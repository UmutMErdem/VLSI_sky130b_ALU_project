* NGSPICE file created from xor3_pex.ext - technology: sky130B

.subckt xor3 C OUT A VDD VSS B
X0 a_338_n478.t9 a_n89_215.t4 a_456_n478.t3 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1 a_692_n1210.t1 A.t0 a_456_n478.t7 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2 a_n89_215.t0 A.t1 VDD.t15 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 a_2236_n478.t11 a_456_n478.t8 VDD.t18 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4 VSS.t2 B.t0 a_692_n1210.t0 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X5 VDD.t1 B.t1 a_338_n478.t1 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X6 a_2648_n504.t3 C.t0 VDD.t4 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7 VDD.t9 C.t1 a_2236_n478.t5 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X8 a_338_n478.t2 B.t2 VDD.t2 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X9 a_2648_n504.t2 C.t2 VDD.t7 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10 VDD.t19 a_456_n478.t9 a_2236_n478.t10 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 a_338_n478.t4 A.t2 VDD.t12 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X12 a_2236_n478.t3 a_1809_215.t4 OUT.t2 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X13 VDD.t3 C.t3 a_2648_n504.t1 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X14 a_2236_n478.t1 a_2648_n504.t4 OUT.t6 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X15 a_456_n1210.t1 a_750_n504.t4 VSS.t4 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X16 VDD.t0 B.t3 a_338_n478.t0 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 a_2236_n478.t9 a_456_n478.t10 VDD.t23 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 a_338_n478.t10 a_750_n504.t5 a_456_n478.t6 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_750_n504.t0 B.t4 VSS.t3 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X20 VDD.t11 A.t3 a_338_n478.t5 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X21 a_338_n478.t3 a_750_n504.t6 a_456_n478.t0 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X22 VSS.t5 A.t4 a_n89_215.t2 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X23 a_338_n478.t11 A.t5 VDD.t10 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X24 OUT.t3 a_1809_215.t5 a_2354_n1210.t0 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X25 VDD.t20 a_456_n478.t11 a_1809_215.t3 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 a_2590_n1210.t1 a_456_n478.t12 OUT.t7 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X27 VDD.t14 A.t6 a_n89_215.t1 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 a_456_n478.t4 a_n89_215.t5 a_338_n478.t8 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X29 a_750_n504.t3 B.t5 VDD.t16 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X30 a_2236_n478.t7 a_2648_n504.t5 OUT.t5 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X31 a_750_n504.t2 B.t6 VDD.t5 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X32 a_456_n478.t2 a_n89_215.t6 a_338_n478.t7 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X33 a_1809_215.t2 a_456_n478.t13 VDD.t21 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X34 VDD.t13 A.t7 a_n89_215.t3 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X35 a_456_n478.t1 a_750_n504.t7 a_338_n478.t6 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X36 VDD.t6 B.t7 a_750_n504.t1 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X37 VDD.t17 C.t4 a_2236_n478.t8 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X38 OUT.t1 a_1809_215.t6 a_2236_n478.t2 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 VSS.t7 a_456_n478.t14 a_1809_215.t0 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X40 VSS.t1 C.t5 a_2590_n1210.t0 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X41 VDD.t22 a_456_n478.t15 a_1809_215.t1 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X42 OUT.t0 a_1809_215.t7 a_2236_n478.t6 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X43 a_2354_n1210.t1 a_2648_n504.t6 VSS.t0 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X44 a_2236_n478.t4 C.t6 VDD.t8 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X45 OUT.t4 a_2648_n504.t7 a_2236_n478.t0 w_n125_153# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X46 a_456_n478.t5 a_n89_215.t7 a_456_n1210.t0 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X47 a_2648_n504.t0 C.t7 VSS.t6 a_647_n1695# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 a_n89_215.n1 a_n89_215.t4 318.922
R1 a_n89_215.n0 a_n89_215.t5 273.935
R2 a_n89_215.n0 a_n89_215.t6 273.935
R3 a_n89_215.n1 a_n89_215.t7 269.116
R4 a_n89_215.n4 a_n89_215.n3 193.227
R5 a_n89_215.t4 a_n89_215.n0 179.142
R6 a_n89_215.n2 a_n89_215.n1 106.999
R7 a_n89_215.n3 a_n89_215.t1 28.568
R8 a_n89_215.n4 a_n89_215.t3 28.565
R9 a_n89_215.t0 a_n89_215.n4 28.565
R10 a_n89_215.n2 a_n89_215.t2 18.149
R11 a_n89_215.n3 a_n89_215.n2 3.726
R12 a_456_n478.n0 a_456_n478.t1 14.282
R13 a_456_n478.t0 a_456_n478.n0 14.282
R14 a_456_n478.n0 a_456_n478.n12 90.436
R15 a_456_n478.n8 a_456_n478.n11 50.575
R16 a_456_n478.n12 a_456_n478.n8 74.302
R17 a_456_n478.n11 a_456_n478.n10 157.665
R18 a_456_n478.n10 a_456_n478.t5 8.7
R19 a_456_n478.n10 a_456_n478.t7 8.7
R20 a_456_n478.n11 a_456_n478.n9 122.999
R21 a_456_n478.n9 a_456_n478.t4 14.282
R22 a_456_n478.n9 a_456_n478.t3 14.282
R23 a_456_n478.n8 a_456_n478.n7 90.416
R24 a_456_n478.n7 a_456_n478.t2 14.282
R25 a_456_n478.n7 a_456_n478.t6 14.282
R26 a_456_n478.n12 a_456_n478.n1 342.688
R27 a_456_n478.n1 a_456_n478.n6 126.566
R28 a_456_n478.n6 a_456_n478.t12 294.653
R29 a_456_n478.n6 a_456_n478.t14 111.663
R30 a_456_n478.n1 a_456_n478.n5 552.333
R31 a_456_n478.n5 a_456_n478.n4 6.615
R32 a_456_n478.n4 a_456_n478.t13 93.989
R33 a_456_n478.n5 a_456_n478.n3 97.816
R34 a_456_n478.n3 a_456_n478.t11 80.333
R35 a_456_n478.n3 a_456_n478.t10 394.151
R36 a_456_n478.t10 a_456_n478.n2 269.523
R37 a_456_n478.n2 a_456_n478.t9 160.666
R38 a_456_n478.n2 a_456_n478.t8 269.523
R39 a_456_n478.n4 a_456_n478.t15 198.043
R40 a_338_n478.n0 a_338_n478.n1 0.001
R41 a_338_n478.n0 a_338_n478.t4 14.282
R42 a_338_n478.t0 a_338_n478.n0 14.282
R43 a_338_n478.n1 a_338_n478.n9 267.767
R44 a_338_n478.n9 a_338_n478.t2 14.282
R45 a_338_n478.n9 a_338_n478.t1 14.282
R46 a_338_n478.n1 a_338_n478.n7 0.669
R47 a_338_n478.n7 a_338_n478.n8 1.511
R48 a_338_n478.n8 a_338_n478.t11 14.282
R49 a_338_n478.n8 a_338_n478.t5 14.282
R50 a_338_n478.n7 a_338_n478.n6 0.227
R51 a_338_n478.n6 a_338_n478.n3 0.575
R52 a_338_n478.n6 a_338_n478.n5 0.2
R53 a_338_n478.n5 a_338_n478.t3 16.058
R54 a_338_n478.n5 a_338_n478.n4 0.999
R55 a_338_n478.n4 a_338_n478.t10 14.282
R56 a_338_n478.n4 a_338_n478.t6 14.282
R57 a_338_n478.n3 a_338_n478.n2 0.999
R58 a_338_n478.n2 a_338_n478.t9 14.282
R59 a_338_n478.n2 a_338_n478.t7 14.282
R60 a_338_n478.n3 a_338_n478.t8 16.058
R61 A A.n4 566.312
R62 A.n1 A.t5 394.151
R63 A.n4 A.t0 294.653
R64 A.n0 A.t2 269.523
R65 A.t5 A.n0 269.523
R66 A.n2 A.t6 198.043
R67 A.n0 A.t3 160.666
R68 A.n4 A.t4 111.663
R69 A.n3 A.n1 97.816
R70 A.n2 A.t1 93.989
R71 A.n1 A.t7 80.333
R72 A A.n3 72.344
R73 A.n3 A.n2 6.615
R74 a_692_n1210.t0 a_692_n1210.t1 17.4
R75 VDD.n12 VDD.t13 28.664
R76 VDD.n17 VDD.t5 28.664
R77 VDD.n1 VDD.t20 28.664
R78 VDD.n6 VDD.t7 28.664
R79 VDD.n13 VDD.t15 28.565
R80 VDD.n13 VDD.t14 28.565
R81 VDD.n18 VDD.t16 28.565
R82 VDD.n18 VDD.t6 28.565
R83 VDD.n2 VDD.t21 28.565
R84 VDD.n2 VDD.t22 28.565
R85 VDD.n7 VDD.t4 28.565
R86 VDD.n7 VDD.t3 28.565
R87 VDD.n12 VDD.t10 14.284
R88 VDD.n17 VDD.t1 14.284
R89 VDD.n1 VDD.t23 14.284
R90 VDD.n6 VDD.t17 14.284
R91 VDD.n11 VDD.t12 14.282
R92 VDD.n11 VDD.t11 14.282
R93 VDD.n16 VDD.t2 14.282
R94 VDD.n16 VDD.t0 14.282
R95 VDD.n0 VDD.t18 14.282
R96 VDD.n0 VDD.t19 14.282
R97 VDD.n5 VDD.t8 14.282
R98 VDD.n5 VDD.t9 14.282
R99 VDD.n21 VDD.n15 4.276
R100 VDD.n10 VDD.n4 4.276
R101 VDD.n14 VDD.n13 2.451
R102 VDD.n3 VDD.n2 2.451
R103 VDD.n19 VDD.n18 2.449
R104 VDD.n8 VDD.n7 2.449
R105 VDD.n15 VDD.n11 0.922
R106 VDD.n20 VDD.n16 0.922
R107 VDD.n4 VDD.n0 0.922
R108 VDD.n9 VDD.n5 0.922
R109 VDD.n14 VDD.n12 0.921
R110 VDD.n19 VDD.n17 0.921
R111 VDD.n3 VDD.n1 0.921
R112 VDD.n8 VDD.n6 0.921
R113 VDD VDD.n10 0.721
R114 VDD.n15 VDD.n14 0.686
R115 VDD.n20 VDD.n19 0.686
R116 VDD.n4 VDD.n3 0.686
R117 VDD.n9 VDD.n8 0.686
R118 VDD VDD.n21 0.27
R119 VDD.n21 VDD.n20 0.179
R120 VDD.n10 VDD.n9 0.179
R121 a_2236_n478.n0 a_2236_n478.t1 14.282
R122 a_2236_n478.t0 a_2236_n478.n0 14.282
R123 a_2236_n478.n0 a_2236_n478.n9 0.999
R124 a_2236_n478.n6 a_2236_n478.n8 0.575
R125 a_2236_n478.n9 a_2236_n478.n6 0.2
R126 a_2236_n478.n9 a_2236_n478.t7 16.058
R127 a_2236_n478.n8 a_2236_n478.n7 0.999
R128 a_2236_n478.n7 a_2236_n478.t3 14.282
R129 a_2236_n478.n7 a_2236_n478.t6 14.282
R130 a_2236_n478.n8 a_2236_n478.t2 16.058
R131 a_2236_n478.n6 a_2236_n478.n4 0.227
R132 a_2236_n478.n4 a_2236_n478.n5 1.511
R133 a_2236_n478.n5 a_2236_n478.t9 14.282
R134 a_2236_n478.n5 a_2236_n478.t10 14.282
R135 a_2236_n478.n4 a_2236_n478.n1 0.669
R136 a_2236_n478.n1 a_2236_n478.n2 0.001
R137 a_2236_n478.n1 a_2236_n478.n3 267.767
R138 a_2236_n478.n3 a_2236_n478.t4 14.282
R139 a_2236_n478.n3 a_2236_n478.t8 14.282
R140 a_2236_n478.n2 a_2236_n478.t11 14.282
R141 a_2236_n478.n2 a_2236_n478.t5 14.282
R142 B B.n3 567.558
R143 B.t6 B.n1 313.873
R144 B.n3 B.t0 294.986
R145 B.n0 B.t3 272.288
R146 B.n2 B.t6 190.152
R147 B.n2 B.t5 190.152
R148 B B.t7 183.395
R149 B.n0 B.t2 160.666
R150 B.n1 B.t1 160.666
R151 B.n3 B.t4 110.859
R152 B.n1 B.n0 96.129
R153 B.t7 B.n2 80.333
R154 VSS.n4 VSS.t3 20.763
R155 VSS.n1 VSS.t6 20.763
R156 VSS.n5 VSS.t5 20.606
R157 VSS.n2 VSS.t7 20.606
R158 VSS.n3 VSS.t4 8.7
R159 VSS.n3 VSS.t2 8.7
R160 VSS.n0 VSS.t0 8.7
R161 VSS.n0 VSS.t1 8.7
R162 VSS.n4 VSS.n3 0.948
R163 VSS.n1 VSS.n0 0.948
R164 VSS VSS.n2 0.389
R165 VSS VSS.n5 0.232
R166 VSS.n5 VSS.n4 0.125
R167 VSS.n2 VSS.n1 0.125
R168 C C.n3 567.558
R169 C.t2 C.n1 313.873
R170 C.n3 C.t5 294.986
R171 C.n0 C.t1 272.288
R172 C.n2 C.t2 190.152
R173 C.n2 C.t0 190.152
R174 C C.t3 183.395
R175 C.n0 C.t6 160.666
R176 C.n1 C.t4 160.666
R177 C.n3 C.t7 110.859
R178 C.n1 C.n0 96.129
R179 C.t3 C.n2 80.333
R180 a_2648_n504.n1 a_2648_n504.t7 318.922
R181 a_2648_n504.n0 a_2648_n504.t4 274.739
R182 a_2648_n504.n0 a_2648_n504.t5 274.739
R183 a_2648_n504.n1 a_2648_n504.t6 269.116
R184 a_2648_n504.t7 a_2648_n504.n0 179.946
R185 a_2648_n504.n2 a_2648_n504.n1 107.263
R186 a_2648_n504.t3 a_2648_n504.n4 29.444
R187 a_2648_n504.n3 a_2648_n504.t1 28.565
R188 a_2648_n504.n3 a_2648_n504.t2 28.565
R189 a_2648_n504.n2 a_2648_n504.t0 18.145
R190 a_2648_n504.n4 a_2648_n504.n2 2.878
R191 a_2648_n504.n4 a_2648_n504.n3 0.764
R192 a_1809_215.n1 a_1809_215.t4 318.922
R193 a_1809_215.n0 a_1809_215.t6 273.935
R194 a_1809_215.n0 a_1809_215.t7 273.935
R195 a_1809_215.n1 a_1809_215.t5 269.116
R196 a_1809_215.n4 a_1809_215.n3 193.227
R197 a_1809_215.t4 a_1809_215.n0 179.142
R198 a_1809_215.n2 a_1809_215.n1 106.999
R199 a_1809_215.n3 a_1809_215.t1 28.568
R200 a_1809_215.t3 a_1809_215.n4 28.565
R201 a_1809_215.n4 a_1809_215.t2 28.565
R202 a_1809_215.n2 a_1809_215.t0 18.149
R203 a_1809_215.n3 a_1809_215.n2 3.726
R204 OUT.n7 OUT.n6 188.878
R205 OUT.n4 OUT.n2 157.665
R206 OUT.n4 OUT.n3 122.999
R207 OUT.n6 OUT.n0 90.436
R208 OUT.n5 OUT.n1 90.416
R209 OUT.n6 OUT.n5 74.302
R210 OUT.n5 OUT.n4 50.575
R211 OUT.n0 OUT.t5 14.282
R212 OUT.n0 OUT.t4 14.282
R213 OUT.n1 OUT.t6 14.282
R214 OUT.n1 OUT.t0 14.282
R215 OUT.n3 OUT.t2 14.282
R216 OUT.n3 OUT.t1 14.282
R217 OUT.n2 OUT.t7 8.7
R218 OUT.n2 OUT.t3 8.7
R219 OUT OUT.n7 5.504
R220 OUT.n7 OUT 5.248
R221 a_750_n504.n1 a_750_n504.t7 318.922
R222 a_750_n504.n0 a_750_n504.t5 274.739
R223 a_750_n504.n0 a_750_n504.t6 274.739
R224 a_750_n504.n1 a_750_n504.t4 269.116
R225 a_750_n504.t7 a_750_n504.n0 179.946
R226 a_750_n504.n2 a_750_n504.n1 107.263
R227 a_750_n504.t3 a_750_n504.n4 29.444
R228 a_750_n504.n3 a_750_n504.t1 28.565
R229 a_750_n504.n3 a_750_n504.t2 28.565
R230 a_750_n504.n2 a_750_n504.t0 18.145
R231 a_750_n504.n4 a_750_n504.n2 2.878
R232 a_750_n504.n4 a_750_n504.n3 0.764
R233 a_456_n1210.t0 a_456_n1210.t1 380.209
R234 a_2354_n1210.t0 a_2354_n1210.t1 380.209
R235 a_2590_n1210.t0 a_2590_n1210.t1 17.4
C0 OUT w_n125_153# 0.15fF
C1 B VSS 0.20fF
C2 VSS A 0.10fF
C3 VDD OUT 0.07fF
C4 B C 0.00fF
C5 w_n125_153# VSS 0.10fF
C6 B A 0.12fF
C7 VDD VSS 0.00fF
C8 C w_n125_153# 0.36fF
C9 B w_n125_153# 0.38fF
C10 w_n125_153# A 0.37fF
C11 VDD C 0.11fF
C12 VDD B 0.15fF
C13 VDD A 0.11fF
C14 OUT VSS 0.11fF
C15 VDD w_n125_153# 0.86fF
C16 OUT C 0.10fF
C17 OUT B 0.01fF
C18 C VSS 0.19fF
C19 VSS a_647_n1695# 2.91fF
C20 OUT a_647_n1695# 0.26fF
C21 VDD a_647_n1695# 3.12fF
C22 C a_647_n1695# 1.30fF
C23 B a_647_n1695# 1.12fF
C24 A a_647_n1695# 1.21fF
C25 w_n125_153# a_647_n1695# 8.59fF
C26 OUT.t5 a_647_n1695# 0.05fF
C27 OUT.t4 a_647_n1695# 0.05fF
C28 OUT.n0 a_647_n1695# 0.33fF $ **FLOATING
C29 OUT.t6 a_647_n1695# 0.05fF
C30 OUT.t0 a_647_n1695# 0.05fF
C31 OUT.n1 a_647_n1695# 0.33fF $ **FLOATING
C32 OUT.t7 a_647_n1695# 0.05fF
C33 OUT.t3 a_647_n1695# 0.05fF
C34 OUT.n2 a_647_n1695# 0.37fF $ **FLOATING
C35 OUT.t2 a_647_n1695# 0.05fF
C36 OUT.t1 a_647_n1695# 0.05fF
C37 OUT.n3 a_647_n1695# 0.33fF $ **FLOATING
C38 OUT.n4 a_647_n1695# 0.15fF $ **FLOATING
C39 OUT.n5 a_647_n1695# 0.10fF $ **FLOATING
C40 OUT.n6 a_647_n1695# 0.17fF $ **FLOATING
C41 OUT.n7 a_647_n1695# 0.13fF $ **FLOATING
C42 VSS.t7 a_647_n1695# 0.02fF
C43 VSS.t6 a_647_n1695# 0.02fF
C44 VSS.t0 a_647_n1695# 0.01fF
C45 VSS.t1 a_647_n1695# 0.01fF
C46 VSS.n0 a_647_n1695# 0.09fF $ **FLOATING
C47 VSS.n1 a_647_n1695# 0.11fF $ **FLOATING
C48 VSS.n2 a_647_n1695# 0.37fF $ **FLOATING
C49 VSS.t5 a_647_n1695# 0.02fF
C50 VSS.t3 a_647_n1695# 0.02fF
C51 VSS.t4 a_647_n1695# 0.01fF
C52 VSS.t2 a_647_n1695# 0.01fF
C53 VSS.n3 a_647_n1695# 0.09fF $ **FLOATING
C54 VSS.n4 a_647_n1695# 0.11fF $ **FLOATING
C55 VSS.n5 a_647_n1695# 0.25fF $ **FLOATING
C56 a_2236_n478.t0 a_647_n1695# 0.06fF
C57 a_2236_n478.n0 a_647_n1695# 0.45fF $ **FLOATING
C58 a_2236_n478.n1 a_647_n1695# 0.37fF $ **FLOATING
C59 a_2236_n478.n2 a_647_n1695# 0.12fF $ **FLOATING
C60 a_2236_n478.t11 a_647_n1695# 0.06fF
C61 a_2236_n478.t5 a_647_n1695# 0.06fF
C62 a_2236_n478.n3 a_647_n1695# 0.53fF $ **FLOATING
C63 a_2236_n478.t4 a_647_n1695# 0.06fF
C64 a_2236_n478.t8 a_647_n1695# 0.06fF
C65 a_2236_n478.n4 a_647_n1695# 0.16fF $ **FLOATING
C66 a_2236_n478.n5 a_647_n1695# 0.48fF $ **FLOATING
C67 a_2236_n478.t9 a_647_n1695# 0.06fF
C68 a_2236_n478.t10 a_647_n1695# 0.06fF
C69 a_2236_n478.n6 a_647_n1695# 0.06fF $ **FLOATING
C70 a_2236_n478.t2 a_647_n1695# 0.12fF
C71 a_2236_n478.n7 a_647_n1695# 0.45fF $ **FLOATING
C72 a_2236_n478.t3 a_647_n1695# 0.06fF
C73 a_2236_n478.t6 a_647_n1695# 0.06fF
C74 a_2236_n478.n8 a_647_n1695# 0.71fF $ **FLOATING
C75 a_2236_n478.t7 a_647_n1695# 0.12fF
C76 a_2236_n478.n9 a_647_n1695# 0.68fF $ **FLOATING
C77 a_2236_n478.t1 a_647_n1695# 0.06fF
C78 VDD.t18 a_647_n1695# 0.02fF
C79 VDD.t19 a_647_n1695# 0.02fF
C80 VDD.n0 a_647_n1695# 0.13fF $ **FLOATING
C81 VDD.t23 a_647_n1695# 0.02fF
C82 VDD.t20 a_647_n1695# 0.01fF
C83 VDD.n1 a_647_n1695# 0.26fF $ **FLOATING
C84 VDD.t21 a_647_n1695# 0.01fF
C85 VDD.t22 a_647_n1695# 0.01fF
C86 VDD.n2 a_647_n1695# 0.10fF $ **FLOATING
C87 VDD.n3 a_647_n1695# 0.09fF $ **FLOATING
C88 VDD.n4 a_647_n1695# 0.04fF $ **FLOATING
C89 VDD.t8 a_647_n1695# 0.02fF
C90 VDD.t9 a_647_n1695# 0.02fF
C91 VDD.n5 a_647_n1695# 0.13fF $ **FLOATING
C92 VDD.t17 a_647_n1695# 0.02fF
C93 VDD.t7 a_647_n1695# 0.01fF
C94 VDD.n6 a_647_n1695# 0.26fF $ **FLOATING
C95 VDD.t4 a_647_n1695# 0.01fF
C96 VDD.t3 a_647_n1695# 0.01fF
C97 VDD.n7 a_647_n1695# 0.10fF $ **FLOATING
C98 VDD.n8 a_647_n1695# 0.08fF $ **FLOATING
C99 VDD.n9 a_647_n1695# 0.04fF $ **FLOATING
C100 VDD.n10 a_647_n1695# 0.50fF $ **FLOATING
C101 VDD.t12 a_647_n1695# 0.02fF
C102 VDD.t11 a_647_n1695# 0.02fF
C103 VDD.n11 a_647_n1695# 0.13fF $ **FLOATING
C104 VDD.t10 a_647_n1695# 0.02fF
C105 VDD.t13 a_647_n1695# 0.01fF
C106 VDD.n12 a_647_n1695# 0.26fF $ **FLOATING
C107 VDD.t15 a_647_n1695# 0.01fF
C108 VDD.t14 a_647_n1695# 0.01fF
C109 VDD.n13 a_647_n1695# 0.10fF $ **FLOATING
C110 VDD.n14 a_647_n1695# 0.09fF $ **FLOATING
C111 VDD.n15 a_647_n1695# 0.04fF $ **FLOATING
C112 VDD.t2 a_647_n1695# 0.02fF
C113 VDD.t0 a_647_n1695# 0.02fF
C114 VDD.n16 a_647_n1695# 0.13fF $ **FLOATING
C115 VDD.t1 a_647_n1695# 0.02fF
C116 VDD.t5 a_647_n1695# 0.01fF
C117 VDD.n17 a_647_n1695# 0.26fF $ **FLOATING
C118 VDD.t16 a_647_n1695# 0.01fF
C119 VDD.t6 a_647_n1695# 0.01fF
C120 VDD.n18 a_647_n1695# 0.10fF $ **FLOATING
C121 VDD.n19 a_647_n1695# 0.08fF $ **FLOATING
C122 VDD.n20 a_647_n1695# 0.04fF $ **FLOATING
C123 VDD.n21 a_647_n1695# 0.28fF $ **FLOATING
C124 a_338_n478.t0 a_647_n1695# 0.06fF
C125 a_338_n478.n0 a_647_n1695# 0.12fF $ **FLOATING
C126 a_338_n478.n1 a_647_n1695# 0.37fF $ **FLOATING
C127 a_338_n478.t8 a_647_n1695# 0.12fF
C128 a_338_n478.n2 a_647_n1695# 0.45fF $ **FLOATING
C129 a_338_n478.t9 a_647_n1695# 0.06fF
C130 a_338_n478.t7 a_647_n1695# 0.06fF
C131 a_338_n478.n3 a_647_n1695# 0.71fF $ **FLOATING
C132 a_338_n478.n4 a_647_n1695# 0.45fF $ **FLOATING
C133 a_338_n478.t10 a_647_n1695# 0.06fF
C134 a_338_n478.t6 a_647_n1695# 0.06fF
C135 a_338_n478.n5 a_647_n1695# 0.68fF $ **FLOATING
C136 a_338_n478.t3 a_647_n1695# 0.12fF
C137 a_338_n478.n6 a_647_n1695# 0.06fF $ **FLOATING
C138 a_338_n478.n7 a_647_n1695# 0.16fF $ **FLOATING
C139 a_338_n478.n8 a_647_n1695# 0.48fF $ **FLOATING
C140 a_338_n478.t11 a_647_n1695# 0.06fF
C141 a_338_n478.t5 a_647_n1695# 0.06fF
C142 a_338_n478.n9 a_647_n1695# 0.53fF $ **FLOATING
C143 a_338_n478.t2 a_647_n1695# 0.06fF
C144 a_338_n478.t1 a_647_n1695# 0.06fF
C145 a_338_n478.t4 a_647_n1695# 0.06fF
C146 a_456_n478.t0 a_647_n1695# 0.02fF
C147 a_456_n478.n0 a_647_n1695# 0.16fF $ **FLOATING
C148 a_456_n478.n1 a_647_n1695# 0.23fF $ **FLOATING
C149 a_456_n478.t15 a_647_n1695# 0.05fF
C150 a_456_n478.t10 a_647_n1695# 0.10fF
C151 a_456_n478.t8 a_647_n1695# 0.08fF
C152 a_456_n478.t9 a_647_n1695# 0.06fF
C153 a_456_n478.n2 a_647_n1695# 0.11fF $ **FLOATING
C154 a_456_n478.t11 a_647_n1695# 0.03fF
C155 a_456_n478.n3 a_647_n1695# 0.08fF $ **FLOATING
C156 a_456_n478.t13 a_647_n1695# 0.03fF
C157 a_456_n478.n4 a_647_n1695# 0.04fF $ **FLOATING
C158 a_456_n478.n5 a_647_n1695# 0.09fF $ **FLOATING
C159 a_456_n478.t14 a_647_n1695# 0.03fF
C160 a_456_n478.n6 a_647_n1695# 0.18fF $ **FLOATING
C161 a_456_n478.t12 a_647_n1695# 0.12fF
C162 a_456_n478.n7 a_647_n1695# 0.16fF $ **FLOATING
C163 a_456_n478.t2 a_647_n1695# 0.02fF
C164 a_456_n478.t6 a_647_n1695# 0.02fF
C165 a_456_n478.n8 a_647_n1695# 0.05fF $ **FLOATING
C166 a_456_n478.n9 a_647_n1695# 0.16fF $ **FLOATING
C167 a_456_n478.t4 a_647_n1695# 0.02fF
C168 a_456_n478.t3 a_647_n1695# 0.02fF
C169 a_456_n478.n10 a_647_n1695# 0.18fF $ **FLOATING
C170 a_456_n478.t5 a_647_n1695# 0.02fF
C171 a_456_n478.t7 a_647_n1695# 0.02fF
C172 a_456_n478.n11 a_647_n1695# 0.07fF $ **FLOATING
C173 a_456_n478.n12 a_647_n1695# 0.15fF $ **FLOATING
C174 a_456_n478.t1 a_647_n1695# 0.02fF
.ends

