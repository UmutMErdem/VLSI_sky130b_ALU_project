magic
tech sky130B
magscale 1 2
timestamp 1736713522
<< nwell >>
rect 6634 5705 7826 5951
rect 6634 5693 7827 5705
rect 6635 5381 7827 5693
rect 13183 5704 14375 5950
rect 19837 5725 21029 5971
rect 19837 5713 21030 5725
rect 13183 5692 14376 5704
rect 13184 5380 14376 5692
rect 19838 5401 21030 5713
rect 28490 5558 29682 5804
rect 28490 5546 29683 5558
rect 28491 5234 29683 5546
rect 30945 5396 31442 5853
rect 30299 5150 33283 5396
rect 30299 4829 33284 5150
rect 30726 4136 31564 4829
rect 32092 4826 33284 4829
rect 12333 4095 12620 4096
rect 13480 4095 13715 4096
rect 25612 4095 25899 4096
rect 26759 4095 26994 4096
rect -30 3805 1162 4051
rect 9851 4041 10091 4042
rect 5784 4007 6071 4008
rect 6931 4007 7166 4008
rect 3302 3953 3542 3954
rect -30 3793 1163 3805
rect -29 3481 1163 3793
rect 3299 3720 3542 3953
rect 3299 3538 3543 3720
rect 5781 3610 6071 4007
rect 6758 3614 7240 4007
rect 9848 3808 10091 4041
rect 9848 3626 10092 3808
rect 12330 3698 12620 4095
rect 13307 3702 13789 4095
rect 23130 4041 23370 4042
rect 18987 4027 19274 4028
rect 20134 4027 20369 4028
rect 16505 3973 16745 3974
rect 2861 3214 4053 3538
rect 5186 3143 6071 3610
rect 5186 3090 6072 3143
rect 6328 3090 7240 3614
rect 9410 3302 10602 3626
rect 11735 3231 12620 3698
rect 11735 3178 12621 3231
rect 12877 3178 13789 3702
rect 16502 3740 16745 3973
rect 16502 3558 16746 3740
rect 18984 3630 19274 4027
rect 19961 3634 20443 4027
rect 16064 3234 17256 3558
rect 11735 3174 12622 3178
rect 5186 3086 6073 3090
rect 5615 2801 6073 3086
rect 6758 2831 7240 3090
rect 12164 2889 12622 3174
rect 13307 2919 13789 3178
rect 18389 3163 19274 3630
rect 18389 3110 19275 3163
rect 19531 3110 20443 3634
rect 23127 3808 23370 4041
rect 23127 3626 23371 3808
rect 25609 3698 25899 4095
rect 26586 3702 27068 4095
rect 22689 3302 23881 3626
rect 25014 3231 25899 3698
rect 25014 3178 25900 3231
rect 26156 3178 27068 3702
rect 25014 3174 25901 3178
rect 18389 3106 19276 3110
rect 5615 2503 6099 2801
rect 6757 2507 7241 2831
rect 12164 2591 12648 2889
rect 13306 2595 13790 2919
rect 18818 2821 19276 3106
rect 19961 2851 20443 3110
rect 25443 2889 25901 3174
rect 26586 2919 27068 3178
rect 28485 2987 29677 3233
rect 28485 2975 29678 2987
rect 18818 2523 19302 2821
rect 19960 2527 20444 2851
rect 25443 2591 25927 2889
rect 26585 2595 27069 2919
rect 28486 2663 29678 2975
rect 9865 2391 10105 2392
rect 23144 2391 23384 2392
rect 3316 2303 3556 2304
rect 3313 2070 3556 2303
rect 9862 2158 10105 2391
rect 16519 2323 16759 2324
rect 3313 1888 3557 2070
rect 9862 1976 10106 2158
rect 16516 2090 16759 2323
rect 23141 2158 23384 2391
rect 2875 1564 4067 1888
rect 7027 1471 7255 1961
rect 9424 1652 10616 1976
rect 13576 1559 13804 2049
rect 16516 1908 16760 2090
rect 16078 1584 17270 1908
rect -38 1220 1154 1466
rect 4338 1271 5661 1471
rect 6721 1271 7559 1471
rect 10887 1359 12210 1559
rect 13270 1359 14108 1559
rect 20230 1491 20458 1981
rect 23141 1976 23385 2158
rect 22703 1652 23895 1976
rect 26855 1559 27083 2049
rect -38 1208 1155 1220
rect -37 896 1155 1208
rect 4338 947 8042 1271
rect 10887 1035 14591 1359
rect 17541 1291 18864 1491
rect 19924 1291 20762 1491
rect 24166 1359 25489 1559
rect 26549 1359 27387 1559
rect 3311 699 3551 700
rect 3308 466 3551 699
rect 3308 284 3552 466
rect 2870 -40 4062 284
rect 4766 254 5604 947
rect 6664 254 7502 947
rect 9860 787 10100 788
rect 9857 554 10100 787
rect 9857 372 10101 554
rect 9419 48 10611 372
rect 11315 342 12153 1035
rect 13213 342 14051 1035
rect 17541 967 21245 1291
rect 24166 1035 27870 1359
rect 30947 1305 31444 1762
rect 30301 1059 33285 1305
rect 16514 719 16754 720
rect 16511 486 16754 719
rect 16511 304 16755 486
rect 16073 -20 17265 304
rect 17969 274 18807 967
rect 19867 274 20705 967
rect 23139 787 23379 788
rect 23136 554 23379 787
rect 23136 372 23380 554
rect 22698 48 23890 372
rect 24594 342 25432 1035
rect 26492 342 27330 1035
rect 30301 738 33286 1059
rect 28485 -46 29677 200
rect 30728 45 31566 738
rect 32094 735 33286 738
rect 28485 -58 29678 -46
rect 28486 -370 29678 -58
rect 5776 -1773 6063 -1772
rect 6923 -1773 7158 -1772
rect 25604 -1773 25891 -1772
rect 26751 -1773 26986 -1772
rect -57 -2058 1135 -1812
rect 3294 -1827 3534 -1826
rect -57 -2070 1136 -2058
rect -56 -2382 1136 -2070
rect 3291 -2060 3534 -1827
rect 3291 -2242 3535 -2060
rect 5773 -2170 6063 -1773
rect 6750 -2166 7232 -1773
rect 18982 -1774 19269 -1773
rect 20129 -1774 20364 -1773
rect 12327 -1775 12614 -1774
rect 13474 -1775 13709 -1774
rect 9845 -1829 10085 -1828
rect 2853 -2566 4045 -2242
rect 5178 -2637 6063 -2170
rect 5178 -2690 6064 -2637
rect 6320 -2690 7232 -2166
rect 9842 -2062 10085 -1829
rect 9842 -2244 10086 -2062
rect 12324 -2172 12614 -1775
rect 13301 -2168 13783 -1775
rect 16500 -1828 16740 -1827
rect 9404 -2568 10596 -2244
rect 5178 -2694 6065 -2690
rect 5607 -2979 6065 -2694
rect 6750 -2949 7232 -2690
rect 11729 -2639 12614 -2172
rect 11729 -2692 12615 -2639
rect 12871 -2692 13783 -2168
rect 16497 -2061 16740 -1828
rect 16497 -2243 16741 -2061
rect 18979 -2171 19269 -1774
rect 19956 -2167 20438 -1774
rect 23122 -1827 23362 -1826
rect 16059 -2567 17251 -2243
rect 11729 -2696 12616 -2692
rect 5607 -3277 6091 -2979
rect 6749 -3273 7233 -2949
rect 12158 -2981 12616 -2696
rect 13301 -2951 13783 -2692
rect 18384 -2638 19269 -2171
rect 18384 -2691 19270 -2638
rect 19526 -2691 20438 -2167
rect 23119 -2060 23362 -1827
rect 23119 -2242 23363 -2060
rect 25601 -2170 25891 -1773
rect 26578 -2166 27060 -1773
rect 28556 -1966 29748 -1720
rect 28556 -1978 29749 -1966
rect 22681 -2566 23873 -2242
rect 18384 -2695 19271 -2691
rect 12158 -3279 12642 -2981
rect 13300 -3275 13784 -2951
rect 18813 -2980 19271 -2695
rect 19956 -2950 20438 -2691
rect 25006 -2637 25891 -2170
rect 25006 -2690 25892 -2637
rect 26148 -2690 27060 -2166
rect 28557 -2290 29749 -1978
rect 30947 -2190 31444 -1733
rect 25006 -2694 25893 -2690
rect 18813 -3278 19297 -2980
rect 19955 -3274 20439 -2950
rect 25435 -2979 25893 -2694
rect 26578 -2949 27060 -2690
rect 30301 -2436 33285 -2190
rect 30301 -2757 33286 -2436
rect 25435 -3277 25919 -2979
rect 26577 -3273 27061 -2949
rect 30728 -3450 31566 -2757
rect 32094 -2760 33286 -2757
rect 3308 -3477 3548 -3476
rect 23136 -3477 23376 -3476
rect 3305 -3710 3548 -3477
rect 16514 -3478 16754 -3477
rect 9859 -3479 10099 -3478
rect 3305 -3892 3549 -3710
rect 9856 -3712 10099 -3479
rect 16511 -3711 16754 -3478
rect 23133 -3710 23376 -3477
rect 2867 -4216 4059 -3892
rect 7019 -4309 7247 -3819
rect 9856 -3894 10100 -3712
rect 9418 -4218 10610 -3894
rect 4330 -4509 5653 -4309
rect 6713 -4509 7551 -4309
rect 13570 -4311 13798 -3821
rect 16511 -3893 16755 -3711
rect 16073 -4217 17265 -3893
rect 20225 -4310 20453 -3820
rect 23133 -3892 23377 -3710
rect 22695 -4216 23887 -3892
rect 26847 -4309 27075 -3819
rect -41 -4818 1151 -4572
rect -41 -4830 1152 -4818
rect -40 -5142 1152 -4830
rect 4330 -4833 8034 -4509
rect 10881 -4511 12204 -4311
rect 13264 -4511 14102 -4311
rect 17536 -4510 18859 -4310
rect 19919 -4510 20757 -4310
rect 24158 -4509 25481 -4309
rect 26541 -4509 27379 -4309
rect 3303 -5081 3543 -5080
rect 3300 -5314 3543 -5081
rect 3300 -5496 3544 -5314
rect 2862 -5820 4054 -5496
rect 4758 -5526 5596 -4833
rect 6656 -5526 7494 -4833
rect 10881 -4835 14585 -4511
rect 17536 -4834 21240 -4510
rect 24158 -4833 27862 -4509
rect 9854 -5083 10094 -5082
rect 9851 -5316 10094 -5083
rect 9851 -5498 10095 -5316
rect 9413 -5822 10605 -5498
rect 11309 -5528 12147 -4835
rect 13207 -5528 14045 -4835
rect 16509 -5082 16749 -5081
rect 16506 -5315 16749 -5082
rect 16506 -5497 16750 -5315
rect 16068 -5821 17260 -5497
rect 17964 -5527 18802 -4834
rect 19862 -5527 20700 -4834
rect 23131 -5081 23371 -5080
rect 23128 -5314 23371 -5081
rect 23128 -5496 23372 -5314
rect 22690 -5820 23882 -5496
rect 24586 -5526 25424 -4833
rect 26484 -5526 27322 -4833
rect 28553 -5036 29745 -4790
rect 28553 -5048 29746 -5036
rect 28554 -5360 29746 -5048
rect 30947 -6538 31444 -6081
rect 30301 -6784 33285 -6538
rect 30301 -7105 33286 -6784
rect 28560 -7881 29752 -7635
rect 30728 -7798 31566 -7105
rect 32094 -7108 33286 -7105
rect 28560 -7893 29753 -7881
rect 6670 -8311 7862 -7999
rect 13224 -8306 14416 -7994
rect 6669 -8323 7862 -8311
rect 13223 -8318 14416 -8306
rect 19873 -8318 21065 -8006
rect 28561 -8205 29753 -7893
rect 6669 -8569 7861 -8323
rect 13223 -8564 14415 -8318
rect 19872 -8330 21065 -8318
rect 19872 -8576 21064 -8330
<< nmos >>
rect 6966 4806 7026 5206
rect 7084 4806 7144 5206
rect 7319 5006 7379 5206
rect 13515 4805 13575 5205
rect 13633 4805 13693 5205
rect 13868 5005 13928 5205
rect 20169 4826 20229 5226
rect 20287 4826 20347 5226
rect 20522 5026 20582 5226
rect 28822 4659 28882 5059
rect 28940 4659 29000 5059
rect 29175 4859 29235 5059
rect 32423 4251 32483 4651
rect 32541 4251 32601 4651
rect 32776 4451 32836 4651
rect 302 2906 362 3306
rect 420 2906 480 3306
rect 655 3106 715 3306
rect 3192 2639 3252 3039
rect 3310 2639 3370 3039
rect 3545 2839 3605 3039
rect 30518 3666 30578 3866
rect 5190 2565 5250 2765
rect 5308 2565 5368 2765
rect 5426 2565 5486 2765
rect 6332 2569 6392 2769
rect 6450 2569 6510 2769
rect 6568 2569 6628 2769
rect 9741 2727 9801 3127
rect 9859 2727 9919 3127
rect 10094 2927 10154 3127
rect 11739 2653 11799 2853
rect 11857 2653 11917 2853
rect 11975 2653 12035 2853
rect 12881 2657 12941 2857
rect 12999 2657 13059 2857
rect 13117 2657 13177 2857
rect 16395 2659 16455 3059
rect 16513 2659 16573 3059
rect 16748 2859 16808 3059
rect 30938 3466 30998 3866
rect 31056 3466 31116 3866
rect 31174 3466 31234 3866
rect 31292 3466 31352 3866
rect 31816 3666 31876 3866
rect 18393 2585 18453 2785
rect 18511 2585 18571 2785
rect 18629 2585 18689 2785
rect 19535 2589 19595 2789
rect 19653 2589 19713 2789
rect 19771 2589 19831 2789
rect 23020 2727 23080 3127
rect 23138 2727 23198 3127
rect 23373 2927 23433 3127
rect 25018 2653 25078 2853
rect 25136 2653 25196 2853
rect 25254 2653 25314 2853
rect 26160 2657 26220 2857
rect 26278 2657 26338 2857
rect 26396 2657 26456 2857
rect 28817 2088 28877 2488
rect 28935 2088 28995 2488
rect 29170 2288 29230 2488
rect 3206 989 3266 1389
rect 3324 989 3384 1389
rect 3559 1189 3619 1389
rect 9755 1077 9815 1477
rect 9873 1077 9933 1477
rect 10108 1277 10168 1477
rect 294 321 354 721
rect 412 321 472 721
rect 647 521 707 721
rect 3201 -615 3261 -215
rect 3319 -615 3379 -215
rect 3554 -415 3614 -215
rect 4558 -216 4618 -16
rect 4978 -416 5038 -16
rect 5096 -416 5156 -16
rect 5214 -416 5274 -16
rect 5332 -416 5392 -16
rect 5856 -216 5916 -16
rect 6456 -216 6516 -16
rect 6876 -416 6936 -16
rect 6994 -416 7054 -16
rect 7112 -416 7172 -16
rect 7230 -416 7290 -16
rect 7754 -216 7814 -16
rect 16409 1009 16469 1409
rect 16527 1009 16587 1409
rect 16762 1209 16822 1409
rect 23034 1077 23094 1477
rect 23152 1077 23212 1477
rect 23387 1277 23447 1477
rect 9750 -527 9810 -127
rect 9868 -527 9928 -127
rect 10103 -327 10163 -127
rect 11107 -128 11167 72
rect 11527 -328 11587 72
rect 11645 -328 11705 72
rect 11763 -328 11823 72
rect 11881 -328 11941 72
rect 12405 -128 12465 72
rect 13005 -128 13065 72
rect 13425 -328 13485 72
rect 13543 -328 13603 72
rect 13661 -328 13721 72
rect 13779 -328 13839 72
rect 14303 -128 14363 72
rect 16404 -595 16464 -195
rect 16522 -595 16582 -195
rect 16757 -395 16817 -195
rect 17761 -196 17821 4
rect 18181 -396 18241 4
rect 18299 -396 18359 4
rect 18417 -396 18477 4
rect 18535 -396 18595 4
rect 19059 -196 19119 4
rect 19659 -196 19719 4
rect 20079 -396 20139 4
rect 20197 -396 20257 4
rect 20315 -396 20375 4
rect 20433 -396 20493 4
rect 20957 -196 21017 4
rect 23029 -527 23089 -127
rect 23147 -527 23207 -127
rect 23382 -327 23442 -127
rect 24386 -128 24446 72
rect 24806 -328 24866 72
rect 24924 -328 24984 72
rect 25042 -328 25102 72
rect 25160 -328 25220 72
rect 25684 -128 25744 72
rect 26284 -128 26344 72
rect 26704 -328 26764 72
rect 26822 -328 26882 72
rect 26940 -328 27000 72
rect 27058 -328 27118 72
rect 27582 -128 27642 72
rect 32425 160 32485 560
rect 32543 160 32603 560
rect 32778 360 32838 560
rect 30520 -425 30580 -225
rect 28817 -945 28877 -545
rect 28935 -945 28995 -545
rect 29170 -745 29230 -545
rect 30940 -625 31000 -225
rect 31058 -625 31118 -225
rect 31176 -625 31236 -225
rect 31294 -625 31354 -225
rect 31818 -425 31878 -225
rect 275 -2957 335 -2557
rect 393 -2957 453 -2557
rect 628 -2757 688 -2557
rect 3184 -3141 3244 -2741
rect 3302 -3141 3362 -2741
rect 3537 -2941 3597 -2741
rect 5182 -3215 5242 -3015
rect 5300 -3215 5360 -3015
rect 5418 -3215 5478 -3015
rect 6324 -3211 6384 -3011
rect 6442 -3211 6502 -3011
rect 6560 -3211 6620 -3011
rect 9735 -3143 9795 -2743
rect 9853 -3143 9913 -2743
rect 10088 -2943 10148 -2743
rect 11733 -3217 11793 -3017
rect 11851 -3217 11911 -3017
rect 11969 -3217 12029 -3017
rect 12875 -3213 12935 -3013
rect 12993 -3213 13053 -3013
rect 13111 -3213 13171 -3013
rect 16390 -3142 16450 -2742
rect 16508 -3142 16568 -2742
rect 16743 -2942 16803 -2742
rect 18388 -3216 18448 -3016
rect 18506 -3216 18566 -3016
rect 18624 -3216 18684 -3016
rect 19530 -3212 19590 -3012
rect 19648 -3212 19708 -3012
rect 19766 -3212 19826 -3012
rect 23012 -3141 23072 -2741
rect 23130 -3141 23190 -2741
rect 23365 -2941 23425 -2741
rect 28888 -2865 28948 -2465
rect 29006 -2865 29066 -2465
rect 29241 -2665 29301 -2465
rect 25010 -3215 25070 -3015
rect 25128 -3215 25188 -3015
rect 25246 -3215 25306 -3015
rect 26152 -3211 26212 -3011
rect 26270 -3211 26330 -3011
rect 26388 -3211 26448 -3011
rect 32425 -3335 32485 -2935
rect 32543 -3335 32603 -2935
rect 32778 -3135 32838 -2935
rect 30520 -3920 30580 -3720
rect 30940 -4120 31000 -3720
rect 31058 -4120 31118 -3720
rect 31176 -4120 31236 -3720
rect 31294 -4120 31354 -3720
rect 31818 -3920 31878 -3720
rect 3198 -4791 3258 -4391
rect 3316 -4791 3376 -4391
rect 3551 -4591 3611 -4391
rect 291 -5717 351 -5317
rect 409 -5717 469 -5317
rect 644 -5517 704 -5317
rect 9749 -4793 9809 -4393
rect 9867 -4793 9927 -4393
rect 10102 -4593 10162 -4393
rect 3193 -6395 3253 -5995
rect 3311 -6395 3371 -5995
rect 3546 -6195 3606 -5995
rect 4550 -5996 4610 -5796
rect 4970 -6196 5030 -5796
rect 5088 -6196 5148 -5796
rect 5206 -6196 5266 -5796
rect 5324 -6196 5384 -5796
rect 5848 -5996 5908 -5796
rect 6448 -5996 6508 -5796
rect 6868 -6196 6928 -5796
rect 6986 -6196 7046 -5796
rect 7104 -6196 7164 -5796
rect 7222 -6196 7282 -5796
rect 7746 -5996 7806 -5796
rect 16404 -4792 16464 -4392
rect 16522 -4792 16582 -4392
rect 16757 -4592 16817 -4392
rect 9744 -6397 9804 -5997
rect 9862 -6397 9922 -5997
rect 10097 -6197 10157 -5997
rect 11101 -5998 11161 -5798
rect 11521 -6198 11581 -5798
rect 11639 -6198 11699 -5798
rect 11757 -6198 11817 -5798
rect 11875 -6198 11935 -5798
rect 12399 -5998 12459 -5798
rect 12999 -5998 13059 -5798
rect 13419 -6198 13479 -5798
rect 13537 -6198 13597 -5798
rect 13655 -6198 13715 -5798
rect 13773 -6198 13833 -5798
rect 14297 -5998 14357 -5798
rect 23026 -4791 23086 -4391
rect 23144 -4791 23204 -4391
rect 23379 -4591 23439 -4391
rect 16399 -6396 16459 -5996
rect 16517 -6396 16577 -5996
rect 16752 -6196 16812 -5996
rect 17756 -5997 17816 -5797
rect 18176 -6197 18236 -5797
rect 18294 -6197 18354 -5797
rect 18412 -6197 18472 -5797
rect 18530 -6197 18590 -5797
rect 19054 -5997 19114 -5797
rect 19654 -5997 19714 -5797
rect 20074 -6197 20134 -5797
rect 20192 -6197 20252 -5797
rect 20310 -6197 20370 -5797
rect 20428 -6197 20488 -5797
rect 20952 -5997 21012 -5797
rect 23021 -6395 23081 -5995
rect 23139 -6395 23199 -5995
rect 23374 -6195 23434 -5995
rect 24378 -5996 24438 -5796
rect 24798 -6196 24858 -5796
rect 24916 -6196 24976 -5796
rect 25034 -6196 25094 -5796
rect 25152 -6196 25212 -5796
rect 25676 -5996 25736 -5796
rect 26276 -5996 26336 -5796
rect 26696 -6196 26756 -5796
rect 26814 -6196 26874 -5796
rect 26932 -6196 26992 -5796
rect 27050 -6196 27110 -5796
rect 27574 -5996 27634 -5796
rect 28885 -5935 28945 -5535
rect 29003 -5935 29063 -5535
rect 29238 -5735 29298 -5535
rect 7001 -7824 7061 -7424
rect 7119 -7824 7179 -7424
rect 7354 -7824 7414 -7624
rect 13555 -7819 13615 -7419
rect 13673 -7819 13733 -7419
rect 13908 -7819 13968 -7619
rect 20204 -7831 20264 -7431
rect 20322 -7831 20382 -7431
rect 20557 -7831 20617 -7631
rect 32425 -7683 32485 -7283
rect 32543 -7683 32603 -7283
rect 32778 -7483 32838 -7283
rect 30520 -8268 30580 -8068
rect 28892 -8780 28952 -8380
rect 29010 -8780 29070 -8380
rect 29245 -8580 29305 -8380
rect 30940 -8468 31000 -8068
rect 31058 -8468 31118 -8068
rect 31176 -8468 31236 -8068
rect 31294 -8468 31354 -8068
rect 31818 -8268 31878 -8068
<< pmos >>
rect 6729 5443 6789 5643
rect 6847 5443 6907 5643
rect 6965 5443 7025 5643
rect 7083 5443 7143 5643
rect 7201 5443 7261 5643
rect 7319 5443 7379 5643
rect 7437 5443 7497 5643
rect 7555 5443 7615 5643
rect 7673 5443 7733 5643
rect 13278 5442 13338 5642
rect 13396 5442 13456 5642
rect 13514 5442 13574 5642
rect 13632 5442 13692 5642
rect 13750 5442 13810 5642
rect 13868 5442 13928 5642
rect 13986 5442 14046 5642
rect 14104 5442 14164 5642
rect 14222 5442 14282 5642
rect 19932 5463 19992 5663
rect 20050 5463 20110 5663
rect 20168 5463 20228 5663
rect 20286 5463 20346 5663
rect 20404 5463 20464 5663
rect 20522 5463 20582 5663
rect 20640 5463 20700 5663
rect 20758 5463 20818 5663
rect 20876 5463 20936 5663
rect 28585 5296 28645 5496
rect 28703 5296 28763 5496
rect 28821 5296 28881 5496
rect 28939 5296 28999 5496
rect 29057 5296 29117 5496
rect 29175 5296 29235 5496
rect 29293 5296 29353 5496
rect 29411 5296 29471 5496
rect 29529 5296 29589 5496
rect 30393 4891 30453 5091
rect 30511 4891 30571 5091
rect 30629 4891 30689 5091
rect 30877 4891 30937 5291
rect 30995 4891 31055 5291
rect 31113 4891 31173 5291
rect 31231 4891 31291 5291
rect 31349 4891 31409 5291
rect 31467 4891 31527 5291
rect 31714 4891 31774 5091
rect 31832 4891 31892 5091
rect 31950 4891 32010 5091
rect 32186 4888 32246 5088
rect 32304 4888 32364 5088
rect 32422 4888 32482 5088
rect 32540 4888 32600 5088
rect 32658 4888 32718 5088
rect 32776 4888 32836 5088
rect 32894 4888 32954 5088
rect 33012 4888 33072 5088
rect 33130 4888 33190 5088
rect 65 3543 125 3743
rect 183 3543 243 3743
rect 301 3543 361 3743
rect 419 3543 479 3743
rect 537 3543 597 3743
rect 655 3543 715 3743
rect 773 3543 833 3743
rect 891 3543 951 3743
rect 1009 3543 1069 3743
rect 30820 4198 30880 4598
rect 30938 4198 30998 4598
rect 31056 4198 31116 4598
rect 31174 4198 31234 4598
rect 31292 4198 31352 4598
rect 31410 4198 31470 4598
rect 2955 3276 3015 3476
rect 3073 3276 3133 3476
rect 3191 3276 3251 3476
rect 3309 3276 3369 3476
rect 3427 3276 3487 3476
rect 3545 3276 3605 3476
rect 3663 3276 3723 3476
rect 3781 3276 3841 3476
rect 3899 3276 3959 3476
rect 5280 3148 5340 3548
rect 5398 3148 5458 3548
rect 5516 3148 5576 3548
rect 5634 3148 5694 3548
rect 5752 3148 5812 3548
rect 5870 3148 5930 3548
rect 6422 3152 6482 3552
rect 6540 3152 6600 3552
rect 6658 3152 6718 3552
rect 6776 3152 6836 3552
rect 6894 3152 6954 3552
rect 7012 3152 7072 3552
rect 9504 3364 9564 3564
rect 9622 3364 9682 3564
rect 9740 3364 9800 3564
rect 9858 3364 9918 3564
rect 9976 3364 10036 3564
rect 10094 3364 10154 3564
rect 10212 3364 10272 3564
rect 10330 3364 10390 3564
rect 10448 3364 10508 3564
rect 11829 3236 11889 3636
rect 11947 3236 12007 3636
rect 12065 3236 12125 3636
rect 12183 3236 12243 3636
rect 12301 3236 12361 3636
rect 12419 3236 12479 3636
rect 12971 3240 13031 3640
rect 13089 3240 13149 3640
rect 13207 3240 13267 3640
rect 13325 3240 13385 3640
rect 13443 3240 13503 3640
rect 13561 3240 13621 3640
rect 16158 3296 16218 3496
rect 16276 3296 16336 3496
rect 16394 3296 16454 3496
rect 16512 3296 16572 3496
rect 16630 3296 16690 3496
rect 16748 3296 16808 3496
rect 16866 3296 16926 3496
rect 16984 3296 17044 3496
rect 17102 3296 17162 3496
rect 5709 2565 5769 2765
rect 5827 2565 5887 2765
rect 5945 2565 6005 2765
rect 6851 2569 6911 2769
rect 6969 2569 7029 2769
rect 7087 2569 7147 2769
rect 18483 3168 18543 3568
rect 18601 3168 18661 3568
rect 18719 3168 18779 3568
rect 18837 3168 18897 3568
rect 18955 3168 19015 3568
rect 19073 3168 19133 3568
rect 19625 3172 19685 3572
rect 19743 3172 19803 3572
rect 19861 3172 19921 3572
rect 19979 3172 20039 3572
rect 20097 3172 20157 3572
rect 20215 3172 20275 3572
rect 22783 3364 22843 3564
rect 22901 3364 22961 3564
rect 23019 3364 23079 3564
rect 23137 3364 23197 3564
rect 23255 3364 23315 3564
rect 23373 3364 23433 3564
rect 23491 3364 23551 3564
rect 23609 3364 23669 3564
rect 23727 3364 23787 3564
rect 12258 2653 12318 2853
rect 12376 2653 12436 2853
rect 12494 2653 12554 2853
rect 13400 2657 13460 2857
rect 13518 2657 13578 2857
rect 13636 2657 13696 2857
rect 25108 3236 25168 3636
rect 25226 3236 25286 3636
rect 25344 3236 25404 3636
rect 25462 3236 25522 3636
rect 25580 3236 25640 3636
rect 25698 3236 25758 3636
rect 26250 3240 26310 3640
rect 26368 3240 26428 3640
rect 26486 3240 26546 3640
rect 26604 3240 26664 3640
rect 26722 3240 26782 3640
rect 26840 3240 26900 3640
rect 18912 2585 18972 2785
rect 19030 2585 19090 2785
rect 19148 2585 19208 2785
rect 20054 2589 20114 2789
rect 20172 2589 20232 2789
rect 20290 2589 20350 2789
rect 25537 2653 25597 2853
rect 25655 2653 25715 2853
rect 25773 2653 25833 2853
rect 26679 2657 26739 2857
rect 26797 2657 26857 2857
rect 26915 2657 26975 2857
rect 28580 2725 28640 2925
rect 28698 2725 28758 2925
rect 28816 2725 28876 2925
rect 28934 2725 28994 2925
rect 29052 2725 29112 2925
rect 29170 2725 29230 2925
rect 29288 2725 29348 2925
rect 29406 2725 29466 2925
rect 29524 2725 29584 2925
rect 2969 1626 3029 1826
rect 3087 1626 3147 1826
rect 3205 1626 3265 1826
rect 3323 1626 3383 1826
rect 3441 1626 3501 1826
rect 3559 1626 3619 1826
rect 3677 1626 3737 1826
rect 3795 1626 3855 1826
rect 3913 1626 3973 1826
rect 9518 1714 9578 1914
rect 9636 1714 9696 1914
rect 9754 1714 9814 1914
rect 9872 1714 9932 1914
rect 9990 1714 10050 1914
rect 10108 1714 10168 1914
rect 10226 1714 10286 1914
rect 10344 1714 10404 1914
rect 10462 1714 10522 1914
rect 16172 1646 16232 1846
rect 16290 1646 16350 1846
rect 16408 1646 16468 1846
rect 16526 1646 16586 1846
rect 16644 1646 16704 1846
rect 16762 1646 16822 1846
rect 16880 1646 16940 1846
rect 16998 1646 17058 1846
rect 17116 1646 17176 1846
rect 22797 1714 22857 1914
rect 22915 1714 22975 1914
rect 23033 1714 23093 1914
rect 23151 1714 23211 1914
rect 23269 1714 23329 1914
rect 23387 1714 23447 1914
rect 23505 1714 23565 1914
rect 23623 1714 23683 1914
rect 23741 1714 23801 1914
rect 57 958 117 1158
rect 175 958 235 1158
rect 293 958 353 1158
rect 411 958 471 1158
rect 529 958 589 1158
rect 647 958 707 1158
rect 765 958 825 1158
rect 883 958 943 1158
rect 1001 958 1061 1158
rect 4433 1009 4493 1209
rect 4551 1009 4611 1209
rect 4669 1009 4729 1209
rect 4917 1009 4977 1409
rect 5035 1009 5095 1409
rect 5153 1009 5213 1409
rect 5271 1009 5331 1409
rect 5389 1009 5449 1409
rect 5507 1009 5567 1409
rect 5754 1009 5814 1209
rect 5872 1009 5932 1209
rect 5990 1009 6050 1209
rect 6331 1009 6391 1209
rect 6449 1009 6509 1209
rect 6567 1009 6627 1209
rect 6815 1009 6875 1409
rect 6933 1009 6993 1409
rect 7051 1009 7111 1409
rect 7169 1009 7229 1409
rect 7287 1009 7347 1409
rect 7405 1009 7465 1409
rect 7652 1009 7712 1209
rect 7770 1009 7830 1209
rect 7888 1009 7948 1209
rect 2964 22 3024 222
rect 3082 22 3142 222
rect 3200 22 3260 222
rect 3318 22 3378 222
rect 3436 22 3496 222
rect 3554 22 3614 222
rect 3672 22 3732 222
rect 3790 22 3850 222
rect 3908 22 3968 222
rect 4860 316 4920 716
rect 4978 316 5038 716
rect 5096 316 5156 716
rect 5214 316 5274 716
rect 5332 316 5392 716
rect 5450 316 5510 716
rect 10982 1097 11042 1297
rect 11100 1097 11160 1297
rect 11218 1097 11278 1297
rect 11466 1097 11526 1497
rect 11584 1097 11644 1497
rect 11702 1097 11762 1497
rect 11820 1097 11880 1497
rect 11938 1097 11998 1497
rect 12056 1097 12116 1497
rect 12303 1097 12363 1297
rect 12421 1097 12481 1297
rect 12539 1097 12599 1297
rect 12880 1097 12940 1297
rect 12998 1097 13058 1297
rect 13116 1097 13176 1297
rect 13364 1097 13424 1497
rect 13482 1097 13542 1497
rect 13600 1097 13660 1497
rect 13718 1097 13778 1497
rect 13836 1097 13896 1497
rect 13954 1097 14014 1497
rect 14201 1097 14261 1297
rect 14319 1097 14379 1297
rect 14437 1097 14497 1297
rect 6758 316 6818 716
rect 6876 316 6936 716
rect 6994 316 7054 716
rect 7112 316 7172 716
rect 7230 316 7290 716
rect 7348 316 7408 716
rect 9513 110 9573 310
rect 9631 110 9691 310
rect 9749 110 9809 310
rect 9867 110 9927 310
rect 9985 110 10045 310
rect 10103 110 10163 310
rect 10221 110 10281 310
rect 10339 110 10399 310
rect 10457 110 10517 310
rect 11409 404 11469 804
rect 11527 404 11587 804
rect 11645 404 11705 804
rect 11763 404 11823 804
rect 11881 404 11941 804
rect 11999 404 12059 804
rect 17636 1029 17696 1229
rect 17754 1029 17814 1229
rect 17872 1029 17932 1229
rect 18120 1029 18180 1429
rect 18238 1029 18298 1429
rect 18356 1029 18416 1429
rect 18474 1029 18534 1429
rect 18592 1029 18652 1429
rect 18710 1029 18770 1429
rect 18957 1029 19017 1229
rect 19075 1029 19135 1229
rect 19193 1029 19253 1229
rect 19534 1029 19594 1229
rect 19652 1029 19712 1229
rect 19770 1029 19830 1229
rect 20018 1029 20078 1429
rect 20136 1029 20196 1429
rect 20254 1029 20314 1429
rect 20372 1029 20432 1429
rect 20490 1029 20550 1429
rect 20608 1029 20668 1429
rect 20855 1029 20915 1229
rect 20973 1029 21033 1229
rect 21091 1029 21151 1229
rect 13307 404 13367 804
rect 13425 404 13485 804
rect 13543 404 13603 804
rect 13661 404 13721 804
rect 13779 404 13839 804
rect 13897 404 13957 804
rect 16167 42 16227 242
rect 16285 42 16345 242
rect 16403 42 16463 242
rect 16521 42 16581 242
rect 16639 42 16699 242
rect 16757 42 16817 242
rect 16875 42 16935 242
rect 16993 42 17053 242
rect 17111 42 17171 242
rect 18063 336 18123 736
rect 18181 336 18241 736
rect 18299 336 18359 736
rect 18417 336 18477 736
rect 18535 336 18595 736
rect 18653 336 18713 736
rect 24261 1097 24321 1297
rect 24379 1097 24439 1297
rect 24497 1097 24557 1297
rect 24745 1097 24805 1497
rect 24863 1097 24923 1497
rect 24981 1097 25041 1497
rect 25099 1097 25159 1497
rect 25217 1097 25277 1497
rect 25335 1097 25395 1497
rect 25582 1097 25642 1297
rect 25700 1097 25760 1297
rect 25818 1097 25878 1297
rect 26159 1097 26219 1297
rect 26277 1097 26337 1297
rect 26395 1097 26455 1297
rect 26643 1097 26703 1497
rect 26761 1097 26821 1497
rect 26879 1097 26939 1497
rect 26997 1097 27057 1497
rect 27115 1097 27175 1497
rect 27233 1097 27293 1497
rect 27480 1097 27540 1297
rect 27598 1097 27658 1297
rect 27716 1097 27776 1297
rect 19961 336 20021 736
rect 20079 336 20139 736
rect 20197 336 20257 736
rect 20315 336 20375 736
rect 20433 336 20493 736
rect 20551 336 20611 736
rect 22792 110 22852 310
rect 22910 110 22970 310
rect 23028 110 23088 310
rect 23146 110 23206 310
rect 23264 110 23324 310
rect 23382 110 23442 310
rect 23500 110 23560 310
rect 23618 110 23678 310
rect 23736 110 23796 310
rect 24688 404 24748 804
rect 24806 404 24866 804
rect 24924 404 24984 804
rect 25042 404 25102 804
rect 25160 404 25220 804
rect 25278 404 25338 804
rect 26586 404 26646 804
rect 26704 404 26764 804
rect 26822 404 26882 804
rect 26940 404 27000 804
rect 27058 404 27118 804
rect 27176 404 27236 804
rect 30395 800 30455 1000
rect 30513 800 30573 1000
rect 30631 800 30691 1000
rect 30879 800 30939 1200
rect 30997 800 31057 1200
rect 31115 800 31175 1200
rect 31233 800 31293 1200
rect 31351 800 31411 1200
rect 31469 800 31529 1200
rect 31716 800 31776 1000
rect 31834 800 31894 1000
rect 31952 800 32012 1000
rect 32188 797 32248 997
rect 32306 797 32366 997
rect 32424 797 32484 997
rect 32542 797 32602 997
rect 32660 797 32720 997
rect 32778 797 32838 997
rect 32896 797 32956 997
rect 33014 797 33074 997
rect 33132 797 33192 997
rect 28580 -308 28640 -108
rect 28698 -308 28758 -108
rect 28816 -308 28876 -108
rect 28934 -308 28994 -108
rect 29052 -308 29112 -108
rect 29170 -308 29230 -108
rect 29288 -308 29348 -108
rect 29406 -308 29466 -108
rect 29524 -308 29584 -108
rect 30822 107 30882 507
rect 30940 107 31000 507
rect 31058 107 31118 507
rect 31176 107 31236 507
rect 31294 107 31354 507
rect 31412 107 31472 507
rect 38 -2320 98 -2120
rect 156 -2320 216 -2120
rect 274 -2320 334 -2120
rect 392 -2320 452 -2120
rect 510 -2320 570 -2120
rect 628 -2320 688 -2120
rect 746 -2320 806 -2120
rect 864 -2320 924 -2120
rect 982 -2320 1042 -2120
rect 2947 -2504 3007 -2304
rect 3065 -2504 3125 -2304
rect 3183 -2504 3243 -2304
rect 3301 -2504 3361 -2304
rect 3419 -2504 3479 -2304
rect 3537 -2504 3597 -2304
rect 3655 -2504 3715 -2304
rect 3773 -2504 3833 -2304
rect 3891 -2504 3951 -2304
rect 5272 -2632 5332 -2232
rect 5390 -2632 5450 -2232
rect 5508 -2632 5568 -2232
rect 5626 -2632 5686 -2232
rect 5744 -2632 5804 -2232
rect 5862 -2632 5922 -2232
rect 6414 -2628 6474 -2228
rect 6532 -2628 6592 -2228
rect 6650 -2628 6710 -2228
rect 6768 -2628 6828 -2228
rect 6886 -2628 6946 -2228
rect 7004 -2628 7064 -2228
rect 9498 -2506 9558 -2306
rect 9616 -2506 9676 -2306
rect 9734 -2506 9794 -2306
rect 9852 -2506 9912 -2306
rect 9970 -2506 10030 -2306
rect 10088 -2506 10148 -2306
rect 10206 -2506 10266 -2306
rect 10324 -2506 10384 -2306
rect 10442 -2506 10502 -2306
rect 11823 -2634 11883 -2234
rect 11941 -2634 12001 -2234
rect 12059 -2634 12119 -2234
rect 12177 -2634 12237 -2234
rect 12295 -2634 12355 -2234
rect 12413 -2634 12473 -2234
rect 12965 -2630 13025 -2230
rect 13083 -2630 13143 -2230
rect 13201 -2630 13261 -2230
rect 13319 -2630 13379 -2230
rect 13437 -2630 13497 -2230
rect 13555 -2630 13615 -2230
rect 16153 -2505 16213 -2305
rect 16271 -2505 16331 -2305
rect 16389 -2505 16449 -2305
rect 16507 -2505 16567 -2305
rect 16625 -2505 16685 -2305
rect 16743 -2505 16803 -2305
rect 16861 -2505 16921 -2305
rect 16979 -2505 17039 -2305
rect 17097 -2505 17157 -2305
rect 5701 -3215 5761 -3015
rect 5819 -3215 5879 -3015
rect 5937 -3215 5997 -3015
rect 6843 -3211 6903 -3011
rect 6961 -3211 7021 -3011
rect 7079 -3211 7139 -3011
rect 18478 -2633 18538 -2233
rect 18596 -2633 18656 -2233
rect 18714 -2633 18774 -2233
rect 18832 -2633 18892 -2233
rect 18950 -2633 19010 -2233
rect 19068 -2633 19128 -2233
rect 19620 -2629 19680 -2229
rect 19738 -2629 19798 -2229
rect 19856 -2629 19916 -2229
rect 19974 -2629 20034 -2229
rect 20092 -2629 20152 -2229
rect 20210 -2629 20270 -2229
rect 28651 -2228 28711 -2028
rect 28769 -2228 28829 -2028
rect 28887 -2228 28947 -2028
rect 29005 -2228 29065 -2028
rect 29123 -2228 29183 -2028
rect 29241 -2228 29301 -2028
rect 29359 -2228 29419 -2028
rect 29477 -2228 29537 -2028
rect 29595 -2228 29655 -2028
rect 22775 -2504 22835 -2304
rect 22893 -2504 22953 -2304
rect 23011 -2504 23071 -2304
rect 23129 -2504 23189 -2304
rect 23247 -2504 23307 -2304
rect 23365 -2504 23425 -2304
rect 23483 -2504 23543 -2304
rect 23601 -2504 23661 -2304
rect 23719 -2504 23779 -2304
rect 12252 -3217 12312 -3017
rect 12370 -3217 12430 -3017
rect 12488 -3217 12548 -3017
rect 13394 -3213 13454 -3013
rect 13512 -3213 13572 -3013
rect 13630 -3213 13690 -3013
rect 25100 -2632 25160 -2232
rect 25218 -2632 25278 -2232
rect 25336 -2632 25396 -2232
rect 25454 -2632 25514 -2232
rect 25572 -2632 25632 -2232
rect 25690 -2632 25750 -2232
rect 26242 -2628 26302 -2228
rect 26360 -2628 26420 -2228
rect 26478 -2628 26538 -2228
rect 26596 -2628 26656 -2228
rect 26714 -2628 26774 -2228
rect 26832 -2628 26892 -2228
rect 18907 -3216 18967 -3016
rect 19025 -3216 19085 -3016
rect 19143 -3216 19203 -3016
rect 20049 -3212 20109 -3012
rect 20167 -3212 20227 -3012
rect 20285 -3212 20345 -3012
rect 30395 -2695 30455 -2495
rect 30513 -2695 30573 -2495
rect 30631 -2695 30691 -2495
rect 30879 -2695 30939 -2295
rect 30997 -2695 31057 -2295
rect 31115 -2695 31175 -2295
rect 31233 -2695 31293 -2295
rect 31351 -2695 31411 -2295
rect 31469 -2695 31529 -2295
rect 31716 -2695 31776 -2495
rect 31834 -2695 31894 -2495
rect 31952 -2695 32012 -2495
rect 32188 -2698 32248 -2498
rect 32306 -2698 32366 -2498
rect 32424 -2698 32484 -2498
rect 32542 -2698 32602 -2498
rect 32660 -2698 32720 -2498
rect 32778 -2698 32838 -2498
rect 32896 -2698 32956 -2498
rect 33014 -2698 33074 -2498
rect 33132 -2698 33192 -2498
rect 25529 -3215 25589 -3015
rect 25647 -3215 25707 -3015
rect 25765 -3215 25825 -3015
rect 26671 -3211 26731 -3011
rect 26789 -3211 26849 -3011
rect 26907 -3211 26967 -3011
rect 30822 -3388 30882 -2988
rect 30940 -3388 31000 -2988
rect 31058 -3388 31118 -2988
rect 31176 -3388 31236 -2988
rect 31294 -3388 31354 -2988
rect 31412 -3388 31472 -2988
rect 2961 -4154 3021 -3954
rect 3079 -4154 3139 -3954
rect 3197 -4154 3257 -3954
rect 3315 -4154 3375 -3954
rect 3433 -4154 3493 -3954
rect 3551 -4154 3611 -3954
rect 3669 -4154 3729 -3954
rect 3787 -4154 3847 -3954
rect 3905 -4154 3965 -3954
rect 9512 -4156 9572 -3956
rect 9630 -4156 9690 -3956
rect 9748 -4156 9808 -3956
rect 9866 -4156 9926 -3956
rect 9984 -4156 10044 -3956
rect 10102 -4156 10162 -3956
rect 10220 -4156 10280 -3956
rect 10338 -4156 10398 -3956
rect 10456 -4156 10516 -3956
rect 16167 -4155 16227 -3955
rect 16285 -4155 16345 -3955
rect 16403 -4155 16463 -3955
rect 16521 -4155 16581 -3955
rect 16639 -4155 16699 -3955
rect 16757 -4155 16817 -3955
rect 16875 -4155 16935 -3955
rect 16993 -4155 17053 -3955
rect 17111 -4155 17171 -3955
rect 22789 -4154 22849 -3954
rect 22907 -4154 22967 -3954
rect 23025 -4154 23085 -3954
rect 23143 -4154 23203 -3954
rect 23261 -4154 23321 -3954
rect 23379 -4154 23439 -3954
rect 23497 -4154 23557 -3954
rect 23615 -4154 23675 -3954
rect 23733 -4154 23793 -3954
rect 4425 -4771 4485 -4571
rect 4543 -4771 4603 -4571
rect 4661 -4771 4721 -4571
rect 4909 -4771 4969 -4371
rect 5027 -4771 5087 -4371
rect 5145 -4771 5205 -4371
rect 5263 -4771 5323 -4371
rect 5381 -4771 5441 -4371
rect 5499 -4771 5559 -4371
rect 5746 -4771 5806 -4571
rect 5864 -4771 5924 -4571
rect 5982 -4771 6042 -4571
rect 6323 -4771 6383 -4571
rect 6441 -4771 6501 -4571
rect 6559 -4771 6619 -4571
rect 6807 -4771 6867 -4371
rect 6925 -4771 6985 -4371
rect 7043 -4771 7103 -4371
rect 7161 -4771 7221 -4371
rect 7279 -4771 7339 -4371
rect 7397 -4771 7457 -4371
rect 7644 -4771 7704 -4571
rect 7762 -4771 7822 -4571
rect 7880 -4771 7940 -4571
rect 54 -5080 114 -4880
rect 172 -5080 232 -4880
rect 290 -5080 350 -4880
rect 408 -5080 468 -4880
rect 526 -5080 586 -4880
rect 644 -5080 704 -4880
rect 762 -5080 822 -4880
rect 880 -5080 940 -4880
rect 998 -5080 1058 -4880
rect 2956 -5758 3016 -5558
rect 3074 -5758 3134 -5558
rect 3192 -5758 3252 -5558
rect 3310 -5758 3370 -5558
rect 3428 -5758 3488 -5558
rect 3546 -5758 3606 -5558
rect 3664 -5758 3724 -5558
rect 3782 -5758 3842 -5558
rect 3900 -5758 3960 -5558
rect 4852 -5464 4912 -5064
rect 4970 -5464 5030 -5064
rect 5088 -5464 5148 -5064
rect 5206 -5464 5266 -5064
rect 5324 -5464 5384 -5064
rect 5442 -5464 5502 -5064
rect 10976 -4773 11036 -4573
rect 11094 -4773 11154 -4573
rect 11212 -4773 11272 -4573
rect 11460 -4773 11520 -4373
rect 11578 -4773 11638 -4373
rect 11696 -4773 11756 -4373
rect 11814 -4773 11874 -4373
rect 11932 -4773 11992 -4373
rect 12050 -4773 12110 -4373
rect 12297 -4773 12357 -4573
rect 12415 -4773 12475 -4573
rect 12533 -4773 12593 -4573
rect 12874 -4773 12934 -4573
rect 12992 -4773 13052 -4573
rect 13110 -4773 13170 -4573
rect 13358 -4773 13418 -4373
rect 13476 -4773 13536 -4373
rect 13594 -4773 13654 -4373
rect 13712 -4773 13772 -4373
rect 13830 -4773 13890 -4373
rect 13948 -4773 14008 -4373
rect 14195 -4773 14255 -4573
rect 14313 -4773 14373 -4573
rect 14431 -4773 14491 -4573
rect 6750 -5464 6810 -5064
rect 6868 -5464 6928 -5064
rect 6986 -5464 7046 -5064
rect 7104 -5464 7164 -5064
rect 7222 -5464 7282 -5064
rect 7340 -5464 7400 -5064
rect 9507 -5760 9567 -5560
rect 9625 -5760 9685 -5560
rect 9743 -5760 9803 -5560
rect 9861 -5760 9921 -5560
rect 9979 -5760 10039 -5560
rect 10097 -5760 10157 -5560
rect 10215 -5760 10275 -5560
rect 10333 -5760 10393 -5560
rect 10451 -5760 10511 -5560
rect 11403 -5466 11463 -5066
rect 11521 -5466 11581 -5066
rect 11639 -5466 11699 -5066
rect 11757 -5466 11817 -5066
rect 11875 -5466 11935 -5066
rect 11993 -5466 12053 -5066
rect 17631 -4772 17691 -4572
rect 17749 -4772 17809 -4572
rect 17867 -4772 17927 -4572
rect 18115 -4772 18175 -4372
rect 18233 -4772 18293 -4372
rect 18351 -4772 18411 -4372
rect 18469 -4772 18529 -4372
rect 18587 -4772 18647 -4372
rect 18705 -4772 18765 -4372
rect 18952 -4772 19012 -4572
rect 19070 -4772 19130 -4572
rect 19188 -4772 19248 -4572
rect 19529 -4772 19589 -4572
rect 19647 -4772 19707 -4572
rect 19765 -4772 19825 -4572
rect 20013 -4772 20073 -4372
rect 20131 -4772 20191 -4372
rect 20249 -4772 20309 -4372
rect 20367 -4772 20427 -4372
rect 20485 -4772 20545 -4372
rect 20603 -4772 20663 -4372
rect 20850 -4772 20910 -4572
rect 20968 -4772 21028 -4572
rect 21086 -4772 21146 -4572
rect 13301 -5466 13361 -5066
rect 13419 -5466 13479 -5066
rect 13537 -5466 13597 -5066
rect 13655 -5466 13715 -5066
rect 13773 -5466 13833 -5066
rect 13891 -5466 13951 -5066
rect 16162 -5759 16222 -5559
rect 16280 -5759 16340 -5559
rect 16398 -5759 16458 -5559
rect 16516 -5759 16576 -5559
rect 16634 -5759 16694 -5559
rect 16752 -5759 16812 -5559
rect 16870 -5759 16930 -5559
rect 16988 -5759 17048 -5559
rect 17106 -5759 17166 -5559
rect 18058 -5465 18118 -5065
rect 18176 -5465 18236 -5065
rect 18294 -5465 18354 -5065
rect 18412 -5465 18472 -5065
rect 18530 -5465 18590 -5065
rect 18648 -5465 18708 -5065
rect 24253 -4771 24313 -4571
rect 24371 -4771 24431 -4571
rect 24489 -4771 24549 -4571
rect 24737 -4771 24797 -4371
rect 24855 -4771 24915 -4371
rect 24973 -4771 25033 -4371
rect 25091 -4771 25151 -4371
rect 25209 -4771 25269 -4371
rect 25327 -4771 25387 -4371
rect 25574 -4771 25634 -4571
rect 25692 -4771 25752 -4571
rect 25810 -4771 25870 -4571
rect 26151 -4771 26211 -4571
rect 26269 -4771 26329 -4571
rect 26387 -4771 26447 -4571
rect 26635 -4771 26695 -4371
rect 26753 -4771 26813 -4371
rect 26871 -4771 26931 -4371
rect 26989 -4771 27049 -4371
rect 27107 -4771 27167 -4371
rect 27225 -4771 27285 -4371
rect 27472 -4771 27532 -4571
rect 27590 -4771 27650 -4571
rect 27708 -4771 27768 -4571
rect 19956 -5465 20016 -5065
rect 20074 -5465 20134 -5065
rect 20192 -5465 20252 -5065
rect 20310 -5465 20370 -5065
rect 20428 -5465 20488 -5065
rect 20546 -5465 20606 -5065
rect 22784 -5758 22844 -5558
rect 22902 -5758 22962 -5558
rect 23020 -5758 23080 -5558
rect 23138 -5758 23198 -5558
rect 23256 -5758 23316 -5558
rect 23374 -5758 23434 -5558
rect 23492 -5758 23552 -5558
rect 23610 -5758 23670 -5558
rect 23728 -5758 23788 -5558
rect 24680 -5464 24740 -5064
rect 24798 -5464 24858 -5064
rect 24916 -5464 24976 -5064
rect 25034 -5464 25094 -5064
rect 25152 -5464 25212 -5064
rect 25270 -5464 25330 -5064
rect 26578 -5464 26638 -5064
rect 26696 -5464 26756 -5064
rect 26814 -5464 26874 -5064
rect 26932 -5464 26992 -5064
rect 27050 -5464 27110 -5064
rect 27168 -5464 27228 -5064
rect 28648 -5298 28708 -5098
rect 28766 -5298 28826 -5098
rect 28884 -5298 28944 -5098
rect 29002 -5298 29062 -5098
rect 29120 -5298 29180 -5098
rect 29238 -5298 29298 -5098
rect 29356 -5298 29416 -5098
rect 29474 -5298 29534 -5098
rect 29592 -5298 29652 -5098
rect 30395 -7043 30455 -6843
rect 30513 -7043 30573 -6843
rect 30631 -7043 30691 -6843
rect 30879 -7043 30939 -6643
rect 30997 -7043 31057 -6643
rect 31115 -7043 31175 -6643
rect 31233 -7043 31293 -6643
rect 31351 -7043 31411 -6643
rect 31469 -7043 31529 -6643
rect 31716 -7043 31776 -6843
rect 31834 -7043 31894 -6843
rect 31952 -7043 32012 -6843
rect 32188 -7046 32248 -6846
rect 32306 -7046 32366 -6846
rect 32424 -7046 32484 -6846
rect 32542 -7046 32602 -6846
rect 32660 -7046 32720 -6846
rect 32778 -7046 32838 -6846
rect 32896 -7046 32956 -6846
rect 33014 -7046 33074 -6846
rect 33132 -7046 33192 -6846
rect 6764 -8261 6824 -8061
rect 6882 -8261 6942 -8061
rect 7000 -8261 7060 -8061
rect 7118 -8261 7178 -8061
rect 7236 -8261 7296 -8061
rect 7354 -8261 7414 -8061
rect 7472 -8261 7532 -8061
rect 7590 -8261 7650 -8061
rect 7708 -8261 7768 -8061
rect 13318 -8256 13378 -8056
rect 13436 -8256 13496 -8056
rect 13554 -8256 13614 -8056
rect 13672 -8256 13732 -8056
rect 13790 -8256 13850 -8056
rect 13908 -8256 13968 -8056
rect 14026 -8256 14086 -8056
rect 14144 -8256 14204 -8056
rect 14262 -8256 14322 -8056
rect 19967 -8268 20027 -8068
rect 20085 -8268 20145 -8068
rect 20203 -8268 20263 -8068
rect 20321 -8268 20381 -8068
rect 20439 -8268 20499 -8068
rect 20557 -8268 20617 -8068
rect 20675 -8268 20735 -8068
rect 20793 -8268 20853 -8068
rect 20911 -8268 20971 -8068
rect 28655 -8143 28715 -7943
rect 28773 -8143 28833 -7943
rect 28891 -8143 28951 -7943
rect 29009 -8143 29069 -7943
rect 29127 -8143 29187 -7943
rect 29245 -8143 29305 -7943
rect 29363 -8143 29423 -7943
rect 29481 -8143 29541 -7943
rect 29599 -8143 29659 -7943
rect 30822 -7736 30882 -7336
rect 30940 -7736 31000 -7336
rect 31058 -7736 31118 -7336
rect 31176 -7736 31236 -7336
rect 31294 -7736 31354 -7336
rect 31412 -7736 31472 -7336
<< ndiff >>
rect 6908 5194 6966 5206
rect 6908 4818 6920 5194
rect 6954 4818 6966 5194
rect 6908 4806 6966 4818
rect 7026 5194 7084 5206
rect 7026 4818 7038 5194
rect 7072 4818 7084 5194
rect 7026 4806 7084 4818
rect 7144 5194 7202 5206
rect 7144 4818 7156 5194
rect 7190 4818 7202 5194
rect 7261 5194 7319 5206
rect 7261 5018 7273 5194
rect 7307 5018 7319 5194
rect 7261 5006 7319 5018
rect 7379 5194 7437 5206
rect 20111 5214 20169 5226
rect 7379 5018 7391 5194
rect 7425 5018 7437 5194
rect 7379 5006 7437 5018
rect 13457 5193 13515 5205
rect 7144 4806 7202 4818
rect 13457 4817 13469 5193
rect 13503 4817 13515 5193
rect 13457 4805 13515 4817
rect 13575 5193 13633 5205
rect 13575 4817 13587 5193
rect 13621 4817 13633 5193
rect 13575 4805 13633 4817
rect 13693 5193 13751 5205
rect 13693 4817 13705 5193
rect 13739 4817 13751 5193
rect 13810 5193 13868 5205
rect 13810 5017 13822 5193
rect 13856 5017 13868 5193
rect 13810 5005 13868 5017
rect 13928 5193 13986 5205
rect 13928 5017 13940 5193
rect 13974 5017 13986 5193
rect 13928 5005 13986 5017
rect 20111 4838 20123 5214
rect 20157 4838 20169 5214
rect 20111 4826 20169 4838
rect 20229 5214 20287 5226
rect 20229 4838 20241 5214
rect 20275 4838 20287 5214
rect 20229 4826 20287 4838
rect 20347 5214 20405 5226
rect 20347 4838 20359 5214
rect 20393 4838 20405 5214
rect 20464 5214 20522 5226
rect 20464 5038 20476 5214
rect 20510 5038 20522 5214
rect 20464 5026 20522 5038
rect 20582 5214 20640 5226
rect 20582 5038 20594 5214
rect 20628 5038 20640 5214
rect 20582 5026 20640 5038
rect 28764 5047 28822 5059
rect 20347 4826 20405 4838
rect 13693 4805 13751 4817
rect 28764 4671 28776 5047
rect 28810 4671 28822 5047
rect 28764 4659 28822 4671
rect 28882 5047 28940 5059
rect 28882 4671 28894 5047
rect 28928 4671 28940 5047
rect 28882 4659 28940 4671
rect 29000 5047 29058 5059
rect 29000 4671 29012 5047
rect 29046 4671 29058 5047
rect 29117 5047 29175 5059
rect 29117 4871 29129 5047
rect 29163 4871 29175 5047
rect 29117 4859 29175 4871
rect 29235 5047 29293 5059
rect 29235 4871 29247 5047
rect 29281 4871 29293 5047
rect 29235 4859 29293 4871
rect 29000 4659 29058 4671
rect 32365 4639 32423 4651
rect 32365 4263 32377 4639
rect 32411 4263 32423 4639
rect 32365 4251 32423 4263
rect 32483 4639 32541 4651
rect 32483 4263 32495 4639
rect 32529 4263 32541 4639
rect 32483 4251 32541 4263
rect 32601 4639 32659 4651
rect 32601 4263 32613 4639
rect 32647 4263 32659 4639
rect 32718 4639 32776 4651
rect 32718 4463 32730 4639
rect 32764 4463 32776 4639
rect 32718 4451 32776 4463
rect 32836 4639 32894 4651
rect 32836 4463 32848 4639
rect 32882 4463 32894 4639
rect 32836 4451 32894 4463
rect 32601 4251 32659 4263
rect 30460 3854 30518 3866
rect 244 3294 302 3306
rect 244 2918 256 3294
rect 290 2918 302 3294
rect 244 2906 302 2918
rect 362 3294 420 3306
rect 362 2918 374 3294
rect 408 2918 420 3294
rect 362 2906 420 2918
rect 480 3294 538 3306
rect 480 2918 492 3294
rect 526 2918 538 3294
rect 597 3294 655 3306
rect 597 3118 609 3294
rect 643 3118 655 3294
rect 597 3106 655 3118
rect 715 3294 773 3306
rect 715 3118 727 3294
rect 761 3118 773 3294
rect 715 3106 773 3118
rect 480 2906 538 2918
rect 3134 3027 3192 3039
rect 3134 2651 3146 3027
rect 3180 2651 3192 3027
rect 3134 2639 3192 2651
rect 3252 3027 3310 3039
rect 3252 2651 3264 3027
rect 3298 2651 3310 3027
rect 3252 2639 3310 2651
rect 3370 3027 3428 3039
rect 3370 2651 3382 3027
rect 3416 2651 3428 3027
rect 3487 3027 3545 3039
rect 3487 2851 3499 3027
rect 3533 2851 3545 3027
rect 3487 2839 3545 2851
rect 3605 3027 3663 3039
rect 3605 2851 3617 3027
rect 3651 2851 3663 3027
rect 3605 2839 3663 2851
rect 30460 3678 30472 3854
rect 30506 3678 30518 3854
rect 30460 3666 30518 3678
rect 30578 3854 30636 3866
rect 30578 3678 30590 3854
rect 30624 3678 30636 3854
rect 30578 3666 30636 3678
rect 30880 3854 30938 3866
rect 9683 3115 9741 3127
rect 5132 2753 5190 2765
rect 3370 2639 3428 2651
rect 5132 2577 5144 2753
rect 5178 2577 5190 2753
rect 5132 2565 5190 2577
rect 5250 2753 5308 2765
rect 5250 2577 5262 2753
rect 5296 2577 5308 2753
rect 5250 2565 5308 2577
rect 5368 2753 5426 2765
rect 5368 2577 5380 2753
rect 5414 2577 5426 2753
rect 5368 2565 5426 2577
rect 5486 2753 5544 2765
rect 5486 2577 5498 2753
rect 5532 2577 5544 2753
rect 5486 2565 5544 2577
rect 6274 2757 6332 2769
rect 6274 2581 6286 2757
rect 6320 2581 6332 2757
rect 6274 2569 6332 2581
rect 6392 2757 6450 2769
rect 6392 2581 6404 2757
rect 6438 2581 6450 2757
rect 6392 2569 6450 2581
rect 6510 2757 6568 2769
rect 6510 2581 6522 2757
rect 6556 2581 6568 2757
rect 6510 2569 6568 2581
rect 6628 2757 6686 2769
rect 6628 2581 6640 2757
rect 6674 2581 6686 2757
rect 6628 2569 6686 2581
rect 9683 2739 9695 3115
rect 9729 2739 9741 3115
rect 9683 2727 9741 2739
rect 9801 3115 9859 3127
rect 9801 2739 9813 3115
rect 9847 2739 9859 3115
rect 9801 2727 9859 2739
rect 9919 3115 9977 3127
rect 9919 2739 9931 3115
rect 9965 2739 9977 3115
rect 10036 3115 10094 3127
rect 10036 2939 10048 3115
rect 10082 2939 10094 3115
rect 10036 2927 10094 2939
rect 10154 3115 10212 3127
rect 10154 2939 10166 3115
rect 10200 2939 10212 3115
rect 10154 2927 10212 2939
rect 16337 3047 16395 3059
rect 11681 2841 11739 2853
rect 9919 2727 9977 2739
rect 11681 2665 11693 2841
rect 11727 2665 11739 2841
rect 11681 2653 11739 2665
rect 11799 2841 11857 2853
rect 11799 2665 11811 2841
rect 11845 2665 11857 2841
rect 11799 2653 11857 2665
rect 11917 2841 11975 2853
rect 11917 2665 11929 2841
rect 11963 2665 11975 2841
rect 11917 2653 11975 2665
rect 12035 2841 12093 2853
rect 12035 2665 12047 2841
rect 12081 2665 12093 2841
rect 12035 2653 12093 2665
rect 12823 2845 12881 2857
rect 12823 2669 12835 2845
rect 12869 2669 12881 2845
rect 12823 2657 12881 2669
rect 12941 2845 12999 2857
rect 12941 2669 12953 2845
rect 12987 2669 12999 2845
rect 12941 2657 12999 2669
rect 13059 2845 13117 2857
rect 13059 2669 13071 2845
rect 13105 2669 13117 2845
rect 13059 2657 13117 2669
rect 13177 2845 13235 2857
rect 13177 2669 13189 2845
rect 13223 2669 13235 2845
rect 13177 2657 13235 2669
rect 16337 2671 16349 3047
rect 16383 2671 16395 3047
rect 16337 2659 16395 2671
rect 16455 3047 16513 3059
rect 16455 2671 16467 3047
rect 16501 2671 16513 3047
rect 16455 2659 16513 2671
rect 16573 3047 16631 3059
rect 16573 2671 16585 3047
rect 16619 2671 16631 3047
rect 16690 3047 16748 3059
rect 16690 2871 16702 3047
rect 16736 2871 16748 3047
rect 16690 2859 16748 2871
rect 16808 3047 16866 3059
rect 16808 2871 16820 3047
rect 16854 2871 16866 3047
rect 16808 2859 16866 2871
rect 30880 3478 30892 3854
rect 30926 3478 30938 3854
rect 30880 3466 30938 3478
rect 30998 3854 31056 3866
rect 30998 3478 31010 3854
rect 31044 3478 31056 3854
rect 30998 3466 31056 3478
rect 31116 3854 31174 3866
rect 31116 3478 31128 3854
rect 31162 3478 31174 3854
rect 31116 3466 31174 3478
rect 31234 3854 31292 3866
rect 31234 3478 31246 3854
rect 31280 3478 31292 3854
rect 31234 3466 31292 3478
rect 31352 3854 31410 3866
rect 31352 3478 31364 3854
rect 31398 3478 31410 3854
rect 31758 3854 31816 3866
rect 31758 3678 31770 3854
rect 31804 3678 31816 3854
rect 31758 3666 31816 3678
rect 31876 3854 31934 3866
rect 31876 3678 31888 3854
rect 31922 3678 31934 3854
rect 31876 3666 31934 3678
rect 31352 3466 31410 3478
rect 22962 3115 23020 3127
rect 18335 2773 18393 2785
rect 16573 2659 16631 2671
rect 18335 2597 18347 2773
rect 18381 2597 18393 2773
rect 18335 2585 18393 2597
rect 18453 2773 18511 2785
rect 18453 2597 18465 2773
rect 18499 2597 18511 2773
rect 18453 2585 18511 2597
rect 18571 2773 18629 2785
rect 18571 2597 18583 2773
rect 18617 2597 18629 2773
rect 18571 2585 18629 2597
rect 18689 2773 18747 2785
rect 18689 2597 18701 2773
rect 18735 2597 18747 2773
rect 18689 2585 18747 2597
rect 19477 2777 19535 2789
rect 19477 2601 19489 2777
rect 19523 2601 19535 2777
rect 19477 2589 19535 2601
rect 19595 2777 19653 2789
rect 19595 2601 19607 2777
rect 19641 2601 19653 2777
rect 19595 2589 19653 2601
rect 19713 2777 19771 2789
rect 19713 2601 19725 2777
rect 19759 2601 19771 2777
rect 19713 2589 19771 2601
rect 19831 2777 19889 2789
rect 19831 2601 19843 2777
rect 19877 2601 19889 2777
rect 19831 2589 19889 2601
rect 22962 2739 22974 3115
rect 23008 2739 23020 3115
rect 22962 2727 23020 2739
rect 23080 3115 23138 3127
rect 23080 2739 23092 3115
rect 23126 2739 23138 3115
rect 23080 2727 23138 2739
rect 23198 3115 23256 3127
rect 23198 2739 23210 3115
rect 23244 2739 23256 3115
rect 23315 3115 23373 3127
rect 23315 2939 23327 3115
rect 23361 2939 23373 3115
rect 23315 2927 23373 2939
rect 23433 3115 23491 3127
rect 23433 2939 23445 3115
rect 23479 2939 23491 3115
rect 23433 2927 23491 2939
rect 24960 2841 25018 2853
rect 23198 2727 23256 2739
rect 24960 2665 24972 2841
rect 25006 2665 25018 2841
rect 24960 2653 25018 2665
rect 25078 2841 25136 2853
rect 25078 2665 25090 2841
rect 25124 2665 25136 2841
rect 25078 2653 25136 2665
rect 25196 2841 25254 2853
rect 25196 2665 25208 2841
rect 25242 2665 25254 2841
rect 25196 2653 25254 2665
rect 25314 2841 25372 2853
rect 25314 2665 25326 2841
rect 25360 2665 25372 2841
rect 25314 2653 25372 2665
rect 26102 2845 26160 2857
rect 26102 2669 26114 2845
rect 26148 2669 26160 2845
rect 26102 2657 26160 2669
rect 26220 2845 26278 2857
rect 26220 2669 26232 2845
rect 26266 2669 26278 2845
rect 26220 2657 26278 2669
rect 26338 2845 26396 2857
rect 26338 2669 26350 2845
rect 26384 2669 26396 2845
rect 26338 2657 26396 2669
rect 26456 2845 26514 2857
rect 26456 2669 26468 2845
rect 26502 2669 26514 2845
rect 26456 2657 26514 2669
rect 28759 2476 28817 2488
rect 28759 2100 28771 2476
rect 28805 2100 28817 2476
rect 28759 2088 28817 2100
rect 28877 2476 28935 2488
rect 28877 2100 28889 2476
rect 28923 2100 28935 2476
rect 28877 2088 28935 2100
rect 28995 2476 29053 2488
rect 28995 2100 29007 2476
rect 29041 2100 29053 2476
rect 29112 2476 29170 2488
rect 29112 2300 29124 2476
rect 29158 2300 29170 2476
rect 29112 2288 29170 2300
rect 29230 2476 29288 2488
rect 29230 2300 29242 2476
rect 29276 2300 29288 2476
rect 29230 2288 29288 2300
rect 28995 2088 29053 2100
rect 9697 1465 9755 1477
rect 3148 1377 3206 1389
rect 3148 1001 3160 1377
rect 3194 1001 3206 1377
rect 3148 989 3206 1001
rect 3266 1377 3324 1389
rect 3266 1001 3278 1377
rect 3312 1001 3324 1377
rect 3266 989 3324 1001
rect 3384 1377 3442 1389
rect 3384 1001 3396 1377
rect 3430 1001 3442 1377
rect 3501 1377 3559 1389
rect 3501 1201 3513 1377
rect 3547 1201 3559 1377
rect 3501 1189 3559 1201
rect 3619 1377 3677 1389
rect 3619 1201 3631 1377
rect 3665 1201 3677 1377
rect 3619 1189 3677 1201
rect 3384 989 3442 1001
rect 9697 1089 9709 1465
rect 9743 1089 9755 1465
rect 9697 1077 9755 1089
rect 9815 1465 9873 1477
rect 9815 1089 9827 1465
rect 9861 1089 9873 1465
rect 9815 1077 9873 1089
rect 9933 1465 9991 1477
rect 9933 1089 9945 1465
rect 9979 1089 9991 1465
rect 10050 1465 10108 1477
rect 10050 1289 10062 1465
rect 10096 1289 10108 1465
rect 10050 1277 10108 1289
rect 10168 1465 10226 1477
rect 10168 1289 10180 1465
rect 10214 1289 10226 1465
rect 10168 1277 10226 1289
rect 9933 1077 9991 1089
rect 236 709 294 721
rect 236 333 248 709
rect 282 333 294 709
rect 236 321 294 333
rect 354 709 412 721
rect 354 333 366 709
rect 400 333 412 709
rect 354 321 412 333
rect 472 709 530 721
rect 472 333 484 709
rect 518 333 530 709
rect 589 709 647 721
rect 589 533 601 709
rect 635 533 647 709
rect 589 521 647 533
rect 707 709 765 721
rect 707 533 719 709
rect 753 533 765 709
rect 707 521 765 533
rect 472 321 530 333
rect 22976 1465 23034 1477
rect 16351 1397 16409 1409
rect 4500 -28 4558 -16
rect 4500 -204 4512 -28
rect 4546 -204 4558 -28
rect 3143 -227 3201 -215
rect 3143 -603 3155 -227
rect 3189 -603 3201 -227
rect 3143 -615 3201 -603
rect 3261 -227 3319 -215
rect 3261 -603 3273 -227
rect 3307 -603 3319 -227
rect 3261 -615 3319 -603
rect 3379 -227 3437 -215
rect 3379 -603 3391 -227
rect 3425 -603 3437 -227
rect 3496 -227 3554 -215
rect 3496 -403 3508 -227
rect 3542 -403 3554 -227
rect 3496 -415 3554 -403
rect 3614 -227 3672 -215
rect 4500 -216 4558 -204
rect 4618 -28 4676 -16
rect 4618 -204 4630 -28
rect 4664 -204 4676 -28
rect 4618 -216 4676 -204
rect 4920 -28 4978 -16
rect 3614 -403 3626 -227
rect 3660 -403 3672 -227
rect 3614 -415 3672 -403
rect 4920 -404 4932 -28
rect 4966 -404 4978 -28
rect 4920 -416 4978 -404
rect 5038 -28 5096 -16
rect 5038 -404 5050 -28
rect 5084 -404 5096 -28
rect 5038 -416 5096 -404
rect 5156 -28 5214 -16
rect 5156 -404 5168 -28
rect 5202 -404 5214 -28
rect 5156 -416 5214 -404
rect 5274 -28 5332 -16
rect 5274 -404 5286 -28
rect 5320 -404 5332 -28
rect 5274 -416 5332 -404
rect 5392 -28 5450 -16
rect 5392 -404 5404 -28
rect 5438 -404 5450 -28
rect 5798 -28 5856 -16
rect 5798 -204 5810 -28
rect 5844 -204 5856 -28
rect 5798 -216 5856 -204
rect 5916 -28 5974 -16
rect 5916 -204 5928 -28
rect 5962 -204 5974 -28
rect 5916 -216 5974 -204
rect 6398 -28 6456 -16
rect 6398 -204 6410 -28
rect 6444 -204 6456 -28
rect 6398 -216 6456 -204
rect 6516 -28 6574 -16
rect 6516 -204 6528 -28
rect 6562 -204 6574 -28
rect 6516 -216 6574 -204
rect 6818 -28 6876 -16
rect 5392 -416 5450 -404
rect 6818 -404 6830 -28
rect 6864 -404 6876 -28
rect 6818 -416 6876 -404
rect 6936 -28 6994 -16
rect 6936 -404 6948 -28
rect 6982 -404 6994 -28
rect 6936 -416 6994 -404
rect 7054 -28 7112 -16
rect 7054 -404 7066 -28
rect 7100 -404 7112 -28
rect 7054 -416 7112 -404
rect 7172 -28 7230 -16
rect 7172 -404 7184 -28
rect 7218 -404 7230 -28
rect 7172 -416 7230 -404
rect 7290 -28 7348 -16
rect 7290 -404 7302 -28
rect 7336 -404 7348 -28
rect 7696 -28 7754 -16
rect 7696 -204 7708 -28
rect 7742 -204 7754 -28
rect 7696 -216 7754 -204
rect 7814 -28 7872 -16
rect 7814 -204 7826 -28
rect 7860 -204 7872 -28
rect 16351 1021 16363 1397
rect 16397 1021 16409 1397
rect 16351 1009 16409 1021
rect 16469 1397 16527 1409
rect 16469 1021 16481 1397
rect 16515 1021 16527 1397
rect 16469 1009 16527 1021
rect 16587 1397 16645 1409
rect 16587 1021 16599 1397
rect 16633 1021 16645 1397
rect 16704 1397 16762 1409
rect 16704 1221 16716 1397
rect 16750 1221 16762 1397
rect 16704 1209 16762 1221
rect 16822 1397 16880 1409
rect 16822 1221 16834 1397
rect 16868 1221 16880 1397
rect 16822 1209 16880 1221
rect 16587 1009 16645 1021
rect 22976 1089 22988 1465
rect 23022 1089 23034 1465
rect 22976 1077 23034 1089
rect 23094 1465 23152 1477
rect 23094 1089 23106 1465
rect 23140 1089 23152 1465
rect 23094 1077 23152 1089
rect 23212 1465 23270 1477
rect 23212 1089 23224 1465
rect 23258 1089 23270 1465
rect 23329 1465 23387 1477
rect 23329 1289 23341 1465
rect 23375 1289 23387 1465
rect 23329 1277 23387 1289
rect 23447 1465 23505 1477
rect 23447 1289 23459 1465
rect 23493 1289 23505 1465
rect 23447 1277 23505 1289
rect 23212 1077 23270 1089
rect 11049 60 11107 72
rect 11049 -116 11061 60
rect 11095 -116 11107 60
rect 7814 -216 7872 -204
rect 9692 -139 9750 -127
rect 7290 -416 7348 -404
rect 9692 -515 9704 -139
rect 9738 -515 9750 -139
rect 3379 -615 3437 -603
rect 9692 -527 9750 -515
rect 9810 -139 9868 -127
rect 9810 -515 9822 -139
rect 9856 -515 9868 -139
rect 9810 -527 9868 -515
rect 9928 -139 9986 -127
rect 9928 -515 9940 -139
rect 9974 -515 9986 -139
rect 10045 -139 10103 -127
rect 10045 -315 10057 -139
rect 10091 -315 10103 -139
rect 10045 -327 10103 -315
rect 10163 -139 10221 -127
rect 11049 -128 11107 -116
rect 11167 60 11225 72
rect 11167 -116 11179 60
rect 11213 -116 11225 60
rect 11167 -128 11225 -116
rect 11469 60 11527 72
rect 10163 -315 10175 -139
rect 10209 -315 10221 -139
rect 10163 -327 10221 -315
rect 11469 -316 11481 60
rect 11515 -316 11527 60
rect 11469 -328 11527 -316
rect 11587 60 11645 72
rect 11587 -316 11599 60
rect 11633 -316 11645 60
rect 11587 -328 11645 -316
rect 11705 60 11763 72
rect 11705 -316 11717 60
rect 11751 -316 11763 60
rect 11705 -328 11763 -316
rect 11823 60 11881 72
rect 11823 -316 11835 60
rect 11869 -316 11881 60
rect 11823 -328 11881 -316
rect 11941 60 11999 72
rect 11941 -316 11953 60
rect 11987 -316 11999 60
rect 12347 60 12405 72
rect 12347 -116 12359 60
rect 12393 -116 12405 60
rect 12347 -128 12405 -116
rect 12465 60 12523 72
rect 12465 -116 12477 60
rect 12511 -116 12523 60
rect 12465 -128 12523 -116
rect 12947 60 13005 72
rect 12947 -116 12959 60
rect 12993 -116 13005 60
rect 12947 -128 13005 -116
rect 13065 60 13123 72
rect 13065 -116 13077 60
rect 13111 -116 13123 60
rect 13065 -128 13123 -116
rect 13367 60 13425 72
rect 11941 -328 11999 -316
rect 13367 -316 13379 60
rect 13413 -316 13425 60
rect 13367 -328 13425 -316
rect 13485 60 13543 72
rect 13485 -316 13497 60
rect 13531 -316 13543 60
rect 13485 -328 13543 -316
rect 13603 60 13661 72
rect 13603 -316 13615 60
rect 13649 -316 13661 60
rect 13603 -328 13661 -316
rect 13721 60 13779 72
rect 13721 -316 13733 60
rect 13767 -316 13779 60
rect 13721 -328 13779 -316
rect 13839 60 13897 72
rect 13839 -316 13851 60
rect 13885 -316 13897 60
rect 14245 60 14303 72
rect 14245 -116 14257 60
rect 14291 -116 14303 60
rect 14245 -128 14303 -116
rect 14363 60 14421 72
rect 14363 -116 14375 60
rect 14409 -116 14421 60
rect 14363 -128 14421 -116
rect 17703 -8 17761 4
rect 17703 -184 17715 -8
rect 17749 -184 17761 -8
rect 13839 -328 13897 -316
rect 16346 -207 16404 -195
rect 9928 -527 9986 -515
rect 16346 -583 16358 -207
rect 16392 -583 16404 -207
rect 16346 -595 16404 -583
rect 16464 -207 16522 -195
rect 16464 -583 16476 -207
rect 16510 -583 16522 -207
rect 16464 -595 16522 -583
rect 16582 -207 16640 -195
rect 16582 -583 16594 -207
rect 16628 -583 16640 -207
rect 16699 -207 16757 -195
rect 16699 -383 16711 -207
rect 16745 -383 16757 -207
rect 16699 -395 16757 -383
rect 16817 -207 16875 -195
rect 17703 -196 17761 -184
rect 17821 -8 17879 4
rect 17821 -184 17833 -8
rect 17867 -184 17879 -8
rect 17821 -196 17879 -184
rect 18123 -8 18181 4
rect 16817 -383 16829 -207
rect 16863 -383 16875 -207
rect 16817 -395 16875 -383
rect 18123 -384 18135 -8
rect 18169 -384 18181 -8
rect 18123 -396 18181 -384
rect 18241 -8 18299 4
rect 18241 -384 18253 -8
rect 18287 -384 18299 -8
rect 18241 -396 18299 -384
rect 18359 -8 18417 4
rect 18359 -384 18371 -8
rect 18405 -384 18417 -8
rect 18359 -396 18417 -384
rect 18477 -8 18535 4
rect 18477 -384 18489 -8
rect 18523 -384 18535 -8
rect 18477 -396 18535 -384
rect 18595 -8 18653 4
rect 18595 -384 18607 -8
rect 18641 -384 18653 -8
rect 19001 -8 19059 4
rect 19001 -184 19013 -8
rect 19047 -184 19059 -8
rect 19001 -196 19059 -184
rect 19119 -8 19177 4
rect 19119 -184 19131 -8
rect 19165 -184 19177 -8
rect 19119 -196 19177 -184
rect 19601 -8 19659 4
rect 19601 -184 19613 -8
rect 19647 -184 19659 -8
rect 19601 -196 19659 -184
rect 19719 -8 19777 4
rect 19719 -184 19731 -8
rect 19765 -184 19777 -8
rect 19719 -196 19777 -184
rect 20021 -8 20079 4
rect 18595 -396 18653 -384
rect 20021 -384 20033 -8
rect 20067 -384 20079 -8
rect 20021 -396 20079 -384
rect 20139 -8 20197 4
rect 20139 -384 20151 -8
rect 20185 -384 20197 -8
rect 20139 -396 20197 -384
rect 20257 -8 20315 4
rect 20257 -384 20269 -8
rect 20303 -384 20315 -8
rect 20257 -396 20315 -384
rect 20375 -8 20433 4
rect 20375 -384 20387 -8
rect 20421 -384 20433 -8
rect 20375 -396 20433 -384
rect 20493 -8 20551 4
rect 20493 -384 20505 -8
rect 20539 -384 20551 -8
rect 20899 -8 20957 4
rect 20899 -184 20911 -8
rect 20945 -184 20957 -8
rect 20899 -196 20957 -184
rect 21017 -8 21075 4
rect 21017 -184 21029 -8
rect 21063 -184 21075 -8
rect 24328 60 24386 72
rect 24328 -116 24340 60
rect 24374 -116 24386 60
rect 21017 -196 21075 -184
rect 22971 -139 23029 -127
rect 20493 -396 20551 -384
rect 16582 -595 16640 -583
rect 22971 -515 22983 -139
rect 23017 -515 23029 -139
rect 22971 -527 23029 -515
rect 23089 -139 23147 -127
rect 23089 -515 23101 -139
rect 23135 -515 23147 -139
rect 23089 -527 23147 -515
rect 23207 -139 23265 -127
rect 23207 -515 23219 -139
rect 23253 -515 23265 -139
rect 23324 -139 23382 -127
rect 23324 -315 23336 -139
rect 23370 -315 23382 -139
rect 23324 -327 23382 -315
rect 23442 -139 23500 -127
rect 24328 -128 24386 -116
rect 24446 60 24504 72
rect 24446 -116 24458 60
rect 24492 -116 24504 60
rect 24446 -128 24504 -116
rect 24748 60 24806 72
rect 23442 -315 23454 -139
rect 23488 -315 23500 -139
rect 23442 -327 23500 -315
rect 24748 -316 24760 60
rect 24794 -316 24806 60
rect 24748 -328 24806 -316
rect 24866 60 24924 72
rect 24866 -316 24878 60
rect 24912 -316 24924 60
rect 24866 -328 24924 -316
rect 24984 60 25042 72
rect 24984 -316 24996 60
rect 25030 -316 25042 60
rect 24984 -328 25042 -316
rect 25102 60 25160 72
rect 25102 -316 25114 60
rect 25148 -316 25160 60
rect 25102 -328 25160 -316
rect 25220 60 25278 72
rect 25220 -316 25232 60
rect 25266 -316 25278 60
rect 25626 60 25684 72
rect 25626 -116 25638 60
rect 25672 -116 25684 60
rect 25626 -128 25684 -116
rect 25744 60 25802 72
rect 25744 -116 25756 60
rect 25790 -116 25802 60
rect 25744 -128 25802 -116
rect 26226 60 26284 72
rect 26226 -116 26238 60
rect 26272 -116 26284 60
rect 26226 -128 26284 -116
rect 26344 60 26402 72
rect 26344 -116 26356 60
rect 26390 -116 26402 60
rect 26344 -128 26402 -116
rect 26646 60 26704 72
rect 25220 -328 25278 -316
rect 26646 -316 26658 60
rect 26692 -316 26704 60
rect 26646 -328 26704 -316
rect 26764 60 26822 72
rect 26764 -316 26776 60
rect 26810 -316 26822 60
rect 26764 -328 26822 -316
rect 26882 60 26940 72
rect 26882 -316 26894 60
rect 26928 -316 26940 60
rect 26882 -328 26940 -316
rect 27000 60 27058 72
rect 27000 -316 27012 60
rect 27046 -316 27058 60
rect 27000 -328 27058 -316
rect 27118 60 27176 72
rect 27118 -316 27130 60
rect 27164 -316 27176 60
rect 27524 60 27582 72
rect 27524 -116 27536 60
rect 27570 -116 27582 60
rect 27524 -128 27582 -116
rect 27642 60 27700 72
rect 27642 -116 27654 60
rect 27688 -116 27700 60
rect 27642 -128 27700 -116
rect 32367 548 32425 560
rect 32367 172 32379 548
rect 32413 172 32425 548
rect 32367 160 32425 172
rect 32485 548 32543 560
rect 32485 172 32497 548
rect 32531 172 32543 548
rect 32485 160 32543 172
rect 32603 548 32661 560
rect 32603 172 32615 548
rect 32649 172 32661 548
rect 32720 548 32778 560
rect 32720 372 32732 548
rect 32766 372 32778 548
rect 32720 360 32778 372
rect 32838 548 32896 560
rect 32838 372 32850 548
rect 32884 372 32896 548
rect 32838 360 32896 372
rect 32603 160 32661 172
rect 30462 -237 30520 -225
rect 27118 -328 27176 -316
rect 23207 -527 23265 -515
rect 30462 -413 30474 -237
rect 30508 -413 30520 -237
rect 30462 -425 30520 -413
rect 30580 -237 30638 -225
rect 30580 -413 30592 -237
rect 30626 -413 30638 -237
rect 30580 -425 30638 -413
rect 30882 -237 30940 -225
rect 28759 -557 28817 -545
rect 28759 -933 28771 -557
rect 28805 -933 28817 -557
rect 28759 -945 28817 -933
rect 28877 -557 28935 -545
rect 28877 -933 28889 -557
rect 28923 -933 28935 -557
rect 28877 -945 28935 -933
rect 28995 -557 29053 -545
rect 28995 -933 29007 -557
rect 29041 -933 29053 -557
rect 29112 -557 29170 -545
rect 29112 -733 29124 -557
rect 29158 -733 29170 -557
rect 29112 -745 29170 -733
rect 29230 -557 29288 -545
rect 29230 -733 29242 -557
rect 29276 -733 29288 -557
rect 30882 -613 30894 -237
rect 30928 -613 30940 -237
rect 30882 -625 30940 -613
rect 31000 -237 31058 -225
rect 31000 -613 31012 -237
rect 31046 -613 31058 -237
rect 31000 -625 31058 -613
rect 31118 -237 31176 -225
rect 31118 -613 31130 -237
rect 31164 -613 31176 -237
rect 31118 -625 31176 -613
rect 31236 -237 31294 -225
rect 31236 -613 31248 -237
rect 31282 -613 31294 -237
rect 31236 -625 31294 -613
rect 31354 -237 31412 -225
rect 31354 -613 31366 -237
rect 31400 -613 31412 -237
rect 31760 -237 31818 -225
rect 31760 -413 31772 -237
rect 31806 -413 31818 -237
rect 31760 -425 31818 -413
rect 31878 -237 31936 -225
rect 31878 -413 31890 -237
rect 31924 -413 31936 -237
rect 31878 -425 31936 -413
rect 31354 -625 31412 -613
rect 29230 -745 29288 -733
rect 28995 -945 29053 -933
rect 217 -2569 275 -2557
rect 217 -2945 229 -2569
rect 263 -2945 275 -2569
rect 217 -2957 275 -2945
rect 335 -2569 393 -2557
rect 335 -2945 347 -2569
rect 381 -2945 393 -2569
rect 335 -2957 393 -2945
rect 453 -2569 511 -2557
rect 453 -2945 465 -2569
rect 499 -2945 511 -2569
rect 570 -2569 628 -2557
rect 570 -2745 582 -2569
rect 616 -2745 628 -2569
rect 570 -2757 628 -2745
rect 688 -2569 746 -2557
rect 688 -2745 700 -2569
rect 734 -2745 746 -2569
rect 688 -2757 746 -2745
rect 3126 -2753 3184 -2741
rect 453 -2957 511 -2945
rect 3126 -3129 3138 -2753
rect 3172 -3129 3184 -2753
rect 3126 -3141 3184 -3129
rect 3244 -2753 3302 -2741
rect 3244 -3129 3256 -2753
rect 3290 -3129 3302 -2753
rect 3244 -3141 3302 -3129
rect 3362 -2753 3420 -2741
rect 3362 -3129 3374 -2753
rect 3408 -3129 3420 -2753
rect 3479 -2753 3537 -2741
rect 3479 -2929 3491 -2753
rect 3525 -2929 3537 -2753
rect 3479 -2941 3537 -2929
rect 3597 -2753 3655 -2741
rect 3597 -2929 3609 -2753
rect 3643 -2929 3655 -2753
rect 3597 -2941 3655 -2929
rect 9677 -2755 9735 -2743
rect 5124 -3027 5182 -3015
rect 3362 -3141 3420 -3129
rect 5124 -3203 5136 -3027
rect 5170 -3203 5182 -3027
rect 5124 -3215 5182 -3203
rect 5242 -3027 5300 -3015
rect 5242 -3203 5254 -3027
rect 5288 -3203 5300 -3027
rect 5242 -3215 5300 -3203
rect 5360 -3027 5418 -3015
rect 5360 -3203 5372 -3027
rect 5406 -3203 5418 -3027
rect 5360 -3215 5418 -3203
rect 5478 -3027 5536 -3015
rect 5478 -3203 5490 -3027
rect 5524 -3203 5536 -3027
rect 5478 -3215 5536 -3203
rect 6266 -3023 6324 -3011
rect 6266 -3199 6278 -3023
rect 6312 -3199 6324 -3023
rect 6266 -3211 6324 -3199
rect 6384 -3023 6442 -3011
rect 6384 -3199 6396 -3023
rect 6430 -3199 6442 -3023
rect 6384 -3211 6442 -3199
rect 6502 -3023 6560 -3011
rect 6502 -3199 6514 -3023
rect 6548 -3199 6560 -3023
rect 6502 -3211 6560 -3199
rect 6620 -3023 6678 -3011
rect 6620 -3199 6632 -3023
rect 6666 -3199 6678 -3023
rect 6620 -3211 6678 -3199
rect 9677 -3131 9689 -2755
rect 9723 -3131 9735 -2755
rect 9677 -3143 9735 -3131
rect 9795 -2755 9853 -2743
rect 9795 -3131 9807 -2755
rect 9841 -3131 9853 -2755
rect 9795 -3143 9853 -3131
rect 9913 -2755 9971 -2743
rect 9913 -3131 9925 -2755
rect 9959 -3131 9971 -2755
rect 10030 -2755 10088 -2743
rect 10030 -2931 10042 -2755
rect 10076 -2931 10088 -2755
rect 10030 -2943 10088 -2931
rect 10148 -2755 10206 -2743
rect 10148 -2931 10160 -2755
rect 10194 -2931 10206 -2755
rect 10148 -2943 10206 -2931
rect 16332 -2754 16390 -2742
rect 11675 -3029 11733 -3017
rect 9913 -3143 9971 -3131
rect 11675 -3205 11687 -3029
rect 11721 -3205 11733 -3029
rect 11675 -3217 11733 -3205
rect 11793 -3029 11851 -3017
rect 11793 -3205 11805 -3029
rect 11839 -3205 11851 -3029
rect 11793 -3217 11851 -3205
rect 11911 -3029 11969 -3017
rect 11911 -3205 11923 -3029
rect 11957 -3205 11969 -3029
rect 11911 -3217 11969 -3205
rect 12029 -3029 12087 -3017
rect 12029 -3205 12041 -3029
rect 12075 -3205 12087 -3029
rect 12029 -3217 12087 -3205
rect 12817 -3025 12875 -3013
rect 12817 -3201 12829 -3025
rect 12863 -3201 12875 -3025
rect 12817 -3213 12875 -3201
rect 12935 -3025 12993 -3013
rect 12935 -3201 12947 -3025
rect 12981 -3201 12993 -3025
rect 12935 -3213 12993 -3201
rect 13053 -3025 13111 -3013
rect 13053 -3201 13065 -3025
rect 13099 -3201 13111 -3025
rect 13053 -3213 13111 -3201
rect 13171 -3025 13229 -3013
rect 13171 -3201 13183 -3025
rect 13217 -3201 13229 -3025
rect 13171 -3213 13229 -3201
rect 16332 -3130 16344 -2754
rect 16378 -3130 16390 -2754
rect 16332 -3142 16390 -3130
rect 16450 -2754 16508 -2742
rect 16450 -3130 16462 -2754
rect 16496 -3130 16508 -2754
rect 16450 -3142 16508 -3130
rect 16568 -2754 16626 -2742
rect 16568 -3130 16580 -2754
rect 16614 -3130 16626 -2754
rect 16685 -2754 16743 -2742
rect 16685 -2930 16697 -2754
rect 16731 -2930 16743 -2754
rect 16685 -2942 16743 -2930
rect 16803 -2754 16861 -2742
rect 16803 -2930 16815 -2754
rect 16849 -2930 16861 -2754
rect 16803 -2942 16861 -2930
rect 28830 -2477 28888 -2465
rect 22954 -2753 23012 -2741
rect 18330 -3028 18388 -3016
rect 16568 -3142 16626 -3130
rect 18330 -3204 18342 -3028
rect 18376 -3204 18388 -3028
rect 18330 -3216 18388 -3204
rect 18448 -3028 18506 -3016
rect 18448 -3204 18460 -3028
rect 18494 -3204 18506 -3028
rect 18448 -3216 18506 -3204
rect 18566 -3028 18624 -3016
rect 18566 -3204 18578 -3028
rect 18612 -3204 18624 -3028
rect 18566 -3216 18624 -3204
rect 18684 -3028 18742 -3016
rect 18684 -3204 18696 -3028
rect 18730 -3204 18742 -3028
rect 18684 -3216 18742 -3204
rect 19472 -3024 19530 -3012
rect 19472 -3200 19484 -3024
rect 19518 -3200 19530 -3024
rect 19472 -3212 19530 -3200
rect 19590 -3024 19648 -3012
rect 19590 -3200 19602 -3024
rect 19636 -3200 19648 -3024
rect 19590 -3212 19648 -3200
rect 19708 -3024 19766 -3012
rect 19708 -3200 19720 -3024
rect 19754 -3200 19766 -3024
rect 19708 -3212 19766 -3200
rect 19826 -3024 19884 -3012
rect 19826 -3200 19838 -3024
rect 19872 -3200 19884 -3024
rect 19826 -3212 19884 -3200
rect 22954 -3129 22966 -2753
rect 23000 -3129 23012 -2753
rect 22954 -3141 23012 -3129
rect 23072 -2753 23130 -2741
rect 23072 -3129 23084 -2753
rect 23118 -3129 23130 -2753
rect 23072 -3141 23130 -3129
rect 23190 -2753 23248 -2741
rect 23190 -3129 23202 -2753
rect 23236 -3129 23248 -2753
rect 23307 -2753 23365 -2741
rect 23307 -2929 23319 -2753
rect 23353 -2929 23365 -2753
rect 23307 -2941 23365 -2929
rect 23425 -2753 23483 -2741
rect 23425 -2929 23437 -2753
rect 23471 -2929 23483 -2753
rect 23425 -2941 23483 -2929
rect 28830 -2853 28842 -2477
rect 28876 -2853 28888 -2477
rect 28830 -2865 28888 -2853
rect 28948 -2477 29006 -2465
rect 28948 -2853 28960 -2477
rect 28994 -2853 29006 -2477
rect 28948 -2865 29006 -2853
rect 29066 -2477 29124 -2465
rect 29066 -2853 29078 -2477
rect 29112 -2853 29124 -2477
rect 29183 -2477 29241 -2465
rect 29183 -2653 29195 -2477
rect 29229 -2653 29241 -2477
rect 29183 -2665 29241 -2653
rect 29301 -2477 29359 -2465
rect 29301 -2653 29313 -2477
rect 29347 -2653 29359 -2477
rect 29301 -2665 29359 -2653
rect 29066 -2865 29124 -2853
rect 24952 -3027 25010 -3015
rect 23190 -3141 23248 -3129
rect 24952 -3203 24964 -3027
rect 24998 -3203 25010 -3027
rect 24952 -3215 25010 -3203
rect 25070 -3027 25128 -3015
rect 25070 -3203 25082 -3027
rect 25116 -3203 25128 -3027
rect 25070 -3215 25128 -3203
rect 25188 -3027 25246 -3015
rect 25188 -3203 25200 -3027
rect 25234 -3203 25246 -3027
rect 25188 -3215 25246 -3203
rect 25306 -3027 25364 -3015
rect 25306 -3203 25318 -3027
rect 25352 -3203 25364 -3027
rect 25306 -3215 25364 -3203
rect 26094 -3023 26152 -3011
rect 26094 -3199 26106 -3023
rect 26140 -3199 26152 -3023
rect 26094 -3211 26152 -3199
rect 26212 -3023 26270 -3011
rect 26212 -3199 26224 -3023
rect 26258 -3199 26270 -3023
rect 26212 -3211 26270 -3199
rect 26330 -3023 26388 -3011
rect 26330 -3199 26342 -3023
rect 26376 -3199 26388 -3023
rect 26330 -3211 26388 -3199
rect 26448 -3023 26506 -3011
rect 26448 -3199 26460 -3023
rect 26494 -3199 26506 -3023
rect 26448 -3211 26506 -3199
rect 32367 -2947 32425 -2935
rect 32367 -3323 32379 -2947
rect 32413 -3323 32425 -2947
rect 32367 -3335 32425 -3323
rect 32485 -2947 32543 -2935
rect 32485 -3323 32497 -2947
rect 32531 -3323 32543 -2947
rect 32485 -3335 32543 -3323
rect 32603 -2947 32661 -2935
rect 32603 -3323 32615 -2947
rect 32649 -3323 32661 -2947
rect 32720 -2947 32778 -2935
rect 32720 -3123 32732 -2947
rect 32766 -3123 32778 -2947
rect 32720 -3135 32778 -3123
rect 32838 -2947 32896 -2935
rect 32838 -3123 32850 -2947
rect 32884 -3123 32896 -2947
rect 32838 -3135 32896 -3123
rect 32603 -3335 32661 -3323
rect 30462 -3732 30520 -3720
rect 30462 -3908 30474 -3732
rect 30508 -3908 30520 -3732
rect 30462 -3920 30520 -3908
rect 30580 -3732 30638 -3720
rect 30580 -3908 30592 -3732
rect 30626 -3908 30638 -3732
rect 30580 -3920 30638 -3908
rect 30882 -3732 30940 -3720
rect 30882 -4108 30894 -3732
rect 30928 -4108 30940 -3732
rect 30882 -4120 30940 -4108
rect 31000 -3732 31058 -3720
rect 31000 -4108 31012 -3732
rect 31046 -4108 31058 -3732
rect 31000 -4120 31058 -4108
rect 31118 -3732 31176 -3720
rect 31118 -4108 31130 -3732
rect 31164 -4108 31176 -3732
rect 31118 -4120 31176 -4108
rect 31236 -3732 31294 -3720
rect 31236 -4108 31248 -3732
rect 31282 -4108 31294 -3732
rect 31236 -4120 31294 -4108
rect 31354 -3732 31412 -3720
rect 31354 -4108 31366 -3732
rect 31400 -4108 31412 -3732
rect 31760 -3732 31818 -3720
rect 31760 -3908 31772 -3732
rect 31806 -3908 31818 -3732
rect 31760 -3920 31818 -3908
rect 31878 -3732 31936 -3720
rect 31878 -3908 31890 -3732
rect 31924 -3908 31936 -3732
rect 31878 -3920 31936 -3908
rect 31354 -4120 31412 -4108
rect 3140 -4403 3198 -4391
rect 3140 -4779 3152 -4403
rect 3186 -4779 3198 -4403
rect 3140 -4791 3198 -4779
rect 3258 -4403 3316 -4391
rect 3258 -4779 3270 -4403
rect 3304 -4779 3316 -4403
rect 3258 -4791 3316 -4779
rect 3376 -4403 3434 -4391
rect 3376 -4779 3388 -4403
rect 3422 -4779 3434 -4403
rect 3493 -4403 3551 -4391
rect 3493 -4579 3505 -4403
rect 3539 -4579 3551 -4403
rect 3493 -4591 3551 -4579
rect 3611 -4403 3669 -4391
rect 3611 -4579 3623 -4403
rect 3657 -4579 3669 -4403
rect 3611 -4591 3669 -4579
rect 3376 -4791 3434 -4779
rect 9691 -4405 9749 -4393
rect 233 -5329 291 -5317
rect 233 -5705 245 -5329
rect 279 -5705 291 -5329
rect 233 -5717 291 -5705
rect 351 -5329 409 -5317
rect 351 -5705 363 -5329
rect 397 -5705 409 -5329
rect 351 -5717 409 -5705
rect 469 -5329 527 -5317
rect 469 -5705 481 -5329
rect 515 -5705 527 -5329
rect 586 -5329 644 -5317
rect 586 -5505 598 -5329
rect 632 -5505 644 -5329
rect 586 -5517 644 -5505
rect 704 -5329 762 -5317
rect 704 -5505 716 -5329
rect 750 -5505 762 -5329
rect 704 -5517 762 -5505
rect 469 -5717 527 -5705
rect 9691 -4781 9703 -4405
rect 9737 -4781 9749 -4405
rect 9691 -4793 9749 -4781
rect 9809 -4405 9867 -4393
rect 9809 -4781 9821 -4405
rect 9855 -4781 9867 -4405
rect 9809 -4793 9867 -4781
rect 9927 -4405 9985 -4393
rect 9927 -4781 9939 -4405
rect 9973 -4781 9985 -4405
rect 10044 -4405 10102 -4393
rect 10044 -4581 10056 -4405
rect 10090 -4581 10102 -4405
rect 10044 -4593 10102 -4581
rect 10162 -4405 10220 -4393
rect 10162 -4581 10174 -4405
rect 10208 -4581 10220 -4405
rect 10162 -4593 10220 -4581
rect 9927 -4793 9985 -4781
rect 16346 -4404 16404 -4392
rect 4492 -5808 4550 -5796
rect 4492 -5984 4504 -5808
rect 4538 -5984 4550 -5808
rect 3135 -6007 3193 -5995
rect 3135 -6383 3147 -6007
rect 3181 -6383 3193 -6007
rect 3135 -6395 3193 -6383
rect 3253 -6007 3311 -5995
rect 3253 -6383 3265 -6007
rect 3299 -6383 3311 -6007
rect 3253 -6395 3311 -6383
rect 3371 -6007 3429 -5995
rect 3371 -6383 3383 -6007
rect 3417 -6383 3429 -6007
rect 3488 -6007 3546 -5995
rect 3488 -6183 3500 -6007
rect 3534 -6183 3546 -6007
rect 3488 -6195 3546 -6183
rect 3606 -6007 3664 -5995
rect 4492 -5996 4550 -5984
rect 4610 -5808 4668 -5796
rect 4610 -5984 4622 -5808
rect 4656 -5984 4668 -5808
rect 4610 -5996 4668 -5984
rect 4912 -5808 4970 -5796
rect 3606 -6183 3618 -6007
rect 3652 -6183 3664 -6007
rect 3606 -6195 3664 -6183
rect 4912 -6184 4924 -5808
rect 4958 -6184 4970 -5808
rect 4912 -6196 4970 -6184
rect 5030 -5808 5088 -5796
rect 5030 -6184 5042 -5808
rect 5076 -6184 5088 -5808
rect 5030 -6196 5088 -6184
rect 5148 -5808 5206 -5796
rect 5148 -6184 5160 -5808
rect 5194 -6184 5206 -5808
rect 5148 -6196 5206 -6184
rect 5266 -5808 5324 -5796
rect 5266 -6184 5278 -5808
rect 5312 -6184 5324 -5808
rect 5266 -6196 5324 -6184
rect 5384 -5808 5442 -5796
rect 5384 -6184 5396 -5808
rect 5430 -6184 5442 -5808
rect 5790 -5808 5848 -5796
rect 5790 -5984 5802 -5808
rect 5836 -5984 5848 -5808
rect 5790 -5996 5848 -5984
rect 5908 -5808 5966 -5796
rect 5908 -5984 5920 -5808
rect 5954 -5984 5966 -5808
rect 5908 -5996 5966 -5984
rect 6390 -5808 6448 -5796
rect 6390 -5984 6402 -5808
rect 6436 -5984 6448 -5808
rect 6390 -5996 6448 -5984
rect 6508 -5808 6566 -5796
rect 6508 -5984 6520 -5808
rect 6554 -5984 6566 -5808
rect 6508 -5996 6566 -5984
rect 6810 -5808 6868 -5796
rect 5384 -6196 5442 -6184
rect 6810 -6184 6822 -5808
rect 6856 -6184 6868 -5808
rect 6810 -6196 6868 -6184
rect 6928 -5808 6986 -5796
rect 6928 -6184 6940 -5808
rect 6974 -6184 6986 -5808
rect 6928 -6196 6986 -6184
rect 7046 -5808 7104 -5796
rect 7046 -6184 7058 -5808
rect 7092 -6184 7104 -5808
rect 7046 -6196 7104 -6184
rect 7164 -5808 7222 -5796
rect 7164 -6184 7176 -5808
rect 7210 -6184 7222 -5808
rect 7164 -6196 7222 -6184
rect 7282 -5808 7340 -5796
rect 7282 -6184 7294 -5808
rect 7328 -6184 7340 -5808
rect 7688 -5808 7746 -5796
rect 7688 -5984 7700 -5808
rect 7734 -5984 7746 -5808
rect 7688 -5996 7746 -5984
rect 7806 -5808 7864 -5796
rect 7806 -5984 7818 -5808
rect 7852 -5984 7864 -5808
rect 7806 -5996 7864 -5984
rect 16346 -4780 16358 -4404
rect 16392 -4780 16404 -4404
rect 16346 -4792 16404 -4780
rect 16464 -4404 16522 -4392
rect 16464 -4780 16476 -4404
rect 16510 -4780 16522 -4404
rect 16464 -4792 16522 -4780
rect 16582 -4404 16640 -4392
rect 16582 -4780 16594 -4404
rect 16628 -4780 16640 -4404
rect 16699 -4404 16757 -4392
rect 16699 -4580 16711 -4404
rect 16745 -4580 16757 -4404
rect 16699 -4592 16757 -4580
rect 16817 -4404 16875 -4392
rect 16817 -4580 16829 -4404
rect 16863 -4580 16875 -4404
rect 16817 -4592 16875 -4580
rect 16582 -4792 16640 -4780
rect 22968 -4403 23026 -4391
rect 11043 -5810 11101 -5798
rect 11043 -5986 11055 -5810
rect 11089 -5986 11101 -5810
rect 9686 -6009 9744 -5997
rect 7282 -6196 7340 -6184
rect 3371 -6395 3429 -6383
rect 9686 -6385 9698 -6009
rect 9732 -6385 9744 -6009
rect 9686 -6397 9744 -6385
rect 9804 -6009 9862 -5997
rect 9804 -6385 9816 -6009
rect 9850 -6385 9862 -6009
rect 9804 -6397 9862 -6385
rect 9922 -6009 9980 -5997
rect 9922 -6385 9934 -6009
rect 9968 -6385 9980 -6009
rect 10039 -6009 10097 -5997
rect 10039 -6185 10051 -6009
rect 10085 -6185 10097 -6009
rect 10039 -6197 10097 -6185
rect 10157 -6009 10215 -5997
rect 11043 -5998 11101 -5986
rect 11161 -5810 11219 -5798
rect 11161 -5986 11173 -5810
rect 11207 -5986 11219 -5810
rect 11161 -5998 11219 -5986
rect 11463 -5810 11521 -5798
rect 10157 -6185 10169 -6009
rect 10203 -6185 10215 -6009
rect 10157 -6197 10215 -6185
rect 11463 -6186 11475 -5810
rect 11509 -6186 11521 -5810
rect 11463 -6198 11521 -6186
rect 11581 -5810 11639 -5798
rect 11581 -6186 11593 -5810
rect 11627 -6186 11639 -5810
rect 11581 -6198 11639 -6186
rect 11699 -5810 11757 -5798
rect 11699 -6186 11711 -5810
rect 11745 -6186 11757 -5810
rect 11699 -6198 11757 -6186
rect 11817 -5810 11875 -5798
rect 11817 -6186 11829 -5810
rect 11863 -6186 11875 -5810
rect 11817 -6198 11875 -6186
rect 11935 -5810 11993 -5798
rect 11935 -6186 11947 -5810
rect 11981 -6186 11993 -5810
rect 12341 -5810 12399 -5798
rect 12341 -5986 12353 -5810
rect 12387 -5986 12399 -5810
rect 12341 -5998 12399 -5986
rect 12459 -5810 12517 -5798
rect 12459 -5986 12471 -5810
rect 12505 -5986 12517 -5810
rect 12459 -5998 12517 -5986
rect 12941 -5810 12999 -5798
rect 12941 -5986 12953 -5810
rect 12987 -5986 12999 -5810
rect 12941 -5998 12999 -5986
rect 13059 -5810 13117 -5798
rect 13059 -5986 13071 -5810
rect 13105 -5986 13117 -5810
rect 13059 -5998 13117 -5986
rect 13361 -5810 13419 -5798
rect 11935 -6198 11993 -6186
rect 13361 -6186 13373 -5810
rect 13407 -6186 13419 -5810
rect 13361 -6198 13419 -6186
rect 13479 -5810 13537 -5798
rect 13479 -6186 13491 -5810
rect 13525 -6186 13537 -5810
rect 13479 -6198 13537 -6186
rect 13597 -5810 13655 -5798
rect 13597 -6186 13609 -5810
rect 13643 -6186 13655 -5810
rect 13597 -6198 13655 -6186
rect 13715 -5810 13773 -5798
rect 13715 -6186 13727 -5810
rect 13761 -6186 13773 -5810
rect 13715 -6198 13773 -6186
rect 13833 -5810 13891 -5798
rect 13833 -6186 13845 -5810
rect 13879 -6186 13891 -5810
rect 14239 -5810 14297 -5798
rect 14239 -5986 14251 -5810
rect 14285 -5986 14297 -5810
rect 14239 -5998 14297 -5986
rect 14357 -5810 14415 -5798
rect 14357 -5986 14369 -5810
rect 14403 -5986 14415 -5810
rect 14357 -5998 14415 -5986
rect 22968 -4779 22980 -4403
rect 23014 -4779 23026 -4403
rect 22968 -4791 23026 -4779
rect 23086 -4403 23144 -4391
rect 23086 -4779 23098 -4403
rect 23132 -4779 23144 -4403
rect 23086 -4791 23144 -4779
rect 23204 -4403 23262 -4391
rect 23204 -4779 23216 -4403
rect 23250 -4779 23262 -4403
rect 23321 -4403 23379 -4391
rect 23321 -4579 23333 -4403
rect 23367 -4579 23379 -4403
rect 23321 -4591 23379 -4579
rect 23439 -4403 23497 -4391
rect 23439 -4579 23451 -4403
rect 23485 -4579 23497 -4403
rect 23439 -4591 23497 -4579
rect 23204 -4791 23262 -4779
rect 17698 -5809 17756 -5797
rect 17698 -5985 17710 -5809
rect 17744 -5985 17756 -5809
rect 16341 -6008 16399 -5996
rect 13833 -6198 13891 -6186
rect 9922 -6397 9980 -6385
rect 16341 -6384 16353 -6008
rect 16387 -6384 16399 -6008
rect 16341 -6396 16399 -6384
rect 16459 -6008 16517 -5996
rect 16459 -6384 16471 -6008
rect 16505 -6384 16517 -6008
rect 16459 -6396 16517 -6384
rect 16577 -6008 16635 -5996
rect 16577 -6384 16589 -6008
rect 16623 -6384 16635 -6008
rect 16694 -6008 16752 -5996
rect 16694 -6184 16706 -6008
rect 16740 -6184 16752 -6008
rect 16694 -6196 16752 -6184
rect 16812 -6008 16870 -5996
rect 17698 -5997 17756 -5985
rect 17816 -5809 17874 -5797
rect 17816 -5985 17828 -5809
rect 17862 -5985 17874 -5809
rect 17816 -5997 17874 -5985
rect 18118 -5809 18176 -5797
rect 16812 -6184 16824 -6008
rect 16858 -6184 16870 -6008
rect 16812 -6196 16870 -6184
rect 18118 -6185 18130 -5809
rect 18164 -6185 18176 -5809
rect 18118 -6197 18176 -6185
rect 18236 -5809 18294 -5797
rect 18236 -6185 18248 -5809
rect 18282 -6185 18294 -5809
rect 18236 -6197 18294 -6185
rect 18354 -5809 18412 -5797
rect 18354 -6185 18366 -5809
rect 18400 -6185 18412 -5809
rect 18354 -6197 18412 -6185
rect 18472 -5809 18530 -5797
rect 18472 -6185 18484 -5809
rect 18518 -6185 18530 -5809
rect 18472 -6197 18530 -6185
rect 18590 -5809 18648 -5797
rect 18590 -6185 18602 -5809
rect 18636 -6185 18648 -5809
rect 18996 -5809 19054 -5797
rect 18996 -5985 19008 -5809
rect 19042 -5985 19054 -5809
rect 18996 -5997 19054 -5985
rect 19114 -5809 19172 -5797
rect 19114 -5985 19126 -5809
rect 19160 -5985 19172 -5809
rect 19114 -5997 19172 -5985
rect 19596 -5809 19654 -5797
rect 19596 -5985 19608 -5809
rect 19642 -5985 19654 -5809
rect 19596 -5997 19654 -5985
rect 19714 -5809 19772 -5797
rect 19714 -5985 19726 -5809
rect 19760 -5985 19772 -5809
rect 19714 -5997 19772 -5985
rect 20016 -5809 20074 -5797
rect 18590 -6197 18648 -6185
rect 20016 -6185 20028 -5809
rect 20062 -6185 20074 -5809
rect 20016 -6197 20074 -6185
rect 20134 -5809 20192 -5797
rect 20134 -6185 20146 -5809
rect 20180 -6185 20192 -5809
rect 20134 -6197 20192 -6185
rect 20252 -5809 20310 -5797
rect 20252 -6185 20264 -5809
rect 20298 -6185 20310 -5809
rect 20252 -6197 20310 -6185
rect 20370 -5809 20428 -5797
rect 20370 -6185 20382 -5809
rect 20416 -6185 20428 -5809
rect 20370 -6197 20428 -6185
rect 20488 -5809 20546 -5797
rect 20488 -6185 20500 -5809
rect 20534 -6185 20546 -5809
rect 20894 -5809 20952 -5797
rect 20894 -5985 20906 -5809
rect 20940 -5985 20952 -5809
rect 20894 -5997 20952 -5985
rect 21012 -5809 21070 -5797
rect 21012 -5985 21024 -5809
rect 21058 -5985 21070 -5809
rect 21012 -5997 21070 -5985
rect 28827 -5547 28885 -5535
rect 24320 -5808 24378 -5796
rect 24320 -5984 24332 -5808
rect 24366 -5984 24378 -5808
rect 22963 -6007 23021 -5995
rect 20488 -6197 20546 -6185
rect 16577 -6396 16635 -6384
rect 22963 -6383 22975 -6007
rect 23009 -6383 23021 -6007
rect 22963 -6395 23021 -6383
rect 23081 -6007 23139 -5995
rect 23081 -6383 23093 -6007
rect 23127 -6383 23139 -6007
rect 23081 -6395 23139 -6383
rect 23199 -6007 23257 -5995
rect 23199 -6383 23211 -6007
rect 23245 -6383 23257 -6007
rect 23316 -6007 23374 -5995
rect 23316 -6183 23328 -6007
rect 23362 -6183 23374 -6007
rect 23316 -6195 23374 -6183
rect 23434 -6007 23492 -5995
rect 24320 -5996 24378 -5984
rect 24438 -5808 24496 -5796
rect 24438 -5984 24450 -5808
rect 24484 -5984 24496 -5808
rect 24438 -5996 24496 -5984
rect 24740 -5808 24798 -5796
rect 23434 -6183 23446 -6007
rect 23480 -6183 23492 -6007
rect 23434 -6195 23492 -6183
rect 24740 -6184 24752 -5808
rect 24786 -6184 24798 -5808
rect 24740 -6196 24798 -6184
rect 24858 -5808 24916 -5796
rect 24858 -6184 24870 -5808
rect 24904 -6184 24916 -5808
rect 24858 -6196 24916 -6184
rect 24976 -5808 25034 -5796
rect 24976 -6184 24988 -5808
rect 25022 -6184 25034 -5808
rect 24976 -6196 25034 -6184
rect 25094 -5808 25152 -5796
rect 25094 -6184 25106 -5808
rect 25140 -6184 25152 -5808
rect 25094 -6196 25152 -6184
rect 25212 -5808 25270 -5796
rect 25212 -6184 25224 -5808
rect 25258 -6184 25270 -5808
rect 25618 -5808 25676 -5796
rect 25618 -5984 25630 -5808
rect 25664 -5984 25676 -5808
rect 25618 -5996 25676 -5984
rect 25736 -5808 25794 -5796
rect 25736 -5984 25748 -5808
rect 25782 -5984 25794 -5808
rect 25736 -5996 25794 -5984
rect 26218 -5808 26276 -5796
rect 26218 -5984 26230 -5808
rect 26264 -5984 26276 -5808
rect 26218 -5996 26276 -5984
rect 26336 -5808 26394 -5796
rect 26336 -5984 26348 -5808
rect 26382 -5984 26394 -5808
rect 26336 -5996 26394 -5984
rect 26638 -5808 26696 -5796
rect 25212 -6196 25270 -6184
rect 26638 -6184 26650 -5808
rect 26684 -6184 26696 -5808
rect 26638 -6196 26696 -6184
rect 26756 -5808 26814 -5796
rect 26756 -6184 26768 -5808
rect 26802 -6184 26814 -5808
rect 26756 -6196 26814 -6184
rect 26874 -5808 26932 -5796
rect 26874 -6184 26886 -5808
rect 26920 -6184 26932 -5808
rect 26874 -6196 26932 -6184
rect 26992 -5808 27050 -5796
rect 26992 -6184 27004 -5808
rect 27038 -6184 27050 -5808
rect 26992 -6196 27050 -6184
rect 27110 -5808 27168 -5796
rect 27110 -6184 27122 -5808
rect 27156 -6184 27168 -5808
rect 27516 -5808 27574 -5796
rect 27516 -5984 27528 -5808
rect 27562 -5984 27574 -5808
rect 27516 -5996 27574 -5984
rect 27634 -5808 27692 -5796
rect 27634 -5984 27646 -5808
rect 27680 -5984 27692 -5808
rect 28827 -5923 28839 -5547
rect 28873 -5923 28885 -5547
rect 28827 -5935 28885 -5923
rect 28945 -5547 29003 -5535
rect 28945 -5923 28957 -5547
rect 28991 -5923 29003 -5547
rect 28945 -5935 29003 -5923
rect 29063 -5547 29121 -5535
rect 29063 -5923 29075 -5547
rect 29109 -5923 29121 -5547
rect 29180 -5547 29238 -5535
rect 29180 -5723 29192 -5547
rect 29226 -5723 29238 -5547
rect 29180 -5735 29238 -5723
rect 29298 -5547 29356 -5535
rect 29298 -5723 29310 -5547
rect 29344 -5723 29356 -5547
rect 29298 -5735 29356 -5723
rect 29063 -5935 29121 -5923
rect 27634 -5996 27692 -5984
rect 27110 -6196 27168 -6184
rect 23199 -6395 23257 -6383
rect 6943 -7436 7001 -7424
rect 6943 -7812 6955 -7436
rect 6989 -7812 7001 -7436
rect 6943 -7824 7001 -7812
rect 7061 -7436 7119 -7424
rect 7061 -7812 7073 -7436
rect 7107 -7812 7119 -7436
rect 7061 -7824 7119 -7812
rect 7179 -7436 7237 -7424
rect 7179 -7812 7191 -7436
rect 7225 -7812 7237 -7436
rect 13497 -7431 13555 -7419
rect 7179 -7824 7237 -7812
rect 7296 -7636 7354 -7624
rect 7296 -7812 7308 -7636
rect 7342 -7812 7354 -7636
rect 7296 -7824 7354 -7812
rect 7414 -7636 7472 -7624
rect 7414 -7812 7426 -7636
rect 7460 -7812 7472 -7636
rect 7414 -7824 7472 -7812
rect 13497 -7807 13509 -7431
rect 13543 -7807 13555 -7431
rect 13497 -7819 13555 -7807
rect 13615 -7431 13673 -7419
rect 13615 -7807 13627 -7431
rect 13661 -7807 13673 -7431
rect 13615 -7819 13673 -7807
rect 13733 -7431 13791 -7419
rect 13733 -7807 13745 -7431
rect 13779 -7807 13791 -7431
rect 20146 -7443 20204 -7431
rect 13733 -7819 13791 -7807
rect 13850 -7631 13908 -7619
rect 13850 -7807 13862 -7631
rect 13896 -7807 13908 -7631
rect 13850 -7819 13908 -7807
rect 13968 -7631 14026 -7619
rect 13968 -7807 13980 -7631
rect 14014 -7807 14026 -7631
rect 13968 -7819 14026 -7807
rect 20146 -7819 20158 -7443
rect 20192 -7819 20204 -7443
rect 20146 -7831 20204 -7819
rect 20264 -7443 20322 -7431
rect 20264 -7819 20276 -7443
rect 20310 -7819 20322 -7443
rect 20264 -7831 20322 -7819
rect 20382 -7443 20440 -7431
rect 20382 -7819 20394 -7443
rect 20428 -7819 20440 -7443
rect 20382 -7831 20440 -7819
rect 20499 -7643 20557 -7631
rect 20499 -7819 20511 -7643
rect 20545 -7819 20557 -7643
rect 20499 -7831 20557 -7819
rect 20617 -7643 20675 -7631
rect 20617 -7819 20629 -7643
rect 20663 -7819 20675 -7643
rect 20617 -7831 20675 -7819
rect 32367 -7295 32425 -7283
rect 32367 -7671 32379 -7295
rect 32413 -7671 32425 -7295
rect 32367 -7683 32425 -7671
rect 32485 -7295 32543 -7283
rect 32485 -7671 32497 -7295
rect 32531 -7671 32543 -7295
rect 32485 -7683 32543 -7671
rect 32603 -7295 32661 -7283
rect 32603 -7671 32615 -7295
rect 32649 -7671 32661 -7295
rect 32720 -7295 32778 -7283
rect 32720 -7471 32732 -7295
rect 32766 -7471 32778 -7295
rect 32720 -7483 32778 -7471
rect 32838 -7295 32896 -7283
rect 32838 -7471 32850 -7295
rect 32884 -7471 32896 -7295
rect 32838 -7483 32896 -7471
rect 32603 -7683 32661 -7671
rect 30462 -8080 30520 -8068
rect 30462 -8256 30474 -8080
rect 30508 -8256 30520 -8080
rect 30462 -8268 30520 -8256
rect 30580 -8080 30638 -8068
rect 30580 -8256 30592 -8080
rect 30626 -8256 30638 -8080
rect 30580 -8268 30638 -8256
rect 30882 -8080 30940 -8068
rect 28834 -8392 28892 -8380
rect 28834 -8768 28846 -8392
rect 28880 -8768 28892 -8392
rect 28834 -8780 28892 -8768
rect 28952 -8392 29010 -8380
rect 28952 -8768 28964 -8392
rect 28998 -8768 29010 -8392
rect 28952 -8780 29010 -8768
rect 29070 -8392 29128 -8380
rect 29070 -8768 29082 -8392
rect 29116 -8768 29128 -8392
rect 29187 -8392 29245 -8380
rect 29187 -8568 29199 -8392
rect 29233 -8568 29245 -8392
rect 29187 -8580 29245 -8568
rect 29305 -8392 29363 -8380
rect 29305 -8568 29317 -8392
rect 29351 -8568 29363 -8392
rect 30882 -8456 30894 -8080
rect 30928 -8456 30940 -8080
rect 30882 -8468 30940 -8456
rect 31000 -8080 31058 -8068
rect 31000 -8456 31012 -8080
rect 31046 -8456 31058 -8080
rect 31000 -8468 31058 -8456
rect 31118 -8080 31176 -8068
rect 31118 -8456 31130 -8080
rect 31164 -8456 31176 -8080
rect 31118 -8468 31176 -8456
rect 31236 -8080 31294 -8068
rect 31236 -8456 31248 -8080
rect 31282 -8456 31294 -8080
rect 31236 -8468 31294 -8456
rect 31354 -8080 31412 -8068
rect 31354 -8456 31366 -8080
rect 31400 -8456 31412 -8080
rect 31760 -8080 31818 -8068
rect 31760 -8256 31772 -8080
rect 31806 -8256 31818 -8080
rect 31760 -8268 31818 -8256
rect 31878 -8080 31936 -8068
rect 31878 -8256 31890 -8080
rect 31924 -8256 31936 -8080
rect 31878 -8268 31936 -8256
rect 31354 -8468 31412 -8456
rect 29305 -8580 29363 -8568
rect 29070 -8780 29128 -8768
<< pdiff >>
rect 6671 5631 6729 5643
rect 6671 5455 6683 5631
rect 6717 5455 6729 5631
rect 6671 5443 6729 5455
rect 6789 5631 6847 5643
rect 6789 5455 6801 5631
rect 6835 5455 6847 5631
rect 6789 5443 6847 5455
rect 6907 5631 6965 5643
rect 6907 5455 6919 5631
rect 6953 5455 6965 5631
rect 6907 5443 6965 5455
rect 7025 5631 7083 5643
rect 7025 5455 7037 5631
rect 7071 5455 7083 5631
rect 7025 5443 7083 5455
rect 7143 5631 7201 5643
rect 7143 5455 7155 5631
rect 7189 5455 7201 5631
rect 7143 5443 7201 5455
rect 7261 5631 7319 5643
rect 7261 5455 7273 5631
rect 7307 5455 7319 5631
rect 7261 5443 7319 5455
rect 7379 5631 7437 5643
rect 7379 5455 7391 5631
rect 7425 5455 7437 5631
rect 7379 5443 7437 5455
rect 7497 5631 7555 5643
rect 7497 5455 7509 5631
rect 7543 5455 7555 5631
rect 7497 5443 7555 5455
rect 7615 5631 7673 5643
rect 7615 5455 7627 5631
rect 7661 5455 7673 5631
rect 7615 5443 7673 5455
rect 7733 5631 7791 5643
rect 19874 5651 19932 5663
rect 7733 5455 7745 5631
rect 7779 5455 7791 5631
rect 7733 5443 7791 5455
rect 13220 5630 13278 5642
rect 13220 5454 13232 5630
rect 13266 5454 13278 5630
rect 13220 5442 13278 5454
rect 13338 5630 13396 5642
rect 13338 5454 13350 5630
rect 13384 5454 13396 5630
rect 13338 5442 13396 5454
rect 13456 5630 13514 5642
rect 13456 5454 13468 5630
rect 13502 5454 13514 5630
rect 13456 5442 13514 5454
rect 13574 5630 13632 5642
rect 13574 5454 13586 5630
rect 13620 5454 13632 5630
rect 13574 5442 13632 5454
rect 13692 5630 13750 5642
rect 13692 5454 13704 5630
rect 13738 5454 13750 5630
rect 13692 5442 13750 5454
rect 13810 5630 13868 5642
rect 13810 5454 13822 5630
rect 13856 5454 13868 5630
rect 13810 5442 13868 5454
rect 13928 5630 13986 5642
rect 13928 5454 13940 5630
rect 13974 5454 13986 5630
rect 13928 5442 13986 5454
rect 14046 5630 14104 5642
rect 14046 5454 14058 5630
rect 14092 5454 14104 5630
rect 14046 5442 14104 5454
rect 14164 5630 14222 5642
rect 14164 5454 14176 5630
rect 14210 5454 14222 5630
rect 14164 5442 14222 5454
rect 14282 5630 14340 5642
rect 14282 5454 14294 5630
rect 14328 5454 14340 5630
rect 19874 5475 19886 5651
rect 19920 5475 19932 5651
rect 19874 5463 19932 5475
rect 19992 5651 20050 5663
rect 19992 5475 20004 5651
rect 20038 5475 20050 5651
rect 19992 5463 20050 5475
rect 20110 5651 20168 5663
rect 20110 5475 20122 5651
rect 20156 5475 20168 5651
rect 20110 5463 20168 5475
rect 20228 5651 20286 5663
rect 20228 5475 20240 5651
rect 20274 5475 20286 5651
rect 20228 5463 20286 5475
rect 20346 5651 20404 5663
rect 20346 5475 20358 5651
rect 20392 5475 20404 5651
rect 20346 5463 20404 5475
rect 20464 5651 20522 5663
rect 20464 5475 20476 5651
rect 20510 5475 20522 5651
rect 20464 5463 20522 5475
rect 20582 5651 20640 5663
rect 20582 5475 20594 5651
rect 20628 5475 20640 5651
rect 20582 5463 20640 5475
rect 20700 5651 20758 5663
rect 20700 5475 20712 5651
rect 20746 5475 20758 5651
rect 20700 5463 20758 5475
rect 20818 5651 20876 5663
rect 20818 5475 20830 5651
rect 20864 5475 20876 5651
rect 20818 5463 20876 5475
rect 20936 5651 20994 5663
rect 20936 5475 20948 5651
rect 20982 5475 20994 5651
rect 20936 5463 20994 5475
rect 28527 5484 28585 5496
rect 14282 5442 14340 5454
rect 28527 5308 28539 5484
rect 28573 5308 28585 5484
rect 28527 5296 28585 5308
rect 28645 5484 28703 5496
rect 28645 5308 28657 5484
rect 28691 5308 28703 5484
rect 28645 5296 28703 5308
rect 28763 5484 28821 5496
rect 28763 5308 28775 5484
rect 28809 5308 28821 5484
rect 28763 5296 28821 5308
rect 28881 5484 28939 5496
rect 28881 5308 28893 5484
rect 28927 5308 28939 5484
rect 28881 5296 28939 5308
rect 28999 5484 29057 5496
rect 28999 5308 29011 5484
rect 29045 5308 29057 5484
rect 28999 5296 29057 5308
rect 29117 5484 29175 5496
rect 29117 5308 29129 5484
rect 29163 5308 29175 5484
rect 29117 5296 29175 5308
rect 29235 5484 29293 5496
rect 29235 5308 29247 5484
rect 29281 5308 29293 5484
rect 29235 5296 29293 5308
rect 29353 5484 29411 5496
rect 29353 5308 29365 5484
rect 29399 5308 29411 5484
rect 29353 5296 29411 5308
rect 29471 5484 29529 5496
rect 29471 5308 29483 5484
rect 29517 5308 29529 5484
rect 29471 5296 29529 5308
rect 29589 5484 29647 5496
rect 29589 5308 29601 5484
rect 29635 5308 29647 5484
rect 29589 5296 29647 5308
rect 30819 5279 30877 5291
rect 30335 5079 30393 5091
rect 30335 4903 30347 5079
rect 30381 4903 30393 5079
rect 30335 4891 30393 4903
rect 30453 5079 30511 5091
rect 30453 4903 30465 5079
rect 30499 4903 30511 5079
rect 30453 4891 30511 4903
rect 30571 5079 30629 5091
rect 30571 4903 30583 5079
rect 30617 4903 30629 5079
rect 30571 4891 30629 4903
rect 30689 5079 30747 5091
rect 30689 4903 30701 5079
rect 30735 4903 30747 5079
rect 30689 4891 30747 4903
rect 30819 4903 30831 5279
rect 30865 4903 30877 5279
rect 30819 4891 30877 4903
rect 30937 5279 30995 5291
rect 30937 4903 30949 5279
rect 30983 4903 30995 5279
rect 30937 4891 30995 4903
rect 31055 5279 31113 5291
rect 31055 4903 31067 5279
rect 31101 4903 31113 5279
rect 31055 4891 31113 4903
rect 31173 5279 31231 5291
rect 31173 4903 31185 5279
rect 31219 4903 31231 5279
rect 31173 4891 31231 4903
rect 31291 5279 31349 5291
rect 31291 4903 31303 5279
rect 31337 4903 31349 5279
rect 31291 4891 31349 4903
rect 31409 5279 31467 5291
rect 31409 4903 31421 5279
rect 31455 4903 31467 5279
rect 31409 4891 31467 4903
rect 31527 5279 31585 5291
rect 31527 4903 31539 5279
rect 31573 4903 31585 5279
rect 31527 4891 31585 4903
rect 31656 5079 31714 5091
rect 31656 4903 31668 5079
rect 31702 4903 31714 5079
rect 31656 4891 31714 4903
rect 31774 5079 31832 5091
rect 31774 4903 31786 5079
rect 31820 4903 31832 5079
rect 31774 4891 31832 4903
rect 31892 5079 31950 5091
rect 31892 4903 31904 5079
rect 31938 4903 31950 5079
rect 31892 4891 31950 4903
rect 32010 5079 32068 5091
rect 32010 4903 32022 5079
rect 32056 4903 32068 5079
rect 32010 4891 32068 4903
rect 32128 5076 32186 5088
rect 32128 4900 32140 5076
rect 32174 4900 32186 5076
rect 32128 4888 32186 4900
rect 32246 5076 32304 5088
rect 32246 4900 32258 5076
rect 32292 4900 32304 5076
rect 32246 4888 32304 4900
rect 32364 5076 32422 5088
rect 32364 4900 32376 5076
rect 32410 4900 32422 5076
rect 32364 4888 32422 4900
rect 32482 5076 32540 5088
rect 32482 4900 32494 5076
rect 32528 4900 32540 5076
rect 32482 4888 32540 4900
rect 32600 5076 32658 5088
rect 32600 4900 32612 5076
rect 32646 4900 32658 5076
rect 32600 4888 32658 4900
rect 32718 5076 32776 5088
rect 32718 4900 32730 5076
rect 32764 4900 32776 5076
rect 32718 4888 32776 4900
rect 32836 5076 32894 5088
rect 32836 4900 32848 5076
rect 32882 4900 32894 5076
rect 32836 4888 32894 4900
rect 32954 5076 33012 5088
rect 32954 4900 32966 5076
rect 33000 4900 33012 5076
rect 32954 4888 33012 4900
rect 33072 5076 33130 5088
rect 33072 4900 33084 5076
rect 33118 4900 33130 5076
rect 33072 4888 33130 4900
rect 33190 5076 33248 5088
rect 33190 4900 33202 5076
rect 33236 4900 33248 5076
rect 33190 4888 33248 4900
rect 30762 4586 30820 4598
rect 7 3731 65 3743
rect 7 3555 19 3731
rect 53 3555 65 3731
rect 7 3543 65 3555
rect 125 3731 183 3743
rect 125 3555 137 3731
rect 171 3555 183 3731
rect 125 3543 183 3555
rect 243 3731 301 3743
rect 243 3555 255 3731
rect 289 3555 301 3731
rect 243 3543 301 3555
rect 361 3731 419 3743
rect 361 3555 373 3731
rect 407 3555 419 3731
rect 361 3543 419 3555
rect 479 3731 537 3743
rect 479 3555 491 3731
rect 525 3555 537 3731
rect 479 3543 537 3555
rect 597 3731 655 3743
rect 597 3555 609 3731
rect 643 3555 655 3731
rect 597 3543 655 3555
rect 715 3731 773 3743
rect 715 3555 727 3731
rect 761 3555 773 3731
rect 715 3543 773 3555
rect 833 3731 891 3743
rect 833 3555 845 3731
rect 879 3555 891 3731
rect 833 3543 891 3555
rect 951 3731 1009 3743
rect 951 3555 963 3731
rect 997 3555 1009 3731
rect 951 3543 1009 3555
rect 1069 3731 1127 3743
rect 1069 3555 1081 3731
rect 1115 3555 1127 3731
rect 30762 4210 30774 4586
rect 30808 4210 30820 4586
rect 30762 4198 30820 4210
rect 30880 4586 30938 4598
rect 30880 4210 30892 4586
rect 30926 4210 30938 4586
rect 30880 4198 30938 4210
rect 30998 4586 31056 4598
rect 30998 4210 31010 4586
rect 31044 4210 31056 4586
rect 30998 4198 31056 4210
rect 31116 4586 31174 4598
rect 31116 4210 31128 4586
rect 31162 4210 31174 4586
rect 31116 4198 31174 4210
rect 31234 4586 31292 4598
rect 31234 4210 31246 4586
rect 31280 4210 31292 4586
rect 31234 4198 31292 4210
rect 31352 4586 31410 4598
rect 31352 4210 31364 4586
rect 31398 4210 31410 4586
rect 31352 4198 31410 4210
rect 31470 4586 31528 4598
rect 31470 4210 31482 4586
rect 31516 4210 31528 4586
rect 31470 4198 31528 4210
rect 11771 3624 11829 3636
rect 1069 3543 1127 3555
rect 9446 3552 9504 3564
rect 5222 3536 5280 3548
rect 2897 3464 2955 3476
rect 2897 3288 2909 3464
rect 2943 3288 2955 3464
rect 2897 3276 2955 3288
rect 3015 3464 3073 3476
rect 3015 3288 3027 3464
rect 3061 3288 3073 3464
rect 3015 3276 3073 3288
rect 3133 3464 3191 3476
rect 3133 3288 3145 3464
rect 3179 3288 3191 3464
rect 3133 3276 3191 3288
rect 3251 3464 3309 3476
rect 3251 3288 3263 3464
rect 3297 3288 3309 3464
rect 3251 3276 3309 3288
rect 3369 3464 3427 3476
rect 3369 3288 3381 3464
rect 3415 3288 3427 3464
rect 3369 3276 3427 3288
rect 3487 3464 3545 3476
rect 3487 3288 3499 3464
rect 3533 3288 3545 3464
rect 3487 3276 3545 3288
rect 3605 3464 3663 3476
rect 3605 3288 3617 3464
rect 3651 3288 3663 3464
rect 3605 3276 3663 3288
rect 3723 3464 3781 3476
rect 3723 3288 3735 3464
rect 3769 3288 3781 3464
rect 3723 3276 3781 3288
rect 3841 3464 3899 3476
rect 3841 3288 3853 3464
rect 3887 3288 3899 3464
rect 3841 3276 3899 3288
rect 3959 3464 4017 3476
rect 3959 3288 3971 3464
rect 4005 3288 4017 3464
rect 3959 3276 4017 3288
rect 5222 3160 5234 3536
rect 5268 3160 5280 3536
rect 5222 3148 5280 3160
rect 5340 3536 5398 3548
rect 5340 3160 5352 3536
rect 5386 3160 5398 3536
rect 5340 3148 5398 3160
rect 5458 3536 5516 3548
rect 5458 3160 5470 3536
rect 5504 3160 5516 3536
rect 5458 3148 5516 3160
rect 5576 3536 5634 3548
rect 5576 3160 5588 3536
rect 5622 3160 5634 3536
rect 5576 3148 5634 3160
rect 5694 3536 5752 3548
rect 5694 3160 5706 3536
rect 5740 3160 5752 3536
rect 5694 3148 5752 3160
rect 5812 3536 5870 3548
rect 5812 3160 5824 3536
rect 5858 3160 5870 3536
rect 5812 3148 5870 3160
rect 5930 3536 5988 3548
rect 5930 3160 5942 3536
rect 5976 3160 5988 3536
rect 5930 3148 5988 3160
rect 6364 3540 6422 3552
rect 6364 3164 6376 3540
rect 6410 3164 6422 3540
rect 6364 3152 6422 3164
rect 6482 3540 6540 3552
rect 6482 3164 6494 3540
rect 6528 3164 6540 3540
rect 6482 3152 6540 3164
rect 6600 3540 6658 3552
rect 6600 3164 6612 3540
rect 6646 3164 6658 3540
rect 6600 3152 6658 3164
rect 6718 3540 6776 3552
rect 6718 3164 6730 3540
rect 6764 3164 6776 3540
rect 6718 3152 6776 3164
rect 6836 3540 6894 3552
rect 6836 3164 6848 3540
rect 6882 3164 6894 3540
rect 6836 3152 6894 3164
rect 6954 3540 7012 3552
rect 6954 3164 6966 3540
rect 7000 3164 7012 3540
rect 6954 3152 7012 3164
rect 7072 3540 7130 3552
rect 7072 3164 7084 3540
rect 7118 3164 7130 3540
rect 9446 3376 9458 3552
rect 9492 3376 9504 3552
rect 9446 3364 9504 3376
rect 9564 3552 9622 3564
rect 9564 3376 9576 3552
rect 9610 3376 9622 3552
rect 9564 3364 9622 3376
rect 9682 3552 9740 3564
rect 9682 3376 9694 3552
rect 9728 3376 9740 3552
rect 9682 3364 9740 3376
rect 9800 3552 9858 3564
rect 9800 3376 9812 3552
rect 9846 3376 9858 3552
rect 9800 3364 9858 3376
rect 9918 3552 9976 3564
rect 9918 3376 9930 3552
rect 9964 3376 9976 3552
rect 9918 3364 9976 3376
rect 10036 3552 10094 3564
rect 10036 3376 10048 3552
rect 10082 3376 10094 3552
rect 10036 3364 10094 3376
rect 10154 3552 10212 3564
rect 10154 3376 10166 3552
rect 10200 3376 10212 3552
rect 10154 3364 10212 3376
rect 10272 3552 10330 3564
rect 10272 3376 10284 3552
rect 10318 3376 10330 3552
rect 10272 3364 10330 3376
rect 10390 3552 10448 3564
rect 10390 3376 10402 3552
rect 10436 3376 10448 3552
rect 10390 3364 10448 3376
rect 10508 3552 10566 3564
rect 10508 3376 10520 3552
rect 10554 3376 10566 3552
rect 10508 3364 10566 3376
rect 7072 3152 7130 3164
rect 11771 3248 11783 3624
rect 11817 3248 11829 3624
rect 11771 3236 11829 3248
rect 11889 3624 11947 3636
rect 11889 3248 11901 3624
rect 11935 3248 11947 3624
rect 11889 3236 11947 3248
rect 12007 3624 12065 3636
rect 12007 3248 12019 3624
rect 12053 3248 12065 3624
rect 12007 3236 12065 3248
rect 12125 3624 12183 3636
rect 12125 3248 12137 3624
rect 12171 3248 12183 3624
rect 12125 3236 12183 3248
rect 12243 3624 12301 3636
rect 12243 3248 12255 3624
rect 12289 3248 12301 3624
rect 12243 3236 12301 3248
rect 12361 3624 12419 3636
rect 12361 3248 12373 3624
rect 12407 3248 12419 3624
rect 12361 3236 12419 3248
rect 12479 3624 12537 3636
rect 12479 3248 12491 3624
rect 12525 3248 12537 3624
rect 12479 3236 12537 3248
rect 12913 3628 12971 3640
rect 12913 3252 12925 3628
rect 12959 3252 12971 3628
rect 12913 3240 12971 3252
rect 13031 3628 13089 3640
rect 13031 3252 13043 3628
rect 13077 3252 13089 3628
rect 13031 3240 13089 3252
rect 13149 3628 13207 3640
rect 13149 3252 13161 3628
rect 13195 3252 13207 3628
rect 13149 3240 13207 3252
rect 13267 3628 13325 3640
rect 13267 3252 13279 3628
rect 13313 3252 13325 3628
rect 13267 3240 13325 3252
rect 13385 3628 13443 3640
rect 13385 3252 13397 3628
rect 13431 3252 13443 3628
rect 13385 3240 13443 3252
rect 13503 3628 13561 3640
rect 13503 3252 13515 3628
rect 13549 3252 13561 3628
rect 13503 3240 13561 3252
rect 13621 3628 13679 3640
rect 13621 3252 13633 3628
rect 13667 3252 13679 3628
rect 25050 3624 25108 3636
rect 18425 3556 18483 3568
rect 16100 3484 16158 3496
rect 16100 3308 16112 3484
rect 16146 3308 16158 3484
rect 16100 3296 16158 3308
rect 16218 3484 16276 3496
rect 16218 3308 16230 3484
rect 16264 3308 16276 3484
rect 16218 3296 16276 3308
rect 16336 3484 16394 3496
rect 16336 3308 16348 3484
rect 16382 3308 16394 3484
rect 16336 3296 16394 3308
rect 16454 3484 16512 3496
rect 16454 3308 16466 3484
rect 16500 3308 16512 3484
rect 16454 3296 16512 3308
rect 16572 3484 16630 3496
rect 16572 3308 16584 3484
rect 16618 3308 16630 3484
rect 16572 3296 16630 3308
rect 16690 3484 16748 3496
rect 16690 3308 16702 3484
rect 16736 3308 16748 3484
rect 16690 3296 16748 3308
rect 16808 3484 16866 3496
rect 16808 3308 16820 3484
rect 16854 3308 16866 3484
rect 16808 3296 16866 3308
rect 16926 3484 16984 3496
rect 16926 3308 16938 3484
rect 16972 3308 16984 3484
rect 16926 3296 16984 3308
rect 17044 3484 17102 3496
rect 17044 3308 17056 3484
rect 17090 3308 17102 3484
rect 17044 3296 17102 3308
rect 17162 3484 17220 3496
rect 17162 3308 17174 3484
rect 17208 3308 17220 3484
rect 17162 3296 17220 3308
rect 13621 3240 13679 3252
rect 5651 2753 5709 2765
rect 5651 2577 5663 2753
rect 5697 2577 5709 2753
rect 5651 2565 5709 2577
rect 5769 2753 5827 2765
rect 5769 2577 5781 2753
rect 5815 2577 5827 2753
rect 5769 2565 5827 2577
rect 5887 2753 5945 2765
rect 5887 2577 5899 2753
rect 5933 2577 5945 2753
rect 5887 2565 5945 2577
rect 6005 2753 6063 2765
rect 6005 2577 6017 2753
rect 6051 2577 6063 2753
rect 6005 2565 6063 2577
rect 6793 2757 6851 2769
rect 6793 2581 6805 2757
rect 6839 2581 6851 2757
rect 6793 2569 6851 2581
rect 6911 2757 6969 2769
rect 6911 2581 6923 2757
rect 6957 2581 6969 2757
rect 6911 2569 6969 2581
rect 7029 2757 7087 2769
rect 7029 2581 7041 2757
rect 7075 2581 7087 2757
rect 7029 2569 7087 2581
rect 7147 2757 7205 2769
rect 7147 2581 7159 2757
rect 7193 2581 7205 2757
rect 18425 3180 18437 3556
rect 18471 3180 18483 3556
rect 18425 3168 18483 3180
rect 18543 3556 18601 3568
rect 18543 3180 18555 3556
rect 18589 3180 18601 3556
rect 18543 3168 18601 3180
rect 18661 3556 18719 3568
rect 18661 3180 18673 3556
rect 18707 3180 18719 3556
rect 18661 3168 18719 3180
rect 18779 3556 18837 3568
rect 18779 3180 18791 3556
rect 18825 3180 18837 3556
rect 18779 3168 18837 3180
rect 18897 3556 18955 3568
rect 18897 3180 18909 3556
rect 18943 3180 18955 3556
rect 18897 3168 18955 3180
rect 19015 3556 19073 3568
rect 19015 3180 19027 3556
rect 19061 3180 19073 3556
rect 19015 3168 19073 3180
rect 19133 3556 19191 3568
rect 19133 3180 19145 3556
rect 19179 3180 19191 3556
rect 19133 3168 19191 3180
rect 19567 3560 19625 3572
rect 19567 3184 19579 3560
rect 19613 3184 19625 3560
rect 19567 3172 19625 3184
rect 19685 3560 19743 3572
rect 19685 3184 19697 3560
rect 19731 3184 19743 3560
rect 19685 3172 19743 3184
rect 19803 3560 19861 3572
rect 19803 3184 19815 3560
rect 19849 3184 19861 3560
rect 19803 3172 19861 3184
rect 19921 3560 19979 3572
rect 19921 3184 19933 3560
rect 19967 3184 19979 3560
rect 19921 3172 19979 3184
rect 20039 3560 20097 3572
rect 20039 3184 20051 3560
rect 20085 3184 20097 3560
rect 20039 3172 20097 3184
rect 20157 3560 20215 3572
rect 20157 3184 20169 3560
rect 20203 3184 20215 3560
rect 20157 3172 20215 3184
rect 20275 3560 20333 3572
rect 20275 3184 20287 3560
rect 20321 3184 20333 3560
rect 22725 3552 22783 3564
rect 22725 3376 22737 3552
rect 22771 3376 22783 3552
rect 22725 3364 22783 3376
rect 22843 3552 22901 3564
rect 22843 3376 22855 3552
rect 22889 3376 22901 3552
rect 22843 3364 22901 3376
rect 22961 3552 23019 3564
rect 22961 3376 22973 3552
rect 23007 3376 23019 3552
rect 22961 3364 23019 3376
rect 23079 3552 23137 3564
rect 23079 3376 23091 3552
rect 23125 3376 23137 3552
rect 23079 3364 23137 3376
rect 23197 3552 23255 3564
rect 23197 3376 23209 3552
rect 23243 3376 23255 3552
rect 23197 3364 23255 3376
rect 23315 3552 23373 3564
rect 23315 3376 23327 3552
rect 23361 3376 23373 3552
rect 23315 3364 23373 3376
rect 23433 3552 23491 3564
rect 23433 3376 23445 3552
rect 23479 3376 23491 3552
rect 23433 3364 23491 3376
rect 23551 3552 23609 3564
rect 23551 3376 23563 3552
rect 23597 3376 23609 3552
rect 23551 3364 23609 3376
rect 23669 3552 23727 3564
rect 23669 3376 23681 3552
rect 23715 3376 23727 3552
rect 23669 3364 23727 3376
rect 23787 3552 23845 3564
rect 23787 3376 23799 3552
rect 23833 3376 23845 3552
rect 23787 3364 23845 3376
rect 20275 3172 20333 3184
rect 12200 2841 12258 2853
rect 12200 2665 12212 2841
rect 12246 2665 12258 2841
rect 12200 2653 12258 2665
rect 12318 2841 12376 2853
rect 12318 2665 12330 2841
rect 12364 2665 12376 2841
rect 12318 2653 12376 2665
rect 12436 2841 12494 2853
rect 12436 2665 12448 2841
rect 12482 2665 12494 2841
rect 12436 2653 12494 2665
rect 12554 2841 12612 2853
rect 12554 2665 12566 2841
rect 12600 2665 12612 2841
rect 12554 2653 12612 2665
rect 13342 2845 13400 2857
rect 13342 2669 13354 2845
rect 13388 2669 13400 2845
rect 13342 2657 13400 2669
rect 13460 2845 13518 2857
rect 13460 2669 13472 2845
rect 13506 2669 13518 2845
rect 13460 2657 13518 2669
rect 13578 2845 13636 2857
rect 13578 2669 13590 2845
rect 13624 2669 13636 2845
rect 13578 2657 13636 2669
rect 13696 2845 13754 2857
rect 13696 2669 13708 2845
rect 13742 2669 13754 2845
rect 13696 2657 13754 2669
rect 25050 3248 25062 3624
rect 25096 3248 25108 3624
rect 25050 3236 25108 3248
rect 25168 3624 25226 3636
rect 25168 3248 25180 3624
rect 25214 3248 25226 3624
rect 25168 3236 25226 3248
rect 25286 3624 25344 3636
rect 25286 3248 25298 3624
rect 25332 3248 25344 3624
rect 25286 3236 25344 3248
rect 25404 3624 25462 3636
rect 25404 3248 25416 3624
rect 25450 3248 25462 3624
rect 25404 3236 25462 3248
rect 25522 3624 25580 3636
rect 25522 3248 25534 3624
rect 25568 3248 25580 3624
rect 25522 3236 25580 3248
rect 25640 3624 25698 3636
rect 25640 3248 25652 3624
rect 25686 3248 25698 3624
rect 25640 3236 25698 3248
rect 25758 3624 25816 3636
rect 25758 3248 25770 3624
rect 25804 3248 25816 3624
rect 25758 3236 25816 3248
rect 26192 3628 26250 3640
rect 26192 3252 26204 3628
rect 26238 3252 26250 3628
rect 26192 3240 26250 3252
rect 26310 3628 26368 3640
rect 26310 3252 26322 3628
rect 26356 3252 26368 3628
rect 26310 3240 26368 3252
rect 26428 3628 26486 3640
rect 26428 3252 26440 3628
rect 26474 3252 26486 3628
rect 26428 3240 26486 3252
rect 26546 3628 26604 3640
rect 26546 3252 26558 3628
rect 26592 3252 26604 3628
rect 26546 3240 26604 3252
rect 26664 3628 26722 3640
rect 26664 3252 26676 3628
rect 26710 3252 26722 3628
rect 26664 3240 26722 3252
rect 26782 3628 26840 3640
rect 26782 3252 26794 3628
rect 26828 3252 26840 3628
rect 26782 3240 26840 3252
rect 26900 3628 26958 3640
rect 26900 3252 26912 3628
rect 26946 3252 26958 3628
rect 26900 3240 26958 3252
rect 7147 2569 7205 2581
rect 18854 2773 18912 2785
rect 18854 2597 18866 2773
rect 18900 2597 18912 2773
rect 18854 2585 18912 2597
rect 18972 2773 19030 2785
rect 18972 2597 18984 2773
rect 19018 2597 19030 2773
rect 18972 2585 19030 2597
rect 19090 2773 19148 2785
rect 19090 2597 19102 2773
rect 19136 2597 19148 2773
rect 19090 2585 19148 2597
rect 19208 2773 19266 2785
rect 19208 2597 19220 2773
rect 19254 2597 19266 2773
rect 19208 2585 19266 2597
rect 19996 2777 20054 2789
rect 19996 2601 20008 2777
rect 20042 2601 20054 2777
rect 19996 2589 20054 2601
rect 20114 2777 20172 2789
rect 20114 2601 20126 2777
rect 20160 2601 20172 2777
rect 20114 2589 20172 2601
rect 20232 2777 20290 2789
rect 20232 2601 20244 2777
rect 20278 2601 20290 2777
rect 20232 2589 20290 2601
rect 20350 2777 20408 2789
rect 20350 2601 20362 2777
rect 20396 2601 20408 2777
rect 28522 2913 28580 2925
rect 25479 2841 25537 2853
rect 25479 2665 25491 2841
rect 25525 2665 25537 2841
rect 25479 2653 25537 2665
rect 25597 2841 25655 2853
rect 25597 2665 25609 2841
rect 25643 2665 25655 2841
rect 25597 2653 25655 2665
rect 25715 2841 25773 2853
rect 25715 2665 25727 2841
rect 25761 2665 25773 2841
rect 25715 2653 25773 2665
rect 25833 2841 25891 2853
rect 25833 2665 25845 2841
rect 25879 2665 25891 2841
rect 25833 2653 25891 2665
rect 26621 2845 26679 2857
rect 26621 2669 26633 2845
rect 26667 2669 26679 2845
rect 26621 2657 26679 2669
rect 26739 2845 26797 2857
rect 26739 2669 26751 2845
rect 26785 2669 26797 2845
rect 26739 2657 26797 2669
rect 26857 2845 26915 2857
rect 26857 2669 26869 2845
rect 26903 2669 26915 2845
rect 26857 2657 26915 2669
rect 26975 2845 27033 2857
rect 26975 2669 26987 2845
rect 27021 2669 27033 2845
rect 28522 2737 28534 2913
rect 28568 2737 28580 2913
rect 28522 2725 28580 2737
rect 28640 2913 28698 2925
rect 28640 2737 28652 2913
rect 28686 2737 28698 2913
rect 28640 2725 28698 2737
rect 28758 2913 28816 2925
rect 28758 2737 28770 2913
rect 28804 2737 28816 2913
rect 28758 2725 28816 2737
rect 28876 2913 28934 2925
rect 28876 2737 28888 2913
rect 28922 2737 28934 2913
rect 28876 2725 28934 2737
rect 28994 2913 29052 2925
rect 28994 2737 29006 2913
rect 29040 2737 29052 2913
rect 28994 2725 29052 2737
rect 29112 2913 29170 2925
rect 29112 2737 29124 2913
rect 29158 2737 29170 2913
rect 29112 2725 29170 2737
rect 29230 2913 29288 2925
rect 29230 2737 29242 2913
rect 29276 2737 29288 2913
rect 29230 2725 29288 2737
rect 29348 2913 29406 2925
rect 29348 2737 29360 2913
rect 29394 2737 29406 2913
rect 29348 2725 29406 2737
rect 29466 2913 29524 2925
rect 29466 2737 29478 2913
rect 29512 2737 29524 2913
rect 29466 2725 29524 2737
rect 29584 2913 29642 2925
rect 29584 2737 29596 2913
rect 29630 2737 29642 2913
rect 29584 2725 29642 2737
rect 26975 2657 27033 2669
rect 20350 2589 20408 2601
rect 2911 1814 2969 1826
rect 2911 1638 2923 1814
rect 2957 1638 2969 1814
rect 2911 1626 2969 1638
rect 3029 1814 3087 1826
rect 3029 1638 3041 1814
rect 3075 1638 3087 1814
rect 3029 1626 3087 1638
rect 3147 1814 3205 1826
rect 3147 1638 3159 1814
rect 3193 1638 3205 1814
rect 3147 1626 3205 1638
rect 3265 1814 3323 1826
rect 3265 1638 3277 1814
rect 3311 1638 3323 1814
rect 3265 1626 3323 1638
rect 3383 1814 3441 1826
rect 3383 1638 3395 1814
rect 3429 1638 3441 1814
rect 3383 1626 3441 1638
rect 3501 1814 3559 1826
rect 3501 1638 3513 1814
rect 3547 1638 3559 1814
rect 3501 1626 3559 1638
rect 3619 1814 3677 1826
rect 3619 1638 3631 1814
rect 3665 1638 3677 1814
rect 3619 1626 3677 1638
rect 3737 1814 3795 1826
rect 3737 1638 3749 1814
rect 3783 1638 3795 1814
rect 3737 1626 3795 1638
rect 3855 1814 3913 1826
rect 3855 1638 3867 1814
rect 3901 1638 3913 1814
rect 3855 1626 3913 1638
rect 3973 1814 4031 1826
rect 3973 1638 3985 1814
rect 4019 1638 4031 1814
rect 9460 1902 9518 1914
rect 9460 1726 9472 1902
rect 9506 1726 9518 1902
rect 9460 1714 9518 1726
rect 9578 1902 9636 1914
rect 9578 1726 9590 1902
rect 9624 1726 9636 1902
rect 9578 1714 9636 1726
rect 9696 1902 9754 1914
rect 9696 1726 9708 1902
rect 9742 1726 9754 1902
rect 9696 1714 9754 1726
rect 9814 1902 9872 1914
rect 9814 1726 9826 1902
rect 9860 1726 9872 1902
rect 9814 1714 9872 1726
rect 9932 1902 9990 1914
rect 9932 1726 9944 1902
rect 9978 1726 9990 1902
rect 9932 1714 9990 1726
rect 10050 1902 10108 1914
rect 10050 1726 10062 1902
rect 10096 1726 10108 1902
rect 10050 1714 10108 1726
rect 10168 1902 10226 1914
rect 10168 1726 10180 1902
rect 10214 1726 10226 1902
rect 10168 1714 10226 1726
rect 10286 1902 10344 1914
rect 10286 1726 10298 1902
rect 10332 1726 10344 1902
rect 10286 1714 10344 1726
rect 10404 1902 10462 1914
rect 10404 1726 10416 1902
rect 10450 1726 10462 1902
rect 10404 1714 10462 1726
rect 10522 1902 10580 1914
rect 10522 1726 10534 1902
rect 10568 1726 10580 1902
rect 16114 1834 16172 1846
rect 10522 1714 10580 1726
rect 3973 1626 4031 1638
rect 16114 1658 16126 1834
rect 16160 1658 16172 1834
rect 16114 1646 16172 1658
rect 16232 1834 16290 1846
rect 16232 1658 16244 1834
rect 16278 1658 16290 1834
rect 16232 1646 16290 1658
rect 16350 1834 16408 1846
rect 16350 1658 16362 1834
rect 16396 1658 16408 1834
rect 16350 1646 16408 1658
rect 16468 1834 16526 1846
rect 16468 1658 16480 1834
rect 16514 1658 16526 1834
rect 16468 1646 16526 1658
rect 16586 1834 16644 1846
rect 16586 1658 16598 1834
rect 16632 1658 16644 1834
rect 16586 1646 16644 1658
rect 16704 1834 16762 1846
rect 16704 1658 16716 1834
rect 16750 1658 16762 1834
rect 16704 1646 16762 1658
rect 16822 1834 16880 1846
rect 16822 1658 16834 1834
rect 16868 1658 16880 1834
rect 16822 1646 16880 1658
rect 16940 1834 16998 1846
rect 16940 1658 16952 1834
rect 16986 1658 16998 1834
rect 16940 1646 16998 1658
rect 17058 1834 17116 1846
rect 17058 1658 17070 1834
rect 17104 1658 17116 1834
rect 17058 1646 17116 1658
rect 17176 1834 17234 1846
rect 17176 1658 17188 1834
rect 17222 1658 17234 1834
rect 22739 1902 22797 1914
rect 22739 1726 22751 1902
rect 22785 1726 22797 1902
rect 22739 1714 22797 1726
rect 22857 1902 22915 1914
rect 22857 1726 22869 1902
rect 22903 1726 22915 1902
rect 22857 1714 22915 1726
rect 22975 1902 23033 1914
rect 22975 1726 22987 1902
rect 23021 1726 23033 1902
rect 22975 1714 23033 1726
rect 23093 1902 23151 1914
rect 23093 1726 23105 1902
rect 23139 1726 23151 1902
rect 23093 1714 23151 1726
rect 23211 1902 23269 1914
rect 23211 1726 23223 1902
rect 23257 1726 23269 1902
rect 23211 1714 23269 1726
rect 23329 1902 23387 1914
rect 23329 1726 23341 1902
rect 23375 1726 23387 1902
rect 23329 1714 23387 1726
rect 23447 1902 23505 1914
rect 23447 1726 23459 1902
rect 23493 1726 23505 1902
rect 23447 1714 23505 1726
rect 23565 1902 23623 1914
rect 23565 1726 23577 1902
rect 23611 1726 23623 1902
rect 23565 1714 23623 1726
rect 23683 1902 23741 1914
rect 23683 1726 23695 1902
rect 23729 1726 23741 1902
rect 23683 1714 23741 1726
rect 23801 1902 23859 1914
rect 23801 1726 23813 1902
rect 23847 1726 23859 1902
rect 23801 1714 23859 1726
rect 17176 1646 17234 1658
rect 11408 1485 11466 1497
rect 4859 1397 4917 1409
rect -1 1146 57 1158
rect -1 970 11 1146
rect 45 970 57 1146
rect -1 958 57 970
rect 117 1146 175 1158
rect 117 970 129 1146
rect 163 970 175 1146
rect 117 958 175 970
rect 235 1146 293 1158
rect 235 970 247 1146
rect 281 970 293 1146
rect 235 958 293 970
rect 353 1146 411 1158
rect 353 970 365 1146
rect 399 970 411 1146
rect 353 958 411 970
rect 471 1146 529 1158
rect 471 970 483 1146
rect 517 970 529 1146
rect 471 958 529 970
rect 589 1146 647 1158
rect 589 970 601 1146
rect 635 970 647 1146
rect 589 958 647 970
rect 707 1146 765 1158
rect 707 970 719 1146
rect 753 970 765 1146
rect 707 958 765 970
rect 825 1146 883 1158
rect 825 970 837 1146
rect 871 970 883 1146
rect 825 958 883 970
rect 943 1146 1001 1158
rect 943 970 955 1146
rect 989 970 1001 1146
rect 943 958 1001 970
rect 1061 1146 1119 1158
rect 1061 970 1073 1146
rect 1107 970 1119 1146
rect 4375 1197 4433 1209
rect 1061 958 1119 970
rect 4375 1021 4387 1197
rect 4421 1021 4433 1197
rect 4375 1009 4433 1021
rect 4493 1197 4551 1209
rect 4493 1021 4505 1197
rect 4539 1021 4551 1197
rect 4493 1009 4551 1021
rect 4611 1197 4669 1209
rect 4611 1021 4623 1197
rect 4657 1021 4669 1197
rect 4611 1009 4669 1021
rect 4729 1197 4787 1209
rect 4729 1021 4741 1197
rect 4775 1021 4787 1197
rect 4729 1009 4787 1021
rect 4859 1021 4871 1397
rect 4905 1021 4917 1397
rect 4859 1009 4917 1021
rect 4977 1397 5035 1409
rect 4977 1021 4989 1397
rect 5023 1021 5035 1397
rect 4977 1009 5035 1021
rect 5095 1397 5153 1409
rect 5095 1021 5107 1397
rect 5141 1021 5153 1397
rect 5095 1009 5153 1021
rect 5213 1397 5271 1409
rect 5213 1021 5225 1397
rect 5259 1021 5271 1397
rect 5213 1009 5271 1021
rect 5331 1397 5389 1409
rect 5331 1021 5343 1397
rect 5377 1021 5389 1397
rect 5331 1009 5389 1021
rect 5449 1397 5507 1409
rect 5449 1021 5461 1397
rect 5495 1021 5507 1397
rect 5449 1009 5507 1021
rect 5567 1397 5625 1409
rect 5567 1021 5579 1397
rect 5613 1021 5625 1397
rect 6757 1397 6815 1409
rect 5567 1009 5625 1021
rect 5696 1197 5754 1209
rect 5696 1021 5708 1197
rect 5742 1021 5754 1197
rect 5696 1009 5754 1021
rect 5814 1197 5872 1209
rect 5814 1021 5826 1197
rect 5860 1021 5872 1197
rect 5814 1009 5872 1021
rect 5932 1197 5990 1209
rect 5932 1021 5944 1197
rect 5978 1021 5990 1197
rect 5932 1009 5990 1021
rect 6050 1197 6108 1209
rect 6050 1021 6062 1197
rect 6096 1021 6108 1197
rect 6050 1009 6108 1021
rect 6273 1197 6331 1209
rect 6273 1021 6285 1197
rect 6319 1021 6331 1197
rect 6273 1009 6331 1021
rect 6391 1197 6449 1209
rect 6391 1021 6403 1197
rect 6437 1021 6449 1197
rect 6391 1009 6449 1021
rect 6509 1197 6567 1209
rect 6509 1021 6521 1197
rect 6555 1021 6567 1197
rect 6509 1009 6567 1021
rect 6627 1197 6685 1209
rect 6627 1021 6639 1197
rect 6673 1021 6685 1197
rect 6627 1009 6685 1021
rect 6757 1021 6769 1397
rect 6803 1021 6815 1397
rect 6757 1009 6815 1021
rect 6875 1397 6933 1409
rect 6875 1021 6887 1397
rect 6921 1021 6933 1397
rect 6875 1009 6933 1021
rect 6993 1397 7051 1409
rect 6993 1021 7005 1397
rect 7039 1021 7051 1397
rect 6993 1009 7051 1021
rect 7111 1397 7169 1409
rect 7111 1021 7123 1397
rect 7157 1021 7169 1397
rect 7111 1009 7169 1021
rect 7229 1397 7287 1409
rect 7229 1021 7241 1397
rect 7275 1021 7287 1397
rect 7229 1009 7287 1021
rect 7347 1397 7405 1409
rect 7347 1021 7359 1397
rect 7393 1021 7405 1397
rect 7347 1009 7405 1021
rect 7465 1397 7523 1409
rect 7465 1021 7477 1397
rect 7511 1021 7523 1397
rect 7465 1009 7523 1021
rect 7594 1197 7652 1209
rect 7594 1021 7606 1197
rect 7640 1021 7652 1197
rect 7594 1009 7652 1021
rect 7712 1197 7770 1209
rect 7712 1021 7724 1197
rect 7758 1021 7770 1197
rect 7712 1009 7770 1021
rect 7830 1197 7888 1209
rect 7830 1021 7842 1197
rect 7876 1021 7888 1197
rect 7830 1009 7888 1021
rect 7948 1197 8006 1209
rect 7948 1021 7960 1197
rect 7994 1021 8006 1197
rect 10924 1285 10982 1297
rect 7948 1009 8006 1021
rect 2906 210 2964 222
rect 2906 34 2918 210
rect 2952 34 2964 210
rect 2906 22 2964 34
rect 3024 210 3082 222
rect 3024 34 3036 210
rect 3070 34 3082 210
rect 3024 22 3082 34
rect 3142 210 3200 222
rect 3142 34 3154 210
rect 3188 34 3200 210
rect 3142 22 3200 34
rect 3260 210 3318 222
rect 3260 34 3272 210
rect 3306 34 3318 210
rect 3260 22 3318 34
rect 3378 210 3436 222
rect 3378 34 3390 210
rect 3424 34 3436 210
rect 3378 22 3436 34
rect 3496 210 3554 222
rect 3496 34 3508 210
rect 3542 34 3554 210
rect 3496 22 3554 34
rect 3614 210 3672 222
rect 3614 34 3626 210
rect 3660 34 3672 210
rect 3614 22 3672 34
rect 3732 210 3790 222
rect 3732 34 3744 210
rect 3778 34 3790 210
rect 3732 22 3790 34
rect 3850 210 3908 222
rect 3850 34 3862 210
rect 3896 34 3908 210
rect 3850 22 3908 34
rect 3968 210 4026 222
rect 3968 34 3980 210
rect 4014 34 4026 210
rect 3968 22 4026 34
rect 4802 704 4860 716
rect 4802 328 4814 704
rect 4848 328 4860 704
rect 4802 316 4860 328
rect 4920 704 4978 716
rect 4920 328 4932 704
rect 4966 328 4978 704
rect 4920 316 4978 328
rect 5038 704 5096 716
rect 5038 328 5050 704
rect 5084 328 5096 704
rect 5038 316 5096 328
rect 5156 704 5214 716
rect 5156 328 5168 704
rect 5202 328 5214 704
rect 5156 316 5214 328
rect 5274 704 5332 716
rect 5274 328 5286 704
rect 5320 328 5332 704
rect 5274 316 5332 328
rect 5392 704 5450 716
rect 5392 328 5404 704
rect 5438 328 5450 704
rect 5392 316 5450 328
rect 5510 704 5568 716
rect 5510 328 5522 704
rect 5556 328 5568 704
rect 5510 316 5568 328
rect 10924 1109 10936 1285
rect 10970 1109 10982 1285
rect 10924 1097 10982 1109
rect 11042 1285 11100 1297
rect 11042 1109 11054 1285
rect 11088 1109 11100 1285
rect 11042 1097 11100 1109
rect 11160 1285 11218 1297
rect 11160 1109 11172 1285
rect 11206 1109 11218 1285
rect 11160 1097 11218 1109
rect 11278 1285 11336 1297
rect 11278 1109 11290 1285
rect 11324 1109 11336 1285
rect 11278 1097 11336 1109
rect 11408 1109 11420 1485
rect 11454 1109 11466 1485
rect 11408 1097 11466 1109
rect 11526 1485 11584 1497
rect 11526 1109 11538 1485
rect 11572 1109 11584 1485
rect 11526 1097 11584 1109
rect 11644 1485 11702 1497
rect 11644 1109 11656 1485
rect 11690 1109 11702 1485
rect 11644 1097 11702 1109
rect 11762 1485 11820 1497
rect 11762 1109 11774 1485
rect 11808 1109 11820 1485
rect 11762 1097 11820 1109
rect 11880 1485 11938 1497
rect 11880 1109 11892 1485
rect 11926 1109 11938 1485
rect 11880 1097 11938 1109
rect 11998 1485 12056 1497
rect 11998 1109 12010 1485
rect 12044 1109 12056 1485
rect 11998 1097 12056 1109
rect 12116 1485 12174 1497
rect 12116 1109 12128 1485
rect 12162 1109 12174 1485
rect 13306 1485 13364 1497
rect 12116 1097 12174 1109
rect 12245 1285 12303 1297
rect 12245 1109 12257 1285
rect 12291 1109 12303 1285
rect 12245 1097 12303 1109
rect 12363 1285 12421 1297
rect 12363 1109 12375 1285
rect 12409 1109 12421 1285
rect 12363 1097 12421 1109
rect 12481 1285 12539 1297
rect 12481 1109 12493 1285
rect 12527 1109 12539 1285
rect 12481 1097 12539 1109
rect 12599 1285 12657 1297
rect 12599 1109 12611 1285
rect 12645 1109 12657 1285
rect 12599 1097 12657 1109
rect 12822 1285 12880 1297
rect 12822 1109 12834 1285
rect 12868 1109 12880 1285
rect 12822 1097 12880 1109
rect 12940 1285 12998 1297
rect 12940 1109 12952 1285
rect 12986 1109 12998 1285
rect 12940 1097 12998 1109
rect 13058 1285 13116 1297
rect 13058 1109 13070 1285
rect 13104 1109 13116 1285
rect 13058 1097 13116 1109
rect 13176 1285 13234 1297
rect 13176 1109 13188 1285
rect 13222 1109 13234 1285
rect 13176 1097 13234 1109
rect 13306 1109 13318 1485
rect 13352 1109 13364 1485
rect 13306 1097 13364 1109
rect 13424 1485 13482 1497
rect 13424 1109 13436 1485
rect 13470 1109 13482 1485
rect 13424 1097 13482 1109
rect 13542 1485 13600 1497
rect 13542 1109 13554 1485
rect 13588 1109 13600 1485
rect 13542 1097 13600 1109
rect 13660 1485 13718 1497
rect 13660 1109 13672 1485
rect 13706 1109 13718 1485
rect 13660 1097 13718 1109
rect 13778 1485 13836 1497
rect 13778 1109 13790 1485
rect 13824 1109 13836 1485
rect 13778 1097 13836 1109
rect 13896 1485 13954 1497
rect 13896 1109 13908 1485
rect 13942 1109 13954 1485
rect 13896 1097 13954 1109
rect 14014 1485 14072 1497
rect 14014 1109 14026 1485
rect 14060 1109 14072 1485
rect 24687 1485 24745 1497
rect 18062 1417 18120 1429
rect 14014 1097 14072 1109
rect 14143 1285 14201 1297
rect 14143 1109 14155 1285
rect 14189 1109 14201 1285
rect 14143 1097 14201 1109
rect 14261 1285 14319 1297
rect 14261 1109 14273 1285
rect 14307 1109 14319 1285
rect 14261 1097 14319 1109
rect 14379 1285 14437 1297
rect 14379 1109 14391 1285
rect 14425 1109 14437 1285
rect 14379 1097 14437 1109
rect 14497 1285 14555 1297
rect 14497 1109 14509 1285
rect 14543 1109 14555 1285
rect 14497 1097 14555 1109
rect 6700 704 6758 716
rect 6700 328 6712 704
rect 6746 328 6758 704
rect 6700 316 6758 328
rect 6818 704 6876 716
rect 6818 328 6830 704
rect 6864 328 6876 704
rect 6818 316 6876 328
rect 6936 704 6994 716
rect 6936 328 6948 704
rect 6982 328 6994 704
rect 6936 316 6994 328
rect 7054 704 7112 716
rect 7054 328 7066 704
rect 7100 328 7112 704
rect 7054 316 7112 328
rect 7172 704 7230 716
rect 7172 328 7184 704
rect 7218 328 7230 704
rect 7172 316 7230 328
rect 7290 704 7348 716
rect 7290 328 7302 704
rect 7336 328 7348 704
rect 7290 316 7348 328
rect 7408 704 7466 716
rect 7408 328 7420 704
rect 7454 328 7466 704
rect 7408 316 7466 328
rect 9455 298 9513 310
rect 9455 122 9467 298
rect 9501 122 9513 298
rect 9455 110 9513 122
rect 9573 298 9631 310
rect 9573 122 9585 298
rect 9619 122 9631 298
rect 9573 110 9631 122
rect 9691 298 9749 310
rect 9691 122 9703 298
rect 9737 122 9749 298
rect 9691 110 9749 122
rect 9809 298 9867 310
rect 9809 122 9821 298
rect 9855 122 9867 298
rect 9809 110 9867 122
rect 9927 298 9985 310
rect 9927 122 9939 298
rect 9973 122 9985 298
rect 9927 110 9985 122
rect 10045 298 10103 310
rect 10045 122 10057 298
rect 10091 122 10103 298
rect 10045 110 10103 122
rect 10163 298 10221 310
rect 10163 122 10175 298
rect 10209 122 10221 298
rect 10163 110 10221 122
rect 10281 298 10339 310
rect 10281 122 10293 298
rect 10327 122 10339 298
rect 10281 110 10339 122
rect 10399 298 10457 310
rect 10399 122 10411 298
rect 10445 122 10457 298
rect 10399 110 10457 122
rect 10517 298 10575 310
rect 10517 122 10529 298
rect 10563 122 10575 298
rect 10517 110 10575 122
rect 11351 792 11409 804
rect 11351 416 11363 792
rect 11397 416 11409 792
rect 11351 404 11409 416
rect 11469 792 11527 804
rect 11469 416 11481 792
rect 11515 416 11527 792
rect 11469 404 11527 416
rect 11587 792 11645 804
rect 11587 416 11599 792
rect 11633 416 11645 792
rect 11587 404 11645 416
rect 11705 792 11763 804
rect 11705 416 11717 792
rect 11751 416 11763 792
rect 11705 404 11763 416
rect 11823 792 11881 804
rect 11823 416 11835 792
rect 11869 416 11881 792
rect 11823 404 11881 416
rect 11941 792 11999 804
rect 11941 416 11953 792
rect 11987 416 11999 792
rect 11941 404 11999 416
rect 12059 792 12117 804
rect 12059 416 12071 792
rect 12105 416 12117 792
rect 12059 404 12117 416
rect 17578 1217 17636 1229
rect 17578 1041 17590 1217
rect 17624 1041 17636 1217
rect 17578 1029 17636 1041
rect 17696 1217 17754 1229
rect 17696 1041 17708 1217
rect 17742 1041 17754 1217
rect 17696 1029 17754 1041
rect 17814 1217 17872 1229
rect 17814 1041 17826 1217
rect 17860 1041 17872 1217
rect 17814 1029 17872 1041
rect 17932 1217 17990 1229
rect 17932 1041 17944 1217
rect 17978 1041 17990 1217
rect 17932 1029 17990 1041
rect 18062 1041 18074 1417
rect 18108 1041 18120 1417
rect 18062 1029 18120 1041
rect 18180 1417 18238 1429
rect 18180 1041 18192 1417
rect 18226 1041 18238 1417
rect 18180 1029 18238 1041
rect 18298 1417 18356 1429
rect 18298 1041 18310 1417
rect 18344 1041 18356 1417
rect 18298 1029 18356 1041
rect 18416 1417 18474 1429
rect 18416 1041 18428 1417
rect 18462 1041 18474 1417
rect 18416 1029 18474 1041
rect 18534 1417 18592 1429
rect 18534 1041 18546 1417
rect 18580 1041 18592 1417
rect 18534 1029 18592 1041
rect 18652 1417 18710 1429
rect 18652 1041 18664 1417
rect 18698 1041 18710 1417
rect 18652 1029 18710 1041
rect 18770 1417 18828 1429
rect 18770 1041 18782 1417
rect 18816 1041 18828 1417
rect 19960 1417 20018 1429
rect 18770 1029 18828 1041
rect 18899 1217 18957 1229
rect 18899 1041 18911 1217
rect 18945 1041 18957 1217
rect 18899 1029 18957 1041
rect 19017 1217 19075 1229
rect 19017 1041 19029 1217
rect 19063 1041 19075 1217
rect 19017 1029 19075 1041
rect 19135 1217 19193 1229
rect 19135 1041 19147 1217
rect 19181 1041 19193 1217
rect 19135 1029 19193 1041
rect 19253 1217 19311 1229
rect 19253 1041 19265 1217
rect 19299 1041 19311 1217
rect 19253 1029 19311 1041
rect 19476 1217 19534 1229
rect 19476 1041 19488 1217
rect 19522 1041 19534 1217
rect 19476 1029 19534 1041
rect 19594 1217 19652 1229
rect 19594 1041 19606 1217
rect 19640 1041 19652 1217
rect 19594 1029 19652 1041
rect 19712 1217 19770 1229
rect 19712 1041 19724 1217
rect 19758 1041 19770 1217
rect 19712 1029 19770 1041
rect 19830 1217 19888 1229
rect 19830 1041 19842 1217
rect 19876 1041 19888 1217
rect 19830 1029 19888 1041
rect 19960 1041 19972 1417
rect 20006 1041 20018 1417
rect 19960 1029 20018 1041
rect 20078 1417 20136 1429
rect 20078 1041 20090 1417
rect 20124 1041 20136 1417
rect 20078 1029 20136 1041
rect 20196 1417 20254 1429
rect 20196 1041 20208 1417
rect 20242 1041 20254 1417
rect 20196 1029 20254 1041
rect 20314 1417 20372 1429
rect 20314 1041 20326 1417
rect 20360 1041 20372 1417
rect 20314 1029 20372 1041
rect 20432 1417 20490 1429
rect 20432 1041 20444 1417
rect 20478 1041 20490 1417
rect 20432 1029 20490 1041
rect 20550 1417 20608 1429
rect 20550 1041 20562 1417
rect 20596 1041 20608 1417
rect 20550 1029 20608 1041
rect 20668 1417 20726 1429
rect 20668 1041 20680 1417
rect 20714 1041 20726 1417
rect 20668 1029 20726 1041
rect 20797 1217 20855 1229
rect 20797 1041 20809 1217
rect 20843 1041 20855 1217
rect 20797 1029 20855 1041
rect 20915 1217 20973 1229
rect 20915 1041 20927 1217
rect 20961 1041 20973 1217
rect 20915 1029 20973 1041
rect 21033 1217 21091 1229
rect 21033 1041 21045 1217
rect 21079 1041 21091 1217
rect 21033 1029 21091 1041
rect 21151 1217 21209 1229
rect 21151 1041 21163 1217
rect 21197 1041 21209 1217
rect 24203 1285 24261 1297
rect 21151 1029 21209 1041
rect 13249 792 13307 804
rect 13249 416 13261 792
rect 13295 416 13307 792
rect 13249 404 13307 416
rect 13367 792 13425 804
rect 13367 416 13379 792
rect 13413 416 13425 792
rect 13367 404 13425 416
rect 13485 792 13543 804
rect 13485 416 13497 792
rect 13531 416 13543 792
rect 13485 404 13543 416
rect 13603 792 13661 804
rect 13603 416 13615 792
rect 13649 416 13661 792
rect 13603 404 13661 416
rect 13721 792 13779 804
rect 13721 416 13733 792
rect 13767 416 13779 792
rect 13721 404 13779 416
rect 13839 792 13897 804
rect 13839 416 13851 792
rect 13885 416 13897 792
rect 13839 404 13897 416
rect 13957 792 14015 804
rect 13957 416 13969 792
rect 14003 416 14015 792
rect 13957 404 14015 416
rect 16109 230 16167 242
rect 16109 54 16121 230
rect 16155 54 16167 230
rect 16109 42 16167 54
rect 16227 230 16285 242
rect 16227 54 16239 230
rect 16273 54 16285 230
rect 16227 42 16285 54
rect 16345 230 16403 242
rect 16345 54 16357 230
rect 16391 54 16403 230
rect 16345 42 16403 54
rect 16463 230 16521 242
rect 16463 54 16475 230
rect 16509 54 16521 230
rect 16463 42 16521 54
rect 16581 230 16639 242
rect 16581 54 16593 230
rect 16627 54 16639 230
rect 16581 42 16639 54
rect 16699 230 16757 242
rect 16699 54 16711 230
rect 16745 54 16757 230
rect 16699 42 16757 54
rect 16817 230 16875 242
rect 16817 54 16829 230
rect 16863 54 16875 230
rect 16817 42 16875 54
rect 16935 230 16993 242
rect 16935 54 16947 230
rect 16981 54 16993 230
rect 16935 42 16993 54
rect 17053 230 17111 242
rect 17053 54 17065 230
rect 17099 54 17111 230
rect 17053 42 17111 54
rect 17171 230 17229 242
rect 17171 54 17183 230
rect 17217 54 17229 230
rect 17171 42 17229 54
rect 18005 724 18063 736
rect 18005 348 18017 724
rect 18051 348 18063 724
rect 18005 336 18063 348
rect 18123 724 18181 736
rect 18123 348 18135 724
rect 18169 348 18181 724
rect 18123 336 18181 348
rect 18241 724 18299 736
rect 18241 348 18253 724
rect 18287 348 18299 724
rect 18241 336 18299 348
rect 18359 724 18417 736
rect 18359 348 18371 724
rect 18405 348 18417 724
rect 18359 336 18417 348
rect 18477 724 18535 736
rect 18477 348 18489 724
rect 18523 348 18535 724
rect 18477 336 18535 348
rect 18595 724 18653 736
rect 18595 348 18607 724
rect 18641 348 18653 724
rect 18595 336 18653 348
rect 18713 724 18771 736
rect 18713 348 18725 724
rect 18759 348 18771 724
rect 18713 336 18771 348
rect 24203 1109 24215 1285
rect 24249 1109 24261 1285
rect 24203 1097 24261 1109
rect 24321 1285 24379 1297
rect 24321 1109 24333 1285
rect 24367 1109 24379 1285
rect 24321 1097 24379 1109
rect 24439 1285 24497 1297
rect 24439 1109 24451 1285
rect 24485 1109 24497 1285
rect 24439 1097 24497 1109
rect 24557 1285 24615 1297
rect 24557 1109 24569 1285
rect 24603 1109 24615 1285
rect 24557 1097 24615 1109
rect 24687 1109 24699 1485
rect 24733 1109 24745 1485
rect 24687 1097 24745 1109
rect 24805 1485 24863 1497
rect 24805 1109 24817 1485
rect 24851 1109 24863 1485
rect 24805 1097 24863 1109
rect 24923 1485 24981 1497
rect 24923 1109 24935 1485
rect 24969 1109 24981 1485
rect 24923 1097 24981 1109
rect 25041 1485 25099 1497
rect 25041 1109 25053 1485
rect 25087 1109 25099 1485
rect 25041 1097 25099 1109
rect 25159 1485 25217 1497
rect 25159 1109 25171 1485
rect 25205 1109 25217 1485
rect 25159 1097 25217 1109
rect 25277 1485 25335 1497
rect 25277 1109 25289 1485
rect 25323 1109 25335 1485
rect 25277 1097 25335 1109
rect 25395 1485 25453 1497
rect 25395 1109 25407 1485
rect 25441 1109 25453 1485
rect 26585 1485 26643 1497
rect 25395 1097 25453 1109
rect 25524 1285 25582 1297
rect 25524 1109 25536 1285
rect 25570 1109 25582 1285
rect 25524 1097 25582 1109
rect 25642 1285 25700 1297
rect 25642 1109 25654 1285
rect 25688 1109 25700 1285
rect 25642 1097 25700 1109
rect 25760 1285 25818 1297
rect 25760 1109 25772 1285
rect 25806 1109 25818 1285
rect 25760 1097 25818 1109
rect 25878 1285 25936 1297
rect 25878 1109 25890 1285
rect 25924 1109 25936 1285
rect 25878 1097 25936 1109
rect 26101 1285 26159 1297
rect 26101 1109 26113 1285
rect 26147 1109 26159 1285
rect 26101 1097 26159 1109
rect 26219 1285 26277 1297
rect 26219 1109 26231 1285
rect 26265 1109 26277 1285
rect 26219 1097 26277 1109
rect 26337 1285 26395 1297
rect 26337 1109 26349 1285
rect 26383 1109 26395 1285
rect 26337 1097 26395 1109
rect 26455 1285 26513 1297
rect 26455 1109 26467 1285
rect 26501 1109 26513 1285
rect 26455 1097 26513 1109
rect 26585 1109 26597 1485
rect 26631 1109 26643 1485
rect 26585 1097 26643 1109
rect 26703 1485 26761 1497
rect 26703 1109 26715 1485
rect 26749 1109 26761 1485
rect 26703 1097 26761 1109
rect 26821 1485 26879 1497
rect 26821 1109 26833 1485
rect 26867 1109 26879 1485
rect 26821 1097 26879 1109
rect 26939 1485 26997 1497
rect 26939 1109 26951 1485
rect 26985 1109 26997 1485
rect 26939 1097 26997 1109
rect 27057 1485 27115 1497
rect 27057 1109 27069 1485
rect 27103 1109 27115 1485
rect 27057 1097 27115 1109
rect 27175 1485 27233 1497
rect 27175 1109 27187 1485
rect 27221 1109 27233 1485
rect 27175 1097 27233 1109
rect 27293 1485 27351 1497
rect 27293 1109 27305 1485
rect 27339 1109 27351 1485
rect 27293 1097 27351 1109
rect 27422 1285 27480 1297
rect 27422 1109 27434 1285
rect 27468 1109 27480 1285
rect 27422 1097 27480 1109
rect 27540 1285 27598 1297
rect 27540 1109 27552 1285
rect 27586 1109 27598 1285
rect 27540 1097 27598 1109
rect 27658 1285 27716 1297
rect 27658 1109 27670 1285
rect 27704 1109 27716 1285
rect 27658 1097 27716 1109
rect 27776 1285 27834 1297
rect 27776 1109 27788 1285
rect 27822 1109 27834 1285
rect 27776 1097 27834 1109
rect 30821 1188 30879 1200
rect 19903 724 19961 736
rect 19903 348 19915 724
rect 19949 348 19961 724
rect 19903 336 19961 348
rect 20021 724 20079 736
rect 20021 348 20033 724
rect 20067 348 20079 724
rect 20021 336 20079 348
rect 20139 724 20197 736
rect 20139 348 20151 724
rect 20185 348 20197 724
rect 20139 336 20197 348
rect 20257 724 20315 736
rect 20257 348 20269 724
rect 20303 348 20315 724
rect 20257 336 20315 348
rect 20375 724 20433 736
rect 20375 348 20387 724
rect 20421 348 20433 724
rect 20375 336 20433 348
rect 20493 724 20551 736
rect 20493 348 20505 724
rect 20539 348 20551 724
rect 20493 336 20551 348
rect 20611 724 20669 736
rect 20611 348 20623 724
rect 20657 348 20669 724
rect 20611 336 20669 348
rect 22734 298 22792 310
rect 22734 122 22746 298
rect 22780 122 22792 298
rect 22734 110 22792 122
rect 22852 298 22910 310
rect 22852 122 22864 298
rect 22898 122 22910 298
rect 22852 110 22910 122
rect 22970 298 23028 310
rect 22970 122 22982 298
rect 23016 122 23028 298
rect 22970 110 23028 122
rect 23088 298 23146 310
rect 23088 122 23100 298
rect 23134 122 23146 298
rect 23088 110 23146 122
rect 23206 298 23264 310
rect 23206 122 23218 298
rect 23252 122 23264 298
rect 23206 110 23264 122
rect 23324 298 23382 310
rect 23324 122 23336 298
rect 23370 122 23382 298
rect 23324 110 23382 122
rect 23442 298 23500 310
rect 23442 122 23454 298
rect 23488 122 23500 298
rect 23442 110 23500 122
rect 23560 298 23618 310
rect 23560 122 23572 298
rect 23606 122 23618 298
rect 23560 110 23618 122
rect 23678 298 23736 310
rect 23678 122 23690 298
rect 23724 122 23736 298
rect 23678 110 23736 122
rect 23796 298 23854 310
rect 23796 122 23808 298
rect 23842 122 23854 298
rect 23796 110 23854 122
rect 24630 792 24688 804
rect 24630 416 24642 792
rect 24676 416 24688 792
rect 24630 404 24688 416
rect 24748 792 24806 804
rect 24748 416 24760 792
rect 24794 416 24806 792
rect 24748 404 24806 416
rect 24866 792 24924 804
rect 24866 416 24878 792
rect 24912 416 24924 792
rect 24866 404 24924 416
rect 24984 792 25042 804
rect 24984 416 24996 792
rect 25030 416 25042 792
rect 24984 404 25042 416
rect 25102 792 25160 804
rect 25102 416 25114 792
rect 25148 416 25160 792
rect 25102 404 25160 416
rect 25220 792 25278 804
rect 25220 416 25232 792
rect 25266 416 25278 792
rect 25220 404 25278 416
rect 25338 792 25396 804
rect 25338 416 25350 792
rect 25384 416 25396 792
rect 25338 404 25396 416
rect 30337 988 30395 1000
rect 26528 792 26586 804
rect 26528 416 26540 792
rect 26574 416 26586 792
rect 26528 404 26586 416
rect 26646 792 26704 804
rect 26646 416 26658 792
rect 26692 416 26704 792
rect 26646 404 26704 416
rect 26764 792 26822 804
rect 26764 416 26776 792
rect 26810 416 26822 792
rect 26764 404 26822 416
rect 26882 792 26940 804
rect 26882 416 26894 792
rect 26928 416 26940 792
rect 26882 404 26940 416
rect 27000 792 27058 804
rect 27000 416 27012 792
rect 27046 416 27058 792
rect 27000 404 27058 416
rect 27118 792 27176 804
rect 27118 416 27130 792
rect 27164 416 27176 792
rect 27118 404 27176 416
rect 27236 792 27294 804
rect 27236 416 27248 792
rect 27282 416 27294 792
rect 27236 404 27294 416
rect 30337 812 30349 988
rect 30383 812 30395 988
rect 30337 800 30395 812
rect 30455 988 30513 1000
rect 30455 812 30467 988
rect 30501 812 30513 988
rect 30455 800 30513 812
rect 30573 988 30631 1000
rect 30573 812 30585 988
rect 30619 812 30631 988
rect 30573 800 30631 812
rect 30691 988 30749 1000
rect 30691 812 30703 988
rect 30737 812 30749 988
rect 30691 800 30749 812
rect 30821 812 30833 1188
rect 30867 812 30879 1188
rect 30821 800 30879 812
rect 30939 1188 30997 1200
rect 30939 812 30951 1188
rect 30985 812 30997 1188
rect 30939 800 30997 812
rect 31057 1188 31115 1200
rect 31057 812 31069 1188
rect 31103 812 31115 1188
rect 31057 800 31115 812
rect 31175 1188 31233 1200
rect 31175 812 31187 1188
rect 31221 812 31233 1188
rect 31175 800 31233 812
rect 31293 1188 31351 1200
rect 31293 812 31305 1188
rect 31339 812 31351 1188
rect 31293 800 31351 812
rect 31411 1188 31469 1200
rect 31411 812 31423 1188
rect 31457 812 31469 1188
rect 31411 800 31469 812
rect 31529 1188 31587 1200
rect 31529 812 31541 1188
rect 31575 812 31587 1188
rect 31529 800 31587 812
rect 31658 988 31716 1000
rect 31658 812 31670 988
rect 31704 812 31716 988
rect 31658 800 31716 812
rect 31776 988 31834 1000
rect 31776 812 31788 988
rect 31822 812 31834 988
rect 31776 800 31834 812
rect 31894 988 31952 1000
rect 31894 812 31906 988
rect 31940 812 31952 988
rect 31894 800 31952 812
rect 32012 988 32070 1000
rect 32012 812 32024 988
rect 32058 812 32070 988
rect 32012 800 32070 812
rect 32130 985 32188 997
rect 32130 809 32142 985
rect 32176 809 32188 985
rect 32130 797 32188 809
rect 32248 985 32306 997
rect 32248 809 32260 985
rect 32294 809 32306 985
rect 32248 797 32306 809
rect 32366 985 32424 997
rect 32366 809 32378 985
rect 32412 809 32424 985
rect 32366 797 32424 809
rect 32484 985 32542 997
rect 32484 809 32496 985
rect 32530 809 32542 985
rect 32484 797 32542 809
rect 32602 985 32660 997
rect 32602 809 32614 985
rect 32648 809 32660 985
rect 32602 797 32660 809
rect 32720 985 32778 997
rect 32720 809 32732 985
rect 32766 809 32778 985
rect 32720 797 32778 809
rect 32838 985 32896 997
rect 32838 809 32850 985
rect 32884 809 32896 985
rect 32838 797 32896 809
rect 32956 985 33014 997
rect 32956 809 32968 985
rect 33002 809 33014 985
rect 32956 797 33014 809
rect 33074 985 33132 997
rect 33074 809 33086 985
rect 33120 809 33132 985
rect 33074 797 33132 809
rect 33192 985 33250 997
rect 33192 809 33204 985
rect 33238 809 33250 985
rect 33192 797 33250 809
rect 30764 495 30822 507
rect 28522 -120 28580 -108
rect 28522 -296 28534 -120
rect 28568 -296 28580 -120
rect 28522 -308 28580 -296
rect 28640 -120 28698 -108
rect 28640 -296 28652 -120
rect 28686 -296 28698 -120
rect 28640 -308 28698 -296
rect 28758 -120 28816 -108
rect 28758 -296 28770 -120
rect 28804 -296 28816 -120
rect 28758 -308 28816 -296
rect 28876 -120 28934 -108
rect 28876 -296 28888 -120
rect 28922 -296 28934 -120
rect 28876 -308 28934 -296
rect 28994 -120 29052 -108
rect 28994 -296 29006 -120
rect 29040 -296 29052 -120
rect 28994 -308 29052 -296
rect 29112 -120 29170 -108
rect 29112 -296 29124 -120
rect 29158 -296 29170 -120
rect 29112 -308 29170 -296
rect 29230 -120 29288 -108
rect 29230 -296 29242 -120
rect 29276 -296 29288 -120
rect 29230 -308 29288 -296
rect 29348 -120 29406 -108
rect 29348 -296 29360 -120
rect 29394 -296 29406 -120
rect 29348 -308 29406 -296
rect 29466 -120 29524 -108
rect 29466 -296 29478 -120
rect 29512 -296 29524 -120
rect 29466 -308 29524 -296
rect 29584 -120 29642 -108
rect 29584 -296 29596 -120
rect 29630 -296 29642 -120
rect 30764 119 30776 495
rect 30810 119 30822 495
rect 30764 107 30822 119
rect 30882 495 30940 507
rect 30882 119 30894 495
rect 30928 119 30940 495
rect 30882 107 30940 119
rect 31000 495 31058 507
rect 31000 119 31012 495
rect 31046 119 31058 495
rect 31000 107 31058 119
rect 31118 495 31176 507
rect 31118 119 31130 495
rect 31164 119 31176 495
rect 31118 107 31176 119
rect 31236 495 31294 507
rect 31236 119 31248 495
rect 31282 119 31294 495
rect 31236 107 31294 119
rect 31354 495 31412 507
rect 31354 119 31366 495
rect 31400 119 31412 495
rect 31354 107 31412 119
rect 31472 495 31530 507
rect 31472 119 31484 495
rect 31518 119 31530 495
rect 31472 107 31530 119
rect 29584 -308 29642 -296
rect -20 -2132 38 -2120
rect -20 -2308 -8 -2132
rect 26 -2308 38 -2132
rect -20 -2320 38 -2308
rect 98 -2132 156 -2120
rect 98 -2308 110 -2132
rect 144 -2308 156 -2132
rect 98 -2320 156 -2308
rect 216 -2132 274 -2120
rect 216 -2308 228 -2132
rect 262 -2308 274 -2132
rect 216 -2320 274 -2308
rect 334 -2132 392 -2120
rect 334 -2308 346 -2132
rect 380 -2308 392 -2132
rect 334 -2320 392 -2308
rect 452 -2132 510 -2120
rect 452 -2308 464 -2132
rect 498 -2308 510 -2132
rect 452 -2320 510 -2308
rect 570 -2132 628 -2120
rect 570 -2308 582 -2132
rect 616 -2308 628 -2132
rect 570 -2320 628 -2308
rect 688 -2132 746 -2120
rect 688 -2308 700 -2132
rect 734 -2308 746 -2132
rect 688 -2320 746 -2308
rect 806 -2132 864 -2120
rect 806 -2308 818 -2132
rect 852 -2308 864 -2132
rect 806 -2320 864 -2308
rect 924 -2132 982 -2120
rect 924 -2308 936 -2132
rect 970 -2308 982 -2132
rect 924 -2320 982 -2308
rect 1042 -2132 1100 -2120
rect 1042 -2308 1054 -2132
rect 1088 -2308 1100 -2132
rect 5214 -2244 5272 -2232
rect 1042 -2320 1100 -2308
rect 2889 -2316 2947 -2304
rect 2889 -2492 2901 -2316
rect 2935 -2492 2947 -2316
rect 2889 -2504 2947 -2492
rect 3007 -2316 3065 -2304
rect 3007 -2492 3019 -2316
rect 3053 -2492 3065 -2316
rect 3007 -2504 3065 -2492
rect 3125 -2316 3183 -2304
rect 3125 -2492 3137 -2316
rect 3171 -2492 3183 -2316
rect 3125 -2504 3183 -2492
rect 3243 -2316 3301 -2304
rect 3243 -2492 3255 -2316
rect 3289 -2492 3301 -2316
rect 3243 -2504 3301 -2492
rect 3361 -2316 3419 -2304
rect 3361 -2492 3373 -2316
rect 3407 -2492 3419 -2316
rect 3361 -2504 3419 -2492
rect 3479 -2316 3537 -2304
rect 3479 -2492 3491 -2316
rect 3525 -2492 3537 -2316
rect 3479 -2504 3537 -2492
rect 3597 -2316 3655 -2304
rect 3597 -2492 3609 -2316
rect 3643 -2492 3655 -2316
rect 3597 -2504 3655 -2492
rect 3715 -2316 3773 -2304
rect 3715 -2492 3727 -2316
rect 3761 -2492 3773 -2316
rect 3715 -2504 3773 -2492
rect 3833 -2316 3891 -2304
rect 3833 -2492 3845 -2316
rect 3879 -2492 3891 -2316
rect 3833 -2504 3891 -2492
rect 3951 -2316 4009 -2304
rect 3951 -2492 3963 -2316
rect 3997 -2492 4009 -2316
rect 3951 -2504 4009 -2492
rect 5214 -2620 5226 -2244
rect 5260 -2620 5272 -2244
rect 5214 -2632 5272 -2620
rect 5332 -2244 5390 -2232
rect 5332 -2620 5344 -2244
rect 5378 -2620 5390 -2244
rect 5332 -2632 5390 -2620
rect 5450 -2244 5508 -2232
rect 5450 -2620 5462 -2244
rect 5496 -2620 5508 -2244
rect 5450 -2632 5508 -2620
rect 5568 -2244 5626 -2232
rect 5568 -2620 5580 -2244
rect 5614 -2620 5626 -2244
rect 5568 -2632 5626 -2620
rect 5686 -2244 5744 -2232
rect 5686 -2620 5698 -2244
rect 5732 -2620 5744 -2244
rect 5686 -2632 5744 -2620
rect 5804 -2244 5862 -2232
rect 5804 -2620 5816 -2244
rect 5850 -2620 5862 -2244
rect 5804 -2632 5862 -2620
rect 5922 -2244 5980 -2232
rect 5922 -2620 5934 -2244
rect 5968 -2620 5980 -2244
rect 5922 -2632 5980 -2620
rect 6356 -2240 6414 -2228
rect 6356 -2616 6368 -2240
rect 6402 -2616 6414 -2240
rect 6356 -2628 6414 -2616
rect 6474 -2240 6532 -2228
rect 6474 -2616 6486 -2240
rect 6520 -2616 6532 -2240
rect 6474 -2628 6532 -2616
rect 6592 -2240 6650 -2228
rect 6592 -2616 6604 -2240
rect 6638 -2616 6650 -2240
rect 6592 -2628 6650 -2616
rect 6710 -2240 6768 -2228
rect 6710 -2616 6722 -2240
rect 6756 -2616 6768 -2240
rect 6710 -2628 6768 -2616
rect 6828 -2240 6886 -2228
rect 6828 -2616 6840 -2240
rect 6874 -2616 6886 -2240
rect 6828 -2628 6886 -2616
rect 6946 -2240 7004 -2228
rect 6946 -2616 6958 -2240
rect 6992 -2616 7004 -2240
rect 6946 -2628 7004 -2616
rect 7064 -2240 7122 -2228
rect 28593 -2040 28651 -2028
rect 7064 -2616 7076 -2240
rect 7110 -2616 7122 -2240
rect 11765 -2246 11823 -2234
rect 9440 -2318 9498 -2306
rect 9440 -2494 9452 -2318
rect 9486 -2494 9498 -2318
rect 9440 -2506 9498 -2494
rect 9558 -2318 9616 -2306
rect 9558 -2494 9570 -2318
rect 9604 -2494 9616 -2318
rect 9558 -2506 9616 -2494
rect 9676 -2318 9734 -2306
rect 9676 -2494 9688 -2318
rect 9722 -2494 9734 -2318
rect 9676 -2506 9734 -2494
rect 9794 -2318 9852 -2306
rect 9794 -2494 9806 -2318
rect 9840 -2494 9852 -2318
rect 9794 -2506 9852 -2494
rect 9912 -2318 9970 -2306
rect 9912 -2494 9924 -2318
rect 9958 -2494 9970 -2318
rect 9912 -2506 9970 -2494
rect 10030 -2318 10088 -2306
rect 10030 -2494 10042 -2318
rect 10076 -2494 10088 -2318
rect 10030 -2506 10088 -2494
rect 10148 -2318 10206 -2306
rect 10148 -2494 10160 -2318
rect 10194 -2494 10206 -2318
rect 10148 -2506 10206 -2494
rect 10266 -2318 10324 -2306
rect 10266 -2494 10278 -2318
rect 10312 -2494 10324 -2318
rect 10266 -2506 10324 -2494
rect 10384 -2318 10442 -2306
rect 10384 -2494 10396 -2318
rect 10430 -2494 10442 -2318
rect 10384 -2506 10442 -2494
rect 10502 -2318 10560 -2306
rect 10502 -2494 10514 -2318
rect 10548 -2494 10560 -2318
rect 10502 -2506 10560 -2494
rect 7064 -2628 7122 -2616
rect 11765 -2622 11777 -2246
rect 11811 -2622 11823 -2246
rect 11765 -2634 11823 -2622
rect 11883 -2246 11941 -2234
rect 11883 -2622 11895 -2246
rect 11929 -2622 11941 -2246
rect 11883 -2634 11941 -2622
rect 12001 -2246 12059 -2234
rect 12001 -2622 12013 -2246
rect 12047 -2622 12059 -2246
rect 12001 -2634 12059 -2622
rect 12119 -2246 12177 -2234
rect 12119 -2622 12131 -2246
rect 12165 -2622 12177 -2246
rect 12119 -2634 12177 -2622
rect 12237 -2246 12295 -2234
rect 12237 -2622 12249 -2246
rect 12283 -2622 12295 -2246
rect 12237 -2634 12295 -2622
rect 12355 -2246 12413 -2234
rect 12355 -2622 12367 -2246
rect 12401 -2622 12413 -2246
rect 12355 -2634 12413 -2622
rect 12473 -2246 12531 -2234
rect 12473 -2622 12485 -2246
rect 12519 -2622 12531 -2246
rect 12473 -2634 12531 -2622
rect 12907 -2242 12965 -2230
rect 12907 -2618 12919 -2242
rect 12953 -2618 12965 -2242
rect 12907 -2630 12965 -2618
rect 13025 -2242 13083 -2230
rect 13025 -2618 13037 -2242
rect 13071 -2618 13083 -2242
rect 13025 -2630 13083 -2618
rect 13143 -2242 13201 -2230
rect 13143 -2618 13155 -2242
rect 13189 -2618 13201 -2242
rect 13143 -2630 13201 -2618
rect 13261 -2242 13319 -2230
rect 13261 -2618 13273 -2242
rect 13307 -2618 13319 -2242
rect 13261 -2630 13319 -2618
rect 13379 -2242 13437 -2230
rect 13379 -2618 13391 -2242
rect 13425 -2618 13437 -2242
rect 13379 -2630 13437 -2618
rect 13497 -2242 13555 -2230
rect 13497 -2618 13509 -2242
rect 13543 -2618 13555 -2242
rect 13497 -2630 13555 -2618
rect 13615 -2242 13673 -2230
rect 13615 -2618 13627 -2242
rect 13661 -2618 13673 -2242
rect 18420 -2245 18478 -2233
rect 16095 -2317 16153 -2305
rect 16095 -2493 16107 -2317
rect 16141 -2493 16153 -2317
rect 16095 -2505 16153 -2493
rect 16213 -2317 16271 -2305
rect 16213 -2493 16225 -2317
rect 16259 -2493 16271 -2317
rect 16213 -2505 16271 -2493
rect 16331 -2317 16389 -2305
rect 16331 -2493 16343 -2317
rect 16377 -2493 16389 -2317
rect 16331 -2505 16389 -2493
rect 16449 -2317 16507 -2305
rect 16449 -2493 16461 -2317
rect 16495 -2493 16507 -2317
rect 16449 -2505 16507 -2493
rect 16567 -2317 16625 -2305
rect 16567 -2493 16579 -2317
rect 16613 -2493 16625 -2317
rect 16567 -2505 16625 -2493
rect 16685 -2317 16743 -2305
rect 16685 -2493 16697 -2317
rect 16731 -2493 16743 -2317
rect 16685 -2505 16743 -2493
rect 16803 -2317 16861 -2305
rect 16803 -2493 16815 -2317
rect 16849 -2493 16861 -2317
rect 16803 -2505 16861 -2493
rect 16921 -2317 16979 -2305
rect 16921 -2493 16933 -2317
rect 16967 -2493 16979 -2317
rect 16921 -2505 16979 -2493
rect 17039 -2317 17097 -2305
rect 17039 -2493 17051 -2317
rect 17085 -2493 17097 -2317
rect 17039 -2505 17097 -2493
rect 17157 -2317 17215 -2305
rect 17157 -2493 17169 -2317
rect 17203 -2493 17215 -2317
rect 17157 -2505 17215 -2493
rect 13615 -2630 13673 -2618
rect 5643 -3027 5701 -3015
rect 5643 -3203 5655 -3027
rect 5689 -3203 5701 -3027
rect 5643 -3215 5701 -3203
rect 5761 -3027 5819 -3015
rect 5761 -3203 5773 -3027
rect 5807 -3203 5819 -3027
rect 5761 -3215 5819 -3203
rect 5879 -3027 5937 -3015
rect 5879 -3203 5891 -3027
rect 5925 -3203 5937 -3027
rect 5879 -3215 5937 -3203
rect 5997 -3027 6055 -3015
rect 5997 -3203 6009 -3027
rect 6043 -3203 6055 -3027
rect 5997 -3215 6055 -3203
rect 6785 -3023 6843 -3011
rect 6785 -3199 6797 -3023
rect 6831 -3199 6843 -3023
rect 6785 -3211 6843 -3199
rect 6903 -3023 6961 -3011
rect 6903 -3199 6915 -3023
rect 6949 -3199 6961 -3023
rect 6903 -3211 6961 -3199
rect 7021 -3023 7079 -3011
rect 7021 -3199 7033 -3023
rect 7067 -3199 7079 -3023
rect 7021 -3211 7079 -3199
rect 7139 -3023 7197 -3011
rect 7139 -3199 7151 -3023
rect 7185 -3199 7197 -3023
rect 18420 -2621 18432 -2245
rect 18466 -2621 18478 -2245
rect 18420 -2633 18478 -2621
rect 18538 -2245 18596 -2233
rect 18538 -2621 18550 -2245
rect 18584 -2621 18596 -2245
rect 18538 -2633 18596 -2621
rect 18656 -2245 18714 -2233
rect 18656 -2621 18668 -2245
rect 18702 -2621 18714 -2245
rect 18656 -2633 18714 -2621
rect 18774 -2245 18832 -2233
rect 18774 -2621 18786 -2245
rect 18820 -2621 18832 -2245
rect 18774 -2633 18832 -2621
rect 18892 -2245 18950 -2233
rect 18892 -2621 18904 -2245
rect 18938 -2621 18950 -2245
rect 18892 -2633 18950 -2621
rect 19010 -2245 19068 -2233
rect 19010 -2621 19022 -2245
rect 19056 -2621 19068 -2245
rect 19010 -2633 19068 -2621
rect 19128 -2245 19186 -2233
rect 19128 -2621 19140 -2245
rect 19174 -2621 19186 -2245
rect 19128 -2633 19186 -2621
rect 19562 -2241 19620 -2229
rect 19562 -2617 19574 -2241
rect 19608 -2617 19620 -2241
rect 19562 -2629 19620 -2617
rect 19680 -2241 19738 -2229
rect 19680 -2617 19692 -2241
rect 19726 -2617 19738 -2241
rect 19680 -2629 19738 -2617
rect 19798 -2241 19856 -2229
rect 19798 -2617 19810 -2241
rect 19844 -2617 19856 -2241
rect 19798 -2629 19856 -2617
rect 19916 -2241 19974 -2229
rect 19916 -2617 19928 -2241
rect 19962 -2617 19974 -2241
rect 19916 -2629 19974 -2617
rect 20034 -2241 20092 -2229
rect 20034 -2617 20046 -2241
rect 20080 -2617 20092 -2241
rect 20034 -2629 20092 -2617
rect 20152 -2241 20210 -2229
rect 20152 -2617 20164 -2241
rect 20198 -2617 20210 -2241
rect 20152 -2629 20210 -2617
rect 20270 -2241 20328 -2229
rect 28593 -2216 28605 -2040
rect 28639 -2216 28651 -2040
rect 28593 -2228 28651 -2216
rect 28711 -2040 28769 -2028
rect 28711 -2216 28723 -2040
rect 28757 -2216 28769 -2040
rect 28711 -2228 28769 -2216
rect 28829 -2040 28887 -2028
rect 28829 -2216 28841 -2040
rect 28875 -2216 28887 -2040
rect 28829 -2228 28887 -2216
rect 28947 -2040 29005 -2028
rect 28947 -2216 28959 -2040
rect 28993 -2216 29005 -2040
rect 28947 -2228 29005 -2216
rect 29065 -2040 29123 -2028
rect 29065 -2216 29077 -2040
rect 29111 -2216 29123 -2040
rect 29065 -2228 29123 -2216
rect 29183 -2040 29241 -2028
rect 29183 -2216 29195 -2040
rect 29229 -2216 29241 -2040
rect 29183 -2228 29241 -2216
rect 29301 -2040 29359 -2028
rect 29301 -2216 29313 -2040
rect 29347 -2216 29359 -2040
rect 29301 -2228 29359 -2216
rect 29419 -2040 29477 -2028
rect 29419 -2216 29431 -2040
rect 29465 -2216 29477 -2040
rect 29419 -2228 29477 -2216
rect 29537 -2040 29595 -2028
rect 29537 -2216 29549 -2040
rect 29583 -2216 29595 -2040
rect 29537 -2228 29595 -2216
rect 29655 -2040 29713 -2028
rect 29655 -2216 29667 -2040
rect 29701 -2216 29713 -2040
rect 29655 -2228 29713 -2216
rect 20270 -2617 20282 -2241
rect 20316 -2617 20328 -2241
rect 25042 -2244 25100 -2232
rect 22717 -2316 22775 -2304
rect 22717 -2492 22729 -2316
rect 22763 -2492 22775 -2316
rect 22717 -2504 22775 -2492
rect 22835 -2316 22893 -2304
rect 22835 -2492 22847 -2316
rect 22881 -2492 22893 -2316
rect 22835 -2504 22893 -2492
rect 22953 -2316 23011 -2304
rect 22953 -2492 22965 -2316
rect 22999 -2492 23011 -2316
rect 22953 -2504 23011 -2492
rect 23071 -2316 23129 -2304
rect 23071 -2492 23083 -2316
rect 23117 -2492 23129 -2316
rect 23071 -2504 23129 -2492
rect 23189 -2316 23247 -2304
rect 23189 -2492 23201 -2316
rect 23235 -2492 23247 -2316
rect 23189 -2504 23247 -2492
rect 23307 -2316 23365 -2304
rect 23307 -2492 23319 -2316
rect 23353 -2492 23365 -2316
rect 23307 -2504 23365 -2492
rect 23425 -2316 23483 -2304
rect 23425 -2492 23437 -2316
rect 23471 -2492 23483 -2316
rect 23425 -2504 23483 -2492
rect 23543 -2316 23601 -2304
rect 23543 -2492 23555 -2316
rect 23589 -2492 23601 -2316
rect 23543 -2504 23601 -2492
rect 23661 -2316 23719 -2304
rect 23661 -2492 23673 -2316
rect 23707 -2492 23719 -2316
rect 23661 -2504 23719 -2492
rect 23779 -2316 23837 -2304
rect 23779 -2492 23791 -2316
rect 23825 -2492 23837 -2316
rect 23779 -2504 23837 -2492
rect 20270 -2629 20328 -2617
rect 7139 -3211 7197 -3199
rect 12194 -3029 12252 -3017
rect 12194 -3205 12206 -3029
rect 12240 -3205 12252 -3029
rect 12194 -3217 12252 -3205
rect 12312 -3029 12370 -3017
rect 12312 -3205 12324 -3029
rect 12358 -3205 12370 -3029
rect 12312 -3217 12370 -3205
rect 12430 -3029 12488 -3017
rect 12430 -3205 12442 -3029
rect 12476 -3205 12488 -3029
rect 12430 -3217 12488 -3205
rect 12548 -3029 12606 -3017
rect 12548 -3205 12560 -3029
rect 12594 -3205 12606 -3029
rect 12548 -3217 12606 -3205
rect 13336 -3025 13394 -3013
rect 13336 -3201 13348 -3025
rect 13382 -3201 13394 -3025
rect 13336 -3213 13394 -3201
rect 13454 -3025 13512 -3013
rect 13454 -3201 13466 -3025
rect 13500 -3201 13512 -3025
rect 13454 -3213 13512 -3201
rect 13572 -3025 13630 -3013
rect 13572 -3201 13584 -3025
rect 13618 -3201 13630 -3025
rect 13572 -3213 13630 -3201
rect 13690 -3025 13748 -3013
rect 13690 -3201 13702 -3025
rect 13736 -3201 13748 -3025
rect 25042 -2620 25054 -2244
rect 25088 -2620 25100 -2244
rect 25042 -2632 25100 -2620
rect 25160 -2244 25218 -2232
rect 25160 -2620 25172 -2244
rect 25206 -2620 25218 -2244
rect 25160 -2632 25218 -2620
rect 25278 -2244 25336 -2232
rect 25278 -2620 25290 -2244
rect 25324 -2620 25336 -2244
rect 25278 -2632 25336 -2620
rect 25396 -2244 25454 -2232
rect 25396 -2620 25408 -2244
rect 25442 -2620 25454 -2244
rect 25396 -2632 25454 -2620
rect 25514 -2244 25572 -2232
rect 25514 -2620 25526 -2244
rect 25560 -2620 25572 -2244
rect 25514 -2632 25572 -2620
rect 25632 -2244 25690 -2232
rect 25632 -2620 25644 -2244
rect 25678 -2620 25690 -2244
rect 25632 -2632 25690 -2620
rect 25750 -2244 25808 -2232
rect 25750 -2620 25762 -2244
rect 25796 -2620 25808 -2244
rect 25750 -2632 25808 -2620
rect 26184 -2240 26242 -2228
rect 26184 -2616 26196 -2240
rect 26230 -2616 26242 -2240
rect 26184 -2628 26242 -2616
rect 26302 -2240 26360 -2228
rect 26302 -2616 26314 -2240
rect 26348 -2616 26360 -2240
rect 26302 -2628 26360 -2616
rect 26420 -2240 26478 -2228
rect 26420 -2616 26432 -2240
rect 26466 -2616 26478 -2240
rect 26420 -2628 26478 -2616
rect 26538 -2240 26596 -2228
rect 26538 -2616 26550 -2240
rect 26584 -2616 26596 -2240
rect 26538 -2628 26596 -2616
rect 26656 -2240 26714 -2228
rect 26656 -2616 26668 -2240
rect 26702 -2616 26714 -2240
rect 26656 -2628 26714 -2616
rect 26774 -2240 26832 -2228
rect 26774 -2616 26786 -2240
rect 26820 -2616 26832 -2240
rect 26774 -2628 26832 -2616
rect 26892 -2240 26950 -2228
rect 26892 -2616 26904 -2240
rect 26938 -2616 26950 -2240
rect 30821 -2307 30879 -2295
rect 26892 -2628 26950 -2616
rect 13690 -3213 13748 -3201
rect 18849 -3028 18907 -3016
rect 18849 -3204 18861 -3028
rect 18895 -3204 18907 -3028
rect 18849 -3216 18907 -3204
rect 18967 -3028 19025 -3016
rect 18967 -3204 18979 -3028
rect 19013 -3204 19025 -3028
rect 18967 -3216 19025 -3204
rect 19085 -3028 19143 -3016
rect 19085 -3204 19097 -3028
rect 19131 -3204 19143 -3028
rect 19085 -3216 19143 -3204
rect 19203 -3028 19261 -3016
rect 19203 -3204 19215 -3028
rect 19249 -3204 19261 -3028
rect 19203 -3216 19261 -3204
rect 19991 -3024 20049 -3012
rect 19991 -3200 20003 -3024
rect 20037 -3200 20049 -3024
rect 19991 -3212 20049 -3200
rect 20109 -3024 20167 -3012
rect 20109 -3200 20121 -3024
rect 20155 -3200 20167 -3024
rect 20109 -3212 20167 -3200
rect 20227 -3024 20285 -3012
rect 20227 -3200 20239 -3024
rect 20273 -3200 20285 -3024
rect 20227 -3212 20285 -3200
rect 20345 -3024 20403 -3012
rect 20345 -3200 20357 -3024
rect 20391 -3200 20403 -3024
rect 30337 -2507 30395 -2495
rect 30337 -2683 30349 -2507
rect 30383 -2683 30395 -2507
rect 30337 -2695 30395 -2683
rect 30455 -2507 30513 -2495
rect 30455 -2683 30467 -2507
rect 30501 -2683 30513 -2507
rect 30455 -2695 30513 -2683
rect 30573 -2507 30631 -2495
rect 30573 -2683 30585 -2507
rect 30619 -2683 30631 -2507
rect 30573 -2695 30631 -2683
rect 30691 -2507 30749 -2495
rect 30691 -2683 30703 -2507
rect 30737 -2683 30749 -2507
rect 30691 -2695 30749 -2683
rect 30821 -2683 30833 -2307
rect 30867 -2683 30879 -2307
rect 30821 -2695 30879 -2683
rect 30939 -2307 30997 -2295
rect 30939 -2683 30951 -2307
rect 30985 -2683 30997 -2307
rect 30939 -2695 30997 -2683
rect 31057 -2307 31115 -2295
rect 31057 -2683 31069 -2307
rect 31103 -2683 31115 -2307
rect 31057 -2695 31115 -2683
rect 31175 -2307 31233 -2295
rect 31175 -2683 31187 -2307
rect 31221 -2683 31233 -2307
rect 31175 -2695 31233 -2683
rect 31293 -2307 31351 -2295
rect 31293 -2683 31305 -2307
rect 31339 -2683 31351 -2307
rect 31293 -2695 31351 -2683
rect 31411 -2307 31469 -2295
rect 31411 -2683 31423 -2307
rect 31457 -2683 31469 -2307
rect 31411 -2695 31469 -2683
rect 31529 -2307 31587 -2295
rect 31529 -2683 31541 -2307
rect 31575 -2683 31587 -2307
rect 31529 -2695 31587 -2683
rect 31658 -2507 31716 -2495
rect 31658 -2683 31670 -2507
rect 31704 -2683 31716 -2507
rect 31658 -2695 31716 -2683
rect 31776 -2507 31834 -2495
rect 31776 -2683 31788 -2507
rect 31822 -2683 31834 -2507
rect 31776 -2695 31834 -2683
rect 31894 -2507 31952 -2495
rect 31894 -2683 31906 -2507
rect 31940 -2683 31952 -2507
rect 31894 -2695 31952 -2683
rect 32012 -2507 32070 -2495
rect 32012 -2683 32024 -2507
rect 32058 -2683 32070 -2507
rect 32012 -2695 32070 -2683
rect 32130 -2510 32188 -2498
rect 32130 -2686 32142 -2510
rect 32176 -2686 32188 -2510
rect 32130 -2698 32188 -2686
rect 32248 -2510 32306 -2498
rect 32248 -2686 32260 -2510
rect 32294 -2686 32306 -2510
rect 32248 -2698 32306 -2686
rect 32366 -2510 32424 -2498
rect 32366 -2686 32378 -2510
rect 32412 -2686 32424 -2510
rect 32366 -2698 32424 -2686
rect 32484 -2510 32542 -2498
rect 32484 -2686 32496 -2510
rect 32530 -2686 32542 -2510
rect 32484 -2698 32542 -2686
rect 32602 -2510 32660 -2498
rect 32602 -2686 32614 -2510
rect 32648 -2686 32660 -2510
rect 32602 -2698 32660 -2686
rect 32720 -2510 32778 -2498
rect 32720 -2686 32732 -2510
rect 32766 -2686 32778 -2510
rect 32720 -2698 32778 -2686
rect 32838 -2510 32896 -2498
rect 32838 -2686 32850 -2510
rect 32884 -2686 32896 -2510
rect 32838 -2698 32896 -2686
rect 32956 -2510 33014 -2498
rect 32956 -2686 32968 -2510
rect 33002 -2686 33014 -2510
rect 32956 -2698 33014 -2686
rect 33074 -2510 33132 -2498
rect 33074 -2686 33086 -2510
rect 33120 -2686 33132 -2510
rect 33074 -2698 33132 -2686
rect 33192 -2510 33250 -2498
rect 33192 -2686 33204 -2510
rect 33238 -2686 33250 -2510
rect 33192 -2698 33250 -2686
rect 20345 -3212 20403 -3200
rect 25471 -3027 25529 -3015
rect 25471 -3203 25483 -3027
rect 25517 -3203 25529 -3027
rect 25471 -3215 25529 -3203
rect 25589 -3027 25647 -3015
rect 25589 -3203 25601 -3027
rect 25635 -3203 25647 -3027
rect 25589 -3215 25647 -3203
rect 25707 -3027 25765 -3015
rect 25707 -3203 25719 -3027
rect 25753 -3203 25765 -3027
rect 25707 -3215 25765 -3203
rect 25825 -3027 25883 -3015
rect 25825 -3203 25837 -3027
rect 25871 -3203 25883 -3027
rect 25825 -3215 25883 -3203
rect 26613 -3023 26671 -3011
rect 26613 -3199 26625 -3023
rect 26659 -3199 26671 -3023
rect 26613 -3211 26671 -3199
rect 26731 -3023 26789 -3011
rect 26731 -3199 26743 -3023
rect 26777 -3199 26789 -3023
rect 26731 -3211 26789 -3199
rect 26849 -3023 26907 -3011
rect 26849 -3199 26861 -3023
rect 26895 -3199 26907 -3023
rect 26849 -3211 26907 -3199
rect 26967 -3023 27025 -3011
rect 26967 -3199 26979 -3023
rect 27013 -3199 27025 -3023
rect 30764 -3000 30822 -2988
rect 26967 -3211 27025 -3199
rect 30764 -3376 30776 -3000
rect 30810 -3376 30822 -3000
rect 30764 -3388 30822 -3376
rect 30882 -3000 30940 -2988
rect 30882 -3376 30894 -3000
rect 30928 -3376 30940 -3000
rect 30882 -3388 30940 -3376
rect 31000 -3000 31058 -2988
rect 31000 -3376 31012 -3000
rect 31046 -3376 31058 -3000
rect 31000 -3388 31058 -3376
rect 31118 -3000 31176 -2988
rect 31118 -3376 31130 -3000
rect 31164 -3376 31176 -3000
rect 31118 -3388 31176 -3376
rect 31236 -3000 31294 -2988
rect 31236 -3376 31248 -3000
rect 31282 -3376 31294 -3000
rect 31236 -3388 31294 -3376
rect 31354 -3000 31412 -2988
rect 31354 -3376 31366 -3000
rect 31400 -3376 31412 -3000
rect 31354 -3388 31412 -3376
rect 31472 -3000 31530 -2988
rect 31472 -3376 31484 -3000
rect 31518 -3376 31530 -3000
rect 31472 -3388 31530 -3376
rect 2903 -3966 2961 -3954
rect 2903 -4142 2915 -3966
rect 2949 -4142 2961 -3966
rect 2903 -4154 2961 -4142
rect 3021 -3966 3079 -3954
rect 3021 -4142 3033 -3966
rect 3067 -4142 3079 -3966
rect 3021 -4154 3079 -4142
rect 3139 -3966 3197 -3954
rect 3139 -4142 3151 -3966
rect 3185 -4142 3197 -3966
rect 3139 -4154 3197 -4142
rect 3257 -3966 3315 -3954
rect 3257 -4142 3269 -3966
rect 3303 -4142 3315 -3966
rect 3257 -4154 3315 -4142
rect 3375 -3966 3433 -3954
rect 3375 -4142 3387 -3966
rect 3421 -4142 3433 -3966
rect 3375 -4154 3433 -4142
rect 3493 -3966 3551 -3954
rect 3493 -4142 3505 -3966
rect 3539 -4142 3551 -3966
rect 3493 -4154 3551 -4142
rect 3611 -3966 3669 -3954
rect 3611 -4142 3623 -3966
rect 3657 -4142 3669 -3966
rect 3611 -4154 3669 -4142
rect 3729 -3966 3787 -3954
rect 3729 -4142 3741 -3966
rect 3775 -4142 3787 -3966
rect 3729 -4154 3787 -4142
rect 3847 -3966 3905 -3954
rect 3847 -4142 3859 -3966
rect 3893 -4142 3905 -3966
rect 3847 -4154 3905 -4142
rect 3965 -3966 4023 -3954
rect 3965 -4142 3977 -3966
rect 4011 -4142 4023 -3966
rect 9454 -3968 9512 -3956
rect 3965 -4154 4023 -4142
rect 9454 -4144 9466 -3968
rect 9500 -4144 9512 -3968
rect 9454 -4156 9512 -4144
rect 9572 -3968 9630 -3956
rect 9572 -4144 9584 -3968
rect 9618 -4144 9630 -3968
rect 9572 -4156 9630 -4144
rect 9690 -3968 9748 -3956
rect 9690 -4144 9702 -3968
rect 9736 -4144 9748 -3968
rect 9690 -4156 9748 -4144
rect 9808 -3968 9866 -3956
rect 9808 -4144 9820 -3968
rect 9854 -4144 9866 -3968
rect 9808 -4156 9866 -4144
rect 9926 -3968 9984 -3956
rect 9926 -4144 9938 -3968
rect 9972 -4144 9984 -3968
rect 9926 -4156 9984 -4144
rect 10044 -3968 10102 -3956
rect 10044 -4144 10056 -3968
rect 10090 -4144 10102 -3968
rect 10044 -4156 10102 -4144
rect 10162 -3968 10220 -3956
rect 10162 -4144 10174 -3968
rect 10208 -4144 10220 -3968
rect 10162 -4156 10220 -4144
rect 10280 -3968 10338 -3956
rect 10280 -4144 10292 -3968
rect 10326 -4144 10338 -3968
rect 10280 -4156 10338 -4144
rect 10398 -3968 10456 -3956
rect 10398 -4144 10410 -3968
rect 10444 -4144 10456 -3968
rect 10398 -4156 10456 -4144
rect 10516 -3968 10574 -3956
rect 10516 -4144 10528 -3968
rect 10562 -4144 10574 -3968
rect 16109 -3967 16167 -3955
rect 10516 -4156 10574 -4144
rect 16109 -4143 16121 -3967
rect 16155 -4143 16167 -3967
rect 16109 -4155 16167 -4143
rect 16227 -3967 16285 -3955
rect 16227 -4143 16239 -3967
rect 16273 -4143 16285 -3967
rect 16227 -4155 16285 -4143
rect 16345 -3967 16403 -3955
rect 16345 -4143 16357 -3967
rect 16391 -4143 16403 -3967
rect 16345 -4155 16403 -4143
rect 16463 -3967 16521 -3955
rect 16463 -4143 16475 -3967
rect 16509 -4143 16521 -3967
rect 16463 -4155 16521 -4143
rect 16581 -3967 16639 -3955
rect 16581 -4143 16593 -3967
rect 16627 -4143 16639 -3967
rect 16581 -4155 16639 -4143
rect 16699 -3967 16757 -3955
rect 16699 -4143 16711 -3967
rect 16745 -4143 16757 -3967
rect 16699 -4155 16757 -4143
rect 16817 -3967 16875 -3955
rect 16817 -4143 16829 -3967
rect 16863 -4143 16875 -3967
rect 16817 -4155 16875 -4143
rect 16935 -3967 16993 -3955
rect 16935 -4143 16947 -3967
rect 16981 -4143 16993 -3967
rect 16935 -4155 16993 -4143
rect 17053 -3967 17111 -3955
rect 17053 -4143 17065 -3967
rect 17099 -4143 17111 -3967
rect 17053 -4155 17111 -4143
rect 17171 -3967 17229 -3955
rect 17171 -4143 17183 -3967
rect 17217 -4143 17229 -3967
rect 22731 -3966 22789 -3954
rect 17171 -4155 17229 -4143
rect 22731 -4142 22743 -3966
rect 22777 -4142 22789 -3966
rect 22731 -4154 22789 -4142
rect 22849 -3966 22907 -3954
rect 22849 -4142 22861 -3966
rect 22895 -4142 22907 -3966
rect 22849 -4154 22907 -4142
rect 22967 -3966 23025 -3954
rect 22967 -4142 22979 -3966
rect 23013 -4142 23025 -3966
rect 22967 -4154 23025 -4142
rect 23085 -3966 23143 -3954
rect 23085 -4142 23097 -3966
rect 23131 -4142 23143 -3966
rect 23085 -4154 23143 -4142
rect 23203 -3966 23261 -3954
rect 23203 -4142 23215 -3966
rect 23249 -4142 23261 -3966
rect 23203 -4154 23261 -4142
rect 23321 -3966 23379 -3954
rect 23321 -4142 23333 -3966
rect 23367 -4142 23379 -3966
rect 23321 -4154 23379 -4142
rect 23439 -3966 23497 -3954
rect 23439 -4142 23451 -3966
rect 23485 -4142 23497 -3966
rect 23439 -4154 23497 -4142
rect 23557 -3966 23615 -3954
rect 23557 -4142 23569 -3966
rect 23603 -4142 23615 -3966
rect 23557 -4154 23615 -4142
rect 23675 -3966 23733 -3954
rect 23675 -4142 23687 -3966
rect 23721 -4142 23733 -3966
rect 23675 -4154 23733 -4142
rect 23793 -3966 23851 -3954
rect 23793 -4142 23805 -3966
rect 23839 -4142 23851 -3966
rect 23793 -4154 23851 -4142
rect 4851 -4383 4909 -4371
rect 4367 -4583 4425 -4571
rect 4367 -4759 4379 -4583
rect 4413 -4759 4425 -4583
rect 4367 -4771 4425 -4759
rect 4485 -4583 4543 -4571
rect 4485 -4759 4497 -4583
rect 4531 -4759 4543 -4583
rect 4485 -4771 4543 -4759
rect 4603 -4583 4661 -4571
rect 4603 -4759 4615 -4583
rect 4649 -4759 4661 -4583
rect 4603 -4771 4661 -4759
rect 4721 -4583 4779 -4571
rect 4721 -4759 4733 -4583
rect 4767 -4759 4779 -4583
rect 4721 -4771 4779 -4759
rect 4851 -4759 4863 -4383
rect 4897 -4759 4909 -4383
rect 4851 -4771 4909 -4759
rect 4969 -4383 5027 -4371
rect 4969 -4759 4981 -4383
rect 5015 -4759 5027 -4383
rect 4969 -4771 5027 -4759
rect 5087 -4383 5145 -4371
rect 5087 -4759 5099 -4383
rect 5133 -4759 5145 -4383
rect 5087 -4771 5145 -4759
rect 5205 -4383 5263 -4371
rect 5205 -4759 5217 -4383
rect 5251 -4759 5263 -4383
rect 5205 -4771 5263 -4759
rect 5323 -4383 5381 -4371
rect 5323 -4759 5335 -4383
rect 5369 -4759 5381 -4383
rect 5323 -4771 5381 -4759
rect 5441 -4383 5499 -4371
rect 5441 -4759 5453 -4383
rect 5487 -4759 5499 -4383
rect 5441 -4771 5499 -4759
rect 5559 -4383 5617 -4371
rect 5559 -4759 5571 -4383
rect 5605 -4759 5617 -4383
rect 6749 -4383 6807 -4371
rect 5559 -4771 5617 -4759
rect 5688 -4583 5746 -4571
rect 5688 -4759 5700 -4583
rect 5734 -4759 5746 -4583
rect 5688 -4771 5746 -4759
rect 5806 -4583 5864 -4571
rect 5806 -4759 5818 -4583
rect 5852 -4759 5864 -4583
rect 5806 -4771 5864 -4759
rect 5924 -4583 5982 -4571
rect 5924 -4759 5936 -4583
rect 5970 -4759 5982 -4583
rect 5924 -4771 5982 -4759
rect 6042 -4583 6100 -4571
rect 6042 -4759 6054 -4583
rect 6088 -4759 6100 -4583
rect 6042 -4771 6100 -4759
rect 6265 -4583 6323 -4571
rect 6265 -4759 6277 -4583
rect 6311 -4759 6323 -4583
rect 6265 -4771 6323 -4759
rect 6383 -4583 6441 -4571
rect 6383 -4759 6395 -4583
rect 6429 -4759 6441 -4583
rect 6383 -4771 6441 -4759
rect 6501 -4583 6559 -4571
rect 6501 -4759 6513 -4583
rect 6547 -4759 6559 -4583
rect 6501 -4771 6559 -4759
rect 6619 -4583 6677 -4571
rect 6619 -4759 6631 -4583
rect 6665 -4759 6677 -4583
rect 6619 -4771 6677 -4759
rect 6749 -4759 6761 -4383
rect 6795 -4759 6807 -4383
rect 6749 -4771 6807 -4759
rect 6867 -4383 6925 -4371
rect 6867 -4759 6879 -4383
rect 6913 -4759 6925 -4383
rect 6867 -4771 6925 -4759
rect 6985 -4383 7043 -4371
rect 6985 -4759 6997 -4383
rect 7031 -4759 7043 -4383
rect 6985 -4771 7043 -4759
rect 7103 -4383 7161 -4371
rect 7103 -4759 7115 -4383
rect 7149 -4759 7161 -4383
rect 7103 -4771 7161 -4759
rect 7221 -4383 7279 -4371
rect 7221 -4759 7233 -4383
rect 7267 -4759 7279 -4383
rect 7221 -4771 7279 -4759
rect 7339 -4383 7397 -4371
rect 7339 -4759 7351 -4383
rect 7385 -4759 7397 -4383
rect 7339 -4771 7397 -4759
rect 7457 -4383 7515 -4371
rect 7457 -4759 7469 -4383
rect 7503 -4759 7515 -4383
rect 11402 -4385 11460 -4373
rect 7457 -4771 7515 -4759
rect 7586 -4583 7644 -4571
rect 7586 -4759 7598 -4583
rect 7632 -4759 7644 -4583
rect 7586 -4771 7644 -4759
rect 7704 -4583 7762 -4571
rect 7704 -4759 7716 -4583
rect 7750 -4759 7762 -4583
rect 7704 -4771 7762 -4759
rect 7822 -4583 7880 -4571
rect 7822 -4759 7834 -4583
rect 7868 -4759 7880 -4583
rect 7822 -4771 7880 -4759
rect 7940 -4583 7998 -4571
rect 7940 -4759 7952 -4583
rect 7986 -4759 7998 -4583
rect 7940 -4771 7998 -4759
rect -4 -4892 54 -4880
rect -4 -5068 8 -4892
rect 42 -5068 54 -4892
rect -4 -5080 54 -5068
rect 114 -4892 172 -4880
rect 114 -5068 126 -4892
rect 160 -5068 172 -4892
rect 114 -5080 172 -5068
rect 232 -4892 290 -4880
rect 232 -5068 244 -4892
rect 278 -5068 290 -4892
rect 232 -5080 290 -5068
rect 350 -4892 408 -4880
rect 350 -5068 362 -4892
rect 396 -5068 408 -4892
rect 350 -5080 408 -5068
rect 468 -4892 526 -4880
rect 468 -5068 480 -4892
rect 514 -5068 526 -4892
rect 468 -5080 526 -5068
rect 586 -4892 644 -4880
rect 586 -5068 598 -4892
rect 632 -5068 644 -4892
rect 586 -5080 644 -5068
rect 704 -4892 762 -4880
rect 704 -5068 716 -4892
rect 750 -5068 762 -4892
rect 704 -5080 762 -5068
rect 822 -4892 880 -4880
rect 822 -5068 834 -4892
rect 868 -5068 880 -4892
rect 822 -5080 880 -5068
rect 940 -4892 998 -4880
rect 940 -5068 952 -4892
rect 986 -5068 998 -4892
rect 940 -5080 998 -5068
rect 1058 -4892 1116 -4880
rect 1058 -5068 1070 -4892
rect 1104 -5068 1116 -4892
rect 1058 -5080 1116 -5068
rect 2898 -5570 2956 -5558
rect 2898 -5746 2910 -5570
rect 2944 -5746 2956 -5570
rect 2898 -5758 2956 -5746
rect 3016 -5570 3074 -5558
rect 3016 -5746 3028 -5570
rect 3062 -5746 3074 -5570
rect 3016 -5758 3074 -5746
rect 3134 -5570 3192 -5558
rect 3134 -5746 3146 -5570
rect 3180 -5746 3192 -5570
rect 3134 -5758 3192 -5746
rect 3252 -5570 3310 -5558
rect 3252 -5746 3264 -5570
rect 3298 -5746 3310 -5570
rect 3252 -5758 3310 -5746
rect 3370 -5570 3428 -5558
rect 3370 -5746 3382 -5570
rect 3416 -5746 3428 -5570
rect 3370 -5758 3428 -5746
rect 3488 -5570 3546 -5558
rect 3488 -5746 3500 -5570
rect 3534 -5746 3546 -5570
rect 3488 -5758 3546 -5746
rect 3606 -5570 3664 -5558
rect 3606 -5746 3618 -5570
rect 3652 -5746 3664 -5570
rect 3606 -5758 3664 -5746
rect 3724 -5570 3782 -5558
rect 3724 -5746 3736 -5570
rect 3770 -5746 3782 -5570
rect 3724 -5758 3782 -5746
rect 3842 -5570 3900 -5558
rect 3842 -5746 3854 -5570
rect 3888 -5746 3900 -5570
rect 3842 -5758 3900 -5746
rect 3960 -5570 4018 -5558
rect 3960 -5746 3972 -5570
rect 4006 -5746 4018 -5570
rect 3960 -5758 4018 -5746
rect 4794 -5076 4852 -5064
rect 4794 -5452 4806 -5076
rect 4840 -5452 4852 -5076
rect 4794 -5464 4852 -5452
rect 4912 -5076 4970 -5064
rect 4912 -5452 4924 -5076
rect 4958 -5452 4970 -5076
rect 4912 -5464 4970 -5452
rect 5030 -5076 5088 -5064
rect 5030 -5452 5042 -5076
rect 5076 -5452 5088 -5076
rect 5030 -5464 5088 -5452
rect 5148 -5076 5206 -5064
rect 5148 -5452 5160 -5076
rect 5194 -5452 5206 -5076
rect 5148 -5464 5206 -5452
rect 5266 -5076 5324 -5064
rect 5266 -5452 5278 -5076
rect 5312 -5452 5324 -5076
rect 5266 -5464 5324 -5452
rect 5384 -5076 5442 -5064
rect 5384 -5452 5396 -5076
rect 5430 -5452 5442 -5076
rect 5384 -5464 5442 -5452
rect 5502 -5076 5560 -5064
rect 5502 -5452 5514 -5076
rect 5548 -5452 5560 -5076
rect 5502 -5464 5560 -5452
rect 10918 -4585 10976 -4573
rect 10918 -4761 10930 -4585
rect 10964 -4761 10976 -4585
rect 10918 -4773 10976 -4761
rect 11036 -4585 11094 -4573
rect 11036 -4761 11048 -4585
rect 11082 -4761 11094 -4585
rect 11036 -4773 11094 -4761
rect 11154 -4585 11212 -4573
rect 11154 -4761 11166 -4585
rect 11200 -4761 11212 -4585
rect 11154 -4773 11212 -4761
rect 11272 -4585 11330 -4573
rect 11272 -4761 11284 -4585
rect 11318 -4761 11330 -4585
rect 11272 -4773 11330 -4761
rect 11402 -4761 11414 -4385
rect 11448 -4761 11460 -4385
rect 11402 -4773 11460 -4761
rect 11520 -4385 11578 -4373
rect 11520 -4761 11532 -4385
rect 11566 -4761 11578 -4385
rect 11520 -4773 11578 -4761
rect 11638 -4385 11696 -4373
rect 11638 -4761 11650 -4385
rect 11684 -4761 11696 -4385
rect 11638 -4773 11696 -4761
rect 11756 -4385 11814 -4373
rect 11756 -4761 11768 -4385
rect 11802 -4761 11814 -4385
rect 11756 -4773 11814 -4761
rect 11874 -4385 11932 -4373
rect 11874 -4761 11886 -4385
rect 11920 -4761 11932 -4385
rect 11874 -4773 11932 -4761
rect 11992 -4385 12050 -4373
rect 11992 -4761 12004 -4385
rect 12038 -4761 12050 -4385
rect 11992 -4773 12050 -4761
rect 12110 -4385 12168 -4373
rect 12110 -4761 12122 -4385
rect 12156 -4761 12168 -4385
rect 13300 -4385 13358 -4373
rect 12110 -4773 12168 -4761
rect 12239 -4585 12297 -4573
rect 12239 -4761 12251 -4585
rect 12285 -4761 12297 -4585
rect 12239 -4773 12297 -4761
rect 12357 -4585 12415 -4573
rect 12357 -4761 12369 -4585
rect 12403 -4761 12415 -4585
rect 12357 -4773 12415 -4761
rect 12475 -4585 12533 -4573
rect 12475 -4761 12487 -4585
rect 12521 -4761 12533 -4585
rect 12475 -4773 12533 -4761
rect 12593 -4585 12651 -4573
rect 12593 -4761 12605 -4585
rect 12639 -4761 12651 -4585
rect 12593 -4773 12651 -4761
rect 12816 -4585 12874 -4573
rect 12816 -4761 12828 -4585
rect 12862 -4761 12874 -4585
rect 12816 -4773 12874 -4761
rect 12934 -4585 12992 -4573
rect 12934 -4761 12946 -4585
rect 12980 -4761 12992 -4585
rect 12934 -4773 12992 -4761
rect 13052 -4585 13110 -4573
rect 13052 -4761 13064 -4585
rect 13098 -4761 13110 -4585
rect 13052 -4773 13110 -4761
rect 13170 -4585 13228 -4573
rect 13170 -4761 13182 -4585
rect 13216 -4761 13228 -4585
rect 13170 -4773 13228 -4761
rect 13300 -4761 13312 -4385
rect 13346 -4761 13358 -4385
rect 13300 -4773 13358 -4761
rect 13418 -4385 13476 -4373
rect 13418 -4761 13430 -4385
rect 13464 -4761 13476 -4385
rect 13418 -4773 13476 -4761
rect 13536 -4385 13594 -4373
rect 13536 -4761 13548 -4385
rect 13582 -4761 13594 -4385
rect 13536 -4773 13594 -4761
rect 13654 -4385 13712 -4373
rect 13654 -4761 13666 -4385
rect 13700 -4761 13712 -4385
rect 13654 -4773 13712 -4761
rect 13772 -4385 13830 -4373
rect 13772 -4761 13784 -4385
rect 13818 -4761 13830 -4385
rect 13772 -4773 13830 -4761
rect 13890 -4385 13948 -4373
rect 13890 -4761 13902 -4385
rect 13936 -4761 13948 -4385
rect 13890 -4773 13948 -4761
rect 14008 -4385 14066 -4373
rect 14008 -4761 14020 -4385
rect 14054 -4761 14066 -4385
rect 18057 -4384 18115 -4372
rect 14008 -4773 14066 -4761
rect 14137 -4585 14195 -4573
rect 14137 -4761 14149 -4585
rect 14183 -4761 14195 -4585
rect 14137 -4773 14195 -4761
rect 14255 -4585 14313 -4573
rect 14255 -4761 14267 -4585
rect 14301 -4761 14313 -4585
rect 14255 -4773 14313 -4761
rect 14373 -4585 14431 -4573
rect 14373 -4761 14385 -4585
rect 14419 -4761 14431 -4585
rect 14373 -4773 14431 -4761
rect 14491 -4585 14549 -4573
rect 14491 -4761 14503 -4585
rect 14537 -4761 14549 -4585
rect 14491 -4773 14549 -4761
rect 6692 -5076 6750 -5064
rect 6692 -5452 6704 -5076
rect 6738 -5452 6750 -5076
rect 6692 -5464 6750 -5452
rect 6810 -5076 6868 -5064
rect 6810 -5452 6822 -5076
rect 6856 -5452 6868 -5076
rect 6810 -5464 6868 -5452
rect 6928 -5076 6986 -5064
rect 6928 -5452 6940 -5076
rect 6974 -5452 6986 -5076
rect 6928 -5464 6986 -5452
rect 7046 -5076 7104 -5064
rect 7046 -5452 7058 -5076
rect 7092 -5452 7104 -5076
rect 7046 -5464 7104 -5452
rect 7164 -5076 7222 -5064
rect 7164 -5452 7176 -5076
rect 7210 -5452 7222 -5076
rect 7164 -5464 7222 -5452
rect 7282 -5076 7340 -5064
rect 7282 -5452 7294 -5076
rect 7328 -5452 7340 -5076
rect 7282 -5464 7340 -5452
rect 7400 -5076 7458 -5064
rect 7400 -5452 7412 -5076
rect 7446 -5452 7458 -5076
rect 7400 -5464 7458 -5452
rect 9449 -5572 9507 -5560
rect 9449 -5748 9461 -5572
rect 9495 -5748 9507 -5572
rect 9449 -5760 9507 -5748
rect 9567 -5572 9625 -5560
rect 9567 -5748 9579 -5572
rect 9613 -5748 9625 -5572
rect 9567 -5760 9625 -5748
rect 9685 -5572 9743 -5560
rect 9685 -5748 9697 -5572
rect 9731 -5748 9743 -5572
rect 9685 -5760 9743 -5748
rect 9803 -5572 9861 -5560
rect 9803 -5748 9815 -5572
rect 9849 -5748 9861 -5572
rect 9803 -5760 9861 -5748
rect 9921 -5572 9979 -5560
rect 9921 -5748 9933 -5572
rect 9967 -5748 9979 -5572
rect 9921 -5760 9979 -5748
rect 10039 -5572 10097 -5560
rect 10039 -5748 10051 -5572
rect 10085 -5748 10097 -5572
rect 10039 -5760 10097 -5748
rect 10157 -5572 10215 -5560
rect 10157 -5748 10169 -5572
rect 10203 -5748 10215 -5572
rect 10157 -5760 10215 -5748
rect 10275 -5572 10333 -5560
rect 10275 -5748 10287 -5572
rect 10321 -5748 10333 -5572
rect 10275 -5760 10333 -5748
rect 10393 -5572 10451 -5560
rect 10393 -5748 10405 -5572
rect 10439 -5748 10451 -5572
rect 10393 -5760 10451 -5748
rect 10511 -5572 10569 -5560
rect 10511 -5748 10523 -5572
rect 10557 -5748 10569 -5572
rect 10511 -5760 10569 -5748
rect 11345 -5078 11403 -5066
rect 11345 -5454 11357 -5078
rect 11391 -5454 11403 -5078
rect 11345 -5466 11403 -5454
rect 11463 -5078 11521 -5066
rect 11463 -5454 11475 -5078
rect 11509 -5454 11521 -5078
rect 11463 -5466 11521 -5454
rect 11581 -5078 11639 -5066
rect 11581 -5454 11593 -5078
rect 11627 -5454 11639 -5078
rect 11581 -5466 11639 -5454
rect 11699 -5078 11757 -5066
rect 11699 -5454 11711 -5078
rect 11745 -5454 11757 -5078
rect 11699 -5466 11757 -5454
rect 11817 -5078 11875 -5066
rect 11817 -5454 11829 -5078
rect 11863 -5454 11875 -5078
rect 11817 -5466 11875 -5454
rect 11935 -5078 11993 -5066
rect 11935 -5454 11947 -5078
rect 11981 -5454 11993 -5078
rect 11935 -5466 11993 -5454
rect 12053 -5078 12111 -5066
rect 12053 -5454 12065 -5078
rect 12099 -5454 12111 -5078
rect 12053 -5466 12111 -5454
rect 17573 -4584 17631 -4572
rect 17573 -4760 17585 -4584
rect 17619 -4760 17631 -4584
rect 17573 -4772 17631 -4760
rect 17691 -4584 17749 -4572
rect 17691 -4760 17703 -4584
rect 17737 -4760 17749 -4584
rect 17691 -4772 17749 -4760
rect 17809 -4584 17867 -4572
rect 17809 -4760 17821 -4584
rect 17855 -4760 17867 -4584
rect 17809 -4772 17867 -4760
rect 17927 -4584 17985 -4572
rect 17927 -4760 17939 -4584
rect 17973 -4760 17985 -4584
rect 17927 -4772 17985 -4760
rect 18057 -4760 18069 -4384
rect 18103 -4760 18115 -4384
rect 18057 -4772 18115 -4760
rect 18175 -4384 18233 -4372
rect 18175 -4760 18187 -4384
rect 18221 -4760 18233 -4384
rect 18175 -4772 18233 -4760
rect 18293 -4384 18351 -4372
rect 18293 -4760 18305 -4384
rect 18339 -4760 18351 -4384
rect 18293 -4772 18351 -4760
rect 18411 -4384 18469 -4372
rect 18411 -4760 18423 -4384
rect 18457 -4760 18469 -4384
rect 18411 -4772 18469 -4760
rect 18529 -4384 18587 -4372
rect 18529 -4760 18541 -4384
rect 18575 -4760 18587 -4384
rect 18529 -4772 18587 -4760
rect 18647 -4384 18705 -4372
rect 18647 -4760 18659 -4384
rect 18693 -4760 18705 -4384
rect 18647 -4772 18705 -4760
rect 18765 -4384 18823 -4372
rect 18765 -4760 18777 -4384
rect 18811 -4760 18823 -4384
rect 19955 -4384 20013 -4372
rect 18765 -4772 18823 -4760
rect 18894 -4584 18952 -4572
rect 18894 -4760 18906 -4584
rect 18940 -4760 18952 -4584
rect 18894 -4772 18952 -4760
rect 19012 -4584 19070 -4572
rect 19012 -4760 19024 -4584
rect 19058 -4760 19070 -4584
rect 19012 -4772 19070 -4760
rect 19130 -4584 19188 -4572
rect 19130 -4760 19142 -4584
rect 19176 -4760 19188 -4584
rect 19130 -4772 19188 -4760
rect 19248 -4584 19306 -4572
rect 19248 -4760 19260 -4584
rect 19294 -4760 19306 -4584
rect 19248 -4772 19306 -4760
rect 19471 -4584 19529 -4572
rect 19471 -4760 19483 -4584
rect 19517 -4760 19529 -4584
rect 19471 -4772 19529 -4760
rect 19589 -4584 19647 -4572
rect 19589 -4760 19601 -4584
rect 19635 -4760 19647 -4584
rect 19589 -4772 19647 -4760
rect 19707 -4584 19765 -4572
rect 19707 -4760 19719 -4584
rect 19753 -4760 19765 -4584
rect 19707 -4772 19765 -4760
rect 19825 -4584 19883 -4572
rect 19825 -4760 19837 -4584
rect 19871 -4760 19883 -4584
rect 19825 -4772 19883 -4760
rect 19955 -4760 19967 -4384
rect 20001 -4760 20013 -4384
rect 19955 -4772 20013 -4760
rect 20073 -4384 20131 -4372
rect 20073 -4760 20085 -4384
rect 20119 -4760 20131 -4384
rect 20073 -4772 20131 -4760
rect 20191 -4384 20249 -4372
rect 20191 -4760 20203 -4384
rect 20237 -4760 20249 -4384
rect 20191 -4772 20249 -4760
rect 20309 -4384 20367 -4372
rect 20309 -4760 20321 -4384
rect 20355 -4760 20367 -4384
rect 20309 -4772 20367 -4760
rect 20427 -4384 20485 -4372
rect 20427 -4760 20439 -4384
rect 20473 -4760 20485 -4384
rect 20427 -4772 20485 -4760
rect 20545 -4384 20603 -4372
rect 20545 -4760 20557 -4384
rect 20591 -4760 20603 -4384
rect 20545 -4772 20603 -4760
rect 20663 -4384 20721 -4372
rect 20663 -4760 20675 -4384
rect 20709 -4760 20721 -4384
rect 24679 -4383 24737 -4371
rect 20663 -4772 20721 -4760
rect 20792 -4584 20850 -4572
rect 20792 -4760 20804 -4584
rect 20838 -4760 20850 -4584
rect 20792 -4772 20850 -4760
rect 20910 -4584 20968 -4572
rect 20910 -4760 20922 -4584
rect 20956 -4760 20968 -4584
rect 20910 -4772 20968 -4760
rect 21028 -4584 21086 -4572
rect 21028 -4760 21040 -4584
rect 21074 -4760 21086 -4584
rect 21028 -4772 21086 -4760
rect 21146 -4584 21204 -4572
rect 21146 -4760 21158 -4584
rect 21192 -4760 21204 -4584
rect 21146 -4772 21204 -4760
rect 13243 -5078 13301 -5066
rect 13243 -5454 13255 -5078
rect 13289 -5454 13301 -5078
rect 13243 -5466 13301 -5454
rect 13361 -5078 13419 -5066
rect 13361 -5454 13373 -5078
rect 13407 -5454 13419 -5078
rect 13361 -5466 13419 -5454
rect 13479 -5078 13537 -5066
rect 13479 -5454 13491 -5078
rect 13525 -5454 13537 -5078
rect 13479 -5466 13537 -5454
rect 13597 -5078 13655 -5066
rect 13597 -5454 13609 -5078
rect 13643 -5454 13655 -5078
rect 13597 -5466 13655 -5454
rect 13715 -5078 13773 -5066
rect 13715 -5454 13727 -5078
rect 13761 -5454 13773 -5078
rect 13715 -5466 13773 -5454
rect 13833 -5078 13891 -5066
rect 13833 -5454 13845 -5078
rect 13879 -5454 13891 -5078
rect 13833 -5466 13891 -5454
rect 13951 -5078 14009 -5066
rect 13951 -5454 13963 -5078
rect 13997 -5454 14009 -5078
rect 13951 -5466 14009 -5454
rect 16104 -5571 16162 -5559
rect 16104 -5747 16116 -5571
rect 16150 -5747 16162 -5571
rect 16104 -5759 16162 -5747
rect 16222 -5571 16280 -5559
rect 16222 -5747 16234 -5571
rect 16268 -5747 16280 -5571
rect 16222 -5759 16280 -5747
rect 16340 -5571 16398 -5559
rect 16340 -5747 16352 -5571
rect 16386 -5747 16398 -5571
rect 16340 -5759 16398 -5747
rect 16458 -5571 16516 -5559
rect 16458 -5747 16470 -5571
rect 16504 -5747 16516 -5571
rect 16458 -5759 16516 -5747
rect 16576 -5571 16634 -5559
rect 16576 -5747 16588 -5571
rect 16622 -5747 16634 -5571
rect 16576 -5759 16634 -5747
rect 16694 -5571 16752 -5559
rect 16694 -5747 16706 -5571
rect 16740 -5747 16752 -5571
rect 16694 -5759 16752 -5747
rect 16812 -5571 16870 -5559
rect 16812 -5747 16824 -5571
rect 16858 -5747 16870 -5571
rect 16812 -5759 16870 -5747
rect 16930 -5571 16988 -5559
rect 16930 -5747 16942 -5571
rect 16976 -5747 16988 -5571
rect 16930 -5759 16988 -5747
rect 17048 -5571 17106 -5559
rect 17048 -5747 17060 -5571
rect 17094 -5747 17106 -5571
rect 17048 -5759 17106 -5747
rect 17166 -5571 17224 -5559
rect 17166 -5747 17178 -5571
rect 17212 -5747 17224 -5571
rect 17166 -5759 17224 -5747
rect 18000 -5077 18058 -5065
rect 18000 -5453 18012 -5077
rect 18046 -5453 18058 -5077
rect 18000 -5465 18058 -5453
rect 18118 -5077 18176 -5065
rect 18118 -5453 18130 -5077
rect 18164 -5453 18176 -5077
rect 18118 -5465 18176 -5453
rect 18236 -5077 18294 -5065
rect 18236 -5453 18248 -5077
rect 18282 -5453 18294 -5077
rect 18236 -5465 18294 -5453
rect 18354 -5077 18412 -5065
rect 18354 -5453 18366 -5077
rect 18400 -5453 18412 -5077
rect 18354 -5465 18412 -5453
rect 18472 -5077 18530 -5065
rect 18472 -5453 18484 -5077
rect 18518 -5453 18530 -5077
rect 18472 -5465 18530 -5453
rect 18590 -5077 18648 -5065
rect 18590 -5453 18602 -5077
rect 18636 -5453 18648 -5077
rect 18590 -5465 18648 -5453
rect 18708 -5077 18766 -5065
rect 18708 -5453 18720 -5077
rect 18754 -5453 18766 -5077
rect 18708 -5465 18766 -5453
rect 24195 -4583 24253 -4571
rect 24195 -4759 24207 -4583
rect 24241 -4759 24253 -4583
rect 24195 -4771 24253 -4759
rect 24313 -4583 24371 -4571
rect 24313 -4759 24325 -4583
rect 24359 -4759 24371 -4583
rect 24313 -4771 24371 -4759
rect 24431 -4583 24489 -4571
rect 24431 -4759 24443 -4583
rect 24477 -4759 24489 -4583
rect 24431 -4771 24489 -4759
rect 24549 -4583 24607 -4571
rect 24549 -4759 24561 -4583
rect 24595 -4759 24607 -4583
rect 24549 -4771 24607 -4759
rect 24679 -4759 24691 -4383
rect 24725 -4759 24737 -4383
rect 24679 -4771 24737 -4759
rect 24797 -4383 24855 -4371
rect 24797 -4759 24809 -4383
rect 24843 -4759 24855 -4383
rect 24797 -4771 24855 -4759
rect 24915 -4383 24973 -4371
rect 24915 -4759 24927 -4383
rect 24961 -4759 24973 -4383
rect 24915 -4771 24973 -4759
rect 25033 -4383 25091 -4371
rect 25033 -4759 25045 -4383
rect 25079 -4759 25091 -4383
rect 25033 -4771 25091 -4759
rect 25151 -4383 25209 -4371
rect 25151 -4759 25163 -4383
rect 25197 -4759 25209 -4383
rect 25151 -4771 25209 -4759
rect 25269 -4383 25327 -4371
rect 25269 -4759 25281 -4383
rect 25315 -4759 25327 -4383
rect 25269 -4771 25327 -4759
rect 25387 -4383 25445 -4371
rect 25387 -4759 25399 -4383
rect 25433 -4759 25445 -4383
rect 26577 -4383 26635 -4371
rect 25387 -4771 25445 -4759
rect 25516 -4583 25574 -4571
rect 25516 -4759 25528 -4583
rect 25562 -4759 25574 -4583
rect 25516 -4771 25574 -4759
rect 25634 -4583 25692 -4571
rect 25634 -4759 25646 -4583
rect 25680 -4759 25692 -4583
rect 25634 -4771 25692 -4759
rect 25752 -4583 25810 -4571
rect 25752 -4759 25764 -4583
rect 25798 -4759 25810 -4583
rect 25752 -4771 25810 -4759
rect 25870 -4583 25928 -4571
rect 25870 -4759 25882 -4583
rect 25916 -4759 25928 -4583
rect 25870 -4771 25928 -4759
rect 26093 -4583 26151 -4571
rect 26093 -4759 26105 -4583
rect 26139 -4759 26151 -4583
rect 26093 -4771 26151 -4759
rect 26211 -4583 26269 -4571
rect 26211 -4759 26223 -4583
rect 26257 -4759 26269 -4583
rect 26211 -4771 26269 -4759
rect 26329 -4583 26387 -4571
rect 26329 -4759 26341 -4583
rect 26375 -4759 26387 -4583
rect 26329 -4771 26387 -4759
rect 26447 -4583 26505 -4571
rect 26447 -4759 26459 -4583
rect 26493 -4759 26505 -4583
rect 26447 -4771 26505 -4759
rect 26577 -4759 26589 -4383
rect 26623 -4759 26635 -4383
rect 26577 -4771 26635 -4759
rect 26695 -4383 26753 -4371
rect 26695 -4759 26707 -4383
rect 26741 -4759 26753 -4383
rect 26695 -4771 26753 -4759
rect 26813 -4383 26871 -4371
rect 26813 -4759 26825 -4383
rect 26859 -4759 26871 -4383
rect 26813 -4771 26871 -4759
rect 26931 -4383 26989 -4371
rect 26931 -4759 26943 -4383
rect 26977 -4759 26989 -4383
rect 26931 -4771 26989 -4759
rect 27049 -4383 27107 -4371
rect 27049 -4759 27061 -4383
rect 27095 -4759 27107 -4383
rect 27049 -4771 27107 -4759
rect 27167 -4383 27225 -4371
rect 27167 -4759 27179 -4383
rect 27213 -4759 27225 -4383
rect 27167 -4771 27225 -4759
rect 27285 -4383 27343 -4371
rect 27285 -4759 27297 -4383
rect 27331 -4759 27343 -4383
rect 27285 -4771 27343 -4759
rect 27414 -4583 27472 -4571
rect 27414 -4759 27426 -4583
rect 27460 -4759 27472 -4583
rect 27414 -4771 27472 -4759
rect 27532 -4583 27590 -4571
rect 27532 -4759 27544 -4583
rect 27578 -4759 27590 -4583
rect 27532 -4771 27590 -4759
rect 27650 -4583 27708 -4571
rect 27650 -4759 27662 -4583
rect 27696 -4759 27708 -4583
rect 27650 -4771 27708 -4759
rect 27768 -4583 27826 -4571
rect 27768 -4759 27780 -4583
rect 27814 -4759 27826 -4583
rect 27768 -4771 27826 -4759
rect 19898 -5077 19956 -5065
rect 19898 -5453 19910 -5077
rect 19944 -5453 19956 -5077
rect 19898 -5465 19956 -5453
rect 20016 -5077 20074 -5065
rect 20016 -5453 20028 -5077
rect 20062 -5453 20074 -5077
rect 20016 -5465 20074 -5453
rect 20134 -5077 20192 -5065
rect 20134 -5453 20146 -5077
rect 20180 -5453 20192 -5077
rect 20134 -5465 20192 -5453
rect 20252 -5077 20310 -5065
rect 20252 -5453 20264 -5077
rect 20298 -5453 20310 -5077
rect 20252 -5465 20310 -5453
rect 20370 -5077 20428 -5065
rect 20370 -5453 20382 -5077
rect 20416 -5453 20428 -5077
rect 20370 -5465 20428 -5453
rect 20488 -5077 20546 -5065
rect 20488 -5453 20500 -5077
rect 20534 -5453 20546 -5077
rect 20488 -5465 20546 -5453
rect 20606 -5077 20664 -5065
rect 20606 -5453 20618 -5077
rect 20652 -5453 20664 -5077
rect 20606 -5465 20664 -5453
rect 22726 -5570 22784 -5558
rect 22726 -5746 22738 -5570
rect 22772 -5746 22784 -5570
rect 22726 -5758 22784 -5746
rect 22844 -5570 22902 -5558
rect 22844 -5746 22856 -5570
rect 22890 -5746 22902 -5570
rect 22844 -5758 22902 -5746
rect 22962 -5570 23020 -5558
rect 22962 -5746 22974 -5570
rect 23008 -5746 23020 -5570
rect 22962 -5758 23020 -5746
rect 23080 -5570 23138 -5558
rect 23080 -5746 23092 -5570
rect 23126 -5746 23138 -5570
rect 23080 -5758 23138 -5746
rect 23198 -5570 23256 -5558
rect 23198 -5746 23210 -5570
rect 23244 -5746 23256 -5570
rect 23198 -5758 23256 -5746
rect 23316 -5570 23374 -5558
rect 23316 -5746 23328 -5570
rect 23362 -5746 23374 -5570
rect 23316 -5758 23374 -5746
rect 23434 -5570 23492 -5558
rect 23434 -5746 23446 -5570
rect 23480 -5746 23492 -5570
rect 23434 -5758 23492 -5746
rect 23552 -5570 23610 -5558
rect 23552 -5746 23564 -5570
rect 23598 -5746 23610 -5570
rect 23552 -5758 23610 -5746
rect 23670 -5570 23728 -5558
rect 23670 -5746 23682 -5570
rect 23716 -5746 23728 -5570
rect 23670 -5758 23728 -5746
rect 23788 -5570 23846 -5558
rect 23788 -5746 23800 -5570
rect 23834 -5746 23846 -5570
rect 23788 -5758 23846 -5746
rect 24622 -5076 24680 -5064
rect 24622 -5452 24634 -5076
rect 24668 -5452 24680 -5076
rect 24622 -5464 24680 -5452
rect 24740 -5076 24798 -5064
rect 24740 -5452 24752 -5076
rect 24786 -5452 24798 -5076
rect 24740 -5464 24798 -5452
rect 24858 -5076 24916 -5064
rect 24858 -5452 24870 -5076
rect 24904 -5452 24916 -5076
rect 24858 -5464 24916 -5452
rect 24976 -5076 25034 -5064
rect 24976 -5452 24988 -5076
rect 25022 -5452 25034 -5076
rect 24976 -5464 25034 -5452
rect 25094 -5076 25152 -5064
rect 25094 -5452 25106 -5076
rect 25140 -5452 25152 -5076
rect 25094 -5464 25152 -5452
rect 25212 -5076 25270 -5064
rect 25212 -5452 25224 -5076
rect 25258 -5452 25270 -5076
rect 25212 -5464 25270 -5452
rect 25330 -5076 25388 -5064
rect 25330 -5452 25342 -5076
rect 25376 -5452 25388 -5076
rect 25330 -5464 25388 -5452
rect 26520 -5076 26578 -5064
rect 26520 -5452 26532 -5076
rect 26566 -5452 26578 -5076
rect 26520 -5464 26578 -5452
rect 26638 -5076 26696 -5064
rect 26638 -5452 26650 -5076
rect 26684 -5452 26696 -5076
rect 26638 -5464 26696 -5452
rect 26756 -5076 26814 -5064
rect 26756 -5452 26768 -5076
rect 26802 -5452 26814 -5076
rect 26756 -5464 26814 -5452
rect 26874 -5076 26932 -5064
rect 26874 -5452 26886 -5076
rect 26920 -5452 26932 -5076
rect 26874 -5464 26932 -5452
rect 26992 -5076 27050 -5064
rect 26992 -5452 27004 -5076
rect 27038 -5452 27050 -5076
rect 26992 -5464 27050 -5452
rect 27110 -5076 27168 -5064
rect 27110 -5452 27122 -5076
rect 27156 -5452 27168 -5076
rect 27110 -5464 27168 -5452
rect 27228 -5076 27286 -5064
rect 27228 -5452 27240 -5076
rect 27274 -5452 27286 -5076
rect 27228 -5464 27286 -5452
rect 28590 -5110 28648 -5098
rect 28590 -5286 28602 -5110
rect 28636 -5286 28648 -5110
rect 28590 -5298 28648 -5286
rect 28708 -5110 28766 -5098
rect 28708 -5286 28720 -5110
rect 28754 -5286 28766 -5110
rect 28708 -5298 28766 -5286
rect 28826 -5110 28884 -5098
rect 28826 -5286 28838 -5110
rect 28872 -5286 28884 -5110
rect 28826 -5298 28884 -5286
rect 28944 -5110 29002 -5098
rect 28944 -5286 28956 -5110
rect 28990 -5286 29002 -5110
rect 28944 -5298 29002 -5286
rect 29062 -5110 29120 -5098
rect 29062 -5286 29074 -5110
rect 29108 -5286 29120 -5110
rect 29062 -5298 29120 -5286
rect 29180 -5110 29238 -5098
rect 29180 -5286 29192 -5110
rect 29226 -5286 29238 -5110
rect 29180 -5298 29238 -5286
rect 29298 -5110 29356 -5098
rect 29298 -5286 29310 -5110
rect 29344 -5286 29356 -5110
rect 29298 -5298 29356 -5286
rect 29416 -5110 29474 -5098
rect 29416 -5286 29428 -5110
rect 29462 -5286 29474 -5110
rect 29416 -5298 29474 -5286
rect 29534 -5110 29592 -5098
rect 29534 -5286 29546 -5110
rect 29580 -5286 29592 -5110
rect 29534 -5298 29592 -5286
rect 29652 -5110 29710 -5098
rect 29652 -5286 29664 -5110
rect 29698 -5286 29710 -5110
rect 29652 -5298 29710 -5286
rect 30821 -6655 30879 -6643
rect 30337 -6855 30395 -6843
rect 30337 -7031 30349 -6855
rect 30383 -7031 30395 -6855
rect 30337 -7043 30395 -7031
rect 30455 -6855 30513 -6843
rect 30455 -7031 30467 -6855
rect 30501 -7031 30513 -6855
rect 30455 -7043 30513 -7031
rect 30573 -6855 30631 -6843
rect 30573 -7031 30585 -6855
rect 30619 -7031 30631 -6855
rect 30573 -7043 30631 -7031
rect 30691 -6855 30749 -6843
rect 30691 -7031 30703 -6855
rect 30737 -7031 30749 -6855
rect 30691 -7043 30749 -7031
rect 30821 -7031 30833 -6655
rect 30867 -7031 30879 -6655
rect 30821 -7043 30879 -7031
rect 30939 -6655 30997 -6643
rect 30939 -7031 30951 -6655
rect 30985 -7031 30997 -6655
rect 30939 -7043 30997 -7031
rect 31057 -6655 31115 -6643
rect 31057 -7031 31069 -6655
rect 31103 -7031 31115 -6655
rect 31057 -7043 31115 -7031
rect 31175 -6655 31233 -6643
rect 31175 -7031 31187 -6655
rect 31221 -7031 31233 -6655
rect 31175 -7043 31233 -7031
rect 31293 -6655 31351 -6643
rect 31293 -7031 31305 -6655
rect 31339 -7031 31351 -6655
rect 31293 -7043 31351 -7031
rect 31411 -6655 31469 -6643
rect 31411 -7031 31423 -6655
rect 31457 -7031 31469 -6655
rect 31411 -7043 31469 -7031
rect 31529 -6655 31587 -6643
rect 31529 -7031 31541 -6655
rect 31575 -7031 31587 -6655
rect 31529 -7043 31587 -7031
rect 31658 -6855 31716 -6843
rect 31658 -7031 31670 -6855
rect 31704 -7031 31716 -6855
rect 31658 -7043 31716 -7031
rect 31776 -6855 31834 -6843
rect 31776 -7031 31788 -6855
rect 31822 -7031 31834 -6855
rect 31776 -7043 31834 -7031
rect 31894 -6855 31952 -6843
rect 31894 -7031 31906 -6855
rect 31940 -7031 31952 -6855
rect 31894 -7043 31952 -7031
rect 32012 -6855 32070 -6843
rect 32012 -7031 32024 -6855
rect 32058 -7031 32070 -6855
rect 32012 -7043 32070 -7031
rect 32130 -6858 32188 -6846
rect 32130 -7034 32142 -6858
rect 32176 -7034 32188 -6858
rect 32130 -7046 32188 -7034
rect 32248 -6858 32306 -6846
rect 32248 -7034 32260 -6858
rect 32294 -7034 32306 -6858
rect 32248 -7046 32306 -7034
rect 32366 -6858 32424 -6846
rect 32366 -7034 32378 -6858
rect 32412 -7034 32424 -6858
rect 32366 -7046 32424 -7034
rect 32484 -6858 32542 -6846
rect 32484 -7034 32496 -6858
rect 32530 -7034 32542 -6858
rect 32484 -7046 32542 -7034
rect 32602 -6858 32660 -6846
rect 32602 -7034 32614 -6858
rect 32648 -7034 32660 -6858
rect 32602 -7046 32660 -7034
rect 32720 -6858 32778 -6846
rect 32720 -7034 32732 -6858
rect 32766 -7034 32778 -6858
rect 32720 -7046 32778 -7034
rect 32838 -6858 32896 -6846
rect 32838 -7034 32850 -6858
rect 32884 -7034 32896 -6858
rect 32838 -7046 32896 -7034
rect 32956 -6858 33014 -6846
rect 32956 -7034 32968 -6858
rect 33002 -7034 33014 -6858
rect 32956 -7046 33014 -7034
rect 33074 -6858 33132 -6846
rect 33074 -7034 33086 -6858
rect 33120 -7034 33132 -6858
rect 33074 -7046 33132 -7034
rect 33192 -6858 33250 -6846
rect 33192 -7034 33204 -6858
rect 33238 -7034 33250 -6858
rect 33192 -7046 33250 -7034
rect 30764 -7348 30822 -7336
rect 28597 -7955 28655 -7943
rect 6706 -8073 6764 -8061
rect 6706 -8249 6718 -8073
rect 6752 -8249 6764 -8073
rect 6706 -8261 6764 -8249
rect 6824 -8073 6882 -8061
rect 6824 -8249 6836 -8073
rect 6870 -8249 6882 -8073
rect 6824 -8261 6882 -8249
rect 6942 -8073 7000 -8061
rect 6942 -8249 6954 -8073
rect 6988 -8249 7000 -8073
rect 6942 -8261 7000 -8249
rect 7060 -8073 7118 -8061
rect 7060 -8249 7072 -8073
rect 7106 -8249 7118 -8073
rect 7060 -8261 7118 -8249
rect 7178 -8073 7236 -8061
rect 7178 -8249 7190 -8073
rect 7224 -8249 7236 -8073
rect 7178 -8261 7236 -8249
rect 7296 -8073 7354 -8061
rect 7296 -8249 7308 -8073
rect 7342 -8249 7354 -8073
rect 7296 -8261 7354 -8249
rect 7414 -8073 7472 -8061
rect 7414 -8249 7426 -8073
rect 7460 -8249 7472 -8073
rect 7414 -8261 7472 -8249
rect 7532 -8073 7590 -8061
rect 7532 -8249 7544 -8073
rect 7578 -8249 7590 -8073
rect 7532 -8261 7590 -8249
rect 7650 -8073 7708 -8061
rect 7650 -8249 7662 -8073
rect 7696 -8249 7708 -8073
rect 7650 -8261 7708 -8249
rect 7768 -8073 7826 -8061
rect 7768 -8249 7780 -8073
rect 7814 -8249 7826 -8073
rect 7768 -8261 7826 -8249
rect 13260 -8068 13318 -8056
rect 13260 -8244 13272 -8068
rect 13306 -8244 13318 -8068
rect 13260 -8256 13318 -8244
rect 13378 -8068 13436 -8056
rect 13378 -8244 13390 -8068
rect 13424 -8244 13436 -8068
rect 13378 -8256 13436 -8244
rect 13496 -8068 13554 -8056
rect 13496 -8244 13508 -8068
rect 13542 -8244 13554 -8068
rect 13496 -8256 13554 -8244
rect 13614 -8068 13672 -8056
rect 13614 -8244 13626 -8068
rect 13660 -8244 13672 -8068
rect 13614 -8256 13672 -8244
rect 13732 -8068 13790 -8056
rect 13732 -8244 13744 -8068
rect 13778 -8244 13790 -8068
rect 13732 -8256 13790 -8244
rect 13850 -8068 13908 -8056
rect 13850 -8244 13862 -8068
rect 13896 -8244 13908 -8068
rect 13850 -8256 13908 -8244
rect 13968 -8068 14026 -8056
rect 13968 -8244 13980 -8068
rect 14014 -8244 14026 -8068
rect 13968 -8256 14026 -8244
rect 14086 -8068 14144 -8056
rect 14086 -8244 14098 -8068
rect 14132 -8244 14144 -8068
rect 14086 -8256 14144 -8244
rect 14204 -8068 14262 -8056
rect 14204 -8244 14216 -8068
rect 14250 -8244 14262 -8068
rect 14204 -8256 14262 -8244
rect 14322 -8068 14380 -8056
rect 14322 -8244 14334 -8068
rect 14368 -8244 14380 -8068
rect 14322 -8256 14380 -8244
rect 19909 -8080 19967 -8068
rect 19909 -8256 19921 -8080
rect 19955 -8256 19967 -8080
rect 19909 -8268 19967 -8256
rect 20027 -8080 20085 -8068
rect 20027 -8256 20039 -8080
rect 20073 -8256 20085 -8080
rect 20027 -8268 20085 -8256
rect 20145 -8080 20203 -8068
rect 20145 -8256 20157 -8080
rect 20191 -8256 20203 -8080
rect 20145 -8268 20203 -8256
rect 20263 -8080 20321 -8068
rect 20263 -8256 20275 -8080
rect 20309 -8256 20321 -8080
rect 20263 -8268 20321 -8256
rect 20381 -8080 20439 -8068
rect 20381 -8256 20393 -8080
rect 20427 -8256 20439 -8080
rect 20381 -8268 20439 -8256
rect 20499 -8080 20557 -8068
rect 20499 -8256 20511 -8080
rect 20545 -8256 20557 -8080
rect 20499 -8268 20557 -8256
rect 20617 -8080 20675 -8068
rect 20617 -8256 20629 -8080
rect 20663 -8256 20675 -8080
rect 20617 -8268 20675 -8256
rect 20735 -8080 20793 -8068
rect 20735 -8256 20747 -8080
rect 20781 -8256 20793 -8080
rect 20735 -8268 20793 -8256
rect 20853 -8080 20911 -8068
rect 20853 -8256 20865 -8080
rect 20899 -8256 20911 -8080
rect 20853 -8268 20911 -8256
rect 20971 -8080 21029 -8068
rect 20971 -8256 20983 -8080
rect 21017 -8256 21029 -8080
rect 28597 -8131 28609 -7955
rect 28643 -8131 28655 -7955
rect 28597 -8143 28655 -8131
rect 28715 -7955 28773 -7943
rect 28715 -8131 28727 -7955
rect 28761 -8131 28773 -7955
rect 28715 -8143 28773 -8131
rect 28833 -7955 28891 -7943
rect 28833 -8131 28845 -7955
rect 28879 -8131 28891 -7955
rect 28833 -8143 28891 -8131
rect 28951 -7955 29009 -7943
rect 28951 -8131 28963 -7955
rect 28997 -8131 29009 -7955
rect 28951 -8143 29009 -8131
rect 29069 -7955 29127 -7943
rect 29069 -8131 29081 -7955
rect 29115 -8131 29127 -7955
rect 29069 -8143 29127 -8131
rect 29187 -7955 29245 -7943
rect 29187 -8131 29199 -7955
rect 29233 -8131 29245 -7955
rect 29187 -8143 29245 -8131
rect 29305 -7955 29363 -7943
rect 29305 -8131 29317 -7955
rect 29351 -8131 29363 -7955
rect 29305 -8143 29363 -8131
rect 29423 -7955 29481 -7943
rect 29423 -8131 29435 -7955
rect 29469 -8131 29481 -7955
rect 29423 -8143 29481 -8131
rect 29541 -7955 29599 -7943
rect 29541 -8131 29553 -7955
rect 29587 -8131 29599 -7955
rect 29541 -8143 29599 -8131
rect 29659 -7955 29717 -7943
rect 29659 -8131 29671 -7955
rect 29705 -8131 29717 -7955
rect 30764 -7724 30776 -7348
rect 30810 -7724 30822 -7348
rect 30764 -7736 30822 -7724
rect 30882 -7348 30940 -7336
rect 30882 -7724 30894 -7348
rect 30928 -7724 30940 -7348
rect 30882 -7736 30940 -7724
rect 31000 -7348 31058 -7336
rect 31000 -7724 31012 -7348
rect 31046 -7724 31058 -7348
rect 31000 -7736 31058 -7724
rect 31118 -7348 31176 -7336
rect 31118 -7724 31130 -7348
rect 31164 -7724 31176 -7348
rect 31118 -7736 31176 -7724
rect 31236 -7348 31294 -7336
rect 31236 -7724 31248 -7348
rect 31282 -7724 31294 -7348
rect 31236 -7736 31294 -7724
rect 31354 -7348 31412 -7336
rect 31354 -7724 31366 -7348
rect 31400 -7724 31412 -7348
rect 31354 -7736 31412 -7724
rect 31472 -7348 31530 -7336
rect 31472 -7724 31484 -7348
rect 31518 -7724 31530 -7348
rect 31472 -7736 31530 -7724
rect 29659 -8143 29717 -8131
rect 20971 -8268 21029 -8256
<< ndiffc >>
rect 6920 4818 6954 5194
rect 7038 4818 7072 5194
rect 7156 4818 7190 5194
rect 7273 5018 7307 5194
rect 7391 5018 7425 5194
rect 13469 4817 13503 5193
rect 13587 4817 13621 5193
rect 13705 4817 13739 5193
rect 13822 5017 13856 5193
rect 13940 5017 13974 5193
rect 20123 4838 20157 5214
rect 20241 4838 20275 5214
rect 20359 4838 20393 5214
rect 20476 5038 20510 5214
rect 20594 5038 20628 5214
rect 28776 4671 28810 5047
rect 28894 4671 28928 5047
rect 29012 4671 29046 5047
rect 29129 4871 29163 5047
rect 29247 4871 29281 5047
rect 32377 4263 32411 4639
rect 32495 4263 32529 4639
rect 32613 4263 32647 4639
rect 32730 4463 32764 4639
rect 32848 4463 32882 4639
rect 256 2918 290 3294
rect 374 2918 408 3294
rect 492 2918 526 3294
rect 609 3118 643 3294
rect 727 3118 761 3294
rect 3146 2651 3180 3027
rect 3264 2651 3298 3027
rect 3382 2651 3416 3027
rect 3499 2851 3533 3027
rect 3617 2851 3651 3027
rect 30472 3678 30506 3854
rect 30590 3678 30624 3854
rect 5144 2577 5178 2753
rect 5262 2577 5296 2753
rect 5380 2577 5414 2753
rect 5498 2577 5532 2753
rect 6286 2581 6320 2757
rect 6404 2581 6438 2757
rect 6522 2581 6556 2757
rect 6640 2581 6674 2757
rect 9695 2739 9729 3115
rect 9813 2739 9847 3115
rect 9931 2739 9965 3115
rect 10048 2939 10082 3115
rect 10166 2939 10200 3115
rect 11693 2665 11727 2841
rect 11811 2665 11845 2841
rect 11929 2665 11963 2841
rect 12047 2665 12081 2841
rect 12835 2669 12869 2845
rect 12953 2669 12987 2845
rect 13071 2669 13105 2845
rect 13189 2669 13223 2845
rect 16349 2671 16383 3047
rect 16467 2671 16501 3047
rect 16585 2671 16619 3047
rect 16702 2871 16736 3047
rect 16820 2871 16854 3047
rect 30892 3478 30926 3854
rect 31010 3478 31044 3854
rect 31128 3478 31162 3854
rect 31246 3478 31280 3854
rect 31364 3478 31398 3854
rect 31770 3678 31804 3854
rect 31888 3678 31922 3854
rect 18347 2597 18381 2773
rect 18465 2597 18499 2773
rect 18583 2597 18617 2773
rect 18701 2597 18735 2773
rect 19489 2601 19523 2777
rect 19607 2601 19641 2777
rect 19725 2601 19759 2777
rect 19843 2601 19877 2777
rect 22974 2739 23008 3115
rect 23092 2739 23126 3115
rect 23210 2739 23244 3115
rect 23327 2939 23361 3115
rect 23445 2939 23479 3115
rect 24972 2665 25006 2841
rect 25090 2665 25124 2841
rect 25208 2665 25242 2841
rect 25326 2665 25360 2841
rect 26114 2669 26148 2845
rect 26232 2669 26266 2845
rect 26350 2669 26384 2845
rect 26468 2669 26502 2845
rect 28771 2100 28805 2476
rect 28889 2100 28923 2476
rect 29007 2100 29041 2476
rect 29124 2300 29158 2476
rect 29242 2300 29276 2476
rect 3160 1001 3194 1377
rect 3278 1001 3312 1377
rect 3396 1001 3430 1377
rect 3513 1201 3547 1377
rect 3631 1201 3665 1377
rect 9709 1089 9743 1465
rect 9827 1089 9861 1465
rect 9945 1089 9979 1465
rect 10062 1289 10096 1465
rect 10180 1289 10214 1465
rect 248 333 282 709
rect 366 333 400 709
rect 484 333 518 709
rect 601 533 635 709
rect 719 533 753 709
rect 4512 -204 4546 -28
rect 3155 -603 3189 -227
rect 3273 -603 3307 -227
rect 3391 -603 3425 -227
rect 3508 -403 3542 -227
rect 4630 -204 4664 -28
rect 3626 -403 3660 -227
rect 4932 -404 4966 -28
rect 5050 -404 5084 -28
rect 5168 -404 5202 -28
rect 5286 -404 5320 -28
rect 5404 -404 5438 -28
rect 5810 -204 5844 -28
rect 5928 -204 5962 -28
rect 6410 -204 6444 -28
rect 6528 -204 6562 -28
rect 6830 -404 6864 -28
rect 6948 -404 6982 -28
rect 7066 -404 7100 -28
rect 7184 -404 7218 -28
rect 7302 -404 7336 -28
rect 7708 -204 7742 -28
rect 7826 -204 7860 -28
rect 16363 1021 16397 1397
rect 16481 1021 16515 1397
rect 16599 1021 16633 1397
rect 16716 1221 16750 1397
rect 16834 1221 16868 1397
rect 22988 1089 23022 1465
rect 23106 1089 23140 1465
rect 23224 1089 23258 1465
rect 23341 1289 23375 1465
rect 23459 1289 23493 1465
rect 11061 -116 11095 60
rect 9704 -515 9738 -139
rect 9822 -515 9856 -139
rect 9940 -515 9974 -139
rect 10057 -315 10091 -139
rect 11179 -116 11213 60
rect 10175 -315 10209 -139
rect 11481 -316 11515 60
rect 11599 -316 11633 60
rect 11717 -316 11751 60
rect 11835 -316 11869 60
rect 11953 -316 11987 60
rect 12359 -116 12393 60
rect 12477 -116 12511 60
rect 12959 -116 12993 60
rect 13077 -116 13111 60
rect 13379 -316 13413 60
rect 13497 -316 13531 60
rect 13615 -316 13649 60
rect 13733 -316 13767 60
rect 13851 -316 13885 60
rect 14257 -116 14291 60
rect 14375 -116 14409 60
rect 17715 -184 17749 -8
rect 16358 -583 16392 -207
rect 16476 -583 16510 -207
rect 16594 -583 16628 -207
rect 16711 -383 16745 -207
rect 17833 -184 17867 -8
rect 16829 -383 16863 -207
rect 18135 -384 18169 -8
rect 18253 -384 18287 -8
rect 18371 -384 18405 -8
rect 18489 -384 18523 -8
rect 18607 -384 18641 -8
rect 19013 -184 19047 -8
rect 19131 -184 19165 -8
rect 19613 -184 19647 -8
rect 19731 -184 19765 -8
rect 20033 -384 20067 -8
rect 20151 -384 20185 -8
rect 20269 -384 20303 -8
rect 20387 -384 20421 -8
rect 20505 -384 20539 -8
rect 20911 -184 20945 -8
rect 21029 -184 21063 -8
rect 24340 -116 24374 60
rect 22983 -515 23017 -139
rect 23101 -515 23135 -139
rect 23219 -515 23253 -139
rect 23336 -315 23370 -139
rect 24458 -116 24492 60
rect 23454 -315 23488 -139
rect 24760 -316 24794 60
rect 24878 -316 24912 60
rect 24996 -316 25030 60
rect 25114 -316 25148 60
rect 25232 -316 25266 60
rect 25638 -116 25672 60
rect 25756 -116 25790 60
rect 26238 -116 26272 60
rect 26356 -116 26390 60
rect 26658 -316 26692 60
rect 26776 -316 26810 60
rect 26894 -316 26928 60
rect 27012 -316 27046 60
rect 27130 -316 27164 60
rect 27536 -116 27570 60
rect 27654 -116 27688 60
rect 32379 172 32413 548
rect 32497 172 32531 548
rect 32615 172 32649 548
rect 32732 372 32766 548
rect 32850 372 32884 548
rect 30474 -413 30508 -237
rect 30592 -413 30626 -237
rect 28771 -933 28805 -557
rect 28889 -933 28923 -557
rect 29007 -933 29041 -557
rect 29124 -733 29158 -557
rect 29242 -733 29276 -557
rect 30894 -613 30928 -237
rect 31012 -613 31046 -237
rect 31130 -613 31164 -237
rect 31248 -613 31282 -237
rect 31366 -613 31400 -237
rect 31772 -413 31806 -237
rect 31890 -413 31924 -237
rect 229 -2945 263 -2569
rect 347 -2945 381 -2569
rect 465 -2945 499 -2569
rect 582 -2745 616 -2569
rect 700 -2745 734 -2569
rect 3138 -3129 3172 -2753
rect 3256 -3129 3290 -2753
rect 3374 -3129 3408 -2753
rect 3491 -2929 3525 -2753
rect 3609 -2929 3643 -2753
rect 5136 -3203 5170 -3027
rect 5254 -3203 5288 -3027
rect 5372 -3203 5406 -3027
rect 5490 -3203 5524 -3027
rect 6278 -3199 6312 -3023
rect 6396 -3199 6430 -3023
rect 6514 -3199 6548 -3023
rect 6632 -3199 6666 -3023
rect 9689 -3131 9723 -2755
rect 9807 -3131 9841 -2755
rect 9925 -3131 9959 -2755
rect 10042 -2931 10076 -2755
rect 10160 -2931 10194 -2755
rect 11687 -3205 11721 -3029
rect 11805 -3205 11839 -3029
rect 11923 -3205 11957 -3029
rect 12041 -3205 12075 -3029
rect 12829 -3201 12863 -3025
rect 12947 -3201 12981 -3025
rect 13065 -3201 13099 -3025
rect 13183 -3201 13217 -3025
rect 16344 -3130 16378 -2754
rect 16462 -3130 16496 -2754
rect 16580 -3130 16614 -2754
rect 16697 -2930 16731 -2754
rect 16815 -2930 16849 -2754
rect 18342 -3204 18376 -3028
rect 18460 -3204 18494 -3028
rect 18578 -3204 18612 -3028
rect 18696 -3204 18730 -3028
rect 19484 -3200 19518 -3024
rect 19602 -3200 19636 -3024
rect 19720 -3200 19754 -3024
rect 19838 -3200 19872 -3024
rect 22966 -3129 23000 -2753
rect 23084 -3129 23118 -2753
rect 23202 -3129 23236 -2753
rect 23319 -2929 23353 -2753
rect 23437 -2929 23471 -2753
rect 28842 -2853 28876 -2477
rect 28960 -2853 28994 -2477
rect 29078 -2853 29112 -2477
rect 29195 -2653 29229 -2477
rect 29313 -2653 29347 -2477
rect 24964 -3203 24998 -3027
rect 25082 -3203 25116 -3027
rect 25200 -3203 25234 -3027
rect 25318 -3203 25352 -3027
rect 26106 -3199 26140 -3023
rect 26224 -3199 26258 -3023
rect 26342 -3199 26376 -3023
rect 26460 -3199 26494 -3023
rect 32379 -3323 32413 -2947
rect 32497 -3323 32531 -2947
rect 32615 -3323 32649 -2947
rect 32732 -3123 32766 -2947
rect 32850 -3123 32884 -2947
rect 30474 -3908 30508 -3732
rect 30592 -3908 30626 -3732
rect 30894 -4108 30928 -3732
rect 31012 -4108 31046 -3732
rect 31130 -4108 31164 -3732
rect 31248 -4108 31282 -3732
rect 31366 -4108 31400 -3732
rect 31772 -3908 31806 -3732
rect 31890 -3908 31924 -3732
rect 3152 -4779 3186 -4403
rect 3270 -4779 3304 -4403
rect 3388 -4779 3422 -4403
rect 3505 -4579 3539 -4403
rect 3623 -4579 3657 -4403
rect 245 -5705 279 -5329
rect 363 -5705 397 -5329
rect 481 -5705 515 -5329
rect 598 -5505 632 -5329
rect 716 -5505 750 -5329
rect 9703 -4781 9737 -4405
rect 9821 -4781 9855 -4405
rect 9939 -4781 9973 -4405
rect 10056 -4581 10090 -4405
rect 10174 -4581 10208 -4405
rect 4504 -5984 4538 -5808
rect 3147 -6383 3181 -6007
rect 3265 -6383 3299 -6007
rect 3383 -6383 3417 -6007
rect 3500 -6183 3534 -6007
rect 4622 -5984 4656 -5808
rect 3618 -6183 3652 -6007
rect 4924 -6184 4958 -5808
rect 5042 -6184 5076 -5808
rect 5160 -6184 5194 -5808
rect 5278 -6184 5312 -5808
rect 5396 -6184 5430 -5808
rect 5802 -5984 5836 -5808
rect 5920 -5984 5954 -5808
rect 6402 -5984 6436 -5808
rect 6520 -5984 6554 -5808
rect 6822 -6184 6856 -5808
rect 6940 -6184 6974 -5808
rect 7058 -6184 7092 -5808
rect 7176 -6184 7210 -5808
rect 7294 -6184 7328 -5808
rect 7700 -5984 7734 -5808
rect 7818 -5984 7852 -5808
rect 16358 -4780 16392 -4404
rect 16476 -4780 16510 -4404
rect 16594 -4780 16628 -4404
rect 16711 -4580 16745 -4404
rect 16829 -4580 16863 -4404
rect 11055 -5986 11089 -5810
rect 9698 -6385 9732 -6009
rect 9816 -6385 9850 -6009
rect 9934 -6385 9968 -6009
rect 10051 -6185 10085 -6009
rect 11173 -5986 11207 -5810
rect 10169 -6185 10203 -6009
rect 11475 -6186 11509 -5810
rect 11593 -6186 11627 -5810
rect 11711 -6186 11745 -5810
rect 11829 -6186 11863 -5810
rect 11947 -6186 11981 -5810
rect 12353 -5986 12387 -5810
rect 12471 -5986 12505 -5810
rect 12953 -5986 12987 -5810
rect 13071 -5986 13105 -5810
rect 13373 -6186 13407 -5810
rect 13491 -6186 13525 -5810
rect 13609 -6186 13643 -5810
rect 13727 -6186 13761 -5810
rect 13845 -6186 13879 -5810
rect 14251 -5986 14285 -5810
rect 14369 -5986 14403 -5810
rect 22980 -4779 23014 -4403
rect 23098 -4779 23132 -4403
rect 23216 -4779 23250 -4403
rect 23333 -4579 23367 -4403
rect 23451 -4579 23485 -4403
rect 17710 -5985 17744 -5809
rect 16353 -6384 16387 -6008
rect 16471 -6384 16505 -6008
rect 16589 -6384 16623 -6008
rect 16706 -6184 16740 -6008
rect 17828 -5985 17862 -5809
rect 16824 -6184 16858 -6008
rect 18130 -6185 18164 -5809
rect 18248 -6185 18282 -5809
rect 18366 -6185 18400 -5809
rect 18484 -6185 18518 -5809
rect 18602 -6185 18636 -5809
rect 19008 -5985 19042 -5809
rect 19126 -5985 19160 -5809
rect 19608 -5985 19642 -5809
rect 19726 -5985 19760 -5809
rect 20028 -6185 20062 -5809
rect 20146 -6185 20180 -5809
rect 20264 -6185 20298 -5809
rect 20382 -6185 20416 -5809
rect 20500 -6185 20534 -5809
rect 20906 -5985 20940 -5809
rect 21024 -5985 21058 -5809
rect 24332 -5984 24366 -5808
rect 22975 -6383 23009 -6007
rect 23093 -6383 23127 -6007
rect 23211 -6383 23245 -6007
rect 23328 -6183 23362 -6007
rect 24450 -5984 24484 -5808
rect 23446 -6183 23480 -6007
rect 24752 -6184 24786 -5808
rect 24870 -6184 24904 -5808
rect 24988 -6184 25022 -5808
rect 25106 -6184 25140 -5808
rect 25224 -6184 25258 -5808
rect 25630 -5984 25664 -5808
rect 25748 -5984 25782 -5808
rect 26230 -5984 26264 -5808
rect 26348 -5984 26382 -5808
rect 26650 -6184 26684 -5808
rect 26768 -6184 26802 -5808
rect 26886 -6184 26920 -5808
rect 27004 -6184 27038 -5808
rect 27122 -6184 27156 -5808
rect 27528 -5984 27562 -5808
rect 27646 -5984 27680 -5808
rect 28839 -5923 28873 -5547
rect 28957 -5923 28991 -5547
rect 29075 -5923 29109 -5547
rect 29192 -5723 29226 -5547
rect 29310 -5723 29344 -5547
rect 6955 -7812 6989 -7436
rect 7073 -7812 7107 -7436
rect 7191 -7812 7225 -7436
rect 7308 -7812 7342 -7636
rect 7426 -7812 7460 -7636
rect 13509 -7807 13543 -7431
rect 13627 -7807 13661 -7431
rect 13745 -7807 13779 -7431
rect 13862 -7807 13896 -7631
rect 13980 -7807 14014 -7631
rect 20158 -7819 20192 -7443
rect 20276 -7819 20310 -7443
rect 20394 -7819 20428 -7443
rect 20511 -7819 20545 -7643
rect 20629 -7819 20663 -7643
rect 32379 -7671 32413 -7295
rect 32497 -7671 32531 -7295
rect 32615 -7671 32649 -7295
rect 32732 -7471 32766 -7295
rect 32850 -7471 32884 -7295
rect 30474 -8256 30508 -8080
rect 30592 -8256 30626 -8080
rect 28846 -8768 28880 -8392
rect 28964 -8768 28998 -8392
rect 29082 -8768 29116 -8392
rect 29199 -8568 29233 -8392
rect 29317 -8568 29351 -8392
rect 30894 -8456 30928 -8080
rect 31012 -8456 31046 -8080
rect 31130 -8456 31164 -8080
rect 31248 -8456 31282 -8080
rect 31366 -8456 31400 -8080
rect 31772 -8256 31806 -8080
rect 31890 -8256 31924 -8080
<< pdiffc >>
rect 6683 5455 6717 5631
rect 6801 5455 6835 5631
rect 6919 5455 6953 5631
rect 7037 5455 7071 5631
rect 7155 5455 7189 5631
rect 7273 5455 7307 5631
rect 7391 5455 7425 5631
rect 7509 5455 7543 5631
rect 7627 5455 7661 5631
rect 7745 5455 7779 5631
rect 13232 5454 13266 5630
rect 13350 5454 13384 5630
rect 13468 5454 13502 5630
rect 13586 5454 13620 5630
rect 13704 5454 13738 5630
rect 13822 5454 13856 5630
rect 13940 5454 13974 5630
rect 14058 5454 14092 5630
rect 14176 5454 14210 5630
rect 14294 5454 14328 5630
rect 19886 5475 19920 5651
rect 20004 5475 20038 5651
rect 20122 5475 20156 5651
rect 20240 5475 20274 5651
rect 20358 5475 20392 5651
rect 20476 5475 20510 5651
rect 20594 5475 20628 5651
rect 20712 5475 20746 5651
rect 20830 5475 20864 5651
rect 20948 5475 20982 5651
rect 28539 5308 28573 5484
rect 28657 5308 28691 5484
rect 28775 5308 28809 5484
rect 28893 5308 28927 5484
rect 29011 5308 29045 5484
rect 29129 5308 29163 5484
rect 29247 5308 29281 5484
rect 29365 5308 29399 5484
rect 29483 5308 29517 5484
rect 29601 5308 29635 5484
rect 30347 4903 30381 5079
rect 30465 4903 30499 5079
rect 30583 4903 30617 5079
rect 30701 4903 30735 5079
rect 30831 4903 30865 5279
rect 30949 4903 30983 5279
rect 31067 4903 31101 5279
rect 31185 4903 31219 5279
rect 31303 4903 31337 5279
rect 31421 4903 31455 5279
rect 31539 4903 31573 5279
rect 31668 4903 31702 5079
rect 31786 4903 31820 5079
rect 31904 4903 31938 5079
rect 32022 4903 32056 5079
rect 32140 4900 32174 5076
rect 32258 4900 32292 5076
rect 32376 4900 32410 5076
rect 32494 4900 32528 5076
rect 32612 4900 32646 5076
rect 32730 4900 32764 5076
rect 32848 4900 32882 5076
rect 32966 4900 33000 5076
rect 33084 4900 33118 5076
rect 33202 4900 33236 5076
rect 19 3555 53 3731
rect 137 3555 171 3731
rect 255 3555 289 3731
rect 373 3555 407 3731
rect 491 3555 525 3731
rect 609 3555 643 3731
rect 727 3555 761 3731
rect 845 3555 879 3731
rect 963 3555 997 3731
rect 1081 3555 1115 3731
rect 30774 4210 30808 4586
rect 30892 4210 30926 4586
rect 31010 4210 31044 4586
rect 31128 4210 31162 4586
rect 31246 4210 31280 4586
rect 31364 4210 31398 4586
rect 31482 4210 31516 4586
rect 2909 3288 2943 3464
rect 3027 3288 3061 3464
rect 3145 3288 3179 3464
rect 3263 3288 3297 3464
rect 3381 3288 3415 3464
rect 3499 3288 3533 3464
rect 3617 3288 3651 3464
rect 3735 3288 3769 3464
rect 3853 3288 3887 3464
rect 3971 3288 4005 3464
rect 5234 3160 5268 3536
rect 5352 3160 5386 3536
rect 5470 3160 5504 3536
rect 5588 3160 5622 3536
rect 5706 3160 5740 3536
rect 5824 3160 5858 3536
rect 5942 3160 5976 3536
rect 6376 3164 6410 3540
rect 6494 3164 6528 3540
rect 6612 3164 6646 3540
rect 6730 3164 6764 3540
rect 6848 3164 6882 3540
rect 6966 3164 7000 3540
rect 7084 3164 7118 3540
rect 9458 3376 9492 3552
rect 9576 3376 9610 3552
rect 9694 3376 9728 3552
rect 9812 3376 9846 3552
rect 9930 3376 9964 3552
rect 10048 3376 10082 3552
rect 10166 3376 10200 3552
rect 10284 3376 10318 3552
rect 10402 3376 10436 3552
rect 10520 3376 10554 3552
rect 11783 3248 11817 3624
rect 11901 3248 11935 3624
rect 12019 3248 12053 3624
rect 12137 3248 12171 3624
rect 12255 3248 12289 3624
rect 12373 3248 12407 3624
rect 12491 3248 12525 3624
rect 12925 3252 12959 3628
rect 13043 3252 13077 3628
rect 13161 3252 13195 3628
rect 13279 3252 13313 3628
rect 13397 3252 13431 3628
rect 13515 3252 13549 3628
rect 13633 3252 13667 3628
rect 16112 3308 16146 3484
rect 16230 3308 16264 3484
rect 16348 3308 16382 3484
rect 16466 3308 16500 3484
rect 16584 3308 16618 3484
rect 16702 3308 16736 3484
rect 16820 3308 16854 3484
rect 16938 3308 16972 3484
rect 17056 3308 17090 3484
rect 17174 3308 17208 3484
rect 5663 2577 5697 2753
rect 5781 2577 5815 2753
rect 5899 2577 5933 2753
rect 6017 2577 6051 2753
rect 6805 2581 6839 2757
rect 6923 2581 6957 2757
rect 7041 2581 7075 2757
rect 7159 2581 7193 2757
rect 18437 3180 18471 3556
rect 18555 3180 18589 3556
rect 18673 3180 18707 3556
rect 18791 3180 18825 3556
rect 18909 3180 18943 3556
rect 19027 3180 19061 3556
rect 19145 3180 19179 3556
rect 19579 3184 19613 3560
rect 19697 3184 19731 3560
rect 19815 3184 19849 3560
rect 19933 3184 19967 3560
rect 20051 3184 20085 3560
rect 20169 3184 20203 3560
rect 20287 3184 20321 3560
rect 22737 3376 22771 3552
rect 22855 3376 22889 3552
rect 22973 3376 23007 3552
rect 23091 3376 23125 3552
rect 23209 3376 23243 3552
rect 23327 3376 23361 3552
rect 23445 3376 23479 3552
rect 23563 3376 23597 3552
rect 23681 3376 23715 3552
rect 23799 3376 23833 3552
rect 12212 2665 12246 2841
rect 12330 2665 12364 2841
rect 12448 2665 12482 2841
rect 12566 2665 12600 2841
rect 13354 2669 13388 2845
rect 13472 2669 13506 2845
rect 13590 2669 13624 2845
rect 13708 2669 13742 2845
rect 25062 3248 25096 3624
rect 25180 3248 25214 3624
rect 25298 3248 25332 3624
rect 25416 3248 25450 3624
rect 25534 3248 25568 3624
rect 25652 3248 25686 3624
rect 25770 3248 25804 3624
rect 26204 3252 26238 3628
rect 26322 3252 26356 3628
rect 26440 3252 26474 3628
rect 26558 3252 26592 3628
rect 26676 3252 26710 3628
rect 26794 3252 26828 3628
rect 26912 3252 26946 3628
rect 18866 2597 18900 2773
rect 18984 2597 19018 2773
rect 19102 2597 19136 2773
rect 19220 2597 19254 2773
rect 20008 2601 20042 2777
rect 20126 2601 20160 2777
rect 20244 2601 20278 2777
rect 20362 2601 20396 2777
rect 25491 2665 25525 2841
rect 25609 2665 25643 2841
rect 25727 2665 25761 2841
rect 25845 2665 25879 2841
rect 26633 2669 26667 2845
rect 26751 2669 26785 2845
rect 26869 2669 26903 2845
rect 26987 2669 27021 2845
rect 28534 2737 28568 2913
rect 28652 2737 28686 2913
rect 28770 2737 28804 2913
rect 28888 2737 28922 2913
rect 29006 2737 29040 2913
rect 29124 2737 29158 2913
rect 29242 2737 29276 2913
rect 29360 2737 29394 2913
rect 29478 2737 29512 2913
rect 29596 2737 29630 2913
rect 2923 1638 2957 1814
rect 3041 1638 3075 1814
rect 3159 1638 3193 1814
rect 3277 1638 3311 1814
rect 3395 1638 3429 1814
rect 3513 1638 3547 1814
rect 3631 1638 3665 1814
rect 3749 1638 3783 1814
rect 3867 1638 3901 1814
rect 3985 1638 4019 1814
rect 9472 1726 9506 1902
rect 9590 1726 9624 1902
rect 9708 1726 9742 1902
rect 9826 1726 9860 1902
rect 9944 1726 9978 1902
rect 10062 1726 10096 1902
rect 10180 1726 10214 1902
rect 10298 1726 10332 1902
rect 10416 1726 10450 1902
rect 10534 1726 10568 1902
rect 16126 1658 16160 1834
rect 16244 1658 16278 1834
rect 16362 1658 16396 1834
rect 16480 1658 16514 1834
rect 16598 1658 16632 1834
rect 16716 1658 16750 1834
rect 16834 1658 16868 1834
rect 16952 1658 16986 1834
rect 17070 1658 17104 1834
rect 17188 1658 17222 1834
rect 22751 1726 22785 1902
rect 22869 1726 22903 1902
rect 22987 1726 23021 1902
rect 23105 1726 23139 1902
rect 23223 1726 23257 1902
rect 23341 1726 23375 1902
rect 23459 1726 23493 1902
rect 23577 1726 23611 1902
rect 23695 1726 23729 1902
rect 23813 1726 23847 1902
rect 11 970 45 1146
rect 129 970 163 1146
rect 247 970 281 1146
rect 365 970 399 1146
rect 483 970 517 1146
rect 601 970 635 1146
rect 719 970 753 1146
rect 837 970 871 1146
rect 955 970 989 1146
rect 1073 970 1107 1146
rect 4387 1021 4421 1197
rect 4505 1021 4539 1197
rect 4623 1021 4657 1197
rect 4741 1021 4775 1197
rect 4871 1021 4905 1397
rect 4989 1021 5023 1397
rect 5107 1021 5141 1397
rect 5225 1021 5259 1397
rect 5343 1021 5377 1397
rect 5461 1021 5495 1397
rect 5579 1021 5613 1397
rect 5708 1021 5742 1197
rect 5826 1021 5860 1197
rect 5944 1021 5978 1197
rect 6062 1021 6096 1197
rect 6285 1021 6319 1197
rect 6403 1021 6437 1197
rect 6521 1021 6555 1197
rect 6639 1021 6673 1197
rect 6769 1021 6803 1397
rect 6887 1021 6921 1397
rect 7005 1021 7039 1397
rect 7123 1021 7157 1397
rect 7241 1021 7275 1397
rect 7359 1021 7393 1397
rect 7477 1021 7511 1397
rect 7606 1021 7640 1197
rect 7724 1021 7758 1197
rect 7842 1021 7876 1197
rect 7960 1021 7994 1197
rect 2918 34 2952 210
rect 3036 34 3070 210
rect 3154 34 3188 210
rect 3272 34 3306 210
rect 3390 34 3424 210
rect 3508 34 3542 210
rect 3626 34 3660 210
rect 3744 34 3778 210
rect 3862 34 3896 210
rect 3980 34 4014 210
rect 4814 328 4848 704
rect 4932 328 4966 704
rect 5050 328 5084 704
rect 5168 328 5202 704
rect 5286 328 5320 704
rect 5404 328 5438 704
rect 5522 328 5556 704
rect 10936 1109 10970 1285
rect 11054 1109 11088 1285
rect 11172 1109 11206 1285
rect 11290 1109 11324 1285
rect 11420 1109 11454 1485
rect 11538 1109 11572 1485
rect 11656 1109 11690 1485
rect 11774 1109 11808 1485
rect 11892 1109 11926 1485
rect 12010 1109 12044 1485
rect 12128 1109 12162 1485
rect 12257 1109 12291 1285
rect 12375 1109 12409 1285
rect 12493 1109 12527 1285
rect 12611 1109 12645 1285
rect 12834 1109 12868 1285
rect 12952 1109 12986 1285
rect 13070 1109 13104 1285
rect 13188 1109 13222 1285
rect 13318 1109 13352 1485
rect 13436 1109 13470 1485
rect 13554 1109 13588 1485
rect 13672 1109 13706 1485
rect 13790 1109 13824 1485
rect 13908 1109 13942 1485
rect 14026 1109 14060 1485
rect 14155 1109 14189 1285
rect 14273 1109 14307 1285
rect 14391 1109 14425 1285
rect 14509 1109 14543 1285
rect 6712 328 6746 704
rect 6830 328 6864 704
rect 6948 328 6982 704
rect 7066 328 7100 704
rect 7184 328 7218 704
rect 7302 328 7336 704
rect 7420 328 7454 704
rect 9467 122 9501 298
rect 9585 122 9619 298
rect 9703 122 9737 298
rect 9821 122 9855 298
rect 9939 122 9973 298
rect 10057 122 10091 298
rect 10175 122 10209 298
rect 10293 122 10327 298
rect 10411 122 10445 298
rect 10529 122 10563 298
rect 11363 416 11397 792
rect 11481 416 11515 792
rect 11599 416 11633 792
rect 11717 416 11751 792
rect 11835 416 11869 792
rect 11953 416 11987 792
rect 12071 416 12105 792
rect 17590 1041 17624 1217
rect 17708 1041 17742 1217
rect 17826 1041 17860 1217
rect 17944 1041 17978 1217
rect 18074 1041 18108 1417
rect 18192 1041 18226 1417
rect 18310 1041 18344 1417
rect 18428 1041 18462 1417
rect 18546 1041 18580 1417
rect 18664 1041 18698 1417
rect 18782 1041 18816 1417
rect 18911 1041 18945 1217
rect 19029 1041 19063 1217
rect 19147 1041 19181 1217
rect 19265 1041 19299 1217
rect 19488 1041 19522 1217
rect 19606 1041 19640 1217
rect 19724 1041 19758 1217
rect 19842 1041 19876 1217
rect 19972 1041 20006 1417
rect 20090 1041 20124 1417
rect 20208 1041 20242 1417
rect 20326 1041 20360 1417
rect 20444 1041 20478 1417
rect 20562 1041 20596 1417
rect 20680 1041 20714 1417
rect 20809 1041 20843 1217
rect 20927 1041 20961 1217
rect 21045 1041 21079 1217
rect 21163 1041 21197 1217
rect 13261 416 13295 792
rect 13379 416 13413 792
rect 13497 416 13531 792
rect 13615 416 13649 792
rect 13733 416 13767 792
rect 13851 416 13885 792
rect 13969 416 14003 792
rect 16121 54 16155 230
rect 16239 54 16273 230
rect 16357 54 16391 230
rect 16475 54 16509 230
rect 16593 54 16627 230
rect 16711 54 16745 230
rect 16829 54 16863 230
rect 16947 54 16981 230
rect 17065 54 17099 230
rect 17183 54 17217 230
rect 18017 348 18051 724
rect 18135 348 18169 724
rect 18253 348 18287 724
rect 18371 348 18405 724
rect 18489 348 18523 724
rect 18607 348 18641 724
rect 18725 348 18759 724
rect 24215 1109 24249 1285
rect 24333 1109 24367 1285
rect 24451 1109 24485 1285
rect 24569 1109 24603 1285
rect 24699 1109 24733 1485
rect 24817 1109 24851 1485
rect 24935 1109 24969 1485
rect 25053 1109 25087 1485
rect 25171 1109 25205 1485
rect 25289 1109 25323 1485
rect 25407 1109 25441 1485
rect 25536 1109 25570 1285
rect 25654 1109 25688 1285
rect 25772 1109 25806 1285
rect 25890 1109 25924 1285
rect 26113 1109 26147 1285
rect 26231 1109 26265 1285
rect 26349 1109 26383 1285
rect 26467 1109 26501 1285
rect 26597 1109 26631 1485
rect 26715 1109 26749 1485
rect 26833 1109 26867 1485
rect 26951 1109 26985 1485
rect 27069 1109 27103 1485
rect 27187 1109 27221 1485
rect 27305 1109 27339 1485
rect 27434 1109 27468 1285
rect 27552 1109 27586 1285
rect 27670 1109 27704 1285
rect 27788 1109 27822 1285
rect 19915 348 19949 724
rect 20033 348 20067 724
rect 20151 348 20185 724
rect 20269 348 20303 724
rect 20387 348 20421 724
rect 20505 348 20539 724
rect 20623 348 20657 724
rect 22746 122 22780 298
rect 22864 122 22898 298
rect 22982 122 23016 298
rect 23100 122 23134 298
rect 23218 122 23252 298
rect 23336 122 23370 298
rect 23454 122 23488 298
rect 23572 122 23606 298
rect 23690 122 23724 298
rect 23808 122 23842 298
rect 24642 416 24676 792
rect 24760 416 24794 792
rect 24878 416 24912 792
rect 24996 416 25030 792
rect 25114 416 25148 792
rect 25232 416 25266 792
rect 25350 416 25384 792
rect 26540 416 26574 792
rect 26658 416 26692 792
rect 26776 416 26810 792
rect 26894 416 26928 792
rect 27012 416 27046 792
rect 27130 416 27164 792
rect 27248 416 27282 792
rect 30349 812 30383 988
rect 30467 812 30501 988
rect 30585 812 30619 988
rect 30703 812 30737 988
rect 30833 812 30867 1188
rect 30951 812 30985 1188
rect 31069 812 31103 1188
rect 31187 812 31221 1188
rect 31305 812 31339 1188
rect 31423 812 31457 1188
rect 31541 812 31575 1188
rect 31670 812 31704 988
rect 31788 812 31822 988
rect 31906 812 31940 988
rect 32024 812 32058 988
rect 32142 809 32176 985
rect 32260 809 32294 985
rect 32378 809 32412 985
rect 32496 809 32530 985
rect 32614 809 32648 985
rect 32732 809 32766 985
rect 32850 809 32884 985
rect 32968 809 33002 985
rect 33086 809 33120 985
rect 33204 809 33238 985
rect 28534 -296 28568 -120
rect 28652 -296 28686 -120
rect 28770 -296 28804 -120
rect 28888 -296 28922 -120
rect 29006 -296 29040 -120
rect 29124 -296 29158 -120
rect 29242 -296 29276 -120
rect 29360 -296 29394 -120
rect 29478 -296 29512 -120
rect 29596 -296 29630 -120
rect 30776 119 30810 495
rect 30894 119 30928 495
rect 31012 119 31046 495
rect 31130 119 31164 495
rect 31248 119 31282 495
rect 31366 119 31400 495
rect 31484 119 31518 495
rect -8 -2308 26 -2132
rect 110 -2308 144 -2132
rect 228 -2308 262 -2132
rect 346 -2308 380 -2132
rect 464 -2308 498 -2132
rect 582 -2308 616 -2132
rect 700 -2308 734 -2132
rect 818 -2308 852 -2132
rect 936 -2308 970 -2132
rect 1054 -2308 1088 -2132
rect 2901 -2492 2935 -2316
rect 3019 -2492 3053 -2316
rect 3137 -2492 3171 -2316
rect 3255 -2492 3289 -2316
rect 3373 -2492 3407 -2316
rect 3491 -2492 3525 -2316
rect 3609 -2492 3643 -2316
rect 3727 -2492 3761 -2316
rect 3845 -2492 3879 -2316
rect 3963 -2492 3997 -2316
rect 5226 -2620 5260 -2244
rect 5344 -2620 5378 -2244
rect 5462 -2620 5496 -2244
rect 5580 -2620 5614 -2244
rect 5698 -2620 5732 -2244
rect 5816 -2620 5850 -2244
rect 5934 -2620 5968 -2244
rect 6368 -2616 6402 -2240
rect 6486 -2616 6520 -2240
rect 6604 -2616 6638 -2240
rect 6722 -2616 6756 -2240
rect 6840 -2616 6874 -2240
rect 6958 -2616 6992 -2240
rect 7076 -2616 7110 -2240
rect 9452 -2494 9486 -2318
rect 9570 -2494 9604 -2318
rect 9688 -2494 9722 -2318
rect 9806 -2494 9840 -2318
rect 9924 -2494 9958 -2318
rect 10042 -2494 10076 -2318
rect 10160 -2494 10194 -2318
rect 10278 -2494 10312 -2318
rect 10396 -2494 10430 -2318
rect 10514 -2494 10548 -2318
rect 11777 -2622 11811 -2246
rect 11895 -2622 11929 -2246
rect 12013 -2622 12047 -2246
rect 12131 -2622 12165 -2246
rect 12249 -2622 12283 -2246
rect 12367 -2622 12401 -2246
rect 12485 -2622 12519 -2246
rect 12919 -2618 12953 -2242
rect 13037 -2618 13071 -2242
rect 13155 -2618 13189 -2242
rect 13273 -2618 13307 -2242
rect 13391 -2618 13425 -2242
rect 13509 -2618 13543 -2242
rect 13627 -2618 13661 -2242
rect 16107 -2493 16141 -2317
rect 16225 -2493 16259 -2317
rect 16343 -2493 16377 -2317
rect 16461 -2493 16495 -2317
rect 16579 -2493 16613 -2317
rect 16697 -2493 16731 -2317
rect 16815 -2493 16849 -2317
rect 16933 -2493 16967 -2317
rect 17051 -2493 17085 -2317
rect 17169 -2493 17203 -2317
rect 5655 -3203 5689 -3027
rect 5773 -3203 5807 -3027
rect 5891 -3203 5925 -3027
rect 6009 -3203 6043 -3027
rect 6797 -3199 6831 -3023
rect 6915 -3199 6949 -3023
rect 7033 -3199 7067 -3023
rect 7151 -3199 7185 -3023
rect 18432 -2621 18466 -2245
rect 18550 -2621 18584 -2245
rect 18668 -2621 18702 -2245
rect 18786 -2621 18820 -2245
rect 18904 -2621 18938 -2245
rect 19022 -2621 19056 -2245
rect 19140 -2621 19174 -2245
rect 19574 -2617 19608 -2241
rect 19692 -2617 19726 -2241
rect 19810 -2617 19844 -2241
rect 19928 -2617 19962 -2241
rect 20046 -2617 20080 -2241
rect 20164 -2617 20198 -2241
rect 28605 -2216 28639 -2040
rect 28723 -2216 28757 -2040
rect 28841 -2216 28875 -2040
rect 28959 -2216 28993 -2040
rect 29077 -2216 29111 -2040
rect 29195 -2216 29229 -2040
rect 29313 -2216 29347 -2040
rect 29431 -2216 29465 -2040
rect 29549 -2216 29583 -2040
rect 29667 -2216 29701 -2040
rect 20282 -2617 20316 -2241
rect 22729 -2492 22763 -2316
rect 22847 -2492 22881 -2316
rect 22965 -2492 22999 -2316
rect 23083 -2492 23117 -2316
rect 23201 -2492 23235 -2316
rect 23319 -2492 23353 -2316
rect 23437 -2492 23471 -2316
rect 23555 -2492 23589 -2316
rect 23673 -2492 23707 -2316
rect 23791 -2492 23825 -2316
rect 12206 -3205 12240 -3029
rect 12324 -3205 12358 -3029
rect 12442 -3205 12476 -3029
rect 12560 -3205 12594 -3029
rect 13348 -3201 13382 -3025
rect 13466 -3201 13500 -3025
rect 13584 -3201 13618 -3025
rect 13702 -3201 13736 -3025
rect 25054 -2620 25088 -2244
rect 25172 -2620 25206 -2244
rect 25290 -2620 25324 -2244
rect 25408 -2620 25442 -2244
rect 25526 -2620 25560 -2244
rect 25644 -2620 25678 -2244
rect 25762 -2620 25796 -2244
rect 26196 -2616 26230 -2240
rect 26314 -2616 26348 -2240
rect 26432 -2616 26466 -2240
rect 26550 -2616 26584 -2240
rect 26668 -2616 26702 -2240
rect 26786 -2616 26820 -2240
rect 26904 -2616 26938 -2240
rect 18861 -3204 18895 -3028
rect 18979 -3204 19013 -3028
rect 19097 -3204 19131 -3028
rect 19215 -3204 19249 -3028
rect 20003 -3200 20037 -3024
rect 20121 -3200 20155 -3024
rect 20239 -3200 20273 -3024
rect 20357 -3200 20391 -3024
rect 30349 -2683 30383 -2507
rect 30467 -2683 30501 -2507
rect 30585 -2683 30619 -2507
rect 30703 -2683 30737 -2507
rect 30833 -2683 30867 -2307
rect 30951 -2683 30985 -2307
rect 31069 -2683 31103 -2307
rect 31187 -2683 31221 -2307
rect 31305 -2683 31339 -2307
rect 31423 -2683 31457 -2307
rect 31541 -2683 31575 -2307
rect 31670 -2683 31704 -2507
rect 31788 -2683 31822 -2507
rect 31906 -2683 31940 -2507
rect 32024 -2683 32058 -2507
rect 32142 -2686 32176 -2510
rect 32260 -2686 32294 -2510
rect 32378 -2686 32412 -2510
rect 32496 -2686 32530 -2510
rect 32614 -2686 32648 -2510
rect 32732 -2686 32766 -2510
rect 32850 -2686 32884 -2510
rect 32968 -2686 33002 -2510
rect 33086 -2686 33120 -2510
rect 33204 -2686 33238 -2510
rect 25483 -3203 25517 -3027
rect 25601 -3203 25635 -3027
rect 25719 -3203 25753 -3027
rect 25837 -3203 25871 -3027
rect 26625 -3199 26659 -3023
rect 26743 -3199 26777 -3023
rect 26861 -3199 26895 -3023
rect 26979 -3199 27013 -3023
rect 30776 -3376 30810 -3000
rect 30894 -3376 30928 -3000
rect 31012 -3376 31046 -3000
rect 31130 -3376 31164 -3000
rect 31248 -3376 31282 -3000
rect 31366 -3376 31400 -3000
rect 31484 -3376 31518 -3000
rect 2915 -4142 2949 -3966
rect 3033 -4142 3067 -3966
rect 3151 -4142 3185 -3966
rect 3269 -4142 3303 -3966
rect 3387 -4142 3421 -3966
rect 3505 -4142 3539 -3966
rect 3623 -4142 3657 -3966
rect 3741 -4142 3775 -3966
rect 3859 -4142 3893 -3966
rect 3977 -4142 4011 -3966
rect 9466 -4144 9500 -3968
rect 9584 -4144 9618 -3968
rect 9702 -4144 9736 -3968
rect 9820 -4144 9854 -3968
rect 9938 -4144 9972 -3968
rect 10056 -4144 10090 -3968
rect 10174 -4144 10208 -3968
rect 10292 -4144 10326 -3968
rect 10410 -4144 10444 -3968
rect 10528 -4144 10562 -3968
rect 16121 -4143 16155 -3967
rect 16239 -4143 16273 -3967
rect 16357 -4143 16391 -3967
rect 16475 -4143 16509 -3967
rect 16593 -4143 16627 -3967
rect 16711 -4143 16745 -3967
rect 16829 -4143 16863 -3967
rect 16947 -4143 16981 -3967
rect 17065 -4143 17099 -3967
rect 17183 -4143 17217 -3967
rect 22743 -4142 22777 -3966
rect 22861 -4142 22895 -3966
rect 22979 -4142 23013 -3966
rect 23097 -4142 23131 -3966
rect 23215 -4142 23249 -3966
rect 23333 -4142 23367 -3966
rect 23451 -4142 23485 -3966
rect 23569 -4142 23603 -3966
rect 23687 -4142 23721 -3966
rect 23805 -4142 23839 -3966
rect 4379 -4759 4413 -4583
rect 4497 -4759 4531 -4583
rect 4615 -4759 4649 -4583
rect 4733 -4759 4767 -4583
rect 4863 -4759 4897 -4383
rect 4981 -4759 5015 -4383
rect 5099 -4759 5133 -4383
rect 5217 -4759 5251 -4383
rect 5335 -4759 5369 -4383
rect 5453 -4759 5487 -4383
rect 5571 -4759 5605 -4383
rect 5700 -4759 5734 -4583
rect 5818 -4759 5852 -4583
rect 5936 -4759 5970 -4583
rect 6054 -4759 6088 -4583
rect 6277 -4759 6311 -4583
rect 6395 -4759 6429 -4583
rect 6513 -4759 6547 -4583
rect 6631 -4759 6665 -4583
rect 6761 -4759 6795 -4383
rect 6879 -4759 6913 -4383
rect 6997 -4759 7031 -4383
rect 7115 -4759 7149 -4383
rect 7233 -4759 7267 -4383
rect 7351 -4759 7385 -4383
rect 7469 -4759 7503 -4383
rect 7598 -4759 7632 -4583
rect 7716 -4759 7750 -4583
rect 7834 -4759 7868 -4583
rect 7952 -4759 7986 -4583
rect 8 -5068 42 -4892
rect 126 -5068 160 -4892
rect 244 -5068 278 -4892
rect 362 -5068 396 -4892
rect 480 -5068 514 -4892
rect 598 -5068 632 -4892
rect 716 -5068 750 -4892
rect 834 -5068 868 -4892
rect 952 -5068 986 -4892
rect 1070 -5068 1104 -4892
rect 2910 -5746 2944 -5570
rect 3028 -5746 3062 -5570
rect 3146 -5746 3180 -5570
rect 3264 -5746 3298 -5570
rect 3382 -5746 3416 -5570
rect 3500 -5746 3534 -5570
rect 3618 -5746 3652 -5570
rect 3736 -5746 3770 -5570
rect 3854 -5746 3888 -5570
rect 3972 -5746 4006 -5570
rect 4806 -5452 4840 -5076
rect 4924 -5452 4958 -5076
rect 5042 -5452 5076 -5076
rect 5160 -5452 5194 -5076
rect 5278 -5452 5312 -5076
rect 5396 -5452 5430 -5076
rect 5514 -5452 5548 -5076
rect 10930 -4761 10964 -4585
rect 11048 -4761 11082 -4585
rect 11166 -4761 11200 -4585
rect 11284 -4761 11318 -4585
rect 11414 -4761 11448 -4385
rect 11532 -4761 11566 -4385
rect 11650 -4761 11684 -4385
rect 11768 -4761 11802 -4385
rect 11886 -4761 11920 -4385
rect 12004 -4761 12038 -4385
rect 12122 -4761 12156 -4385
rect 12251 -4761 12285 -4585
rect 12369 -4761 12403 -4585
rect 12487 -4761 12521 -4585
rect 12605 -4761 12639 -4585
rect 12828 -4761 12862 -4585
rect 12946 -4761 12980 -4585
rect 13064 -4761 13098 -4585
rect 13182 -4761 13216 -4585
rect 13312 -4761 13346 -4385
rect 13430 -4761 13464 -4385
rect 13548 -4761 13582 -4385
rect 13666 -4761 13700 -4385
rect 13784 -4761 13818 -4385
rect 13902 -4761 13936 -4385
rect 14020 -4761 14054 -4385
rect 14149 -4761 14183 -4585
rect 14267 -4761 14301 -4585
rect 14385 -4761 14419 -4585
rect 14503 -4761 14537 -4585
rect 6704 -5452 6738 -5076
rect 6822 -5452 6856 -5076
rect 6940 -5452 6974 -5076
rect 7058 -5452 7092 -5076
rect 7176 -5452 7210 -5076
rect 7294 -5452 7328 -5076
rect 7412 -5452 7446 -5076
rect 9461 -5748 9495 -5572
rect 9579 -5748 9613 -5572
rect 9697 -5748 9731 -5572
rect 9815 -5748 9849 -5572
rect 9933 -5748 9967 -5572
rect 10051 -5748 10085 -5572
rect 10169 -5748 10203 -5572
rect 10287 -5748 10321 -5572
rect 10405 -5748 10439 -5572
rect 10523 -5748 10557 -5572
rect 11357 -5454 11391 -5078
rect 11475 -5454 11509 -5078
rect 11593 -5454 11627 -5078
rect 11711 -5454 11745 -5078
rect 11829 -5454 11863 -5078
rect 11947 -5454 11981 -5078
rect 12065 -5454 12099 -5078
rect 17585 -4760 17619 -4584
rect 17703 -4760 17737 -4584
rect 17821 -4760 17855 -4584
rect 17939 -4760 17973 -4584
rect 18069 -4760 18103 -4384
rect 18187 -4760 18221 -4384
rect 18305 -4760 18339 -4384
rect 18423 -4760 18457 -4384
rect 18541 -4760 18575 -4384
rect 18659 -4760 18693 -4384
rect 18777 -4760 18811 -4384
rect 18906 -4760 18940 -4584
rect 19024 -4760 19058 -4584
rect 19142 -4760 19176 -4584
rect 19260 -4760 19294 -4584
rect 19483 -4760 19517 -4584
rect 19601 -4760 19635 -4584
rect 19719 -4760 19753 -4584
rect 19837 -4760 19871 -4584
rect 19967 -4760 20001 -4384
rect 20085 -4760 20119 -4384
rect 20203 -4760 20237 -4384
rect 20321 -4760 20355 -4384
rect 20439 -4760 20473 -4384
rect 20557 -4760 20591 -4384
rect 20675 -4760 20709 -4384
rect 20804 -4760 20838 -4584
rect 20922 -4760 20956 -4584
rect 21040 -4760 21074 -4584
rect 21158 -4760 21192 -4584
rect 13255 -5454 13289 -5078
rect 13373 -5454 13407 -5078
rect 13491 -5454 13525 -5078
rect 13609 -5454 13643 -5078
rect 13727 -5454 13761 -5078
rect 13845 -5454 13879 -5078
rect 13963 -5454 13997 -5078
rect 16116 -5747 16150 -5571
rect 16234 -5747 16268 -5571
rect 16352 -5747 16386 -5571
rect 16470 -5747 16504 -5571
rect 16588 -5747 16622 -5571
rect 16706 -5747 16740 -5571
rect 16824 -5747 16858 -5571
rect 16942 -5747 16976 -5571
rect 17060 -5747 17094 -5571
rect 17178 -5747 17212 -5571
rect 18012 -5453 18046 -5077
rect 18130 -5453 18164 -5077
rect 18248 -5453 18282 -5077
rect 18366 -5453 18400 -5077
rect 18484 -5453 18518 -5077
rect 18602 -5453 18636 -5077
rect 18720 -5453 18754 -5077
rect 24207 -4759 24241 -4583
rect 24325 -4759 24359 -4583
rect 24443 -4759 24477 -4583
rect 24561 -4759 24595 -4583
rect 24691 -4759 24725 -4383
rect 24809 -4759 24843 -4383
rect 24927 -4759 24961 -4383
rect 25045 -4759 25079 -4383
rect 25163 -4759 25197 -4383
rect 25281 -4759 25315 -4383
rect 25399 -4759 25433 -4383
rect 25528 -4759 25562 -4583
rect 25646 -4759 25680 -4583
rect 25764 -4759 25798 -4583
rect 25882 -4759 25916 -4583
rect 26105 -4759 26139 -4583
rect 26223 -4759 26257 -4583
rect 26341 -4759 26375 -4583
rect 26459 -4759 26493 -4583
rect 26589 -4759 26623 -4383
rect 26707 -4759 26741 -4383
rect 26825 -4759 26859 -4383
rect 26943 -4759 26977 -4383
rect 27061 -4759 27095 -4383
rect 27179 -4759 27213 -4383
rect 27297 -4759 27331 -4383
rect 27426 -4759 27460 -4583
rect 27544 -4759 27578 -4583
rect 27662 -4759 27696 -4583
rect 27780 -4759 27814 -4583
rect 19910 -5453 19944 -5077
rect 20028 -5453 20062 -5077
rect 20146 -5453 20180 -5077
rect 20264 -5453 20298 -5077
rect 20382 -5453 20416 -5077
rect 20500 -5453 20534 -5077
rect 20618 -5453 20652 -5077
rect 22738 -5746 22772 -5570
rect 22856 -5746 22890 -5570
rect 22974 -5746 23008 -5570
rect 23092 -5746 23126 -5570
rect 23210 -5746 23244 -5570
rect 23328 -5746 23362 -5570
rect 23446 -5746 23480 -5570
rect 23564 -5746 23598 -5570
rect 23682 -5746 23716 -5570
rect 23800 -5746 23834 -5570
rect 24634 -5452 24668 -5076
rect 24752 -5452 24786 -5076
rect 24870 -5452 24904 -5076
rect 24988 -5452 25022 -5076
rect 25106 -5452 25140 -5076
rect 25224 -5452 25258 -5076
rect 25342 -5452 25376 -5076
rect 26532 -5452 26566 -5076
rect 26650 -5452 26684 -5076
rect 26768 -5452 26802 -5076
rect 26886 -5452 26920 -5076
rect 27004 -5452 27038 -5076
rect 27122 -5452 27156 -5076
rect 27240 -5452 27274 -5076
rect 28602 -5286 28636 -5110
rect 28720 -5286 28754 -5110
rect 28838 -5286 28872 -5110
rect 28956 -5286 28990 -5110
rect 29074 -5286 29108 -5110
rect 29192 -5286 29226 -5110
rect 29310 -5286 29344 -5110
rect 29428 -5286 29462 -5110
rect 29546 -5286 29580 -5110
rect 29664 -5286 29698 -5110
rect 30349 -7031 30383 -6855
rect 30467 -7031 30501 -6855
rect 30585 -7031 30619 -6855
rect 30703 -7031 30737 -6855
rect 30833 -7031 30867 -6655
rect 30951 -7031 30985 -6655
rect 31069 -7031 31103 -6655
rect 31187 -7031 31221 -6655
rect 31305 -7031 31339 -6655
rect 31423 -7031 31457 -6655
rect 31541 -7031 31575 -6655
rect 31670 -7031 31704 -6855
rect 31788 -7031 31822 -6855
rect 31906 -7031 31940 -6855
rect 32024 -7031 32058 -6855
rect 32142 -7034 32176 -6858
rect 32260 -7034 32294 -6858
rect 32378 -7034 32412 -6858
rect 32496 -7034 32530 -6858
rect 32614 -7034 32648 -6858
rect 32732 -7034 32766 -6858
rect 32850 -7034 32884 -6858
rect 32968 -7034 33002 -6858
rect 33086 -7034 33120 -6858
rect 33204 -7034 33238 -6858
rect 6718 -8249 6752 -8073
rect 6836 -8249 6870 -8073
rect 6954 -8249 6988 -8073
rect 7072 -8249 7106 -8073
rect 7190 -8249 7224 -8073
rect 7308 -8249 7342 -8073
rect 7426 -8249 7460 -8073
rect 7544 -8249 7578 -8073
rect 7662 -8249 7696 -8073
rect 7780 -8249 7814 -8073
rect 13272 -8244 13306 -8068
rect 13390 -8244 13424 -8068
rect 13508 -8244 13542 -8068
rect 13626 -8244 13660 -8068
rect 13744 -8244 13778 -8068
rect 13862 -8244 13896 -8068
rect 13980 -8244 14014 -8068
rect 14098 -8244 14132 -8068
rect 14216 -8244 14250 -8068
rect 14334 -8244 14368 -8068
rect 19921 -8256 19955 -8080
rect 20039 -8256 20073 -8080
rect 20157 -8256 20191 -8080
rect 20275 -8256 20309 -8080
rect 20393 -8256 20427 -8080
rect 20511 -8256 20545 -8080
rect 20629 -8256 20663 -8080
rect 20747 -8256 20781 -8080
rect 20865 -8256 20899 -8080
rect 20983 -8256 21017 -8080
rect 28609 -8131 28643 -7955
rect 28727 -8131 28761 -7955
rect 28845 -8131 28879 -7955
rect 28963 -8131 28997 -7955
rect 29081 -8131 29115 -7955
rect 29199 -8131 29233 -7955
rect 29317 -8131 29351 -7955
rect 29435 -8131 29469 -7955
rect 29553 -8131 29587 -7955
rect 29671 -8131 29705 -7955
rect 30776 -7724 30810 -7348
rect 30894 -7724 30928 -7348
rect 31012 -7724 31046 -7348
rect 31130 -7724 31164 -7348
rect 31248 -7724 31282 -7348
rect 31366 -7724 31400 -7348
rect 31484 -7724 31518 -7348
<< psubdiff >>
rect 7172 4663 7384 4693
rect 7172 4607 7212 4663
rect 7346 4607 7384 4663
rect 7172 4585 7384 4607
rect 13721 4662 13933 4692
rect 13721 4606 13761 4662
rect 13895 4606 13933 4662
rect 13721 4584 13933 4606
rect 20375 4683 20587 4713
rect 20375 4627 20415 4683
rect 20549 4627 20587 4683
rect 20375 4605 20587 4627
rect 29028 4516 29240 4546
rect 29028 4460 29068 4516
rect 29202 4460 29240 4516
rect 29028 4438 29240 4460
rect 32629 4108 32841 4138
rect 32629 4052 32669 4108
rect 32803 4052 32841 4108
rect 32629 4030 32841 4052
rect 508 2763 720 2793
rect 508 2707 548 2763
rect 682 2707 720 2763
rect 508 2685 720 2707
rect 3670 2701 3904 2735
rect 3670 2611 3716 2701
rect 3879 2611 3904 2701
rect 3670 2580 3904 2611
rect 10219 2789 10453 2823
rect 10219 2699 10265 2789
rect 10428 2699 10453 2789
rect 10219 2668 10453 2699
rect 31039 3307 31281 3319
rect 16873 2721 17107 2755
rect 16873 2631 16919 2721
rect 17082 2631 17107 2721
rect 16873 2600 17107 2631
rect 31039 3205 31086 3307
rect 31221 3205 31281 3307
rect 31039 3188 31281 3205
rect 23498 2789 23732 2823
rect 23498 2699 23544 2789
rect 23707 2699 23732 2789
rect 23498 2668 23732 2699
rect 11716 2418 11871 2464
rect 5167 2330 5322 2376
rect 5167 2167 5198 2330
rect 5288 2167 5322 2330
rect 5167 2142 5322 2167
rect 6309 2328 6464 2374
rect 6309 2165 6340 2328
rect 6430 2165 6464 2328
rect 6309 2140 6464 2165
rect 11716 2255 11747 2418
rect 11837 2255 11871 2418
rect 11716 2230 11871 2255
rect 12858 2416 13013 2462
rect 12858 2253 12889 2416
rect 12979 2253 13013 2416
rect 24995 2418 25150 2464
rect 18370 2350 18525 2396
rect 12858 2228 13013 2253
rect 18370 2187 18401 2350
rect 18491 2187 18525 2350
rect 18370 2162 18525 2187
rect 19512 2348 19667 2394
rect 19512 2185 19543 2348
rect 19633 2185 19667 2348
rect 19512 2160 19667 2185
rect 24995 2255 25026 2418
rect 25116 2255 25150 2418
rect 24995 2230 25150 2255
rect 26137 2416 26292 2462
rect 26137 2253 26168 2416
rect 26258 2253 26292 2416
rect 26137 2228 26292 2253
rect 29023 1945 29235 1975
rect 29023 1889 29063 1945
rect 29197 1889 29235 1945
rect 29023 1867 29235 1889
rect 3684 1051 3918 1085
rect 3684 961 3730 1051
rect 3893 961 3918 1051
rect 10233 1139 10467 1173
rect 3684 930 3918 961
rect 500 178 712 208
rect 500 122 540 178
rect 674 122 712 178
rect 500 100 712 122
rect 10233 1049 10279 1139
rect 10442 1049 10467 1139
rect 10233 1018 10467 1049
rect 16887 1071 17121 1105
rect 16887 981 16933 1071
rect 17096 981 17121 1071
rect 23512 1139 23746 1173
rect 16887 950 17121 981
rect 3679 -553 3913 -519
rect 23512 1049 23558 1139
rect 23721 1049 23746 1139
rect 23512 1018 23746 1049
rect 10228 -465 10462 -431
rect 3679 -643 3725 -553
rect 3888 -643 3913 -553
rect 10228 -555 10274 -465
rect 10437 -555 10462 -465
rect 10228 -586 10462 -555
rect 3679 -674 3913 -643
rect 11660 -625 11815 -579
rect 16882 -533 17116 -499
rect 32631 17 32843 47
rect 32631 -39 32671 17
rect 32805 -39 32843 17
rect 32631 -61 32843 -39
rect 23507 -465 23741 -431
rect 5111 -713 5266 -667
rect 5111 -876 5142 -713
rect 5232 -876 5266 -713
rect 11660 -788 11691 -625
rect 11781 -788 11815 -625
rect 16882 -623 16928 -533
rect 17091 -623 17116 -533
rect 23507 -555 23553 -465
rect 23716 -555 23741 -465
rect 23507 -586 23741 -555
rect 16882 -654 17116 -623
rect 24939 -625 25094 -579
rect 11660 -813 11815 -788
rect 18314 -693 18469 -647
rect 5111 -901 5266 -876
rect 18314 -856 18345 -693
rect 18435 -856 18469 -693
rect 24939 -788 24970 -625
rect 25060 -788 25094 -625
rect 24939 -813 25094 -788
rect 18314 -881 18469 -856
rect 31041 -784 31283 -772
rect 31041 -886 31088 -784
rect 31223 -886 31283 -784
rect 31041 -903 31283 -886
rect 29023 -1088 29235 -1058
rect 29023 -1144 29063 -1088
rect 29197 -1144 29235 -1088
rect 29023 -1166 29235 -1144
rect 481 -3100 693 -3070
rect 481 -3156 521 -3100
rect 655 -3156 693 -3100
rect 3662 -3079 3896 -3045
rect 481 -3178 693 -3156
rect 3662 -3169 3708 -3079
rect 3871 -3169 3896 -3079
rect 3662 -3200 3896 -3169
rect 10213 -3081 10447 -3047
rect 10213 -3171 10259 -3081
rect 10422 -3171 10447 -3081
rect 10213 -3202 10447 -3171
rect 16868 -3080 17102 -3046
rect 16868 -3170 16914 -3080
rect 17077 -3170 17102 -3080
rect 16868 -3201 17102 -3170
rect 29094 -3008 29306 -2978
rect 23490 -3079 23724 -3045
rect 23490 -3169 23536 -3079
rect 23699 -3169 23724 -3079
rect 23490 -3200 23724 -3169
rect 29094 -3064 29134 -3008
rect 29268 -3064 29306 -3008
rect 29094 -3086 29306 -3064
rect 5159 -3450 5314 -3404
rect 5159 -3613 5190 -3450
rect 5280 -3613 5314 -3450
rect 5159 -3638 5314 -3613
rect 6301 -3452 6456 -3406
rect 6301 -3615 6332 -3452
rect 6422 -3615 6456 -3452
rect 11710 -3452 11865 -3406
rect 6301 -3640 6456 -3615
rect 11710 -3615 11741 -3452
rect 11831 -3615 11865 -3452
rect 11710 -3640 11865 -3615
rect 12852 -3454 13007 -3408
rect 12852 -3617 12883 -3454
rect 12973 -3617 13007 -3454
rect 18365 -3451 18520 -3405
rect 12852 -3642 13007 -3617
rect 18365 -3614 18396 -3451
rect 18486 -3614 18520 -3451
rect 18365 -3639 18520 -3614
rect 19507 -3453 19662 -3407
rect 19507 -3616 19538 -3453
rect 19628 -3616 19662 -3453
rect 24987 -3450 25142 -3404
rect 19507 -3641 19662 -3616
rect 24987 -3613 25018 -3450
rect 25108 -3613 25142 -3450
rect 24987 -3638 25142 -3613
rect 26129 -3452 26284 -3406
rect 26129 -3615 26160 -3452
rect 26250 -3615 26284 -3452
rect 26129 -3640 26284 -3615
rect 32631 -3478 32843 -3448
rect 32631 -3534 32671 -3478
rect 32805 -3534 32843 -3478
rect 32631 -3556 32843 -3534
rect 3676 -4729 3910 -4695
rect 3676 -4819 3722 -4729
rect 3885 -4819 3910 -4729
rect 3676 -4850 3910 -4819
rect 497 -5860 709 -5830
rect 497 -5916 537 -5860
rect 671 -5916 709 -5860
rect 497 -5938 709 -5916
rect 10227 -4731 10461 -4697
rect 10227 -4821 10273 -4731
rect 10436 -4821 10461 -4731
rect 10227 -4852 10461 -4821
rect 16882 -4730 17116 -4696
rect 16882 -4820 16928 -4730
rect 17091 -4820 17116 -4730
rect 31041 -4279 31283 -4267
rect 16882 -4851 17116 -4820
rect 3671 -6333 3905 -6299
rect 3671 -6423 3717 -6333
rect 3880 -6423 3905 -6333
rect 23504 -4729 23738 -4695
rect 23504 -4819 23550 -4729
rect 23713 -4819 23738 -4729
rect 31041 -4381 31088 -4279
rect 31223 -4381 31283 -4279
rect 31041 -4398 31283 -4381
rect 23504 -4850 23738 -4819
rect 10222 -6335 10456 -6301
rect 3671 -6454 3905 -6423
rect 5103 -6493 5258 -6447
rect 10222 -6425 10268 -6335
rect 10431 -6425 10456 -6335
rect 16877 -6334 17111 -6300
rect 10222 -6456 10456 -6425
rect 5103 -6656 5134 -6493
rect 5224 -6656 5258 -6493
rect 5103 -6681 5258 -6656
rect 11654 -6495 11809 -6449
rect 16877 -6424 16923 -6334
rect 17086 -6424 17111 -6334
rect 29091 -6078 29303 -6048
rect 29091 -6134 29131 -6078
rect 29265 -6134 29303 -6078
rect 29091 -6156 29303 -6134
rect 23499 -6333 23733 -6299
rect 16877 -6455 17111 -6424
rect 11654 -6658 11685 -6495
rect 11775 -6658 11809 -6495
rect 11654 -6683 11809 -6658
rect 18309 -6494 18464 -6448
rect 23499 -6423 23545 -6333
rect 23708 -6423 23733 -6333
rect 23499 -6454 23733 -6423
rect 18309 -6657 18340 -6494
rect 18430 -6657 18464 -6494
rect 18309 -6682 18464 -6657
rect 24931 -6493 25086 -6447
rect 24931 -6656 24962 -6493
rect 25052 -6656 25086 -6493
rect 24931 -6681 25086 -6656
rect 7207 -7225 7419 -7203
rect 7207 -7281 7247 -7225
rect 7381 -7281 7419 -7225
rect 7207 -7311 7419 -7281
rect 13761 -7220 13973 -7198
rect 13761 -7276 13801 -7220
rect 13935 -7276 13973 -7220
rect 13761 -7306 13973 -7276
rect 20410 -7232 20622 -7210
rect 20410 -7288 20450 -7232
rect 20584 -7288 20622 -7232
rect 20410 -7318 20622 -7288
rect 32631 -7826 32843 -7796
rect 32631 -7882 32671 -7826
rect 32805 -7882 32843 -7826
rect 32631 -7904 32843 -7882
rect 31041 -8627 31283 -8615
rect 31041 -8729 31088 -8627
rect 31223 -8729 31283 -8627
rect 31041 -8746 31283 -8729
rect 29098 -8923 29310 -8893
rect 29098 -8979 29138 -8923
rect 29272 -8979 29310 -8923
rect 29098 -9001 29310 -8979
<< nsubdiff >>
rect 6932 5871 7176 5909
rect 6932 5801 6988 5871
rect 7124 5801 7176 5871
rect 6932 5779 7176 5801
rect 13481 5870 13725 5908
rect 13481 5800 13537 5870
rect 13673 5800 13725 5870
rect 13481 5778 13725 5800
rect 20135 5891 20379 5929
rect 20135 5821 20191 5891
rect 20327 5821 20379 5891
rect 20135 5799 20379 5821
rect 30981 5783 31402 5817
rect 28788 5724 29032 5762
rect 28788 5654 28844 5724
rect 28980 5654 29032 5724
rect 28788 5632 29032 5654
rect 30981 5638 31044 5783
rect 31353 5638 31402 5783
rect 30981 5617 31402 5638
rect 32389 5316 32633 5354
rect 32389 5246 32445 5316
rect 32581 5246 32633 5316
rect 32389 5224 32633 5246
rect 12371 4020 12524 4060
rect 268 3971 512 4009
rect 268 3901 324 3971
rect 460 3901 512 3971
rect 5822 3932 5975 3972
rect 268 3879 512 3901
rect 3340 3878 3493 3918
rect 3340 3729 3383 3878
rect 3450 3729 3493 3878
rect 3340 3660 3493 3729
rect 5822 3783 5865 3932
rect 5932 3783 5975 3932
rect 5822 3714 5975 3783
rect 6969 3932 7122 3972
rect 6969 3783 7012 3932
rect 7079 3783 7122 3932
rect 6969 3714 7122 3783
rect 9889 3966 10042 4006
rect 9889 3817 9932 3966
rect 9999 3817 10042 3966
rect 9889 3748 10042 3817
rect 12371 3871 12414 4020
rect 12481 3871 12524 4020
rect 12371 3802 12524 3871
rect 13518 4020 13671 4060
rect 13518 3871 13561 4020
rect 13628 3871 13671 4020
rect 25650 4020 25803 4060
rect 19025 3952 19178 3992
rect 13518 3802 13671 3871
rect 16543 3898 16696 3938
rect 16543 3749 16586 3898
rect 16653 3749 16696 3898
rect 16543 3680 16696 3749
rect 19025 3803 19068 3952
rect 19135 3803 19178 3952
rect 19025 3734 19178 3803
rect 20172 3952 20325 3992
rect 20172 3803 20215 3952
rect 20282 3803 20325 3952
rect 20172 3734 20325 3803
rect 23168 3966 23321 4006
rect 23168 3817 23211 3966
rect 23278 3817 23321 3966
rect 23168 3748 23321 3817
rect 25650 3871 25693 4020
rect 25760 3871 25803 4020
rect 25650 3802 25803 3871
rect 26797 4020 26950 4060
rect 26797 3871 26840 4020
rect 26907 3871 26950 4020
rect 26797 3802 26950 3871
rect 28783 3153 29027 3191
rect 28783 3083 28839 3153
rect 28975 3083 29027 3153
rect 28783 3061 29027 3083
rect 3354 2228 3507 2268
rect 3354 2079 3397 2228
rect 3464 2079 3507 2228
rect 9903 2316 10056 2356
rect 9903 2167 9946 2316
rect 10013 2167 10056 2316
rect 16557 2248 16710 2288
rect 9903 2098 10056 2167
rect 16557 2099 16600 2248
rect 16667 2099 16710 2248
rect 23182 2316 23335 2356
rect 23182 2167 23225 2316
rect 23292 2167 23335 2316
rect 3354 2010 3507 2079
rect 16557 2030 16710 2099
rect 23182 2098 23335 2167
rect 13614 1973 13767 2013
rect 7065 1885 7218 1925
rect 7065 1736 7108 1885
rect 7175 1736 7218 1885
rect 7065 1667 7218 1736
rect 13614 1824 13657 1973
rect 13724 1824 13767 1973
rect 26893 1973 27046 2013
rect 20268 1905 20421 1945
rect 13614 1755 13767 1824
rect 260 1386 504 1424
rect 20268 1756 20311 1905
rect 20378 1756 20421 1905
rect 20268 1687 20421 1756
rect 26893 1824 26936 1973
rect 27003 1824 27046 1973
rect 26893 1755 27046 1824
rect 260 1316 316 1386
rect 452 1316 504 1386
rect 260 1294 504 1316
rect 3349 624 3502 664
rect 3349 475 3392 624
rect 3459 475 3502 624
rect 3349 406 3502 475
rect 30983 1692 31404 1726
rect 30983 1547 31046 1692
rect 31355 1547 31404 1692
rect 30983 1526 31404 1547
rect 9898 712 10051 752
rect 9898 563 9941 712
rect 10008 563 10051 712
rect 9898 494 10051 563
rect 16552 644 16705 684
rect 16552 495 16595 644
rect 16662 495 16705 644
rect 16552 426 16705 495
rect 32391 1225 32635 1263
rect 23177 712 23330 752
rect 23177 563 23220 712
rect 23287 563 23330 712
rect 23177 494 23330 563
rect 32391 1155 32447 1225
rect 32583 1155 32635 1225
rect 32391 1133 32635 1155
rect 28783 120 29027 158
rect 28783 50 28839 120
rect 28975 50 29027 120
rect 28783 28 29027 50
rect 28854 -1800 29098 -1762
rect 5814 -1848 5967 -1808
rect 241 -1892 485 -1854
rect 241 -1962 297 -1892
rect 433 -1962 485 -1892
rect 241 -1984 485 -1962
rect 3332 -1902 3485 -1862
rect 3332 -2051 3375 -1902
rect 3442 -2051 3485 -1902
rect 3332 -2120 3485 -2051
rect 5814 -1997 5857 -1848
rect 5924 -1997 5967 -1848
rect 5814 -2066 5967 -1997
rect 6961 -1848 7114 -1808
rect 6961 -1997 7004 -1848
rect 7071 -1997 7114 -1848
rect 12365 -1850 12518 -1810
rect 6961 -2066 7114 -1997
rect 9883 -1904 10036 -1864
rect 9883 -2053 9926 -1904
rect 9993 -2053 10036 -1904
rect 9883 -2122 10036 -2053
rect 12365 -1999 12408 -1850
rect 12475 -1999 12518 -1850
rect 12365 -2068 12518 -1999
rect 13512 -1850 13665 -1810
rect 13512 -1999 13555 -1850
rect 13622 -1999 13665 -1850
rect 19020 -1849 19173 -1809
rect 13512 -2068 13665 -1999
rect 16538 -1903 16691 -1863
rect 16538 -2052 16581 -1903
rect 16648 -2052 16691 -1903
rect 16538 -2121 16691 -2052
rect 19020 -1998 19063 -1849
rect 19130 -1998 19173 -1849
rect 19020 -2067 19173 -1998
rect 20167 -1849 20320 -1809
rect 20167 -1998 20210 -1849
rect 20277 -1998 20320 -1849
rect 25642 -1848 25795 -1808
rect 20167 -2067 20320 -1998
rect 23160 -1902 23313 -1862
rect 23160 -2051 23203 -1902
rect 23270 -2051 23313 -1902
rect 23160 -2120 23313 -2051
rect 25642 -1997 25685 -1848
rect 25752 -1997 25795 -1848
rect 25642 -2066 25795 -1997
rect 26789 -1848 26942 -1808
rect 26789 -1997 26832 -1848
rect 26899 -1997 26942 -1848
rect 28854 -1870 28910 -1800
rect 29046 -1870 29098 -1800
rect 28854 -1892 29098 -1870
rect 30983 -1803 31404 -1769
rect 30983 -1948 31046 -1803
rect 31355 -1948 31404 -1803
rect 30983 -1969 31404 -1948
rect 26789 -2066 26942 -1997
rect 32391 -2270 32635 -2232
rect 32391 -2340 32447 -2270
rect 32583 -2340 32635 -2270
rect 32391 -2362 32635 -2340
rect 3346 -3552 3499 -3512
rect 3346 -3701 3389 -3552
rect 3456 -3701 3499 -3552
rect 9897 -3554 10050 -3514
rect 3346 -3770 3499 -3701
rect 9897 -3703 9940 -3554
rect 10007 -3703 10050 -3554
rect 16552 -3553 16705 -3513
rect 9897 -3772 10050 -3703
rect 16552 -3702 16595 -3553
rect 16662 -3702 16705 -3553
rect 23174 -3552 23327 -3512
rect 16552 -3771 16705 -3702
rect 23174 -3701 23217 -3552
rect 23284 -3701 23327 -3552
rect 23174 -3770 23327 -3701
rect 7057 -3895 7210 -3855
rect 7057 -4044 7100 -3895
rect 7167 -4044 7210 -3895
rect 13608 -3897 13761 -3857
rect 7057 -4113 7210 -4044
rect 13608 -4046 13651 -3897
rect 13718 -4046 13761 -3897
rect 20263 -3896 20416 -3856
rect 13608 -4115 13761 -4046
rect 20263 -4045 20306 -3896
rect 20373 -4045 20416 -3896
rect 26885 -3895 27038 -3855
rect 20263 -4114 20416 -4045
rect 26885 -4044 26928 -3895
rect 26995 -4044 27038 -3895
rect 26885 -4113 27038 -4044
rect 257 -4652 501 -4614
rect 257 -4722 313 -4652
rect 449 -4722 501 -4652
rect 257 -4744 501 -4722
rect 3341 -5156 3494 -5116
rect 3341 -5305 3384 -5156
rect 3451 -5305 3494 -5156
rect 3341 -5374 3494 -5305
rect 9892 -5158 10045 -5118
rect 9892 -5307 9935 -5158
rect 10002 -5307 10045 -5158
rect 9892 -5376 10045 -5307
rect 16547 -5157 16700 -5117
rect 16547 -5306 16590 -5157
rect 16657 -5306 16700 -5157
rect 16547 -5375 16700 -5306
rect 23169 -5156 23322 -5116
rect 23169 -5305 23212 -5156
rect 23279 -5305 23322 -5156
rect 23169 -5374 23322 -5305
rect 28851 -4870 29095 -4832
rect 28851 -4940 28907 -4870
rect 29043 -4940 29095 -4870
rect 28851 -4962 29095 -4940
rect 30983 -6151 31404 -6117
rect 30983 -6296 31046 -6151
rect 31355 -6296 31404 -6151
rect 30983 -6317 31404 -6296
rect 32391 -6618 32635 -6580
rect 32391 -6688 32447 -6618
rect 32583 -6688 32635 -6618
rect 32391 -6710 32635 -6688
rect 28858 -7715 29102 -7677
rect 28858 -7785 28914 -7715
rect 29050 -7785 29102 -7715
rect 28858 -7807 29102 -7785
rect 6967 -8419 7211 -8397
rect 6967 -8489 7023 -8419
rect 7159 -8489 7211 -8419
rect 6967 -8527 7211 -8489
rect 13521 -8414 13765 -8392
rect 13521 -8484 13577 -8414
rect 13713 -8484 13765 -8414
rect 13521 -8522 13765 -8484
rect 20170 -8426 20414 -8404
rect 20170 -8496 20226 -8426
rect 20362 -8496 20414 -8426
rect 20170 -8534 20414 -8496
<< psubdiffcont >>
rect 7212 4607 7346 4663
rect 13761 4606 13895 4662
rect 20415 4627 20549 4683
rect 29068 4460 29202 4516
rect 32669 4052 32803 4108
rect 548 2707 682 2763
rect 3716 2611 3879 2701
rect 10265 2699 10428 2789
rect 16919 2631 17082 2721
rect 31086 3205 31221 3307
rect 23544 2699 23707 2789
rect 5198 2167 5288 2330
rect 6340 2165 6430 2328
rect 11747 2255 11837 2418
rect 12889 2253 12979 2416
rect 18401 2187 18491 2350
rect 19543 2185 19633 2348
rect 25026 2255 25116 2418
rect 26168 2253 26258 2416
rect 29063 1889 29197 1945
rect 3730 961 3893 1051
rect 540 122 674 178
rect 10279 1049 10442 1139
rect 16933 981 17096 1071
rect 23558 1049 23721 1139
rect 3725 -643 3888 -553
rect 10274 -555 10437 -465
rect 32671 -39 32805 17
rect 5142 -876 5232 -713
rect 11691 -788 11781 -625
rect 16928 -623 17091 -533
rect 23553 -555 23716 -465
rect 18345 -856 18435 -693
rect 24970 -788 25060 -625
rect 31088 -886 31223 -784
rect 29063 -1144 29197 -1088
rect 521 -3156 655 -3100
rect 3708 -3169 3871 -3079
rect 10259 -3171 10422 -3081
rect 16914 -3170 17077 -3080
rect 23536 -3169 23699 -3079
rect 29134 -3064 29268 -3008
rect 5190 -3613 5280 -3450
rect 6332 -3615 6422 -3452
rect 11741 -3615 11831 -3452
rect 12883 -3617 12973 -3454
rect 18396 -3614 18486 -3451
rect 19538 -3616 19628 -3453
rect 25018 -3613 25108 -3450
rect 26160 -3615 26250 -3452
rect 32671 -3534 32805 -3478
rect 3722 -4819 3885 -4729
rect 537 -5916 671 -5860
rect 10273 -4821 10436 -4731
rect 16928 -4820 17091 -4730
rect 3717 -6423 3880 -6333
rect 23550 -4819 23713 -4729
rect 31088 -4381 31223 -4279
rect 10268 -6425 10431 -6335
rect 5134 -6656 5224 -6493
rect 16923 -6424 17086 -6334
rect 29131 -6134 29265 -6078
rect 11685 -6658 11775 -6495
rect 23545 -6423 23708 -6333
rect 18340 -6657 18430 -6494
rect 24962 -6656 25052 -6493
rect 7247 -7281 7381 -7225
rect 13801 -7276 13935 -7220
rect 20450 -7288 20584 -7232
rect 32671 -7882 32805 -7826
rect 31088 -8729 31223 -8627
rect 29138 -8979 29272 -8923
<< nsubdiffcont >>
rect 6988 5801 7124 5871
rect 13537 5800 13673 5870
rect 20191 5821 20327 5891
rect 28844 5654 28980 5724
rect 31044 5638 31353 5783
rect 32445 5246 32581 5316
rect 324 3901 460 3971
rect 3383 3729 3450 3878
rect 5865 3783 5932 3932
rect 7012 3783 7079 3932
rect 9932 3817 9999 3966
rect 12414 3871 12481 4020
rect 13561 3871 13628 4020
rect 16586 3749 16653 3898
rect 19068 3803 19135 3952
rect 20215 3803 20282 3952
rect 23211 3817 23278 3966
rect 25693 3871 25760 4020
rect 26840 3871 26907 4020
rect 28839 3083 28975 3153
rect 3397 2079 3464 2228
rect 9946 2167 10013 2316
rect 16600 2099 16667 2248
rect 23225 2167 23292 2316
rect 7108 1736 7175 1885
rect 13657 1824 13724 1973
rect 20311 1756 20378 1905
rect 26936 1824 27003 1973
rect 316 1316 452 1386
rect 3392 475 3459 624
rect 31046 1547 31355 1692
rect 9941 563 10008 712
rect 16595 495 16662 644
rect 23220 563 23287 712
rect 32447 1155 32583 1225
rect 28839 50 28975 120
rect 297 -1962 433 -1892
rect 3375 -2051 3442 -1902
rect 5857 -1997 5924 -1848
rect 7004 -1997 7071 -1848
rect 9926 -2053 9993 -1904
rect 12408 -1999 12475 -1850
rect 13555 -1999 13622 -1850
rect 16581 -2052 16648 -1903
rect 19063 -1998 19130 -1849
rect 20210 -1998 20277 -1849
rect 23203 -2051 23270 -1902
rect 25685 -1997 25752 -1848
rect 26832 -1997 26899 -1848
rect 28910 -1870 29046 -1800
rect 31046 -1948 31355 -1803
rect 32447 -2340 32583 -2270
rect 3389 -3701 3456 -3552
rect 9940 -3703 10007 -3554
rect 16595 -3702 16662 -3553
rect 23217 -3701 23284 -3552
rect 7100 -4044 7167 -3895
rect 13651 -4046 13718 -3897
rect 20306 -4045 20373 -3896
rect 26928 -4044 26995 -3895
rect 313 -4722 449 -4652
rect 3384 -5305 3451 -5156
rect 9935 -5307 10002 -5158
rect 16590 -5306 16657 -5157
rect 23212 -5305 23279 -5156
rect 28907 -4940 29043 -4870
rect 31046 -6296 31355 -6151
rect 32447 -6688 32583 -6618
rect 28914 -7785 29050 -7715
rect 7023 -8489 7159 -8419
rect 13577 -8484 13713 -8414
rect 20226 -8496 20362 -8426
<< poly >>
rect 6729 5664 7025 5700
rect 6729 5643 6789 5664
rect 6847 5643 6907 5664
rect 6965 5643 7025 5664
rect 7083 5663 7379 5699
rect 7083 5643 7143 5663
rect 7201 5643 7261 5663
rect 7319 5643 7379 5663
rect 7437 5663 7733 5699
rect 7437 5643 7497 5663
rect 7555 5643 7615 5663
rect 7673 5643 7733 5663
rect 13278 5663 13574 5699
rect 13278 5642 13338 5663
rect 13396 5642 13456 5663
rect 13514 5642 13574 5663
rect 13632 5662 13928 5698
rect 13632 5642 13692 5662
rect 13750 5642 13810 5662
rect 13868 5642 13928 5662
rect 13986 5662 14282 5698
rect 19932 5684 20228 5720
rect 19932 5663 19992 5684
rect 20050 5663 20110 5684
rect 20168 5663 20228 5684
rect 20286 5683 20582 5719
rect 20286 5663 20346 5683
rect 20404 5663 20464 5683
rect 20522 5663 20582 5683
rect 20640 5683 20936 5719
rect 20640 5663 20700 5683
rect 20758 5663 20818 5683
rect 20876 5663 20936 5683
rect 13986 5642 14046 5662
rect 14104 5642 14164 5662
rect 14222 5642 14282 5662
rect 6729 5417 6789 5443
rect 6847 5417 6907 5443
rect 6965 5417 7025 5443
rect 7083 5423 7143 5443
rect 7083 5417 7144 5423
rect 7201 5417 7261 5443
rect 7319 5417 7379 5443
rect 6966 5232 7024 5417
rect 6966 5206 7026 5232
rect 7084 5206 7144 5417
rect 7437 5411 7497 5443
rect 7555 5417 7615 5443
rect 7673 5417 7733 5443
rect 28585 5517 28881 5553
rect 28585 5496 28645 5517
rect 28703 5496 28763 5517
rect 28821 5496 28881 5517
rect 28939 5516 29235 5552
rect 28939 5496 28999 5516
rect 29057 5496 29117 5516
rect 29175 5496 29235 5516
rect 29293 5516 29589 5552
rect 29293 5496 29353 5516
rect 29411 5496 29471 5516
rect 29529 5496 29589 5516
rect 13278 5416 13338 5442
rect 13396 5416 13456 5442
rect 13514 5416 13574 5442
rect 13632 5422 13692 5442
rect 13632 5416 13693 5422
rect 13750 5416 13810 5442
rect 13868 5416 13928 5442
rect 7434 5395 7500 5411
rect 7434 5361 7450 5395
rect 7484 5361 7500 5395
rect 7434 5345 7500 5361
rect 7316 5278 7382 5294
rect 7316 5244 7332 5278
rect 7366 5244 7382 5278
rect 7316 5228 7382 5244
rect 13515 5231 13573 5416
rect 7319 5206 7379 5228
rect 13515 5205 13575 5231
rect 13633 5205 13693 5416
rect 13986 5410 14046 5442
rect 14104 5416 14164 5442
rect 14222 5416 14282 5442
rect 19932 5437 19992 5463
rect 20050 5437 20110 5463
rect 20168 5437 20228 5463
rect 20286 5443 20346 5463
rect 20286 5437 20347 5443
rect 20404 5437 20464 5463
rect 20522 5437 20582 5463
rect 13983 5394 14049 5410
rect 13983 5360 13999 5394
rect 14033 5360 14049 5394
rect 13983 5344 14049 5360
rect 13865 5277 13931 5293
rect 13865 5243 13881 5277
rect 13915 5243 13931 5277
rect 13865 5227 13931 5243
rect 20169 5252 20227 5437
rect 13868 5205 13928 5227
rect 20169 5226 20229 5252
rect 20287 5226 20347 5437
rect 20640 5431 20700 5463
rect 20758 5437 20818 5463
rect 20876 5437 20936 5463
rect 20637 5415 20703 5431
rect 20637 5381 20653 5415
rect 20687 5381 20703 5415
rect 20637 5365 20703 5381
rect 20519 5298 20585 5314
rect 20519 5264 20535 5298
rect 20569 5264 20585 5298
rect 30877 5306 31173 5357
rect 28585 5270 28645 5296
rect 28703 5270 28763 5296
rect 28821 5270 28881 5296
rect 28939 5276 28999 5296
rect 28939 5270 29000 5276
rect 29057 5270 29117 5296
rect 29175 5270 29235 5296
rect 20519 5248 20585 5264
rect 20522 5226 20582 5248
rect 7319 4980 7379 5006
rect 6966 4784 7026 4806
rect 7084 4784 7144 4806
rect 13868 4979 13928 5005
rect 28822 5085 28880 5270
rect 28822 5059 28882 5085
rect 28940 5059 29000 5270
rect 29293 5264 29353 5296
rect 29411 5270 29471 5296
rect 29529 5270 29589 5296
rect 30877 5291 30937 5306
rect 30995 5291 31055 5306
rect 31113 5291 31173 5306
rect 31231 5291 31291 5317
rect 31349 5291 31409 5317
rect 31467 5291 31527 5317
rect 29290 5248 29356 5264
rect 29290 5214 29306 5248
rect 29340 5214 29356 5248
rect 29290 5198 29356 5214
rect 29172 5131 29238 5147
rect 29172 5097 29188 5131
rect 29222 5097 29238 5131
rect 29172 5081 29238 5097
rect 30393 5091 30453 5117
rect 30511 5091 30571 5117
rect 30629 5091 30689 5117
rect 29175 5059 29235 5081
rect 20522 5000 20582 5026
rect 6963 4768 7029 4784
rect 6963 4734 6979 4768
rect 7013 4734 7029 4768
rect 6963 4718 7029 4734
rect 7081 4768 7147 4784
rect 13515 4783 13575 4805
rect 13633 4783 13693 4805
rect 20169 4804 20229 4826
rect 20287 4804 20347 4826
rect 20166 4788 20232 4804
rect 7081 4734 7097 4768
rect 7131 4734 7147 4768
rect 7081 4718 7147 4734
rect 13512 4767 13578 4783
rect 13512 4733 13528 4767
rect 13562 4733 13578 4767
rect 13512 4717 13578 4733
rect 13630 4767 13696 4783
rect 13630 4733 13646 4767
rect 13680 4733 13696 4767
rect 20166 4754 20182 4788
rect 20216 4754 20232 4788
rect 20166 4738 20232 4754
rect 20284 4788 20350 4804
rect 20284 4754 20300 4788
rect 20334 4754 20350 4788
rect 20284 4738 20350 4754
rect 13630 4717 13696 4733
rect 31714 5108 32010 5159
rect 31714 5091 31774 5108
rect 31832 5091 31892 5108
rect 31950 5091 32010 5108
rect 32186 5109 32482 5145
rect 32186 5088 32246 5109
rect 32304 5088 32364 5109
rect 32422 5088 32482 5109
rect 32540 5108 32836 5144
rect 32540 5088 32600 5108
rect 32658 5088 32718 5108
rect 32776 5088 32836 5108
rect 32894 5108 33190 5144
rect 32894 5088 32954 5108
rect 33012 5088 33072 5108
rect 33130 5088 33190 5108
rect 30393 4874 30453 4891
rect 30511 4874 30571 4891
rect 30629 4874 30689 4891
rect 30877 4874 30937 4891
rect 29175 4833 29235 4859
rect 30393 4823 30937 4874
rect 30995 4865 31055 4891
rect 31113 4865 31173 4891
rect 31231 4872 31291 4891
rect 31349 4872 31409 4891
rect 31467 4872 31527 4891
rect 31714 4872 31774 4891
rect 31832 4872 31892 4891
rect 28822 4637 28882 4659
rect 28940 4637 29000 4659
rect 28819 4621 28885 4637
rect 28819 4587 28835 4621
rect 28869 4587 28885 4621
rect 28819 4571 28885 4587
rect 28937 4621 29003 4637
rect 28937 4587 28953 4621
rect 28987 4587 29003 4621
rect 28937 4571 29003 4587
rect 30518 4619 30578 4823
rect 31231 4821 31774 4872
rect 31816 4865 31892 4872
rect 31950 4865 32010 4891
rect 31816 4821 31891 4865
rect 32186 4862 32246 4888
rect 32304 4862 32364 4888
rect 32422 4862 32482 4888
rect 32540 4868 32600 4888
rect 32540 4862 32601 4868
rect 32658 4862 32718 4888
rect 32776 4862 32836 4888
rect 31816 4739 31876 4821
rect 31816 4721 32050 4739
rect 31816 4687 31999 4721
rect 32033 4687 32050 4721
rect 30820 4621 31116 4681
rect 30518 4602 30649 4619
rect 30518 4568 30599 4602
rect 30633 4568 30649 4602
rect 30820 4598 30880 4621
rect 30938 4598 30998 4621
rect 31056 4598 31116 4621
rect 31174 4622 31470 4682
rect 31174 4598 31234 4622
rect 31292 4598 31352 4622
rect 31410 4598 31470 4622
rect 31816 4671 32050 4687
rect 32423 4677 32481 4862
rect 30518 4551 30649 4568
rect 65 3764 361 3800
rect 65 3743 125 3764
rect 183 3743 243 3764
rect 301 3743 361 3764
rect 419 3763 715 3799
rect 419 3743 479 3763
rect 537 3743 597 3763
rect 655 3743 715 3763
rect 773 3763 1069 3799
rect 773 3743 833 3763
rect 891 3743 951 3763
rect 1009 3743 1069 3763
rect 5103 3712 5169 3728
rect 6233 3718 6299 3734
rect 5103 3678 5119 3712
rect 5153 3705 5169 3712
rect 5153 3678 5678 3705
rect 5103 3662 5678 3678
rect 6233 3684 6249 3718
rect 6283 3709 6299 3718
rect 11652 3800 11718 3816
rect 12782 3806 12848 3822
rect 11652 3766 11668 3800
rect 11702 3793 11718 3800
rect 11702 3766 12227 3793
rect 11652 3750 12227 3766
rect 12782 3772 12798 3806
rect 12832 3797 12848 3806
rect 12832 3772 13369 3797
rect 12782 3754 13369 3772
rect 6283 3684 6820 3709
rect 12183 3698 12227 3750
rect 13325 3702 13369 3754
rect 6233 3666 6820 3684
rect 5634 3610 5678 3662
rect 6776 3614 6820 3666
rect 11652 3682 12125 3698
rect 11652 3648 11668 3682
rect 11702 3657 12125 3682
rect 11702 3656 11889 3657
rect 11702 3648 11718 3656
rect 11652 3632 11718 3648
rect 11829 3636 11889 3656
rect 11947 3636 12007 3657
rect 12065 3636 12125 3657
rect 12183 3657 12479 3698
rect 12183 3636 12243 3657
rect 12301 3636 12361 3657
rect 12419 3636 12479 3657
rect 12782 3686 13267 3702
rect 12782 3652 12798 3686
rect 12832 3661 13267 3686
rect 12832 3660 13031 3661
rect 12832 3652 12848 3660
rect 12782 3636 12848 3652
rect 12971 3640 13031 3660
rect 13089 3640 13149 3661
rect 13207 3640 13267 3661
rect 13325 3661 13621 3702
rect 18306 3732 18372 3748
rect 19436 3738 19502 3754
rect 18306 3698 18322 3732
rect 18356 3725 18372 3732
rect 18356 3698 18881 3725
rect 18306 3682 18881 3698
rect 19436 3704 19452 3738
rect 19486 3729 19502 3738
rect 24931 3800 24997 3816
rect 26061 3806 26127 3822
rect 24931 3766 24947 3800
rect 24981 3793 24997 3800
rect 24981 3766 25506 3793
rect 24931 3750 25506 3766
rect 26061 3772 26077 3806
rect 26111 3797 26127 3806
rect 30518 3971 30578 4551
rect 30820 4172 30880 4198
rect 30788 4031 30855 4038
rect 30938 4031 30998 4198
rect 31056 4172 31116 4198
rect 31174 4172 31234 4198
rect 30788 4022 30998 4031
rect 30788 3988 30804 4022
rect 30838 3988 30998 4022
rect 30788 3972 30998 3988
rect 30518 3955 30669 3971
rect 30518 3921 30619 3955
rect 30653 3921 30669 3955
rect 30518 3905 30669 3921
rect 30518 3866 30578 3905
rect 30938 3866 30998 3972
rect 31292 4031 31352 4198
rect 31410 4172 31470 4198
rect 31435 4031 31502 4038
rect 31292 4022 31502 4031
rect 31292 3988 31452 4022
rect 31486 3988 31502 4022
rect 31292 3972 31502 3988
rect 31054 3938 31120 3954
rect 31054 3904 31070 3938
rect 31104 3904 31120 3938
rect 31054 3888 31120 3904
rect 31172 3939 31238 3954
rect 31172 3905 31188 3939
rect 31222 3905 31238 3939
rect 31172 3889 31238 3905
rect 31056 3866 31116 3888
rect 31174 3866 31234 3889
rect 31292 3866 31352 3972
rect 31816 3970 31876 4671
rect 32423 4651 32483 4677
rect 32541 4651 32601 4862
rect 32894 4856 32954 4888
rect 33012 4862 33072 4888
rect 33130 4862 33190 4888
rect 32891 4840 32957 4856
rect 32891 4806 32907 4840
rect 32941 4806 32957 4840
rect 32891 4790 32957 4806
rect 32773 4723 32839 4739
rect 32773 4689 32789 4723
rect 32823 4689 32839 4723
rect 32773 4673 32839 4689
rect 32776 4651 32836 4673
rect 32776 4425 32836 4451
rect 32423 4229 32483 4251
rect 32541 4229 32601 4251
rect 32420 4213 32486 4229
rect 32420 4179 32436 4213
rect 32470 4179 32486 4213
rect 32420 4163 32486 4179
rect 32538 4213 32604 4229
rect 32538 4179 32554 4213
rect 32588 4179 32604 4213
rect 32538 4163 32604 4179
rect 31726 3954 31876 3970
rect 31726 3920 31742 3954
rect 31776 3920 31876 3954
rect 31726 3904 31876 3920
rect 31816 3866 31876 3904
rect 26111 3772 26648 3797
rect 26061 3754 26648 3772
rect 19486 3704 20023 3729
rect 19436 3686 20023 3704
rect 25462 3698 25506 3750
rect 26604 3702 26648 3754
rect 13325 3640 13385 3661
rect 13443 3640 13503 3661
rect 13561 3640 13621 3661
rect 5103 3594 5576 3610
rect 5103 3560 5119 3594
rect 5153 3569 5576 3594
rect 5153 3568 5340 3569
rect 5153 3560 5169 3568
rect 5103 3544 5169 3560
rect 5280 3548 5340 3568
rect 5398 3548 5458 3569
rect 5516 3548 5576 3569
rect 5634 3569 5930 3610
rect 5634 3548 5694 3569
rect 5752 3548 5812 3569
rect 5870 3548 5930 3569
rect 6233 3598 6718 3614
rect 6233 3564 6249 3598
rect 6283 3573 6718 3598
rect 6283 3572 6482 3573
rect 6283 3564 6299 3572
rect 6233 3548 6299 3564
rect 6422 3552 6482 3572
rect 6540 3552 6600 3573
rect 6658 3552 6718 3573
rect 6776 3573 7072 3614
rect 6776 3552 6836 3573
rect 6894 3552 6954 3573
rect 7012 3552 7072 3573
rect 9504 3585 9800 3621
rect 9504 3564 9564 3585
rect 9622 3564 9682 3585
rect 9740 3564 9800 3585
rect 9858 3584 10154 3620
rect 9858 3564 9918 3584
rect 9976 3564 10036 3584
rect 10094 3564 10154 3584
rect 10212 3584 10508 3620
rect 10212 3564 10272 3584
rect 10330 3564 10390 3584
rect 10448 3564 10508 3584
rect 65 3517 125 3543
rect 183 3517 243 3543
rect 301 3517 361 3543
rect 419 3523 479 3543
rect 419 3517 480 3523
rect 537 3517 597 3543
rect 655 3517 715 3543
rect 302 3332 360 3517
rect 302 3306 362 3332
rect 420 3306 480 3517
rect 773 3511 833 3543
rect 891 3517 951 3543
rect 1009 3517 1069 3543
rect 770 3495 836 3511
rect 770 3461 786 3495
rect 820 3461 836 3495
rect 2955 3497 3251 3533
rect 2955 3476 3015 3497
rect 3073 3476 3133 3497
rect 3191 3476 3251 3497
rect 3309 3496 3605 3532
rect 3309 3476 3369 3496
rect 3427 3476 3487 3496
rect 3545 3476 3605 3496
rect 3663 3496 3959 3532
rect 3663 3476 3723 3496
rect 3781 3476 3841 3496
rect 3899 3476 3959 3496
rect 770 3445 836 3461
rect 652 3378 718 3394
rect 652 3344 668 3378
rect 702 3344 718 3378
rect 652 3328 718 3344
rect 655 3306 715 3328
rect 2955 3250 3015 3276
rect 3073 3250 3133 3276
rect 3191 3250 3251 3276
rect 3309 3256 3369 3276
rect 3309 3250 3370 3256
rect 3427 3250 3487 3276
rect 3545 3250 3605 3276
rect 655 3080 715 3106
rect 3192 3065 3250 3250
rect 3192 3039 3252 3065
rect 3310 3039 3370 3250
rect 3663 3244 3723 3276
rect 3781 3250 3841 3276
rect 3899 3250 3959 3276
rect 3660 3228 3726 3244
rect 3660 3194 3676 3228
rect 3710 3194 3726 3228
rect 3660 3178 3726 3194
rect 9504 3338 9564 3364
rect 9622 3338 9682 3364
rect 9740 3338 9800 3364
rect 9858 3344 9918 3364
rect 9858 3338 9919 3344
rect 9976 3338 10036 3364
rect 10094 3338 10154 3364
rect 9741 3153 9799 3338
rect 5280 3131 5340 3148
rect 3542 3111 3608 3127
rect 3542 3077 3558 3111
rect 3592 3077 3608 3111
rect 3542 3061 3608 3077
rect 3545 3039 3605 3061
rect 5280 3042 5341 3131
rect 5398 3122 5458 3148
rect 5516 3122 5576 3148
rect 302 2884 362 2906
rect 420 2884 480 2906
rect 299 2868 365 2884
rect 299 2834 315 2868
rect 349 2834 365 2868
rect 299 2818 365 2834
rect 417 2868 483 2884
rect 417 2834 433 2868
rect 467 2834 483 2868
rect 417 2818 483 2834
rect 5190 2989 5341 3042
rect 3545 2813 3605 2839
rect 5190 2765 5250 2989
rect 5634 2947 5694 3148
rect 5752 3122 5812 3148
rect 5870 3122 5930 3148
rect 6422 3135 6482 3152
rect 6422 3046 6483 3135
rect 6540 3126 6600 3152
rect 6658 3126 6718 3152
rect 5308 2896 5694 2947
rect 6332 2993 6483 3046
rect 5308 2765 5368 2896
rect 5423 2838 5489 2854
rect 5423 2804 5439 2838
rect 5473 2804 5489 2838
rect 5423 2788 5489 2804
rect 5426 2765 5486 2788
rect 5709 2765 5769 2791
rect 5827 2765 5887 2791
rect 5945 2765 6005 2791
rect 6332 2769 6392 2993
rect 6776 2951 6836 3152
rect 6894 3126 6954 3152
rect 7012 3126 7072 3152
rect 9741 3127 9801 3153
rect 9859 3127 9919 3338
rect 10212 3332 10272 3364
rect 10330 3338 10390 3364
rect 10448 3338 10508 3364
rect 10209 3316 10275 3332
rect 10209 3282 10225 3316
rect 10259 3282 10275 3316
rect 10209 3266 10275 3282
rect 18837 3630 18881 3682
rect 19979 3634 20023 3686
rect 24931 3682 25404 3698
rect 24931 3648 24947 3682
rect 24981 3657 25404 3682
rect 24981 3656 25168 3657
rect 24981 3648 24997 3656
rect 18306 3614 18779 3630
rect 18306 3580 18322 3614
rect 18356 3589 18779 3614
rect 18356 3588 18543 3589
rect 18356 3580 18372 3588
rect 18306 3564 18372 3580
rect 18483 3568 18543 3588
rect 18601 3568 18661 3589
rect 18719 3568 18779 3589
rect 18837 3589 19133 3630
rect 18837 3568 18897 3589
rect 18955 3568 19015 3589
rect 19073 3568 19133 3589
rect 19436 3618 19921 3634
rect 19436 3584 19452 3618
rect 19486 3593 19921 3618
rect 19486 3592 19685 3593
rect 19486 3584 19502 3592
rect 19436 3568 19502 3584
rect 19625 3572 19685 3592
rect 19743 3572 19803 3593
rect 19861 3572 19921 3593
rect 19979 3593 20275 3634
rect 24931 3632 24997 3648
rect 25108 3636 25168 3656
rect 25226 3636 25286 3657
rect 25344 3636 25404 3657
rect 25462 3657 25758 3698
rect 25462 3636 25522 3657
rect 25580 3636 25640 3657
rect 25698 3636 25758 3657
rect 26061 3686 26546 3702
rect 26061 3652 26077 3686
rect 26111 3661 26546 3686
rect 26111 3660 26310 3661
rect 26111 3652 26127 3660
rect 26061 3636 26127 3652
rect 26250 3640 26310 3660
rect 26368 3640 26428 3661
rect 26486 3640 26546 3661
rect 26604 3661 26900 3702
rect 26604 3640 26664 3661
rect 26722 3640 26782 3661
rect 26840 3640 26900 3661
rect 30518 3640 30578 3666
rect 19979 3572 20039 3593
rect 20097 3572 20157 3593
rect 20215 3572 20275 3593
rect 22783 3585 23079 3621
rect 16158 3517 16454 3553
rect 16158 3496 16218 3517
rect 16276 3496 16336 3517
rect 16394 3496 16454 3517
rect 16512 3516 16808 3552
rect 16512 3496 16572 3516
rect 16630 3496 16690 3516
rect 16748 3496 16808 3516
rect 16866 3516 17162 3552
rect 16866 3496 16926 3516
rect 16984 3496 17044 3516
rect 17102 3496 17162 3516
rect 16158 3270 16218 3296
rect 16276 3270 16336 3296
rect 16394 3270 16454 3296
rect 16512 3276 16572 3296
rect 16512 3270 16573 3276
rect 16630 3270 16690 3296
rect 16748 3270 16808 3296
rect 11829 3219 11889 3236
rect 10091 3199 10157 3215
rect 10091 3165 10107 3199
rect 10141 3165 10157 3199
rect 10091 3149 10157 3165
rect 10094 3127 10154 3149
rect 11829 3130 11890 3219
rect 11947 3210 12007 3236
rect 12065 3210 12125 3236
rect 6450 2900 6836 2951
rect 6450 2769 6510 2900
rect 6565 2842 6631 2858
rect 6565 2808 6581 2842
rect 6615 2808 6631 2842
rect 6565 2792 6631 2808
rect 6568 2769 6628 2792
rect 6851 2769 6911 2795
rect 6969 2769 7029 2795
rect 7087 2769 7147 2795
rect 3192 2617 3252 2639
rect 3310 2617 3370 2639
rect 3189 2601 3255 2617
rect 3189 2567 3205 2601
rect 3239 2567 3255 2601
rect 3189 2551 3255 2567
rect 3307 2601 3373 2617
rect 3307 2567 3323 2601
rect 3357 2567 3373 2601
rect 3307 2551 3373 2567
rect 11739 3077 11890 3130
rect 10094 2901 10154 2927
rect 11739 2853 11799 3077
rect 12183 3035 12243 3236
rect 12301 3210 12361 3236
rect 12419 3210 12479 3236
rect 12971 3223 13031 3240
rect 12971 3134 13032 3223
rect 13089 3214 13149 3240
rect 13207 3214 13267 3240
rect 11857 2984 12243 3035
rect 12881 3081 13032 3134
rect 11857 2853 11917 2984
rect 11972 2926 12038 2942
rect 11972 2892 11988 2926
rect 12022 2892 12038 2926
rect 11972 2876 12038 2892
rect 11975 2853 12035 2876
rect 12258 2853 12318 2879
rect 12376 2853 12436 2879
rect 12494 2853 12554 2879
rect 12881 2857 12941 3081
rect 13325 3039 13385 3240
rect 13443 3214 13503 3240
rect 13561 3214 13621 3240
rect 16395 3085 16453 3270
rect 16395 3059 16455 3085
rect 16513 3059 16573 3270
rect 16866 3264 16926 3296
rect 16984 3270 17044 3296
rect 17102 3270 17162 3296
rect 16863 3248 16929 3264
rect 16863 3214 16879 3248
rect 16913 3214 16929 3248
rect 16863 3198 16929 3214
rect 22783 3564 22843 3585
rect 22901 3564 22961 3585
rect 23019 3564 23079 3585
rect 23137 3584 23433 3620
rect 23137 3564 23197 3584
rect 23255 3564 23315 3584
rect 23373 3564 23433 3584
rect 23491 3584 23787 3620
rect 23491 3564 23551 3584
rect 23609 3564 23669 3584
rect 23727 3564 23787 3584
rect 22783 3338 22843 3364
rect 22901 3338 22961 3364
rect 23019 3338 23079 3364
rect 23137 3344 23197 3364
rect 23137 3338 23198 3344
rect 23255 3338 23315 3364
rect 23373 3338 23433 3364
rect 18483 3151 18543 3168
rect 16745 3131 16811 3147
rect 16745 3097 16761 3131
rect 16795 3097 16811 3131
rect 16745 3081 16811 3097
rect 16748 3059 16808 3081
rect 18483 3062 18544 3151
rect 18601 3142 18661 3168
rect 18719 3142 18779 3168
rect 12999 2988 13385 3039
rect 12999 2857 13059 2988
rect 13114 2930 13180 2946
rect 13114 2896 13130 2930
rect 13164 2896 13180 2930
rect 13114 2880 13180 2896
rect 13117 2857 13177 2880
rect 13400 2857 13460 2883
rect 13518 2857 13578 2883
rect 13636 2857 13696 2883
rect 9741 2705 9801 2727
rect 9859 2705 9919 2727
rect 9738 2689 9804 2705
rect 9738 2655 9754 2689
rect 9788 2655 9804 2689
rect 9738 2639 9804 2655
rect 9856 2689 9922 2705
rect 9856 2655 9872 2689
rect 9906 2655 9922 2689
rect 9856 2639 9922 2655
rect 18393 3009 18544 3062
rect 16748 2833 16808 2859
rect 18393 2785 18453 3009
rect 18837 2967 18897 3168
rect 18955 3142 19015 3168
rect 19073 3142 19133 3168
rect 19625 3155 19685 3172
rect 19625 3066 19686 3155
rect 19743 3146 19803 3172
rect 19861 3146 19921 3172
rect 18511 2916 18897 2967
rect 19535 3013 19686 3066
rect 18511 2785 18571 2916
rect 18626 2858 18692 2874
rect 18626 2824 18642 2858
rect 18676 2824 18692 2858
rect 18626 2808 18692 2824
rect 18629 2785 18689 2808
rect 18912 2785 18972 2811
rect 19030 2785 19090 2811
rect 19148 2785 19208 2811
rect 19535 2789 19595 3013
rect 19979 2971 20039 3172
rect 20097 3146 20157 3172
rect 20215 3146 20275 3172
rect 23020 3153 23078 3338
rect 23020 3127 23080 3153
rect 23138 3127 23198 3338
rect 23491 3332 23551 3364
rect 23609 3338 23669 3364
rect 23727 3338 23787 3364
rect 23488 3316 23554 3332
rect 23488 3282 23504 3316
rect 23538 3282 23554 3316
rect 23488 3266 23554 3282
rect 31816 3640 31876 3666
rect 30938 3440 30998 3466
rect 31056 3440 31116 3466
rect 31174 3440 31234 3466
rect 31292 3440 31352 3466
rect 25108 3219 25168 3236
rect 23370 3199 23436 3215
rect 23370 3165 23386 3199
rect 23420 3165 23436 3199
rect 23370 3149 23436 3165
rect 23373 3127 23433 3149
rect 25108 3130 25169 3219
rect 25226 3210 25286 3236
rect 25344 3210 25404 3236
rect 19653 2920 20039 2971
rect 19653 2789 19713 2920
rect 19768 2862 19834 2878
rect 19768 2828 19784 2862
rect 19818 2828 19834 2862
rect 19768 2812 19834 2828
rect 19771 2789 19831 2812
rect 20054 2789 20114 2815
rect 20172 2789 20232 2815
rect 20290 2789 20350 2815
rect 11739 2627 11799 2653
rect 11857 2627 11917 2653
rect 11975 2621 12035 2653
rect 12258 2621 12318 2653
rect 12376 2621 12436 2653
rect 12494 2621 12554 2653
rect 12881 2631 12941 2657
rect 12999 2631 13059 2657
rect 11975 2580 12554 2621
rect 13117 2625 13177 2657
rect 13400 2625 13460 2657
rect 13518 2625 13578 2657
rect 13636 2625 13696 2657
rect 16395 2637 16455 2659
rect 16513 2637 16573 2659
rect 13117 2584 13696 2625
rect 16392 2621 16458 2637
rect 16392 2587 16408 2621
rect 16442 2587 16458 2621
rect 16392 2571 16458 2587
rect 16510 2621 16576 2637
rect 16510 2587 16526 2621
rect 16560 2587 16576 2621
rect 16510 2571 16576 2587
rect 25018 3077 25169 3130
rect 23373 2901 23433 2927
rect 25018 2853 25078 3077
rect 25462 3035 25522 3236
rect 25580 3210 25640 3236
rect 25698 3210 25758 3236
rect 26250 3223 26310 3240
rect 26250 3134 26311 3223
rect 26368 3214 26428 3240
rect 26486 3214 26546 3240
rect 25136 2984 25522 3035
rect 26160 3081 26311 3134
rect 25136 2853 25196 2984
rect 25251 2926 25317 2942
rect 25251 2892 25267 2926
rect 25301 2892 25317 2926
rect 25251 2876 25317 2892
rect 25254 2853 25314 2876
rect 25537 2853 25597 2879
rect 25655 2853 25715 2879
rect 25773 2853 25833 2879
rect 26160 2857 26220 3081
rect 26604 3039 26664 3240
rect 26722 3214 26782 3240
rect 26840 3214 26900 3240
rect 26278 2988 26664 3039
rect 26278 2857 26338 2988
rect 28580 2946 28876 2982
rect 26393 2930 26459 2946
rect 26393 2896 26409 2930
rect 26443 2896 26459 2930
rect 28580 2925 28640 2946
rect 28698 2925 28758 2946
rect 28816 2925 28876 2946
rect 28934 2945 29230 2981
rect 28934 2925 28994 2945
rect 29052 2925 29112 2945
rect 29170 2925 29230 2945
rect 29288 2945 29584 2981
rect 29288 2925 29348 2945
rect 29406 2925 29466 2945
rect 29524 2925 29584 2945
rect 26393 2880 26459 2896
rect 26396 2857 26456 2880
rect 26679 2857 26739 2883
rect 26797 2857 26857 2883
rect 26915 2857 26975 2883
rect 23020 2705 23080 2727
rect 23138 2705 23198 2727
rect 23017 2689 23083 2705
rect 23017 2655 23033 2689
rect 23067 2655 23083 2689
rect 23017 2639 23083 2655
rect 23135 2689 23201 2705
rect 23135 2655 23151 2689
rect 23185 2655 23201 2689
rect 23135 2639 23201 2655
rect 28580 2699 28640 2725
rect 28698 2699 28758 2725
rect 28816 2699 28876 2725
rect 28934 2705 28994 2725
rect 28934 2699 28995 2705
rect 29052 2699 29112 2725
rect 29170 2699 29230 2725
rect 25018 2627 25078 2653
rect 25136 2627 25196 2653
rect 25254 2621 25314 2653
rect 25537 2621 25597 2653
rect 25655 2621 25715 2653
rect 25773 2621 25833 2653
rect 26160 2631 26220 2657
rect 26278 2631 26338 2657
rect 5190 2539 5250 2565
rect 5308 2539 5368 2565
rect 5426 2533 5486 2565
rect 5709 2533 5769 2565
rect 5827 2533 5887 2565
rect 5945 2533 6005 2565
rect 6332 2543 6392 2569
rect 6450 2543 6510 2569
rect 5426 2492 6005 2533
rect 6568 2537 6628 2569
rect 6851 2537 6911 2569
rect 6969 2537 7029 2569
rect 7087 2537 7147 2569
rect 18393 2559 18453 2585
rect 18511 2559 18571 2585
rect 6568 2496 7147 2537
rect 18629 2553 18689 2585
rect 18912 2553 18972 2585
rect 19030 2553 19090 2585
rect 19148 2553 19208 2585
rect 19535 2563 19595 2589
rect 19653 2563 19713 2589
rect 18629 2512 19208 2553
rect 19771 2557 19831 2589
rect 20054 2557 20114 2589
rect 20172 2557 20232 2589
rect 20290 2557 20350 2589
rect 25254 2580 25833 2621
rect 26396 2625 26456 2657
rect 26679 2625 26739 2657
rect 26797 2625 26857 2657
rect 26915 2625 26975 2657
rect 26396 2584 26975 2625
rect 19771 2516 20350 2557
rect 28817 2514 28875 2699
rect 28817 2488 28877 2514
rect 28935 2488 28995 2699
rect 29288 2693 29348 2725
rect 29406 2699 29466 2725
rect 29524 2699 29584 2725
rect 29285 2677 29351 2693
rect 29285 2643 29301 2677
rect 29335 2643 29351 2677
rect 29285 2627 29351 2643
rect 29167 2560 29233 2576
rect 29167 2526 29183 2560
rect 29217 2526 29233 2560
rect 29167 2510 29233 2526
rect 29170 2488 29230 2510
rect 29170 2262 29230 2288
rect 28817 2066 28877 2088
rect 28935 2066 28995 2088
rect 28814 2050 28880 2066
rect 28814 2016 28830 2050
rect 28864 2016 28880 2050
rect 9518 1935 9814 1971
rect 9518 1914 9578 1935
rect 9636 1914 9696 1935
rect 9754 1914 9814 1935
rect 9872 1934 10168 1970
rect 9872 1914 9932 1934
rect 9990 1914 10050 1934
rect 10108 1914 10168 1934
rect 10226 1934 10522 1970
rect 10226 1914 10286 1934
rect 10344 1914 10404 1934
rect 10462 1914 10522 1934
rect 2969 1847 3265 1883
rect 2969 1826 3029 1847
rect 3087 1826 3147 1847
rect 3205 1826 3265 1847
rect 3323 1846 3619 1882
rect 3323 1826 3383 1846
rect 3441 1826 3501 1846
rect 3559 1826 3619 1846
rect 3677 1846 3973 1882
rect 3677 1826 3737 1846
rect 3795 1826 3855 1846
rect 3913 1826 3973 1846
rect 28814 2000 28880 2016
rect 28932 2050 28998 2066
rect 28932 2016 28948 2050
rect 28982 2016 28998 2050
rect 28932 2000 28998 2016
rect 22797 1935 23093 1971
rect 22797 1914 22857 1935
rect 22915 1914 22975 1935
rect 23033 1914 23093 1935
rect 23151 1934 23447 1970
rect 23151 1914 23211 1934
rect 23269 1914 23329 1934
rect 23387 1914 23447 1934
rect 23505 1934 23801 1970
rect 23505 1914 23565 1934
rect 23623 1914 23683 1934
rect 23741 1914 23801 1934
rect 16172 1867 16468 1903
rect 16172 1846 16232 1867
rect 16290 1846 16350 1867
rect 16408 1846 16468 1867
rect 16526 1866 16822 1902
rect 16526 1846 16586 1866
rect 16644 1846 16704 1866
rect 16762 1846 16822 1866
rect 16880 1866 17176 1902
rect 16880 1846 16940 1866
rect 16998 1846 17058 1866
rect 17116 1846 17176 1866
rect 9518 1688 9578 1714
rect 9636 1688 9696 1714
rect 9754 1688 9814 1714
rect 9872 1694 9932 1714
rect 9872 1688 9933 1694
rect 9990 1688 10050 1714
rect 10108 1688 10168 1714
rect 2969 1600 3029 1626
rect 3087 1600 3147 1626
rect 3205 1600 3265 1626
rect 3323 1606 3383 1626
rect 3323 1600 3384 1606
rect 3441 1600 3501 1626
rect 3559 1600 3619 1626
rect 3206 1415 3264 1600
rect 3206 1389 3266 1415
rect 3324 1389 3384 1600
rect 3677 1594 3737 1626
rect 3795 1600 3855 1626
rect 3913 1600 3973 1626
rect 3674 1578 3740 1594
rect 3674 1544 3690 1578
rect 3724 1544 3740 1578
rect 3674 1528 3740 1544
rect 9755 1503 9813 1688
rect 9755 1477 9815 1503
rect 9873 1477 9933 1688
rect 10226 1682 10286 1714
rect 10344 1688 10404 1714
rect 10462 1688 10522 1714
rect 10223 1666 10289 1682
rect 10223 1632 10239 1666
rect 10273 1632 10289 1666
rect 22797 1688 22857 1714
rect 22915 1688 22975 1714
rect 23033 1688 23093 1714
rect 23151 1694 23211 1714
rect 23151 1688 23212 1694
rect 23269 1688 23329 1714
rect 23387 1688 23447 1714
rect 10223 1616 10289 1632
rect 16172 1620 16232 1646
rect 16290 1620 16350 1646
rect 16408 1620 16468 1646
rect 16526 1626 16586 1646
rect 16526 1620 16587 1626
rect 16644 1620 16704 1646
rect 16762 1620 16822 1646
rect 10105 1549 10171 1565
rect 10105 1515 10121 1549
rect 10155 1515 10171 1549
rect 10105 1499 10171 1515
rect 11466 1512 11762 1563
rect 10108 1477 10168 1499
rect 11466 1497 11526 1512
rect 11584 1497 11644 1512
rect 11702 1497 11762 1512
rect 11820 1497 11880 1523
rect 11938 1497 11998 1523
rect 12056 1497 12116 1523
rect 13364 1512 13660 1563
rect 13364 1497 13424 1512
rect 13482 1497 13542 1512
rect 13600 1497 13660 1512
rect 13718 1497 13778 1523
rect 13836 1497 13896 1523
rect 13954 1497 14014 1523
rect 3556 1461 3622 1477
rect 3556 1427 3572 1461
rect 3606 1427 3622 1461
rect 3556 1411 3622 1427
rect 4917 1424 5213 1475
rect 3559 1389 3619 1411
rect 4917 1409 4977 1424
rect 5035 1409 5095 1424
rect 5153 1409 5213 1424
rect 5271 1409 5331 1435
rect 5389 1409 5449 1435
rect 5507 1409 5567 1435
rect 6815 1424 7111 1475
rect 6815 1409 6875 1424
rect 6933 1409 6993 1424
rect 7051 1409 7111 1424
rect 7169 1409 7229 1435
rect 7287 1409 7347 1435
rect 7405 1409 7465 1435
rect 57 1179 353 1215
rect 57 1158 117 1179
rect 175 1158 235 1179
rect 293 1158 353 1179
rect 411 1178 707 1214
rect 411 1158 471 1178
rect 529 1158 589 1178
rect 647 1158 707 1178
rect 765 1178 1061 1214
rect 765 1158 825 1178
rect 883 1158 943 1178
rect 1001 1158 1061 1178
rect 4433 1209 4493 1235
rect 4551 1209 4611 1235
rect 4669 1209 4729 1235
rect 3559 1163 3619 1189
rect 3206 967 3266 989
rect 3324 973 3384 989
rect 57 932 117 958
rect 175 932 235 958
rect 293 932 353 958
rect 411 938 471 958
rect 411 932 472 938
rect 529 932 589 958
rect 647 932 707 958
rect 294 747 352 932
rect 294 721 354 747
rect 412 721 472 932
rect 765 926 825 958
rect 883 932 943 958
rect 1001 932 1061 958
rect 3203 951 3269 967
rect 762 910 828 926
rect 762 876 778 910
rect 812 876 828 910
rect 3203 917 3219 951
rect 3253 917 3269 951
rect 3203 901 3269 917
rect 3318 951 3392 973
rect 3318 917 3337 951
rect 3371 917 3392 951
rect 5754 1226 6050 1277
rect 5754 1209 5814 1226
rect 5872 1209 5932 1226
rect 5990 1209 6050 1226
rect 6331 1209 6391 1235
rect 6449 1209 6509 1235
rect 6567 1209 6627 1235
rect 7652 1226 7948 1277
rect 7652 1209 7712 1226
rect 7770 1209 7830 1226
rect 7888 1209 7948 1226
rect 10982 1297 11042 1323
rect 11100 1297 11160 1323
rect 11218 1297 11278 1323
rect 10108 1251 10168 1277
rect 9755 1055 9815 1077
rect 9873 1061 9933 1077
rect 9752 1039 9818 1055
rect 4433 992 4493 1009
rect 4551 992 4611 1009
rect 4669 992 4729 1009
rect 4917 992 4977 1009
rect 4433 941 4977 992
rect 5035 983 5095 1009
rect 5153 983 5213 1009
rect 5271 990 5331 1009
rect 5389 990 5449 1009
rect 5507 990 5567 1009
rect 5754 990 5814 1009
rect 5872 990 5932 1009
rect 762 860 828 876
rect 3318 860 3392 917
rect 4558 860 4618 941
rect 5271 939 5814 990
rect 5856 983 5932 990
rect 5990 983 6050 1009
rect 6331 992 6391 1009
rect 6449 992 6509 1009
rect 6567 992 6627 1009
rect 6815 992 6875 1009
rect 5856 939 5931 983
rect 6331 941 6875 992
rect 6933 983 6993 1009
rect 7051 983 7111 1009
rect 7169 990 7229 1009
rect 7287 990 7347 1009
rect 7405 990 7465 1009
rect 7652 990 7712 1009
rect 7770 990 7830 1009
rect 3318 835 4618 860
rect 644 793 710 809
rect 644 759 660 793
rect 694 759 710 793
rect 3317 787 4618 835
rect 5856 819 5916 939
rect 644 743 710 759
rect 647 721 707 743
rect 647 495 707 521
rect 294 299 354 321
rect 412 299 472 321
rect 291 283 357 299
rect 291 249 307 283
rect 341 249 357 283
rect 291 233 357 249
rect 409 283 475 299
rect 409 249 425 283
rect 459 249 475 283
rect 409 233 475 249
rect 2964 243 3260 279
rect 2964 222 3024 243
rect 3082 222 3142 243
rect 3200 222 3260 243
rect 3318 242 3614 278
rect 3318 222 3378 242
rect 3436 222 3496 242
rect 3554 222 3614 242
rect 3672 242 3968 278
rect 3672 222 3732 242
rect 3790 222 3850 242
rect 3908 222 3968 242
rect 4558 89 4618 787
rect 4860 739 5156 799
rect 4860 716 4920 739
rect 4978 716 5038 739
rect 5096 716 5156 739
rect 5214 740 5510 800
rect 5855 799 5916 819
rect 5214 716 5274 740
rect 5332 716 5392 740
rect 5450 716 5510 740
rect 5836 783 5916 799
rect 5836 749 5851 783
rect 5885 749 5916 783
rect 5836 733 5916 749
rect 5855 710 5916 733
rect 5856 564 5916 710
rect 5855 391 5916 564
rect 4860 290 4920 316
rect 4828 149 4895 156
rect 4978 149 5038 316
rect 5096 290 5156 316
rect 5214 290 5274 316
rect 4828 140 5038 149
rect 4828 106 4844 140
rect 4878 106 5038 140
rect 4828 90 5038 106
rect 4558 73 4709 89
rect 4558 39 4659 73
rect 4693 39 4709 73
rect 4558 23 4709 39
rect 2964 -4 3024 22
rect 3082 -4 3142 22
rect 3200 -4 3260 22
rect 3318 2 3378 22
rect 3318 -4 3379 2
rect 3436 -4 3496 22
rect 3554 -4 3614 22
rect 3201 -189 3259 -4
rect 3201 -215 3261 -189
rect 3319 -215 3379 -4
rect 3672 -10 3732 22
rect 3790 -4 3850 22
rect 3908 -4 3968 22
rect 3669 -26 3735 -10
rect 4558 -16 4618 23
rect 4978 -16 5038 90
rect 5332 149 5392 316
rect 5450 290 5510 316
rect 5475 149 5542 156
rect 5332 140 5542 149
rect 5332 106 5492 140
rect 5526 106 5542 140
rect 5332 90 5542 106
rect 5094 56 5160 72
rect 5094 22 5110 56
rect 5144 22 5160 56
rect 5094 6 5160 22
rect 5212 57 5278 72
rect 5212 23 5228 57
rect 5262 23 5278 57
rect 5212 7 5278 23
rect 5096 -16 5156 6
rect 5214 -16 5274 7
rect 5332 -16 5392 90
rect 5856 88 5916 391
rect 5766 72 5916 88
rect 5766 38 5782 72
rect 5816 38 5916 72
rect 5766 22 5916 38
rect 5856 -16 5916 22
rect 6456 283 6516 941
rect 7169 939 7712 990
rect 7754 983 7830 990
rect 7888 983 7948 1009
rect 9752 1005 9768 1039
rect 9802 1005 9818 1039
rect 9752 989 9818 1005
rect 9867 1039 9941 1061
rect 9867 1005 9886 1039
rect 9920 1005 9941 1039
rect 12303 1314 12599 1365
rect 12303 1297 12363 1314
rect 12421 1297 12481 1314
rect 12539 1297 12599 1314
rect 12880 1297 12940 1323
rect 12998 1297 13058 1323
rect 13116 1297 13176 1323
rect 16409 1435 16467 1620
rect 16409 1409 16469 1435
rect 16527 1409 16587 1620
rect 16880 1614 16940 1646
rect 16998 1620 17058 1646
rect 17116 1620 17176 1646
rect 16877 1598 16943 1614
rect 16877 1564 16893 1598
rect 16927 1564 16943 1598
rect 16877 1548 16943 1564
rect 23034 1503 23092 1688
rect 16759 1481 16825 1497
rect 16759 1447 16775 1481
rect 16809 1447 16825 1481
rect 16759 1431 16825 1447
rect 18120 1444 18416 1495
rect 16762 1409 16822 1431
rect 18120 1429 18180 1444
rect 18238 1429 18298 1444
rect 18356 1429 18416 1444
rect 18474 1429 18534 1455
rect 18592 1429 18652 1455
rect 18710 1429 18770 1455
rect 20018 1444 20314 1495
rect 23034 1477 23094 1503
rect 23152 1477 23212 1688
rect 23505 1682 23565 1714
rect 23623 1688 23683 1714
rect 23741 1688 23801 1714
rect 23502 1666 23568 1682
rect 23502 1632 23518 1666
rect 23552 1632 23568 1666
rect 23502 1616 23568 1632
rect 23384 1549 23450 1565
rect 23384 1515 23400 1549
rect 23434 1515 23450 1549
rect 23384 1499 23450 1515
rect 24745 1512 25041 1563
rect 23387 1477 23447 1499
rect 24745 1497 24805 1512
rect 24863 1497 24923 1512
rect 24981 1497 25041 1512
rect 25099 1497 25159 1523
rect 25217 1497 25277 1523
rect 25335 1497 25395 1523
rect 26643 1512 26939 1563
rect 26643 1497 26703 1512
rect 26761 1497 26821 1512
rect 26879 1497 26939 1512
rect 26997 1497 27057 1523
rect 27115 1497 27175 1523
rect 27233 1497 27293 1523
rect 20018 1429 20078 1444
rect 20136 1429 20196 1444
rect 20254 1429 20314 1444
rect 20372 1429 20432 1455
rect 20490 1429 20550 1455
rect 20608 1429 20668 1455
rect 14201 1314 14497 1365
rect 14201 1297 14261 1314
rect 14319 1297 14379 1314
rect 14437 1297 14497 1314
rect 10982 1080 11042 1097
rect 11100 1080 11160 1097
rect 11218 1080 11278 1097
rect 11466 1080 11526 1097
rect 10982 1029 11526 1080
rect 11584 1071 11644 1097
rect 11702 1071 11762 1097
rect 11820 1078 11880 1097
rect 11938 1078 11998 1097
rect 12056 1078 12116 1097
rect 12303 1078 12363 1097
rect 12421 1078 12481 1097
rect 7754 939 7829 983
rect 9867 948 9941 1005
rect 11107 948 11167 1029
rect 11820 1027 12363 1078
rect 12405 1071 12481 1078
rect 12539 1071 12599 1097
rect 12880 1080 12940 1097
rect 12998 1080 13058 1097
rect 13116 1080 13176 1097
rect 13364 1080 13424 1097
rect 12405 1027 12480 1071
rect 12880 1029 13424 1080
rect 13482 1071 13542 1097
rect 13600 1071 13660 1097
rect 13718 1078 13778 1097
rect 13836 1078 13896 1097
rect 13954 1078 14014 1097
rect 14201 1078 14261 1097
rect 14319 1078 14379 1097
rect 6758 739 7054 799
rect 6758 716 6818 739
rect 6876 716 6936 739
rect 6994 716 7054 739
rect 7112 740 7408 800
rect 7112 716 7172 740
rect 7230 716 7290 740
rect 7348 716 7408 740
rect 7754 786 7814 939
rect 9867 923 11167 948
rect 9866 875 11167 923
rect 12405 907 12465 1027
rect 7754 762 8008 786
rect 7754 728 7958 762
rect 7992 728 8008 762
rect 7754 712 8008 728
rect 6758 290 6818 316
rect 6456 267 6523 283
rect 6456 233 6472 267
rect 6506 233 6523 267
rect 6456 217 6523 233
rect 6456 89 6516 217
rect 6726 149 6793 156
rect 6876 149 6936 316
rect 6994 290 7054 316
rect 7112 290 7172 316
rect 6726 140 6936 149
rect 6726 106 6742 140
rect 6776 106 6936 140
rect 6726 90 6936 106
rect 6456 73 6607 89
rect 6456 39 6557 73
rect 6591 39 6607 73
rect 6456 23 6607 39
rect 6456 -16 6516 23
rect 6876 -16 6936 90
rect 7230 149 7290 316
rect 7348 290 7408 316
rect 7371 150 7438 157
rect 7365 149 7438 150
rect 7230 141 7438 149
rect 7230 107 7388 141
rect 7422 107 7438 141
rect 7230 91 7438 107
rect 7230 90 7427 91
rect 6992 56 7058 72
rect 6992 22 7008 56
rect 7042 22 7058 56
rect 6992 6 7058 22
rect 7110 57 7176 72
rect 7110 23 7126 57
rect 7160 23 7176 57
rect 7110 7 7176 23
rect 6994 -16 7054 6
rect 7112 -16 7172 7
rect 7230 -16 7290 90
rect 7754 88 7814 712
rect 9513 331 9809 367
rect 9513 310 9573 331
rect 9631 310 9691 331
rect 9749 310 9809 331
rect 9867 330 10163 366
rect 9867 310 9927 330
rect 9985 310 10045 330
rect 10103 310 10163 330
rect 10221 330 10517 366
rect 10221 310 10281 330
rect 10339 310 10399 330
rect 10457 310 10517 330
rect 11107 177 11167 875
rect 11409 827 11705 887
rect 11409 804 11469 827
rect 11527 804 11587 827
rect 11645 804 11705 827
rect 11763 828 12059 888
rect 12404 887 12465 907
rect 11763 804 11823 828
rect 11881 804 11941 828
rect 11999 804 12059 828
rect 12385 871 12465 887
rect 12385 837 12400 871
rect 12434 837 12465 871
rect 12385 821 12465 837
rect 12404 798 12465 821
rect 12405 652 12465 798
rect 12404 479 12465 652
rect 11409 378 11469 404
rect 11377 237 11444 244
rect 11527 237 11587 404
rect 11645 378 11705 404
rect 11763 378 11823 404
rect 11377 228 11587 237
rect 11377 194 11393 228
rect 11427 194 11587 228
rect 11377 178 11587 194
rect 11107 161 11258 177
rect 11107 127 11208 161
rect 11242 127 11258 161
rect 11107 111 11258 127
rect 7664 72 7814 88
rect 9513 84 9573 110
rect 9631 84 9691 110
rect 9749 84 9809 110
rect 9867 90 9927 110
rect 9867 84 9928 90
rect 9985 84 10045 110
rect 10103 84 10163 110
rect 7664 38 7680 72
rect 7714 38 7814 72
rect 7664 22 7814 38
rect 7754 -16 7814 22
rect 3669 -60 3685 -26
rect 3719 -60 3735 -26
rect 3669 -76 3735 -60
rect 3551 -143 3617 -127
rect 3551 -177 3567 -143
rect 3601 -177 3617 -143
rect 3551 -193 3617 -177
rect 3554 -215 3614 -193
rect 4558 -242 4618 -216
rect 3554 -441 3614 -415
rect 5856 -242 5916 -216
rect 6456 -242 6516 -216
rect 9750 -101 9808 84
rect 9750 -127 9810 -101
rect 9868 -127 9928 84
rect 10221 78 10281 110
rect 10339 84 10399 110
rect 10457 84 10517 110
rect 10218 62 10284 78
rect 11107 72 11167 111
rect 11527 72 11587 178
rect 11881 237 11941 404
rect 11999 378 12059 404
rect 12024 237 12091 244
rect 11881 228 12091 237
rect 11881 194 12041 228
rect 12075 194 12091 228
rect 11881 178 12091 194
rect 11643 144 11709 160
rect 11643 110 11659 144
rect 11693 110 11709 144
rect 11643 94 11709 110
rect 11761 145 11827 160
rect 11761 111 11777 145
rect 11811 111 11827 145
rect 11761 95 11827 111
rect 11645 72 11705 94
rect 11763 72 11823 95
rect 11881 72 11941 178
rect 12405 176 12465 479
rect 12315 160 12465 176
rect 12315 126 12331 160
rect 12365 126 12465 160
rect 12315 110 12465 126
rect 12405 72 12465 110
rect 13005 371 13065 1029
rect 13718 1027 14261 1078
rect 14303 1071 14379 1078
rect 14437 1071 14497 1097
rect 14303 1027 14378 1071
rect 13307 827 13603 887
rect 13307 804 13367 827
rect 13425 804 13485 827
rect 13543 804 13603 827
rect 13661 828 13957 888
rect 13661 804 13721 828
rect 13779 804 13839 828
rect 13897 804 13957 828
rect 14303 874 14363 1027
rect 17636 1229 17696 1255
rect 17754 1229 17814 1255
rect 17872 1229 17932 1255
rect 16762 1183 16822 1209
rect 16409 987 16469 1009
rect 16527 993 16587 1009
rect 16406 971 16472 987
rect 16406 937 16422 971
rect 16456 937 16472 971
rect 16406 921 16472 937
rect 16521 971 16595 993
rect 16521 937 16540 971
rect 16574 937 16595 971
rect 18957 1246 19253 1297
rect 18957 1229 19017 1246
rect 19075 1229 19135 1246
rect 19193 1229 19253 1246
rect 19534 1229 19594 1255
rect 19652 1229 19712 1255
rect 19770 1229 19830 1255
rect 20855 1246 21151 1297
rect 20855 1229 20915 1246
rect 20973 1229 21033 1246
rect 21091 1229 21151 1246
rect 24261 1297 24321 1323
rect 24379 1297 24439 1323
rect 24497 1297 24557 1323
rect 23387 1251 23447 1277
rect 23034 1055 23094 1077
rect 23152 1061 23212 1077
rect 23031 1039 23097 1055
rect 17636 1012 17696 1029
rect 17754 1012 17814 1029
rect 17872 1012 17932 1029
rect 18120 1012 18180 1029
rect 17636 961 18180 1012
rect 18238 1003 18298 1029
rect 18356 1003 18416 1029
rect 18474 1010 18534 1029
rect 18592 1010 18652 1029
rect 18710 1010 18770 1029
rect 18957 1010 19017 1029
rect 19075 1010 19135 1029
rect 16521 880 16595 937
rect 17761 880 17821 961
rect 18474 959 19017 1010
rect 19059 1003 19135 1010
rect 19193 1003 19253 1029
rect 19534 1012 19594 1029
rect 19652 1012 19712 1029
rect 19770 1012 19830 1029
rect 20018 1012 20078 1029
rect 19059 959 19134 1003
rect 19534 961 20078 1012
rect 20136 1003 20196 1029
rect 20254 1003 20314 1029
rect 20372 1010 20432 1029
rect 20490 1010 20550 1029
rect 20608 1010 20668 1029
rect 20855 1010 20915 1029
rect 20973 1010 21033 1029
rect 14303 850 14557 874
rect 16521 855 17821 880
rect 14303 816 14507 850
rect 14541 816 14557 850
rect 14303 800 14557 816
rect 16520 807 17821 855
rect 19059 839 19119 959
rect 13307 378 13367 404
rect 13005 355 13072 371
rect 13005 321 13021 355
rect 13055 321 13072 355
rect 13005 305 13072 321
rect 13005 177 13065 305
rect 13275 237 13342 244
rect 13425 237 13485 404
rect 13543 378 13603 404
rect 13661 378 13721 404
rect 13275 228 13485 237
rect 13275 194 13291 228
rect 13325 194 13485 228
rect 13275 178 13485 194
rect 13005 161 13156 177
rect 13005 127 13106 161
rect 13140 127 13156 161
rect 13005 111 13156 127
rect 13005 72 13065 111
rect 13425 72 13485 178
rect 13779 237 13839 404
rect 13897 378 13957 404
rect 13920 238 13987 245
rect 13914 237 13987 238
rect 13779 229 13987 237
rect 13779 195 13937 229
rect 13971 195 13987 229
rect 13779 179 13987 195
rect 13779 178 13976 179
rect 13541 144 13607 160
rect 13541 110 13557 144
rect 13591 110 13607 144
rect 13541 94 13607 110
rect 13659 145 13725 160
rect 13659 111 13675 145
rect 13709 111 13725 145
rect 13659 95 13725 111
rect 13543 72 13603 94
rect 13661 72 13721 95
rect 13779 72 13839 178
rect 14303 176 14363 800
rect 16167 263 16463 299
rect 16167 242 16227 263
rect 16285 242 16345 263
rect 16403 242 16463 263
rect 16521 262 16817 298
rect 16521 242 16581 262
rect 16639 242 16699 262
rect 16757 242 16817 262
rect 16875 262 17171 298
rect 16875 242 16935 262
rect 16993 242 17053 262
rect 17111 242 17171 262
rect 14213 160 14363 176
rect 14213 126 14229 160
rect 14263 126 14363 160
rect 14213 110 14363 126
rect 14303 72 14363 110
rect 10218 28 10234 62
rect 10268 28 10284 62
rect 10218 12 10284 28
rect 10100 -55 10166 -39
rect 10100 -89 10116 -55
rect 10150 -89 10166 -55
rect 10100 -105 10166 -89
rect 10103 -127 10163 -105
rect 7754 -242 7814 -216
rect 4978 -442 5038 -416
rect 5096 -442 5156 -416
rect 5214 -442 5274 -416
rect 5332 -442 5392 -416
rect 6876 -442 6936 -416
rect 6994 -442 7054 -416
rect 7112 -442 7172 -416
rect 7230 -442 7290 -416
rect 11107 -154 11167 -128
rect 10103 -353 10163 -327
rect 12405 -154 12465 -128
rect 13005 -154 13065 -128
rect 17761 109 17821 807
rect 18063 759 18359 819
rect 18063 736 18123 759
rect 18181 736 18241 759
rect 18299 736 18359 759
rect 18417 760 18713 820
rect 19058 819 19119 839
rect 18417 736 18477 760
rect 18535 736 18595 760
rect 18653 736 18713 760
rect 19039 803 19119 819
rect 19039 769 19054 803
rect 19088 769 19119 803
rect 19039 753 19119 769
rect 19058 730 19119 753
rect 19059 584 19119 730
rect 19058 411 19119 584
rect 18063 310 18123 336
rect 18031 169 18098 176
rect 18181 169 18241 336
rect 18299 310 18359 336
rect 18417 310 18477 336
rect 18031 160 18241 169
rect 18031 126 18047 160
rect 18081 126 18241 160
rect 18031 110 18241 126
rect 17761 93 17912 109
rect 17761 59 17862 93
rect 17896 59 17912 93
rect 17761 43 17912 59
rect 16167 16 16227 42
rect 16285 16 16345 42
rect 16403 16 16463 42
rect 16521 22 16581 42
rect 16521 16 16582 22
rect 16639 16 16699 42
rect 16757 16 16817 42
rect 14303 -154 14363 -128
rect 16404 -169 16462 16
rect 16404 -195 16464 -169
rect 16522 -195 16582 16
rect 16875 10 16935 42
rect 16993 16 17053 42
rect 17111 16 17171 42
rect 16872 -6 16938 10
rect 17761 4 17821 43
rect 18181 4 18241 110
rect 18535 169 18595 336
rect 18653 310 18713 336
rect 18678 169 18745 176
rect 18535 160 18745 169
rect 18535 126 18695 160
rect 18729 126 18745 160
rect 18535 110 18745 126
rect 18297 76 18363 92
rect 18297 42 18313 76
rect 18347 42 18363 76
rect 18297 26 18363 42
rect 18415 77 18481 92
rect 18415 43 18431 77
rect 18465 43 18481 77
rect 18415 27 18481 43
rect 18299 4 18359 26
rect 18417 4 18477 27
rect 18535 4 18595 110
rect 19059 108 19119 411
rect 18969 92 19119 108
rect 18969 58 18985 92
rect 19019 58 19119 92
rect 18969 42 19119 58
rect 19059 4 19119 42
rect 19659 303 19719 961
rect 20372 959 20915 1010
rect 20957 1003 21033 1010
rect 21091 1003 21151 1029
rect 23031 1005 23047 1039
rect 23081 1005 23097 1039
rect 20957 959 21032 1003
rect 23031 989 23097 1005
rect 23146 1039 23220 1061
rect 23146 1005 23165 1039
rect 23199 1005 23220 1039
rect 25582 1314 25878 1365
rect 25582 1297 25642 1314
rect 25700 1297 25760 1314
rect 25818 1297 25878 1314
rect 26159 1297 26219 1323
rect 26277 1297 26337 1323
rect 26395 1297 26455 1323
rect 27480 1314 27776 1365
rect 27480 1297 27540 1314
rect 27598 1297 27658 1314
rect 27716 1297 27776 1314
rect 30879 1215 31175 1266
rect 30879 1200 30939 1215
rect 30997 1200 31057 1215
rect 31115 1200 31175 1215
rect 31233 1200 31293 1226
rect 31351 1200 31411 1226
rect 31469 1200 31529 1226
rect 24261 1080 24321 1097
rect 24379 1080 24439 1097
rect 24497 1080 24557 1097
rect 24745 1080 24805 1097
rect 24261 1029 24805 1080
rect 24863 1071 24923 1097
rect 24981 1071 25041 1097
rect 25099 1078 25159 1097
rect 25217 1078 25277 1097
rect 25335 1078 25395 1097
rect 25582 1078 25642 1097
rect 25700 1078 25760 1097
rect 19961 759 20257 819
rect 19961 736 20021 759
rect 20079 736 20139 759
rect 20197 736 20257 759
rect 20315 760 20611 820
rect 20315 736 20375 760
rect 20433 736 20493 760
rect 20551 736 20611 760
rect 20957 806 21017 959
rect 23146 948 23220 1005
rect 24386 948 24446 1029
rect 25099 1027 25642 1078
rect 25684 1071 25760 1078
rect 25818 1071 25878 1097
rect 26159 1080 26219 1097
rect 26277 1080 26337 1097
rect 26395 1080 26455 1097
rect 26643 1080 26703 1097
rect 25684 1027 25759 1071
rect 26159 1029 26703 1080
rect 26761 1071 26821 1097
rect 26879 1071 26939 1097
rect 26997 1078 27057 1097
rect 27115 1078 27175 1097
rect 27233 1078 27293 1097
rect 27480 1078 27540 1097
rect 27598 1078 27658 1097
rect 23146 923 24446 948
rect 23145 875 24446 923
rect 25684 907 25744 1027
rect 20957 782 21211 806
rect 20957 748 21161 782
rect 21195 748 21211 782
rect 20957 732 21211 748
rect 19961 310 20021 336
rect 19659 287 19726 303
rect 19659 253 19675 287
rect 19709 253 19726 287
rect 19659 237 19726 253
rect 19659 109 19719 237
rect 19929 169 19996 176
rect 20079 169 20139 336
rect 20197 310 20257 336
rect 20315 310 20375 336
rect 19929 160 20139 169
rect 19929 126 19945 160
rect 19979 126 20139 160
rect 19929 110 20139 126
rect 19659 93 19810 109
rect 19659 59 19760 93
rect 19794 59 19810 93
rect 19659 43 19810 59
rect 19659 4 19719 43
rect 20079 4 20139 110
rect 20433 169 20493 336
rect 20551 310 20611 336
rect 20574 170 20641 177
rect 20568 169 20641 170
rect 20433 161 20641 169
rect 20433 127 20591 161
rect 20625 127 20641 161
rect 20433 111 20641 127
rect 20433 110 20630 111
rect 20195 76 20261 92
rect 20195 42 20211 76
rect 20245 42 20261 76
rect 20195 26 20261 42
rect 20313 77 20379 92
rect 20313 43 20329 77
rect 20363 43 20379 77
rect 20313 27 20379 43
rect 20197 4 20257 26
rect 20315 4 20375 27
rect 20433 4 20493 110
rect 20957 108 21017 732
rect 22792 331 23088 367
rect 22792 310 22852 331
rect 22910 310 22970 331
rect 23028 310 23088 331
rect 23146 330 23442 366
rect 23146 310 23206 330
rect 23264 310 23324 330
rect 23382 310 23442 330
rect 23500 330 23796 366
rect 23500 310 23560 330
rect 23618 310 23678 330
rect 23736 310 23796 330
rect 24386 177 24446 875
rect 24688 827 24984 887
rect 24688 804 24748 827
rect 24806 804 24866 827
rect 24924 804 24984 827
rect 25042 828 25338 888
rect 25683 887 25744 907
rect 25042 804 25102 828
rect 25160 804 25220 828
rect 25278 804 25338 828
rect 25664 871 25744 887
rect 25664 837 25679 871
rect 25713 837 25744 871
rect 25664 821 25744 837
rect 25683 798 25744 821
rect 25684 652 25744 798
rect 25683 479 25744 652
rect 24688 378 24748 404
rect 24656 237 24723 244
rect 24806 237 24866 404
rect 24924 378 24984 404
rect 25042 378 25102 404
rect 24656 228 24866 237
rect 24656 194 24672 228
rect 24706 194 24866 228
rect 24656 178 24866 194
rect 24386 161 24537 177
rect 24386 127 24487 161
rect 24521 127 24537 161
rect 24386 111 24537 127
rect 20867 92 21017 108
rect 20867 58 20883 92
rect 20917 58 21017 92
rect 22792 84 22852 110
rect 22910 84 22970 110
rect 23028 84 23088 110
rect 23146 90 23206 110
rect 23146 84 23207 90
rect 23264 84 23324 110
rect 23382 84 23442 110
rect 20867 42 21017 58
rect 20957 4 21017 42
rect 16872 -40 16888 -6
rect 16922 -40 16938 -6
rect 16872 -56 16938 -40
rect 16754 -123 16820 -107
rect 16754 -157 16770 -123
rect 16804 -157 16820 -123
rect 16754 -173 16820 -157
rect 16757 -195 16817 -173
rect 11527 -354 11587 -328
rect 11645 -354 11705 -328
rect 11763 -354 11823 -328
rect 11881 -354 11941 -328
rect 13425 -354 13485 -328
rect 13543 -354 13603 -328
rect 13661 -354 13721 -328
rect 13779 -354 13839 -328
rect 9750 -549 9810 -527
rect 9868 -549 9928 -527
rect 3201 -637 3261 -615
rect 3319 -637 3379 -615
rect 3198 -653 3264 -637
rect 3198 -687 3214 -653
rect 3248 -687 3264 -653
rect 3198 -703 3264 -687
rect 3316 -653 3382 -637
rect 3316 -687 3332 -653
rect 3366 -687 3382 -653
rect 9747 -565 9813 -549
rect 9747 -599 9763 -565
rect 9797 -599 9813 -565
rect 9747 -615 9813 -599
rect 9865 -565 9931 -549
rect 9865 -599 9881 -565
rect 9915 -599 9931 -565
rect 9865 -615 9931 -599
rect 17761 -222 17821 -196
rect 16757 -421 16817 -395
rect 19059 -222 19119 -196
rect 19659 -222 19719 -196
rect 23029 -101 23087 84
rect 23029 -127 23089 -101
rect 23147 -127 23207 84
rect 23500 78 23560 110
rect 23618 84 23678 110
rect 23736 84 23796 110
rect 23497 62 23563 78
rect 24386 72 24446 111
rect 24806 72 24866 178
rect 25160 237 25220 404
rect 25278 378 25338 404
rect 25303 237 25370 244
rect 25160 228 25370 237
rect 25160 194 25320 228
rect 25354 194 25370 228
rect 25160 178 25370 194
rect 24922 144 24988 160
rect 24922 110 24938 144
rect 24972 110 24988 144
rect 24922 94 24988 110
rect 25040 145 25106 160
rect 25040 111 25056 145
rect 25090 111 25106 145
rect 25040 95 25106 111
rect 24924 72 24984 94
rect 25042 72 25102 95
rect 25160 72 25220 178
rect 25684 176 25744 479
rect 25594 160 25744 176
rect 25594 126 25610 160
rect 25644 126 25744 160
rect 25594 110 25744 126
rect 25684 72 25744 110
rect 26284 371 26344 1029
rect 26997 1027 27540 1078
rect 27582 1071 27658 1078
rect 27716 1071 27776 1097
rect 27582 1027 27657 1071
rect 26586 827 26882 887
rect 26586 804 26646 827
rect 26704 804 26764 827
rect 26822 804 26882 827
rect 26940 828 27236 888
rect 26940 804 27000 828
rect 27058 804 27118 828
rect 27176 804 27236 828
rect 27582 874 27642 1027
rect 30395 1000 30455 1026
rect 30513 1000 30573 1026
rect 30631 1000 30691 1026
rect 27582 850 27836 874
rect 27582 816 27786 850
rect 27820 816 27836 850
rect 27582 800 27836 816
rect 31716 1017 32012 1068
rect 31716 1000 31776 1017
rect 31834 1000 31894 1017
rect 31952 1000 32012 1017
rect 32188 1018 32484 1054
rect 32188 997 32248 1018
rect 32306 997 32366 1018
rect 32424 997 32484 1018
rect 32542 1017 32838 1053
rect 32542 997 32602 1017
rect 32660 997 32720 1017
rect 32778 997 32838 1017
rect 32896 1017 33192 1053
rect 32896 997 32956 1017
rect 33014 997 33074 1017
rect 33132 997 33192 1017
rect 26586 378 26646 404
rect 26284 355 26351 371
rect 26284 321 26300 355
rect 26334 321 26351 355
rect 26284 305 26351 321
rect 26284 177 26344 305
rect 26554 237 26621 244
rect 26704 237 26764 404
rect 26822 378 26882 404
rect 26940 378 27000 404
rect 26554 228 26764 237
rect 26554 194 26570 228
rect 26604 194 26764 228
rect 26554 178 26764 194
rect 26284 161 26435 177
rect 26284 127 26385 161
rect 26419 127 26435 161
rect 26284 111 26435 127
rect 26284 72 26344 111
rect 26704 72 26764 178
rect 27058 237 27118 404
rect 27176 378 27236 404
rect 27199 238 27266 245
rect 27193 237 27266 238
rect 27058 229 27266 237
rect 27058 195 27216 229
rect 27250 195 27266 229
rect 27058 179 27266 195
rect 27058 178 27255 179
rect 26820 144 26886 160
rect 26820 110 26836 144
rect 26870 110 26886 144
rect 26820 94 26886 110
rect 26938 145 27004 160
rect 26938 111 26954 145
rect 26988 111 27004 145
rect 26938 95 27004 111
rect 26822 72 26882 94
rect 26940 72 27000 95
rect 27058 72 27118 178
rect 27582 176 27642 800
rect 30395 783 30455 800
rect 30513 783 30573 800
rect 30631 783 30691 800
rect 30879 783 30939 800
rect 30395 732 30939 783
rect 30997 774 31057 800
rect 31115 774 31175 800
rect 31233 781 31293 800
rect 31351 781 31411 800
rect 31469 781 31529 800
rect 31716 781 31776 800
rect 31834 781 31894 800
rect 27492 160 27642 176
rect 27492 126 27508 160
rect 27542 126 27642 160
rect 30520 528 30580 732
rect 31233 730 31776 781
rect 31818 774 31894 781
rect 31952 774 32012 800
rect 31818 730 31893 774
rect 32188 771 32248 797
rect 32306 771 32366 797
rect 32424 771 32484 797
rect 32542 777 32602 797
rect 32542 771 32603 777
rect 32660 771 32720 797
rect 32778 771 32838 797
rect 31818 648 31878 730
rect 31818 630 32052 648
rect 31818 596 32001 630
rect 32035 596 32052 630
rect 30822 530 31118 590
rect 30520 511 30651 528
rect 30520 477 30601 511
rect 30635 477 30651 511
rect 30822 507 30882 530
rect 30940 507 31000 530
rect 31058 507 31118 530
rect 31176 531 31472 591
rect 31176 507 31236 531
rect 31294 507 31354 531
rect 31412 507 31472 531
rect 31818 580 32052 596
rect 32425 586 32483 771
rect 30520 460 30651 477
rect 27492 110 27642 126
rect 27582 72 27642 110
rect 23497 28 23513 62
rect 23547 28 23563 62
rect 23497 12 23563 28
rect 23379 -55 23445 -39
rect 23379 -89 23395 -55
rect 23429 -89 23445 -55
rect 23379 -105 23445 -89
rect 23382 -127 23442 -105
rect 20957 -222 21017 -196
rect 18181 -422 18241 -396
rect 18299 -422 18359 -396
rect 18417 -422 18477 -396
rect 18535 -422 18595 -396
rect 20079 -422 20139 -396
rect 20197 -422 20257 -396
rect 20315 -422 20375 -396
rect 20433 -422 20493 -396
rect 24386 -154 24446 -128
rect 23382 -353 23442 -327
rect 25684 -154 25744 -128
rect 26284 -154 26344 -128
rect 28580 -87 28876 -51
rect 28580 -108 28640 -87
rect 28698 -108 28758 -87
rect 28816 -108 28876 -87
rect 28934 -88 29230 -52
rect 28934 -108 28994 -88
rect 29052 -108 29112 -88
rect 29170 -108 29230 -88
rect 29288 -88 29584 -52
rect 29288 -108 29348 -88
rect 29406 -108 29466 -88
rect 29524 -108 29584 -88
rect 27582 -154 27642 -128
rect 30520 -120 30580 460
rect 30822 81 30882 107
rect 30790 -60 30857 -53
rect 30940 -60 31000 107
rect 31058 81 31118 107
rect 31176 81 31236 107
rect 30790 -69 31000 -60
rect 30790 -103 30806 -69
rect 30840 -103 31000 -69
rect 30790 -119 31000 -103
rect 30520 -136 30671 -120
rect 30520 -170 30621 -136
rect 30655 -170 30671 -136
rect 30520 -186 30671 -170
rect 30520 -225 30580 -186
rect 30940 -225 31000 -119
rect 31294 -60 31354 107
rect 31412 81 31472 107
rect 31437 -60 31504 -53
rect 31294 -69 31504 -60
rect 31294 -103 31454 -69
rect 31488 -103 31504 -69
rect 31294 -119 31504 -103
rect 31056 -153 31122 -137
rect 31056 -187 31072 -153
rect 31106 -187 31122 -153
rect 31056 -203 31122 -187
rect 31174 -152 31240 -137
rect 31174 -186 31190 -152
rect 31224 -186 31240 -152
rect 31174 -202 31240 -186
rect 31058 -225 31118 -203
rect 31176 -225 31236 -202
rect 31294 -225 31354 -119
rect 31818 -121 31878 580
rect 32425 560 32485 586
rect 32543 560 32603 771
rect 32896 765 32956 797
rect 33014 771 33074 797
rect 33132 771 33192 797
rect 32893 749 32959 765
rect 32893 715 32909 749
rect 32943 715 32959 749
rect 32893 699 32959 715
rect 32775 632 32841 648
rect 32775 598 32791 632
rect 32825 598 32841 632
rect 32775 582 32841 598
rect 32778 560 32838 582
rect 32778 334 32838 360
rect 32425 138 32485 160
rect 32543 138 32603 160
rect 32422 122 32488 138
rect 32422 88 32438 122
rect 32472 88 32488 122
rect 32422 72 32488 88
rect 32540 122 32606 138
rect 32540 88 32556 122
rect 32590 88 32606 122
rect 32540 72 32606 88
rect 31728 -137 31878 -121
rect 31728 -171 31744 -137
rect 31778 -171 31878 -137
rect 31728 -187 31878 -171
rect 31818 -225 31878 -187
rect 24806 -354 24866 -328
rect 24924 -354 24984 -328
rect 25042 -354 25102 -328
rect 25160 -354 25220 -328
rect 26704 -354 26764 -328
rect 26822 -354 26882 -328
rect 26940 -354 27000 -328
rect 27058 -354 27118 -328
rect 28580 -334 28640 -308
rect 28698 -334 28758 -308
rect 28816 -334 28876 -308
rect 28934 -328 28994 -308
rect 28934 -334 28995 -328
rect 29052 -334 29112 -308
rect 29170 -334 29230 -308
rect 16404 -617 16464 -595
rect 16522 -617 16582 -595
rect 3316 -703 3382 -687
rect 16401 -633 16467 -617
rect 16401 -667 16417 -633
rect 16451 -667 16467 -633
rect 16401 -683 16467 -667
rect 16519 -633 16585 -617
rect 16519 -667 16535 -633
rect 16569 -667 16585 -633
rect 23029 -549 23089 -527
rect 23147 -549 23207 -527
rect 23026 -565 23092 -549
rect 23026 -599 23042 -565
rect 23076 -599 23092 -565
rect 23026 -615 23092 -599
rect 23144 -565 23210 -549
rect 23144 -599 23160 -565
rect 23194 -599 23210 -565
rect 28817 -519 28875 -334
rect 28817 -545 28877 -519
rect 28935 -545 28995 -334
rect 29288 -340 29348 -308
rect 29406 -334 29466 -308
rect 29524 -334 29584 -308
rect 29285 -356 29351 -340
rect 29285 -390 29301 -356
rect 29335 -390 29351 -356
rect 29285 -406 29351 -390
rect 30520 -451 30580 -425
rect 29167 -473 29233 -457
rect 29167 -507 29183 -473
rect 29217 -507 29233 -473
rect 29167 -523 29233 -507
rect 29170 -545 29230 -523
rect 23144 -615 23210 -599
rect 16519 -683 16585 -667
rect 31818 -451 31878 -425
rect 30940 -651 31000 -625
rect 31058 -651 31118 -625
rect 31176 -651 31236 -625
rect 31294 -651 31354 -625
rect 29170 -771 29230 -745
rect 28817 -967 28877 -945
rect 28935 -967 28995 -945
rect 28814 -983 28880 -967
rect 28814 -1017 28830 -983
rect 28864 -1017 28880 -983
rect 28814 -1033 28880 -1017
rect 28932 -983 28998 -967
rect 28932 -1017 28948 -983
rect 28982 -1017 28998 -983
rect 28932 -1033 28998 -1017
rect 38 -2099 334 -2063
rect 38 -2120 98 -2099
rect 156 -2120 216 -2099
rect 274 -2120 334 -2099
rect 392 -2100 688 -2064
rect 392 -2120 452 -2100
rect 510 -2120 570 -2100
rect 628 -2120 688 -2100
rect 746 -2100 1042 -2064
rect 746 -2120 806 -2100
rect 864 -2120 924 -2100
rect 982 -2120 1042 -2100
rect 5095 -2068 5161 -2052
rect 6225 -2062 6291 -2046
rect 5095 -2102 5111 -2068
rect 5145 -2075 5161 -2068
rect 5145 -2102 5670 -2075
rect 5095 -2118 5670 -2102
rect 6225 -2096 6241 -2062
rect 6275 -2071 6291 -2062
rect 6275 -2096 6812 -2071
rect 6225 -2114 6812 -2096
rect 5626 -2170 5670 -2118
rect 6768 -2166 6812 -2114
rect 11646 -2070 11712 -2054
rect 12776 -2064 12842 -2048
rect 11646 -2104 11662 -2070
rect 11696 -2077 11712 -2070
rect 11696 -2104 12221 -2077
rect 11646 -2120 12221 -2104
rect 12776 -2098 12792 -2064
rect 12826 -2073 12842 -2064
rect 12826 -2098 13363 -2073
rect 12776 -2116 13363 -2098
rect 5095 -2186 5568 -2170
rect 5095 -2220 5111 -2186
rect 5145 -2211 5568 -2186
rect 5145 -2212 5332 -2211
rect 5145 -2220 5161 -2212
rect 5095 -2236 5161 -2220
rect 5272 -2232 5332 -2212
rect 5390 -2232 5450 -2211
rect 5508 -2232 5568 -2211
rect 5626 -2211 5922 -2170
rect 5626 -2232 5686 -2211
rect 5744 -2232 5804 -2211
rect 5862 -2232 5922 -2211
rect 6225 -2182 6710 -2166
rect 6225 -2216 6241 -2182
rect 6275 -2207 6710 -2182
rect 6275 -2208 6474 -2207
rect 6275 -2216 6291 -2208
rect 6225 -2232 6291 -2216
rect 6414 -2228 6474 -2208
rect 6532 -2228 6592 -2207
rect 6650 -2228 6710 -2207
rect 6768 -2207 7064 -2166
rect 12177 -2172 12221 -2120
rect 13319 -2168 13363 -2116
rect 18301 -2069 18367 -2053
rect 19431 -2063 19497 -2047
rect 18301 -2103 18317 -2069
rect 18351 -2076 18367 -2069
rect 18351 -2103 18876 -2076
rect 18301 -2119 18876 -2103
rect 19431 -2097 19447 -2063
rect 19481 -2072 19497 -2063
rect 19481 -2097 20018 -2072
rect 19431 -2115 20018 -2097
rect 6768 -2228 6828 -2207
rect 6886 -2228 6946 -2207
rect 7004 -2228 7064 -2207
rect 11646 -2188 12119 -2172
rect 11646 -2222 11662 -2188
rect 11696 -2213 12119 -2188
rect 11696 -2214 11883 -2213
rect 11696 -2222 11712 -2214
rect 2947 -2283 3243 -2247
rect 2947 -2304 3007 -2283
rect 3065 -2304 3125 -2283
rect 3183 -2304 3243 -2283
rect 3301 -2284 3597 -2248
rect 3301 -2304 3361 -2284
rect 3419 -2304 3479 -2284
rect 3537 -2304 3597 -2284
rect 3655 -2284 3951 -2248
rect 3655 -2304 3715 -2284
rect 3773 -2304 3833 -2284
rect 3891 -2304 3951 -2284
rect 38 -2346 98 -2320
rect 156 -2346 216 -2320
rect 274 -2346 334 -2320
rect 392 -2340 452 -2320
rect 392 -2346 453 -2340
rect 510 -2346 570 -2320
rect 628 -2346 688 -2320
rect 275 -2531 333 -2346
rect 275 -2557 335 -2531
rect 393 -2557 453 -2346
rect 746 -2352 806 -2320
rect 864 -2346 924 -2320
rect 982 -2346 1042 -2320
rect 743 -2368 809 -2352
rect 743 -2402 759 -2368
rect 793 -2402 809 -2368
rect 743 -2418 809 -2402
rect 625 -2485 691 -2469
rect 625 -2519 641 -2485
rect 675 -2519 691 -2485
rect 625 -2535 691 -2519
rect 2947 -2530 3007 -2504
rect 3065 -2530 3125 -2504
rect 3183 -2530 3243 -2504
rect 3301 -2524 3361 -2504
rect 3301 -2530 3362 -2524
rect 3419 -2530 3479 -2504
rect 3537 -2530 3597 -2504
rect 628 -2557 688 -2535
rect 3184 -2715 3242 -2530
rect 3184 -2741 3244 -2715
rect 3302 -2741 3362 -2530
rect 3655 -2536 3715 -2504
rect 3773 -2530 3833 -2504
rect 3891 -2530 3951 -2504
rect 3652 -2552 3718 -2536
rect 3652 -2586 3668 -2552
rect 3702 -2586 3718 -2552
rect 3652 -2602 3718 -2586
rect 11646 -2238 11712 -2222
rect 11823 -2234 11883 -2214
rect 11941 -2234 12001 -2213
rect 12059 -2234 12119 -2213
rect 12177 -2213 12473 -2172
rect 12177 -2234 12237 -2213
rect 12295 -2234 12355 -2213
rect 12413 -2234 12473 -2213
rect 12776 -2184 13261 -2168
rect 12776 -2218 12792 -2184
rect 12826 -2209 13261 -2184
rect 12826 -2210 13025 -2209
rect 12826 -2218 12842 -2210
rect 12776 -2234 12842 -2218
rect 12965 -2230 13025 -2210
rect 13083 -2230 13143 -2209
rect 13201 -2230 13261 -2209
rect 13319 -2209 13615 -2168
rect 18832 -2171 18876 -2119
rect 19974 -2167 20018 -2115
rect 24923 -2068 24989 -2052
rect 26053 -2062 26119 -2046
rect 24923 -2102 24939 -2068
rect 24973 -2075 24989 -2068
rect 24973 -2102 25498 -2075
rect 24923 -2118 25498 -2102
rect 26053 -2096 26069 -2062
rect 26103 -2071 26119 -2062
rect 28651 -2007 28947 -1971
rect 28651 -2028 28711 -2007
rect 28769 -2028 28829 -2007
rect 28887 -2028 28947 -2007
rect 29005 -2008 29301 -1972
rect 29005 -2028 29065 -2008
rect 29123 -2028 29183 -2008
rect 29241 -2028 29301 -2008
rect 29359 -2008 29655 -1972
rect 29359 -2028 29419 -2008
rect 29477 -2028 29537 -2008
rect 29595 -2028 29655 -2008
rect 26103 -2096 26640 -2071
rect 26053 -2114 26640 -2096
rect 13319 -2230 13379 -2209
rect 13437 -2230 13497 -2209
rect 13555 -2230 13615 -2209
rect 18301 -2187 18774 -2171
rect 18301 -2221 18317 -2187
rect 18351 -2212 18774 -2187
rect 18351 -2213 18538 -2212
rect 18351 -2221 18367 -2213
rect 9498 -2285 9794 -2249
rect 9498 -2306 9558 -2285
rect 9616 -2306 9676 -2285
rect 9734 -2306 9794 -2285
rect 9852 -2286 10148 -2250
rect 9852 -2306 9912 -2286
rect 9970 -2306 10030 -2286
rect 10088 -2306 10148 -2286
rect 10206 -2286 10502 -2250
rect 10206 -2306 10266 -2286
rect 10324 -2306 10384 -2286
rect 10442 -2306 10502 -2286
rect 9498 -2532 9558 -2506
rect 9616 -2532 9676 -2506
rect 9734 -2532 9794 -2506
rect 9852 -2526 9912 -2506
rect 9852 -2532 9913 -2526
rect 9970 -2532 10030 -2506
rect 10088 -2532 10148 -2506
rect 5272 -2649 5332 -2632
rect 3534 -2669 3600 -2653
rect 3534 -2703 3550 -2669
rect 3584 -2703 3600 -2669
rect 3534 -2719 3600 -2703
rect 3537 -2741 3597 -2719
rect 5272 -2738 5333 -2649
rect 5390 -2658 5450 -2632
rect 5508 -2658 5568 -2632
rect 628 -2783 688 -2757
rect 275 -2979 335 -2957
rect 393 -2979 453 -2957
rect 272 -2995 338 -2979
rect 272 -3029 288 -2995
rect 322 -3029 338 -2995
rect 272 -3045 338 -3029
rect 390 -2995 456 -2979
rect 390 -3029 406 -2995
rect 440 -3029 456 -2995
rect 390 -3045 456 -3029
rect 5182 -2791 5333 -2738
rect 3537 -2967 3597 -2941
rect 5182 -3015 5242 -2791
rect 5626 -2833 5686 -2632
rect 5744 -2658 5804 -2632
rect 5862 -2658 5922 -2632
rect 6414 -2645 6474 -2628
rect 6414 -2734 6475 -2645
rect 6532 -2654 6592 -2628
rect 6650 -2654 6710 -2628
rect 5300 -2884 5686 -2833
rect 6324 -2787 6475 -2734
rect 5300 -3015 5360 -2884
rect 5415 -2942 5481 -2926
rect 5415 -2976 5431 -2942
rect 5465 -2976 5481 -2942
rect 5415 -2992 5481 -2976
rect 5418 -3015 5478 -2992
rect 5701 -3015 5761 -2989
rect 5819 -3015 5879 -2989
rect 5937 -3015 5997 -2989
rect 6324 -3011 6384 -2787
rect 6768 -2829 6828 -2628
rect 6886 -2654 6946 -2628
rect 7004 -2654 7064 -2628
rect 9735 -2717 9793 -2532
rect 9735 -2743 9795 -2717
rect 9853 -2743 9913 -2532
rect 10206 -2538 10266 -2506
rect 10324 -2532 10384 -2506
rect 10442 -2532 10502 -2506
rect 10203 -2554 10269 -2538
rect 10203 -2588 10219 -2554
rect 10253 -2588 10269 -2554
rect 10203 -2604 10269 -2588
rect 18301 -2237 18367 -2221
rect 18478 -2233 18538 -2213
rect 18596 -2233 18656 -2212
rect 18714 -2233 18774 -2212
rect 18832 -2212 19128 -2171
rect 18832 -2233 18892 -2212
rect 18950 -2233 19010 -2212
rect 19068 -2233 19128 -2212
rect 19431 -2183 19916 -2167
rect 19431 -2217 19447 -2183
rect 19481 -2208 19916 -2183
rect 19481 -2209 19680 -2208
rect 19481 -2217 19497 -2209
rect 19431 -2233 19497 -2217
rect 19620 -2229 19680 -2209
rect 19738 -2229 19798 -2208
rect 19856 -2229 19916 -2208
rect 19974 -2208 20270 -2167
rect 25454 -2170 25498 -2118
rect 26596 -2166 26640 -2114
rect 19974 -2229 20034 -2208
rect 20092 -2229 20152 -2208
rect 20210 -2229 20270 -2208
rect 24923 -2186 25396 -2170
rect 24923 -2220 24939 -2186
rect 24973 -2211 25396 -2186
rect 24973 -2212 25160 -2211
rect 24973 -2220 24989 -2212
rect 16153 -2284 16449 -2248
rect 16153 -2305 16213 -2284
rect 16271 -2305 16331 -2284
rect 16389 -2305 16449 -2284
rect 16507 -2285 16803 -2249
rect 16507 -2305 16567 -2285
rect 16625 -2305 16685 -2285
rect 16743 -2305 16803 -2285
rect 16861 -2285 17157 -2249
rect 16861 -2305 16921 -2285
rect 16979 -2305 17039 -2285
rect 17097 -2305 17157 -2285
rect 16153 -2531 16213 -2505
rect 16271 -2531 16331 -2505
rect 16389 -2531 16449 -2505
rect 16507 -2525 16567 -2505
rect 16507 -2531 16568 -2525
rect 16625 -2531 16685 -2505
rect 16743 -2531 16803 -2505
rect 11823 -2651 11883 -2634
rect 10085 -2671 10151 -2655
rect 10085 -2705 10101 -2671
rect 10135 -2705 10151 -2671
rect 10085 -2721 10151 -2705
rect 10088 -2743 10148 -2721
rect 11823 -2740 11884 -2651
rect 11941 -2660 12001 -2634
rect 12059 -2660 12119 -2634
rect 6442 -2880 6828 -2829
rect 6442 -3011 6502 -2880
rect 6557 -2938 6623 -2922
rect 6557 -2972 6573 -2938
rect 6607 -2972 6623 -2938
rect 6557 -2988 6623 -2972
rect 6560 -3011 6620 -2988
rect 6843 -3011 6903 -2985
rect 6961 -3011 7021 -2985
rect 7079 -3011 7139 -2985
rect 3184 -3163 3244 -3141
rect 3302 -3163 3362 -3141
rect 3181 -3179 3247 -3163
rect 3181 -3213 3197 -3179
rect 3231 -3213 3247 -3179
rect 3181 -3229 3247 -3213
rect 3299 -3179 3365 -3163
rect 3299 -3213 3315 -3179
rect 3349 -3213 3365 -3179
rect 3299 -3229 3365 -3213
rect 11733 -2793 11884 -2740
rect 10088 -2969 10148 -2943
rect 11733 -3017 11793 -2793
rect 12177 -2835 12237 -2634
rect 12295 -2660 12355 -2634
rect 12413 -2660 12473 -2634
rect 12965 -2647 13025 -2630
rect 12965 -2736 13026 -2647
rect 13083 -2656 13143 -2630
rect 13201 -2656 13261 -2630
rect 11851 -2886 12237 -2835
rect 12875 -2789 13026 -2736
rect 11851 -3017 11911 -2886
rect 11966 -2944 12032 -2928
rect 11966 -2978 11982 -2944
rect 12016 -2978 12032 -2944
rect 11966 -2994 12032 -2978
rect 11969 -3017 12029 -2994
rect 12252 -3017 12312 -2991
rect 12370 -3017 12430 -2991
rect 12488 -3017 12548 -2991
rect 12875 -3013 12935 -2789
rect 13319 -2831 13379 -2630
rect 13437 -2656 13497 -2630
rect 13555 -2656 13615 -2630
rect 16390 -2716 16448 -2531
rect 16390 -2742 16450 -2716
rect 16508 -2742 16568 -2531
rect 16861 -2537 16921 -2505
rect 16979 -2531 17039 -2505
rect 17097 -2531 17157 -2505
rect 16858 -2553 16924 -2537
rect 16858 -2587 16874 -2553
rect 16908 -2587 16924 -2553
rect 16858 -2603 16924 -2587
rect 24923 -2236 24989 -2220
rect 25100 -2232 25160 -2212
rect 25218 -2232 25278 -2211
rect 25336 -2232 25396 -2211
rect 25454 -2211 25750 -2170
rect 25454 -2232 25514 -2211
rect 25572 -2232 25632 -2211
rect 25690 -2232 25750 -2211
rect 26053 -2182 26538 -2166
rect 26053 -2216 26069 -2182
rect 26103 -2207 26538 -2182
rect 26103 -2208 26302 -2207
rect 26103 -2216 26119 -2208
rect 26053 -2232 26119 -2216
rect 26242 -2228 26302 -2208
rect 26360 -2228 26420 -2207
rect 26478 -2228 26538 -2207
rect 26596 -2207 26892 -2166
rect 26596 -2228 26656 -2207
rect 26714 -2228 26774 -2207
rect 26832 -2228 26892 -2207
rect 22775 -2283 23071 -2247
rect 22775 -2304 22835 -2283
rect 22893 -2304 22953 -2283
rect 23011 -2304 23071 -2283
rect 23129 -2284 23425 -2248
rect 23129 -2304 23189 -2284
rect 23247 -2304 23307 -2284
rect 23365 -2304 23425 -2284
rect 23483 -2284 23779 -2248
rect 23483 -2304 23543 -2284
rect 23601 -2304 23661 -2284
rect 23719 -2304 23779 -2284
rect 22775 -2530 22835 -2504
rect 22893 -2530 22953 -2504
rect 23011 -2530 23071 -2504
rect 23129 -2524 23189 -2504
rect 23129 -2530 23190 -2524
rect 23247 -2530 23307 -2504
rect 23365 -2530 23425 -2504
rect 18478 -2650 18538 -2633
rect 16740 -2670 16806 -2654
rect 16740 -2704 16756 -2670
rect 16790 -2704 16806 -2670
rect 16740 -2720 16806 -2704
rect 16743 -2742 16803 -2720
rect 18478 -2739 18539 -2650
rect 18596 -2659 18656 -2633
rect 18714 -2659 18774 -2633
rect 12993 -2882 13379 -2831
rect 12993 -3013 13053 -2882
rect 13108 -2940 13174 -2924
rect 13108 -2974 13124 -2940
rect 13158 -2974 13174 -2940
rect 13108 -2990 13174 -2974
rect 13111 -3013 13171 -2990
rect 13394 -3013 13454 -2987
rect 13512 -3013 13572 -2987
rect 13630 -3013 13690 -2987
rect 9735 -3165 9795 -3143
rect 9853 -3165 9913 -3143
rect 9732 -3181 9798 -3165
rect 5182 -3241 5242 -3215
rect 5300 -3241 5360 -3215
rect 5418 -3247 5478 -3215
rect 5701 -3247 5761 -3215
rect 5819 -3247 5879 -3215
rect 5937 -3247 5997 -3215
rect 6324 -3237 6384 -3211
rect 6442 -3237 6502 -3211
rect 5418 -3288 5997 -3247
rect 6560 -3243 6620 -3211
rect 6843 -3243 6903 -3211
rect 6961 -3243 7021 -3211
rect 7079 -3243 7139 -3211
rect 9732 -3215 9748 -3181
rect 9782 -3215 9798 -3181
rect 9732 -3231 9798 -3215
rect 9850 -3181 9916 -3165
rect 9850 -3215 9866 -3181
rect 9900 -3215 9916 -3181
rect 9850 -3231 9916 -3215
rect 18388 -2792 18539 -2739
rect 16743 -2968 16803 -2942
rect 18388 -3016 18448 -2792
rect 18832 -2834 18892 -2633
rect 18950 -2659 19010 -2633
rect 19068 -2659 19128 -2633
rect 19620 -2646 19680 -2629
rect 19620 -2735 19681 -2646
rect 19738 -2655 19798 -2629
rect 19856 -2655 19916 -2629
rect 18506 -2885 18892 -2834
rect 19530 -2788 19681 -2735
rect 18506 -3016 18566 -2885
rect 18621 -2943 18687 -2927
rect 18621 -2977 18637 -2943
rect 18671 -2977 18687 -2943
rect 18621 -2993 18687 -2977
rect 18624 -3016 18684 -2993
rect 18907 -3016 18967 -2990
rect 19025 -3016 19085 -2990
rect 19143 -3016 19203 -2990
rect 19530 -3012 19590 -2788
rect 19974 -2830 20034 -2629
rect 20092 -2655 20152 -2629
rect 20210 -2655 20270 -2629
rect 23012 -2715 23070 -2530
rect 23012 -2741 23072 -2715
rect 23130 -2741 23190 -2530
rect 23483 -2536 23543 -2504
rect 23601 -2530 23661 -2504
rect 23719 -2530 23779 -2504
rect 23480 -2552 23546 -2536
rect 23480 -2586 23496 -2552
rect 23530 -2586 23546 -2552
rect 23480 -2602 23546 -2586
rect 28651 -2254 28711 -2228
rect 28769 -2254 28829 -2228
rect 28887 -2254 28947 -2228
rect 29005 -2248 29065 -2228
rect 29005 -2254 29066 -2248
rect 29123 -2254 29183 -2228
rect 29241 -2254 29301 -2228
rect 28888 -2439 28946 -2254
rect 28888 -2465 28948 -2439
rect 29006 -2465 29066 -2254
rect 29359 -2260 29419 -2228
rect 29477 -2254 29537 -2228
rect 29595 -2254 29655 -2228
rect 29356 -2276 29422 -2260
rect 29356 -2310 29372 -2276
rect 29406 -2310 29422 -2276
rect 30879 -2280 31175 -2229
rect 30879 -2295 30939 -2280
rect 30997 -2295 31057 -2280
rect 31115 -2295 31175 -2280
rect 31233 -2295 31293 -2269
rect 31351 -2295 31411 -2269
rect 31469 -2295 31529 -2269
rect 29356 -2326 29422 -2310
rect 29238 -2393 29304 -2377
rect 29238 -2427 29254 -2393
rect 29288 -2427 29304 -2393
rect 29238 -2443 29304 -2427
rect 29241 -2465 29301 -2443
rect 25100 -2649 25160 -2632
rect 23362 -2669 23428 -2653
rect 23362 -2703 23378 -2669
rect 23412 -2703 23428 -2669
rect 23362 -2719 23428 -2703
rect 23365 -2741 23425 -2719
rect 25100 -2738 25161 -2649
rect 25218 -2658 25278 -2632
rect 25336 -2658 25396 -2632
rect 19648 -2881 20034 -2830
rect 19648 -3012 19708 -2881
rect 19763 -2939 19829 -2923
rect 19763 -2973 19779 -2939
rect 19813 -2973 19829 -2939
rect 19763 -2989 19829 -2973
rect 19766 -3012 19826 -2989
rect 20049 -3012 20109 -2986
rect 20167 -3012 20227 -2986
rect 20285 -3012 20345 -2986
rect 16390 -3164 16450 -3142
rect 16508 -3164 16568 -3142
rect 16387 -3180 16453 -3164
rect 11733 -3243 11793 -3217
rect 11851 -3243 11911 -3217
rect 6560 -3284 7139 -3243
rect 11969 -3249 12029 -3217
rect 12252 -3249 12312 -3217
rect 12370 -3249 12430 -3217
rect 12488 -3249 12548 -3217
rect 12875 -3239 12935 -3213
rect 12993 -3239 13053 -3213
rect 11969 -3290 12548 -3249
rect 13111 -3245 13171 -3213
rect 13394 -3245 13454 -3213
rect 13512 -3245 13572 -3213
rect 13630 -3245 13690 -3213
rect 16387 -3214 16403 -3180
rect 16437 -3214 16453 -3180
rect 16387 -3230 16453 -3214
rect 16505 -3180 16571 -3164
rect 16505 -3214 16521 -3180
rect 16555 -3214 16571 -3180
rect 16505 -3230 16571 -3214
rect 25010 -2791 25161 -2738
rect 23365 -2967 23425 -2941
rect 25010 -3015 25070 -2791
rect 25454 -2833 25514 -2632
rect 25572 -2658 25632 -2632
rect 25690 -2658 25750 -2632
rect 26242 -2645 26302 -2628
rect 26242 -2734 26303 -2645
rect 26360 -2654 26420 -2628
rect 26478 -2654 26538 -2628
rect 25128 -2884 25514 -2833
rect 26152 -2787 26303 -2734
rect 25128 -3015 25188 -2884
rect 25243 -2942 25309 -2926
rect 25243 -2976 25259 -2942
rect 25293 -2976 25309 -2942
rect 25243 -2992 25309 -2976
rect 25246 -3015 25306 -2992
rect 25529 -3015 25589 -2989
rect 25647 -3015 25707 -2989
rect 25765 -3015 25825 -2989
rect 26152 -3011 26212 -2787
rect 26596 -2829 26656 -2628
rect 26714 -2654 26774 -2628
rect 26832 -2654 26892 -2628
rect 26270 -2880 26656 -2829
rect 30395 -2495 30455 -2469
rect 30513 -2495 30573 -2469
rect 30631 -2495 30691 -2469
rect 29241 -2691 29301 -2665
rect 31716 -2478 32012 -2427
rect 31716 -2495 31776 -2478
rect 31834 -2495 31894 -2478
rect 31952 -2495 32012 -2478
rect 32188 -2477 32484 -2441
rect 32188 -2498 32248 -2477
rect 32306 -2498 32366 -2477
rect 32424 -2498 32484 -2477
rect 32542 -2478 32838 -2442
rect 32542 -2498 32602 -2478
rect 32660 -2498 32720 -2478
rect 32778 -2498 32838 -2478
rect 32896 -2478 33192 -2442
rect 32896 -2498 32956 -2478
rect 33014 -2498 33074 -2478
rect 33132 -2498 33192 -2478
rect 30395 -2712 30455 -2695
rect 30513 -2712 30573 -2695
rect 30631 -2712 30691 -2695
rect 30879 -2712 30939 -2695
rect 30395 -2763 30939 -2712
rect 30997 -2721 31057 -2695
rect 31115 -2721 31175 -2695
rect 31233 -2714 31293 -2695
rect 31351 -2714 31411 -2695
rect 31469 -2714 31529 -2695
rect 31716 -2714 31776 -2695
rect 31834 -2714 31894 -2695
rect 26270 -3011 26330 -2880
rect 28888 -2887 28948 -2865
rect 29006 -2887 29066 -2865
rect 28885 -2903 28951 -2887
rect 26385 -2938 26451 -2922
rect 26385 -2972 26401 -2938
rect 26435 -2972 26451 -2938
rect 28885 -2937 28901 -2903
rect 28935 -2937 28951 -2903
rect 28885 -2953 28951 -2937
rect 29003 -2903 29069 -2887
rect 29003 -2937 29019 -2903
rect 29053 -2937 29069 -2903
rect 29003 -2953 29069 -2937
rect 26385 -2988 26451 -2972
rect 30520 -2967 30580 -2763
rect 31233 -2765 31776 -2714
rect 31818 -2721 31894 -2714
rect 31952 -2721 32012 -2695
rect 31818 -2765 31893 -2721
rect 32188 -2724 32248 -2698
rect 32306 -2724 32366 -2698
rect 32424 -2724 32484 -2698
rect 32542 -2718 32602 -2698
rect 32542 -2724 32603 -2718
rect 32660 -2724 32720 -2698
rect 32778 -2724 32838 -2698
rect 31818 -2847 31878 -2765
rect 31818 -2865 32052 -2847
rect 31818 -2899 32001 -2865
rect 32035 -2899 32052 -2865
rect 30822 -2965 31118 -2905
rect 26388 -3011 26448 -2988
rect 26671 -3011 26731 -2985
rect 26789 -3011 26849 -2985
rect 26907 -3011 26967 -2985
rect 23012 -3163 23072 -3141
rect 23130 -3163 23190 -3141
rect 23009 -3179 23075 -3163
rect 18388 -3242 18448 -3216
rect 18506 -3242 18566 -3216
rect 13111 -3286 13690 -3245
rect 18624 -3248 18684 -3216
rect 18907 -3248 18967 -3216
rect 19025 -3248 19085 -3216
rect 19143 -3248 19203 -3216
rect 19530 -3238 19590 -3212
rect 19648 -3238 19708 -3212
rect 18624 -3289 19203 -3248
rect 19766 -3244 19826 -3212
rect 20049 -3244 20109 -3212
rect 20167 -3244 20227 -3212
rect 20285 -3244 20345 -3212
rect 23009 -3213 23025 -3179
rect 23059 -3213 23075 -3179
rect 23009 -3229 23075 -3213
rect 23127 -3179 23193 -3163
rect 23127 -3213 23143 -3179
rect 23177 -3213 23193 -3179
rect 23127 -3229 23193 -3213
rect 30520 -2984 30651 -2967
rect 30520 -3018 30601 -2984
rect 30635 -3018 30651 -2984
rect 30822 -2988 30882 -2965
rect 30940 -2988 31000 -2965
rect 31058 -2988 31118 -2965
rect 31176 -2964 31472 -2904
rect 31176 -2988 31236 -2964
rect 31294 -2988 31354 -2964
rect 31412 -2988 31472 -2964
rect 31818 -2915 32052 -2899
rect 32425 -2909 32483 -2724
rect 30520 -3035 30651 -3018
rect 25010 -3241 25070 -3215
rect 25128 -3241 25188 -3215
rect 19766 -3285 20345 -3244
rect 25246 -3247 25306 -3215
rect 25529 -3247 25589 -3215
rect 25647 -3247 25707 -3215
rect 25765 -3247 25825 -3215
rect 26152 -3237 26212 -3211
rect 26270 -3237 26330 -3211
rect 25246 -3288 25825 -3247
rect 26388 -3243 26448 -3211
rect 26671 -3243 26731 -3211
rect 26789 -3243 26849 -3211
rect 26907 -3243 26967 -3211
rect 26388 -3284 26967 -3243
rect 30520 -3615 30580 -3035
rect 30822 -3414 30882 -3388
rect 30790 -3555 30857 -3548
rect 30940 -3555 31000 -3388
rect 31058 -3414 31118 -3388
rect 31176 -3414 31236 -3388
rect 30790 -3564 31000 -3555
rect 30790 -3598 30806 -3564
rect 30840 -3598 31000 -3564
rect 30790 -3614 31000 -3598
rect 30520 -3631 30671 -3615
rect 30520 -3665 30621 -3631
rect 30655 -3665 30671 -3631
rect 30520 -3681 30671 -3665
rect 30520 -3720 30580 -3681
rect 30940 -3720 31000 -3614
rect 31294 -3555 31354 -3388
rect 31412 -3414 31472 -3388
rect 31437 -3555 31504 -3548
rect 31294 -3564 31504 -3555
rect 31294 -3598 31454 -3564
rect 31488 -3598 31504 -3564
rect 31294 -3614 31504 -3598
rect 31056 -3648 31122 -3632
rect 31056 -3682 31072 -3648
rect 31106 -3682 31122 -3648
rect 31056 -3698 31122 -3682
rect 31174 -3647 31240 -3632
rect 31174 -3681 31190 -3647
rect 31224 -3681 31240 -3647
rect 31174 -3697 31240 -3681
rect 31058 -3720 31118 -3698
rect 31176 -3720 31236 -3697
rect 31294 -3720 31354 -3614
rect 31818 -3616 31878 -2915
rect 32425 -2935 32485 -2909
rect 32543 -2935 32603 -2724
rect 32896 -2730 32956 -2698
rect 33014 -2724 33074 -2698
rect 33132 -2724 33192 -2698
rect 32893 -2746 32959 -2730
rect 32893 -2780 32909 -2746
rect 32943 -2780 32959 -2746
rect 32893 -2796 32959 -2780
rect 32775 -2863 32841 -2847
rect 32775 -2897 32791 -2863
rect 32825 -2897 32841 -2863
rect 32775 -2913 32841 -2897
rect 32778 -2935 32838 -2913
rect 32778 -3161 32838 -3135
rect 32425 -3357 32485 -3335
rect 32543 -3357 32603 -3335
rect 32422 -3373 32488 -3357
rect 32422 -3407 32438 -3373
rect 32472 -3407 32488 -3373
rect 32422 -3423 32488 -3407
rect 32540 -3373 32606 -3357
rect 32540 -3407 32556 -3373
rect 32590 -3407 32606 -3373
rect 32540 -3423 32606 -3407
rect 31728 -3632 31878 -3616
rect 31728 -3666 31744 -3632
rect 31778 -3666 31878 -3632
rect 31728 -3682 31878 -3666
rect 31818 -3720 31878 -3682
rect 2961 -3933 3257 -3897
rect 2961 -3954 3021 -3933
rect 3079 -3954 3139 -3933
rect 3197 -3954 3257 -3933
rect 3315 -3934 3611 -3898
rect 3315 -3954 3375 -3934
rect 3433 -3954 3493 -3934
rect 3551 -3954 3611 -3934
rect 3669 -3934 3965 -3898
rect 3669 -3954 3729 -3934
rect 3787 -3954 3847 -3934
rect 3905 -3954 3965 -3934
rect 9512 -3935 9808 -3899
rect 9512 -3956 9572 -3935
rect 9630 -3956 9690 -3935
rect 9748 -3956 9808 -3935
rect 9866 -3936 10162 -3900
rect 9866 -3956 9926 -3936
rect 9984 -3956 10044 -3936
rect 10102 -3956 10162 -3936
rect 10220 -3936 10516 -3900
rect 10220 -3956 10280 -3936
rect 10338 -3956 10398 -3936
rect 10456 -3956 10516 -3936
rect 2961 -4180 3021 -4154
rect 3079 -4180 3139 -4154
rect 3197 -4180 3257 -4154
rect 3315 -4174 3375 -4154
rect 3315 -4180 3376 -4174
rect 3433 -4180 3493 -4154
rect 3551 -4180 3611 -4154
rect 3198 -4365 3256 -4180
rect 3198 -4391 3258 -4365
rect 3316 -4391 3376 -4180
rect 3669 -4186 3729 -4154
rect 3787 -4180 3847 -4154
rect 3905 -4180 3965 -4154
rect 16167 -3934 16463 -3898
rect 16167 -3955 16227 -3934
rect 16285 -3955 16345 -3934
rect 16403 -3955 16463 -3934
rect 16521 -3935 16817 -3899
rect 16521 -3955 16581 -3935
rect 16639 -3955 16699 -3935
rect 16757 -3955 16817 -3935
rect 16875 -3935 17171 -3899
rect 16875 -3955 16935 -3935
rect 16993 -3955 17053 -3935
rect 17111 -3955 17171 -3935
rect 22789 -3933 23085 -3897
rect 22789 -3954 22849 -3933
rect 22907 -3954 22967 -3933
rect 23025 -3954 23085 -3933
rect 23143 -3934 23439 -3898
rect 23143 -3954 23203 -3934
rect 23261 -3954 23321 -3934
rect 23379 -3954 23439 -3934
rect 23497 -3934 23793 -3898
rect 23497 -3954 23557 -3934
rect 23615 -3954 23675 -3934
rect 23733 -3954 23793 -3934
rect 30520 -3946 30580 -3920
rect 31818 -3946 31878 -3920
rect 30940 -4146 31000 -4120
rect 31058 -4146 31118 -4120
rect 31176 -4146 31236 -4120
rect 31294 -4146 31354 -4120
rect 9512 -4182 9572 -4156
rect 9630 -4182 9690 -4156
rect 9748 -4182 9808 -4156
rect 9866 -4176 9926 -4156
rect 9866 -4182 9927 -4176
rect 9984 -4182 10044 -4156
rect 10102 -4182 10162 -4156
rect 3666 -4202 3732 -4186
rect 3666 -4236 3682 -4202
rect 3716 -4236 3732 -4202
rect 3666 -4252 3732 -4236
rect 3548 -4319 3614 -4303
rect 3548 -4353 3564 -4319
rect 3598 -4353 3614 -4319
rect 3548 -4369 3614 -4353
rect 4909 -4356 5205 -4305
rect 3551 -4391 3611 -4369
rect 4909 -4371 4969 -4356
rect 5027 -4371 5087 -4356
rect 5145 -4371 5205 -4356
rect 5263 -4371 5323 -4345
rect 5381 -4371 5441 -4345
rect 5499 -4371 5559 -4345
rect 6807 -4356 7103 -4305
rect 6807 -4371 6867 -4356
rect 6925 -4371 6985 -4356
rect 7043 -4371 7103 -4356
rect 7161 -4371 7221 -4345
rect 7279 -4371 7339 -4345
rect 7397 -4371 7457 -4345
rect 9749 -4367 9807 -4182
rect 4425 -4571 4485 -4545
rect 4543 -4571 4603 -4545
rect 4661 -4571 4721 -4545
rect 3551 -4617 3611 -4591
rect 3198 -4813 3258 -4791
rect 3316 -4807 3376 -4791
rect 54 -4859 350 -4823
rect 54 -4880 114 -4859
rect 172 -4880 232 -4859
rect 290 -4880 350 -4859
rect 408 -4860 704 -4824
rect 408 -4880 468 -4860
rect 526 -4880 586 -4860
rect 644 -4880 704 -4860
rect 762 -4860 1058 -4824
rect 762 -4880 822 -4860
rect 880 -4880 940 -4860
rect 998 -4880 1058 -4860
rect 3195 -4829 3261 -4813
rect 3195 -4863 3211 -4829
rect 3245 -4863 3261 -4829
rect 3195 -4879 3261 -4863
rect 3310 -4829 3384 -4807
rect 3310 -4863 3329 -4829
rect 3363 -4863 3384 -4829
rect 5746 -4554 6042 -4503
rect 5746 -4571 5806 -4554
rect 5864 -4571 5924 -4554
rect 5982 -4571 6042 -4554
rect 6323 -4571 6383 -4545
rect 6441 -4571 6501 -4545
rect 6559 -4571 6619 -4545
rect 9749 -4393 9809 -4367
rect 9867 -4393 9927 -4182
rect 10220 -4188 10280 -4156
rect 10338 -4182 10398 -4156
rect 10456 -4182 10516 -4156
rect 16167 -4181 16227 -4155
rect 16285 -4181 16345 -4155
rect 16403 -4181 16463 -4155
rect 16521 -4175 16581 -4155
rect 16521 -4181 16582 -4175
rect 16639 -4181 16699 -4155
rect 16757 -4181 16817 -4155
rect 10217 -4204 10283 -4188
rect 10217 -4238 10233 -4204
rect 10267 -4238 10283 -4204
rect 10217 -4254 10283 -4238
rect 10099 -4321 10165 -4305
rect 10099 -4355 10115 -4321
rect 10149 -4355 10165 -4321
rect 10099 -4371 10165 -4355
rect 11460 -4358 11756 -4307
rect 10102 -4393 10162 -4371
rect 11460 -4373 11520 -4358
rect 11578 -4373 11638 -4358
rect 11696 -4373 11756 -4358
rect 11814 -4373 11874 -4347
rect 11932 -4373 11992 -4347
rect 12050 -4373 12110 -4347
rect 13358 -4358 13654 -4307
rect 13358 -4373 13418 -4358
rect 13476 -4373 13536 -4358
rect 13594 -4373 13654 -4358
rect 13712 -4373 13772 -4347
rect 13830 -4373 13890 -4347
rect 13948 -4373 14008 -4347
rect 16404 -4366 16462 -4181
rect 7644 -4554 7940 -4503
rect 7644 -4571 7704 -4554
rect 7762 -4571 7822 -4554
rect 7880 -4571 7940 -4554
rect 4425 -4788 4485 -4771
rect 4543 -4788 4603 -4771
rect 4661 -4788 4721 -4771
rect 4909 -4788 4969 -4771
rect 4425 -4839 4969 -4788
rect 5027 -4797 5087 -4771
rect 5145 -4797 5205 -4771
rect 5263 -4790 5323 -4771
rect 5381 -4790 5441 -4771
rect 5499 -4790 5559 -4771
rect 5746 -4790 5806 -4771
rect 5864 -4790 5924 -4771
rect 3310 -4920 3384 -4863
rect 4550 -4920 4610 -4839
rect 5263 -4841 5806 -4790
rect 5848 -4797 5924 -4790
rect 5982 -4797 6042 -4771
rect 6323 -4788 6383 -4771
rect 6441 -4788 6501 -4771
rect 6559 -4788 6619 -4771
rect 6807 -4788 6867 -4771
rect 5848 -4841 5923 -4797
rect 6323 -4839 6867 -4788
rect 6925 -4797 6985 -4771
rect 7043 -4797 7103 -4771
rect 7161 -4790 7221 -4771
rect 7279 -4790 7339 -4771
rect 7397 -4790 7457 -4771
rect 7644 -4790 7704 -4771
rect 7762 -4790 7822 -4771
rect 3310 -4945 4610 -4920
rect 3309 -4993 4610 -4945
rect 5848 -4961 5908 -4841
rect 54 -5106 114 -5080
rect 172 -5106 232 -5080
rect 290 -5106 350 -5080
rect 408 -5100 468 -5080
rect 408 -5106 469 -5100
rect 526 -5106 586 -5080
rect 644 -5106 704 -5080
rect 291 -5291 349 -5106
rect 291 -5317 351 -5291
rect 409 -5317 469 -5106
rect 762 -5112 822 -5080
rect 880 -5106 940 -5080
rect 998 -5106 1058 -5080
rect 759 -5128 825 -5112
rect 759 -5162 775 -5128
rect 809 -5162 825 -5128
rect 759 -5178 825 -5162
rect 641 -5245 707 -5229
rect 641 -5279 657 -5245
rect 691 -5279 707 -5245
rect 641 -5295 707 -5279
rect 644 -5317 704 -5295
rect 644 -5543 704 -5517
rect 2956 -5537 3252 -5501
rect 2956 -5558 3016 -5537
rect 3074 -5558 3134 -5537
rect 3192 -5558 3252 -5537
rect 3310 -5538 3606 -5502
rect 3310 -5558 3370 -5538
rect 3428 -5558 3488 -5538
rect 3546 -5558 3606 -5538
rect 3664 -5538 3960 -5502
rect 3664 -5558 3724 -5538
rect 3782 -5558 3842 -5538
rect 3900 -5558 3960 -5538
rect 291 -5739 351 -5717
rect 409 -5739 469 -5717
rect 288 -5755 354 -5739
rect 288 -5789 304 -5755
rect 338 -5789 354 -5755
rect 288 -5805 354 -5789
rect 406 -5755 472 -5739
rect 406 -5789 422 -5755
rect 456 -5789 472 -5755
rect 4550 -5691 4610 -4993
rect 4852 -5041 5148 -4981
rect 4852 -5064 4912 -5041
rect 4970 -5064 5030 -5041
rect 5088 -5064 5148 -5041
rect 5206 -5040 5502 -4980
rect 5847 -4981 5908 -4961
rect 5206 -5064 5266 -5040
rect 5324 -5064 5384 -5040
rect 5442 -5064 5502 -5040
rect 5828 -4997 5908 -4981
rect 5828 -5031 5843 -4997
rect 5877 -5031 5908 -4997
rect 5828 -5047 5908 -5031
rect 5847 -5070 5908 -5047
rect 5848 -5216 5908 -5070
rect 5847 -5389 5908 -5216
rect 4852 -5490 4912 -5464
rect 4820 -5631 4887 -5624
rect 4970 -5631 5030 -5464
rect 5088 -5490 5148 -5464
rect 5206 -5490 5266 -5464
rect 4820 -5640 5030 -5631
rect 4820 -5674 4836 -5640
rect 4870 -5674 5030 -5640
rect 4820 -5690 5030 -5674
rect 4550 -5707 4701 -5691
rect 4550 -5741 4651 -5707
rect 4685 -5741 4701 -5707
rect 4550 -5757 4701 -5741
rect 2956 -5784 3016 -5758
rect 3074 -5784 3134 -5758
rect 3192 -5784 3252 -5758
rect 3310 -5778 3370 -5758
rect 3310 -5784 3371 -5778
rect 3428 -5784 3488 -5758
rect 3546 -5784 3606 -5758
rect 406 -5805 472 -5789
rect 3193 -5969 3251 -5784
rect 3193 -5995 3253 -5969
rect 3311 -5995 3371 -5784
rect 3664 -5790 3724 -5758
rect 3782 -5784 3842 -5758
rect 3900 -5784 3960 -5758
rect 3661 -5806 3727 -5790
rect 4550 -5796 4610 -5757
rect 4970 -5796 5030 -5690
rect 5324 -5631 5384 -5464
rect 5442 -5490 5502 -5464
rect 5467 -5631 5534 -5624
rect 5324 -5640 5534 -5631
rect 5324 -5674 5484 -5640
rect 5518 -5674 5534 -5640
rect 5324 -5690 5534 -5674
rect 5086 -5724 5152 -5708
rect 5086 -5758 5102 -5724
rect 5136 -5758 5152 -5724
rect 5086 -5774 5152 -5758
rect 5204 -5723 5270 -5708
rect 5204 -5757 5220 -5723
rect 5254 -5757 5270 -5723
rect 5204 -5773 5270 -5757
rect 5088 -5796 5148 -5774
rect 5206 -5796 5266 -5773
rect 5324 -5796 5384 -5690
rect 5848 -5692 5908 -5389
rect 5758 -5708 5908 -5692
rect 5758 -5742 5774 -5708
rect 5808 -5742 5908 -5708
rect 5758 -5758 5908 -5742
rect 5848 -5796 5908 -5758
rect 6448 -5497 6508 -4839
rect 7161 -4841 7704 -4790
rect 7746 -4797 7822 -4790
rect 7880 -4797 7940 -4771
rect 10976 -4573 11036 -4547
rect 11094 -4573 11154 -4547
rect 11212 -4573 11272 -4547
rect 10102 -4619 10162 -4593
rect 7746 -4841 7821 -4797
rect 9749 -4815 9809 -4793
rect 9867 -4809 9927 -4793
rect 9746 -4831 9812 -4815
rect 6750 -5041 7046 -4981
rect 6750 -5064 6810 -5041
rect 6868 -5064 6928 -5041
rect 6986 -5064 7046 -5041
rect 7104 -5040 7400 -4980
rect 7104 -5064 7164 -5040
rect 7222 -5064 7282 -5040
rect 7340 -5064 7400 -5040
rect 7746 -4994 7806 -4841
rect 9746 -4865 9762 -4831
rect 9796 -4865 9812 -4831
rect 9746 -4881 9812 -4865
rect 9861 -4831 9935 -4809
rect 9861 -4865 9880 -4831
rect 9914 -4865 9935 -4831
rect 12297 -4556 12593 -4505
rect 12297 -4573 12357 -4556
rect 12415 -4573 12475 -4556
rect 12533 -4573 12593 -4556
rect 12874 -4573 12934 -4547
rect 12992 -4573 13052 -4547
rect 13110 -4573 13170 -4547
rect 16404 -4392 16464 -4366
rect 16522 -4392 16582 -4181
rect 16875 -4187 16935 -4155
rect 16993 -4181 17053 -4155
rect 17111 -4181 17171 -4155
rect 22789 -4180 22849 -4154
rect 22907 -4180 22967 -4154
rect 23025 -4180 23085 -4154
rect 23143 -4174 23203 -4154
rect 23143 -4180 23204 -4174
rect 23261 -4180 23321 -4154
rect 23379 -4180 23439 -4154
rect 16872 -4203 16938 -4187
rect 16872 -4237 16888 -4203
rect 16922 -4237 16938 -4203
rect 16872 -4253 16938 -4237
rect 16754 -4320 16820 -4304
rect 16754 -4354 16770 -4320
rect 16804 -4354 16820 -4320
rect 16754 -4370 16820 -4354
rect 18115 -4357 18411 -4306
rect 16757 -4392 16817 -4370
rect 18115 -4372 18175 -4357
rect 18233 -4372 18293 -4357
rect 18351 -4372 18411 -4357
rect 18469 -4372 18529 -4346
rect 18587 -4372 18647 -4346
rect 18705 -4372 18765 -4346
rect 20013 -4357 20309 -4306
rect 20013 -4372 20073 -4357
rect 20131 -4372 20191 -4357
rect 20249 -4372 20309 -4357
rect 20367 -4372 20427 -4346
rect 20485 -4372 20545 -4346
rect 20603 -4372 20663 -4346
rect 23026 -4365 23084 -4180
rect 14195 -4556 14491 -4505
rect 14195 -4573 14255 -4556
rect 14313 -4573 14373 -4556
rect 14431 -4573 14491 -4556
rect 10976 -4790 11036 -4773
rect 11094 -4790 11154 -4773
rect 11212 -4790 11272 -4773
rect 11460 -4790 11520 -4773
rect 10976 -4841 11520 -4790
rect 11578 -4799 11638 -4773
rect 11696 -4799 11756 -4773
rect 11814 -4792 11874 -4773
rect 11932 -4792 11992 -4773
rect 12050 -4792 12110 -4773
rect 12297 -4792 12357 -4773
rect 12415 -4792 12475 -4773
rect 9861 -4922 9935 -4865
rect 11101 -4922 11161 -4841
rect 11814 -4843 12357 -4792
rect 12399 -4799 12475 -4792
rect 12533 -4799 12593 -4773
rect 12874 -4790 12934 -4773
rect 12992 -4790 13052 -4773
rect 13110 -4790 13170 -4773
rect 13358 -4790 13418 -4773
rect 12399 -4843 12474 -4799
rect 12874 -4841 13418 -4790
rect 13476 -4799 13536 -4773
rect 13594 -4799 13654 -4773
rect 13712 -4792 13772 -4773
rect 13830 -4792 13890 -4773
rect 13948 -4792 14008 -4773
rect 14195 -4792 14255 -4773
rect 14313 -4792 14373 -4773
rect 9861 -4947 11161 -4922
rect 7746 -5018 8000 -4994
rect 9860 -4995 11161 -4947
rect 12399 -4963 12459 -4843
rect 7746 -5052 7950 -5018
rect 7984 -5052 8000 -5018
rect 7746 -5068 8000 -5052
rect 6750 -5490 6810 -5464
rect 6448 -5513 6515 -5497
rect 6448 -5547 6464 -5513
rect 6498 -5547 6515 -5513
rect 6448 -5563 6515 -5547
rect 6448 -5691 6508 -5563
rect 6718 -5631 6785 -5624
rect 6868 -5631 6928 -5464
rect 6986 -5490 7046 -5464
rect 7104 -5490 7164 -5464
rect 6718 -5640 6928 -5631
rect 6718 -5674 6734 -5640
rect 6768 -5674 6928 -5640
rect 6718 -5690 6928 -5674
rect 6448 -5707 6599 -5691
rect 6448 -5741 6549 -5707
rect 6583 -5741 6599 -5707
rect 6448 -5757 6599 -5741
rect 6448 -5796 6508 -5757
rect 6868 -5796 6928 -5690
rect 7222 -5631 7282 -5464
rect 7340 -5490 7400 -5464
rect 7363 -5630 7430 -5623
rect 7357 -5631 7430 -5630
rect 7222 -5639 7430 -5631
rect 7222 -5673 7380 -5639
rect 7414 -5673 7430 -5639
rect 7222 -5689 7430 -5673
rect 7222 -5690 7419 -5689
rect 6984 -5724 7050 -5708
rect 6984 -5758 7000 -5724
rect 7034 -5758 7050 -5724
rect 6984 -5774 7050 -5758
rect 7102 -5723 7168 -5708
rect 7102 -5757 7118 -5723
rect 7152 -5757 7168 -5723
rect 7102 -5773 7168 -5757
rect 6986 -5796 7046 -5774
rect 7104 -5796 7164 -5773
rect 7222 -5796 7282 -5690
rect 7746 -5692 7806 -5068
rect 9507 -5539 9803 -5503
rect 9507 -5560 9567 -5539
rect 9625 -5560 9685 -5539
rect 9743 -5560 9803 -5539
rect 9861 -5540 10157 -5504
rect 9861 -5560 9921 -5540
rect 9979 -5560 10039 -5540
rect 10097 -5560 10157 -5540
rect 10215 -5540 10511 -5504
rect 10215 -5560 10275 -5540
rect 10333 -5560 10393 -5540
rect 10451 -5560 10511 -5540
rect 7656 -5708 7806 -5692
rect 7656 -5742 7672 -5708
rect 7706 -5742 7806 -5708
rect 7656 -5758 7806 -5742
rect 7746 -5796 7806 -5758
rect 11101 -5693 11161 -4995
rect 11403 -5043 11699 -4983
rect 11403 -5066 11463 -5043
rect 11521 -5066 11581 -5043
rect 11639 -5066 11699 -5043
rect 11757 -5042 12053 -4982
rect 12398 -4983 12459 -4963
rect 11757 -5066 11817 -5042
rect 11875 -5066 11935 -5042
rect 11993 -5066 12053 -5042
rect 12379 -4999 12459 -4983
rect 12379 -5033 12394 -4999
rect 12428 -5033 12459 -4999
rect 12379 -5049 12459 -5033
rect 12398 -5072 12459 -5049
rect 12399 -5218 12459 -5072
rect 12398 -5391 12459 -5218
rect 11403 -5492 11463 -5466
rect 11371 -5633 11438 -5626
rect 11521 -5633 11581 -5466
rect 11639 -5492 11699 -5466
rect 11757 -5492 11817 -5466
rect 11371 -5642 11581 -5633
rect 11371 -5676 11387 -5642
rect 11421 -5676 11581 -5642
rect 11371 -5692 11581 -5676
rect 11101 -5709 11252 -5693
rect 11101 -5743 11202 -5709
rect 11236 -5743 11252 -5709
rect 11101 -5759 11252 -5743
rect 9507 -5786 9567 -5760
rect 9625 -5786 9685 -5760
rect 9743 -5786 9803 -5760
rect 9861 -5780 9921 -5760
rect 9861 -5786 9922 -5780
rect 9979 -5786 10039 -5760
rect 10097 -5786 10157 -5760
rect 3661 -5840 3677 -5806
rect 3711 -5840 3727 -5806
rect 3661 -5856 3727 -5840
rect 3543 -5923 3609 -5907
rect 3543 -5957 3559 -5923
rect 3593 -5957 3609 -5923
rect 3543 -5973 3609 -5957
rect 3546 -5995 3606 -5973
rect 4550 -6022 4610 -5996
rect 3546 -6221 3606 -6195
rect 5848 -6022 5908 -5996
rect 6448 -6022 6508 -5996
rect 9744 -5971 9802 -5786
rect 7746 -6022 7806 -5996
rect 9744 -5997 9804 -5971
rect 9862 -5997 9922 -5786
rect 10215 -5792 10275 -5760
rect 10333 -5786 10393 -5760
rect 10451 -5786 10511 -5760
rect 10212 -5808 10278 -5792
rect 11101 -5798 11161 -5759
rect 11521 -5798 11581 -5692
rect 11875 -5633 11935 -5466
rect 11993 -5492 12053 -5466
rect 12018 -5633 12085 -5626
rect 11875 -5642 12085 -5633
rect 11875 -5676 12035 -5642
rect 12069 -5676 12085 -5642
rect 11875 -5692 12085 -5676
rect 11637 -5726 11703 -5710
rect 11637 -5760 11653 -5726
rect 11687 -5760 11703 -5726
rect 11637 -5776 11703 -5760
rect 11755 -5725 11821 -5710
rect 11755 -5759 11771 -5725
rect 11805 -5759 11821 -5725
rect 11755 -5775 11821 -5759
rect 11639 -5798 11699 -5776
rect 11757 -5798 11817 -5775
rect 11875 -5798 11935 -5692
rect 12399 -5694 12459 -5391
rect 12309 -5710 12459 -5694
rect 12309 -5744 12325 -5710
rect 12359 -5744 12459 -5710
rect 12309 -5760 12459 -5744
rect 12399 -5798 12459 -5760
rect 12999 -5499 13059 -4841
rect 13712 -4843 14255 -4792
rect 14297 -4799 14373 -4792
rect 14431 -4799 14491 -4773
rect 17631 -4572 17691 -4546
rect 17749 -4572 17809 -4546
rect 17867 -4572 17927 -4546
rect 16757 -4618 16817 -4592
rect 14297 -4843 14372 -4799
rect 16404 -4814 16464 -4792
rect 16522 -4808 16582 -4792
rect 16401 -4830 16467 -4814
rect 13301 -5043 13597 -4983
rect 13301 -5066 13361 -5043
rect 13419 -5066 13479 -5043
rect 13537 -5066 13597 -5043
rect 13655 -5042 13951 -4982
rect 13655 -5066 13715 -5042
rect 13773 -5066 13833 -5042
rect 13891 -5066 13951 -5042
rect 14297 -4996 14357 -4843
rect 16401 -4864 16417 -4830
rect 16451 -4864 16467 -4830
rect 16401 -4880 16467 -4864
rect 16516 -4830 16590 -4808
rect 16516 -4864 16535 -4830
rect 16569 -4864 16590 -4830
rect 18952 -4555 19248 -4504
rect 18952 -4572 19012 -4555
rect 19070 -4572 19130 -4555
rect 19188 -4572 19248 -4555
rect 19529 -4572 19589 -4546
rect 19647 -4572 19707 -4546
rect 19765 -4572 19825 -4546
rect 23026 -4391 23086 -4365
rect 23144 -4391 23204 -4180
rect 23497 -4186 23557 -4154
rect 23615 -4180 23675 -4154
rect 23733 -4180 23793 -4154
rect 23494 -4202 23560 -4186
rect 23494 -4236 23510 -4202
rect 23544 -4236 23560 -4202
rect 23494 -4252 23560 -4236
rect 23376 -4319 23442 -4303
rect 23376 -4353 23392 -4319
rect 23426 -4353 23442 -4319
rect 23376 -4369 23442 -4353
rect 24737 -4356 25033 -4305
rect 23379 -4391 23439 -4369
rect 24737 -4371 24797 -4356
rect 24855 -4371 24915 -4356
rect 24973 -4371 25033 -4356
rect 25091 -4371 25151 -4345
rect 25209 -4371 25269 -4345
rect 25327 -4371 25387 -4345
rect 26635 -4356 26931 -4305
rect 26635 -4371 26695 -4356
rect 26753 -4371 26813 -4356
rect 26871 -4371 26931 -4356
rect 26989 -4371 27049 -4345
rect 27107 -4371 27167 -4345
rect 27225 -4371 27285 -4345
rect 20850 -4555 21146 -4504
rect 20850 -4572 20910 -4555
rect 20968 -4572 21028 -4555
rect 21086 -4572 21146 -4555
rect 17631 -4789 17691 -4772
rect 17749 -4789 17809 -4772
rect 17867 -4789 17927 -4772
rect 18115 -4789 18175 -4772
rect 17631 -4840 18175 -4789
rect 18233 -4798 18293 -4772
rect 18351 -4798 18411 -4772
rect 18469 -4791 18529 -4772
rect 18587 -4791 18647 -4772
rect 18705 -4791 18765 -4772
rect 18952 -4791 19012 -4772
rect 19070 -4791 19130 -4772
rect 16516 -4921 16590 -4864
rect 17756 -4921 17816 -4840
rect 18469 -4842 19012 -4791
rect 19054 -4798 19130 -4791
rect 19188 -4798 19248 -4772
rect 19529 -4789 19589 -4772
rect 19647 -4789 19707 -4772
rect 19765 -4789 19825 -4772
rect 20013 -4789 20073 -4772
rect 19054 -4842 19129 -4798
rect 19529 -4840 20073 -4789
rect 20131 -4798 20191 -4772
rect 20249 -4798 20309 -4772
rect 20367 -4791 20427 -4772
rect 20485 -4791 20545 -4772
rect 20603 -4791 20663 -4772
rect 20850 -4791 20910 -4772
rect 20968 -4791 21028 -4772
rect 16516 -4946 17816 -4921
rect 16515 -4994 17816 -4946
rect 19054 -4962 19114 -4842
rect 14297 -5020 14551 -4996
rect 14297 -5054 14501 -5020
rect 14535 -5054 14551 -5020
rect 14297 -5070 14551 -5054
rect 13301 -5492 13361 -5466
rect 12999 -5515 13066 -5499
rect 12999 -5549 13015 -5515
rect 13049 -5549 13066 -5515
rect 12999 -5565 13066 -5549
rect 12999 -5693 13059 -5565
rect 13269 -5633 13336 -5626
rect 13419 -5633 13479 -5466
rect 13537 -5492 13597 -5466
rect 13655 -5492 13715 -5466
rect 13269 -5642 13479 -5633
rect 13269 -5676 13285 -5642
rect 13319 -5676 13479 -5642
rect 13269 -5692 13479 -5676
rect 12999 -5709 13150 -5693
rect 12999 -5743 13100 -5709
rect 13134 -5743 13150 -5709
rect 12999 -5759 13150 -5743
rect 12999 -5798 13059 -5759
rect 13419 -5798 13479 -5692
rect 13773 -5633 13833 -5466
rect 13891 -5492 13951 -5466
rect 13914 -5632 13981 -5625
rect 13908 -5633 13981 -5632
rect 13773 -5641 13981 -5633
rect 13773 -5675 13931 -5641
rect 13965 -5675 13981 -5641
rect 13773 -5691 13981 -5675
rect 13773 -5692 13970 -5691
rect 13535 -5726 13601 -5710
rect 13535 -5760 13551 -5726
rect 13585 -5760 13601 -5726
rect 13535 -5776 13601 -5760
rect 13653 -5725 13719 -5710
rect 13653 -5759 13669 -5725
rect 13703 -5759 13719 -5725
rect 13653 -5775 13719 -5759
rect 13537 -5798 13597 -5776
rect 13655 -5798 13715 -5775
rect 13773 -5798 13833 -5692
rect 14297 -5694 14357 -5070
rect 16162 -5538 16458 -5502
rect 16162 -5559 16222 -5538
rect 16280 -5559 16340 -5538
rect 16398 -5559 16458 -5538
rect 16516 -5539 16812 -5503
rect 16516 -5559 16576 -5539
rect 16634 -5559 16694 -5539
rect 16752 -5559 16812 -5539
rect 16870 -5539 17166 -5503
rect 16870 -5559 16930 -5539
rect 16988 -5559 17048 -5539
rect 17106 -5559 17166 -5539
rect 14207 -5710 14357 -5694
rect 14207 -5744 14223 -5710
rect 14257 -5744 14357 -5710
rect 14207 -5760 14357 -5744
rect 17756 -5692 17816 -4994
rect 18058 -5042 18354 -4982
rect 18058 -5065 18118 -5042
rect 18176 -5065 18236 -5042
rect 18294 -5065 18354 -5042
rect 18412 -5041 18708 -4981
rect 19053 -4982 19114 -4962
rect 18412 -5065 18472 -5041
rect 18530 -5065 18590 -5041
rect 18648 -5065 18708 -5041
rect 19034 -4998 19114 -4982
rect 19034 -5032 19049 -4998
rect 19083 -5032 19114 -4998
rect 19034 -5048 19114 -5032
rect 19053 -5071 19114 -5048
rect 19054 -5217 19114 -5071
rect 19053 -5390 19114 -5217
rect 18058 -5491 18118 -5465
rect 18026 -5632 18093 -5625
rect 18176 -5632 18236 -5465
rect 18294 -5491 18354 -5465
rect 18412 -5491 18472 -5465
rect 18026 -5641 18236 -5632
rect 18026 -5675 18042 -5641
rect 18076 -5675 18236 -5641
rect 18026 -5691 18236 -5675
rect 17756 -5708 17907 -5692
rect 17756 -5742 17857 -5708
rect 17891 -5742 17907 -5708
rect 17756 -5758 17907 -5742
rect 14297 -5798 14357 -5760
rect 16162 -5785 16222 -5759
rect 16280 -5785 16340 -5759
rect 16398 -5785 16458 -5759
rect 16516 -5779 16576 -5759
rect 16516 -5785 16577 -5779
rect 16634 -5785 16694 -5759
rect 16752 -5785 16812 -5759
rect 10212 -5842 10228 -5808
rect 10262 -5842 10278 -5808
rect 10212 -5858 10278 -5842
rect 10094 -5925 10160 -5909
rect 10094 -5959 10110 -5925
rect 10144 -5959 10160 -5925
rect 10094 -5975 10160 -5959
rect 10097 -5997 10157 -5975
rect 4970 -6222 5030 -6196
rect 5088 -6222 5148 -6196
rect 5206 -6222 5266 -6196
rect 5324 -6222 5384 -6196
rect 6868 -6222 6928 -6196
rect 6986 -6222 7046 -6196
rect 7104 -6222 7164 -6196
rect 7222 -6222 7282 -6196
rect 3193 -6417 3253 -6395
rect 3311 -6417 3371 -6395
rect 3190 -6433 3256 -6417
rect 3190 -6467 3206 -6433
rect 3240 -6467 3256 -6433
rect 3190 -6483 3256 -6467
rect 3308 -6433 3374 -6417
rect 3308 -6467 3324 -6433
rect 3358 -6467 3374 -6433
rect 11101 -6024 11161 -5998
rect 10097 -6223 10157 -6197
rect 12399 -6024 12459 -5998
rect 12999 -6024 13059 -5998
rect 16399 -5970 16457 -5785
rect 16399 -5996 16459 -5970
rect 16517 -5996 16577 -5785
rect 16870 -5791 16930 -5759
rect 16988 -5785 17048 -5759
rect 17106 -5785 17166 -5759
rect 16867 -5807 16933 -5791
rect 17756 -5797 17816 -5758
rect 18176 -5797 18236 -5691
rect 18530 -5632 18590 -5465
rect 18648 -5491 18708 -5465
rect 18673 -5632 18740 -5625
rect 18530 -5641 18740 -5632
rect 18530 -5675 18690 -5641
rect 18724 -5675 18740 -5641
rect 18530 -5691 18740 -5675
rect 18292 -5725 18358 -5709
rect 18292 -5759 18308 -5725
rect 18342 -5759 18358 -5725
rect 18292 -5775 18358 -5759
rect 18410 -5724 18476 -5709
rect 18410 -5758 18426 -5724
rect 18460 -5758 18476 -5724
rect 18410 -5774 18476 -5758
rect 18294 -5797 18354 -5775
rect 18412 -5797 18472 -5774
rect 18530 -5797 18590 -5691
rect 19054 -5693 19114 -5390
rect 18964 -5709 19114 -5693
rect 18964 -5743 18980 -5709
rect 19014 -5743 19114 -5709
rect 18964 -5759 19114 -5743
rect 19054 -5797 19114 -5759
rect 19654 -5498 19714 -4840
rect 20367 -4842 20910 -4791
rect 20952 -4798 21028 -4791
rect 21086 -4798 21146 -4772
rect 24253 -4571 24313 -4545
rect 24371 -4571 24431 -4545
rect 24489 -4571 24549 -4545
rect 23379 -4617 23439 -4591
rect 20952 -4842 21027 -4798
rect 23026 -4813 23086 -4791
rect 23144 -4807 23204 -4791
rect 23023 -4829 23089 -4813
rect 19956 -5042 20252 -4982
rect 19956 -5065 20016 -5042
rect 20074 -5065 20134 -5042
rect 20192 -5065 20252 -5042
rect 20310 -5041 20606 -4981
rect 20310 -5065 20370 -5041
rect 20428 -5065 20488 -5041
rect 20546 -5065 20606 -5041
rect 20952 -4995 21012 -4842
rect 23023 -4863 23039 -4829
rect 23073 -4863 23089 -4829
rect 23023 -4879 23089 -4863
rect 23138 -4829 23212 -4807
rect 23138 -4863 23157 -4829
rect 23191 -4863 23212 -4829
rect 25574 -4554 25870 -4503
rect 25574 -4571 25634 -4554
rect 25692 -4571 25752 -4554
rect 25810 -4571 25870 -4554
rect 26151 -4571 26211 -4545
rect 26269 -4571 26329 -4545
rect 26387 -4571 26447 -4545
rect 27472 -4554 27768 -4503
rect 27472 -4571 27532 -4554
rect 27590 -4571 27650 -4554
rect 27708 -4571 27768 -4554
rect 24253 -4788 24313 -4771
rect 24371 -4788 24431 -4771
rect 24489 -4788 24549 -4771
rect 24737 -4788 24797 -4771
rect 24253 -4839 24797 -4788
rect 24855 -4797 24915 -4771
rect 24973 -4797 25033 -4771
rect 25091 -4790 25151 -4771
rect 25209 -4790 25269 -4771
rect 25327 -4790 25387 -4771
rect 25574 -4790 25634 -4771
rect 25692 -4790 25752 -4771
rect 23138 -4920 23212 -4863
rect 24378 -4920 24438 -4839
rect 25091 -4841 25634 -4790
rect 25676 -4797 25752 -4790
rect 25810 -4797 25870 -4771
rect 26151 -4788 26211 -4771
rect 26269 -4788 26329 -4771
rect 26387 -4788 26447 -4771
rect 26635 -4788 26695 -4771
rect 25676 -4841 25751 -4797
rect 26151 -4839 26695 -4788
rect 26753 -4797 26813 -4771
rect 26871 -4797 26931 -4771
rect 26989 -4790 27049 -4771
rect 27107 -4790 27167 -4771
rect 27225 -4790 27285 -4771
rect 27472 -4790 27532 -4771
rect 27590 -4790 27650 -4771
rect 23138 -4945 24438 -4920
rect 23137 -4993 24438 -4945
rect 25676 -4961 25736 -4841
rect 20952 -5019 21206 -4995
rect 20952 -5053 21156 -5019
rect 21190 -5053 21206 -5019
rect 20952 -5069 21206 -5053
rect 19956 -5491 20016 -5465
rect 19654 -5514 19721 -5498
rect 19654 -5548 19670 -5514
rect 19704 -5548 19721 -5514
rect 19654 -5564 19721 -5548
rect 19654 -5692 19714 -5564
rect 19924 -5632 19991 -5625
rect 20074 -5632 20134 -5465
rect 20192 -5491 20252 -5465
rect 20310 -5491 20370 -5465
rect 19924 -5641 20134 -5632
rect 19924 -5675 19940 -5641
rect 19974 -5675 20134 -5641
rect 19924 -5691 20134 -5675
rect 19654 -5708 19805 -5692
rect 19654 -5742 19755 -5708
rect 19789 -5742 19805 -5708
rect 19654 -5758 19805 -5742
rect 19654 -5797 19714 -5758
rect 20074 -5797 20134 -5691
rect 20428 -5632 20488 -5465
rect 20546 -5491 20606 -5465
rect 20569 -5631 20636 -5624
rect 20563 -5632 20636 -5631
rect 20428 -5640 20636 -5632
rect 20428 -5674 20586 -5640
rect 20620 -5674 20636 -5640
rect 20428 -5690 20636 -5674
rect 20428 -5691 20625 -5690
rect 20190 -5725 20256 -5709
rect 20190 -5759 20206 -5725
rect 20240 -5759 20256 -5725
rect 20190 -5775 20256 -5759
rect 20308 -5724 20374 -5709
rect 20308 -5758 20324 -5724
rect 20358 -5758 20374 -5724
rect 20308 -5774 20374 -5758
rect 20192 -5797 20252 -5775
rect 20310 -5797 20370 -5774
rect 20428 -5797 20488 -5691
rect 20952 -5693 21012 -5069
rect 22784 -5537 23080 -5501
rect 22784 -5558 22844 -5537
rect 22902 -5558 22962 -5537
rect 23020 -5558 23080 -5537
rect 23138 -5538 23434 -5502
rect 23138 -5558 23198 -5538
rect 23256 -5558 23316 -5538
rect 23374 -5558 23434 -5538
rect 23492 -5538 23788 -5502
rect 23492 -5558 23552 -5538
rect 23610 -5558 23670 -5538
rect 23728 -5558 23788 -5538
rect 20862 -5709 21012 -5693
rect 20862 -5743 20878 -5709
rect 20912 -5743 21012 -5709
rect 20862 -5759 21012 -5743
rect 24378 -5691 24438 -4993
rect 24680 -5041 24976 -4981
rect 24680 -5064 24740 -5041
rect 24798 -5064 24858 -5041
rect 24916 -5064 24976 -5041
rect 25034 -5040 25330 -4980
rect 25675 -4981 25736 -4961
rect 25034 -5064 25094 -5040
rect 25152 -5064 25212 -5040
rect 25270 -5064 25330 -5040
rect 25656 -4997 25736 -4981
rect 25656 -5031 25671 -4997
rect 25705 -5031 25736 -4997
rect 25656 -5047 25736 -5031
rect 25675 -5070 25736 -5047
rect 25676 -5216 25736 -5070
rect 25675 -5389 25736 -5216
rect 24680 -5490 24740 -5464
rect 24648 -5631 24715 -5624
rect 24798 -5631 24858 -5464
rect 24916 -5490 24976 -5464
rect 25034 -5490 25094 -5464
rect 24648 -5640 24858 -5631
rect 24648 -5674 24664 -5640
rect 24698 -5674 24858 -5640
rect 24648 -5690 24858 -5674
rect 24378 -5707 24529 -5691
rect 24378 -5741 24479 -5707
rect 24513 -5741 24529 -5707
rect 24378 -5757 24529 -5741
rect 20952 -5797 21012 -5759
rect 22784 -5784 22844 -5758
rect 22902 -5784 22962 -5758
rect 23020 -5784 23080 -5758
rect 23138 -5778 23198 -5758
rect 23138 -5784 23199 -5778
rect 23256 -5784 23316 -5758
rect 23374 -5784 23434 -5758
rect 16867 -5841 16883 -5807
rect 16917 -5841 16933 -5807
rect 16867 -5857 16933 -5841
rect 16749 -5924 16815 -5908
rect 16749 -5958 16765 -5924
rect 16799 -5958 16815 -5924
rect 16749 -5974 16815 -5958
rect 16752 -5996 16812 -5974
rect 14297 -6024 14357 -5998
rect 11521 -6224 11581 -6198
rect 11639 -6224 11699 -6198
rect 11757 -6224 11817 -6198
rect 11875 -6224 11935 -6198
rect 13419 -6224 13479 -6198
rect 13537 -6224 13597 -6198
rect 13655 -6224 13715 -6198
rect 13773 -6224 13833 -6198
rect 9744 -6419 9804 -6397
rect 9862 -6419 9922 -6397
rect 9741 -6435 9807 -6419
rect 3308 -6483 3374 -6467
rect 9741 -6469 9757 -6435
rect 9791 -6469 9807 -6435
rect 9741 -6485 9807 -6469
rect 9859 -6435 9925 -6419
rect 9859 -6469 9875 -6435
rect 9909 -6469 9925 -6435
rect 17756 -6023 17816 -5997
rect 16752 -6222 16812 -6196
rect 19054 -6023 19114 -5997
rect 19654 -6023 19714 -5997
rect 23021 -5969 23079 -5784
rect 23021 -5995 23081 -5969
rect 23139 -5995 23199 -5784
rect 23492 -5790 23552 -5758
rect 23610 -5784 23670 -5758
rect 23728 -5784 23788 -5758
rect 23489 -5806 23555 -5790
rect 24378 -5796 24438 -5757
rect 24798 -5796 24858 -5690
rect 25152 -5631 25212 -5464
rect 25270 -5490 25330 -5464
rect 25295 -5631 25362 -5624
rect 25152 -5640 25362 -5631
rect 25152 -5674 25312 -5640
rect 25346 -5674 25362 -5640
rect 25152 -5690 25362 -5674
rect 24914 -5724 24980 -5708
rect 24914 -5758 24930 -5724
rect 24964 -5758 24980 -5724
rect 24914 -5774 24980 -5758
rect 25032 -5723 25098 -5708
rect 25032 -5757 25048 -5723
rect 25082 -5757 25098 -5723
rect 25032 -5773 25098 -5757
rect 24916 -5796 24976 -5774
rect 25034 -5796 25094 -5773
rect 25152 -5796 25212 -5690
rect 25676 -5692 25736 -5389
rect 25586 -5708 25736 -5692
rect 25586 -5742 25602 -5708
rect 25636 -5742 25736 -5708
rect 25586 -5758 25736 -5742
rect 25676 -5796 25736 -5758
rect 26276 -5497 26336 -4839
rect 26989 -4841 27532 -4790
rect 27574 -4797 27650 -4790
rect 27708 -4797 27768 -4771
rect 27574 -4841 27649 -4797
rect 26578 -5041 26874 -4981
rect 26578 -5064 26638 -5041
rect 26696 -5064 26756 -5041
rect 26814 -5064 26874 -5041
rect 26932 -5040 27228 -4980
rect 26932 -5064 26992 -5040
rect 27050 -5064 27110 -5040
rect 27168 -5064 27228 -5040
rect 27574 -4994 27634 -4841
rect 27574 -5018 27828 -4994
rect 27574 -5052 27778 -5018
rect 27812 -5052 27828 -5018
rect 27574 -5068 27828 -5052
rect 26578 -5490 26638 -5464
rect 26276 -5513 26343 -5497
rect 26276 -5547 26292 -5513
rect 26326 -5547 26343 -5513
rect 26276 -5563 26343 -5547
rect 26276 -5691 26336 -5563
rect 26546 -5631 26613 -5624
rect 26696 -5631 26756 -5464
rect 26814 -5490 26874 -5464
rect 26932 -5490 26992 -5464
rect 26546 -5640 26756 -5631
rect 26546 -5674 26562 -5640
rect 26596 -5674 26756 -5640
rect 26546 -5690 26756 -5674
rect 26276 -5707 26427 -5691
rect 26276 -5741 26377 -5707
rect 26411 -5741 26427 -5707
rect 26276 -5757 26427 -5741
rect 26276 -5796 26336 -5757
rect 26696 -5796 26756 -5690
rect 27050 -5631 27110 -5464
rect 27168 -5490 27228 -5464
rect 27191 -5630 27258 -5623
rect 27185 -5631 27258 -5630
rect 27050 -5639 27258 -5631
rect 27050 -5673 27208 -5639
rect 27242 -5673 27258 -5639
rect 27050 -5689 27258 -5673
rect 27050 -5690 27247 -5689
rect 26812 -5724 26878 -5708
rect 26812 -5758 26828 -5724
rect 26862 -5758 26878 -5724
rect 26812 -5774 26878 -5758
rect 26930 -5723 26996 -5708
rect 26930 -5757 26946 -5723
rect 26980 -5757 26996 -5723
rect 26930 -5773 26996 -5757
rect 26814 -5796 26874 -5774
rect 26932 -5796 26992 -5773
rect 27050 -5796 27110 -5690
rect 27574 -5692 27634 -5068
rect 28648 -5077 28944 -5041
rect 28648 -5098 28708 -5077
rect 28766 -5098 28826 -5077
rect 28884 -5098 28944 -5077
rect 29002 -5078 29298 -5042
rect 29002 -5098 29062 -5078
rect 29120 -5098 29180 -5078
rect 29238 -5098 29298 -5078
rect 29356 -5078 29652 -5042
rect 29356 -5098 29416 -5078
rect 29474 -5098 29534 -5078
rect 29592 -5098 29652 -5078
rect 28648 -5324 28708 -5298
rect 28766 -5324 28826 -5298
rect 28884 -5324 28944 -5298
rect 29002 -5318 29062 -5298
rect 29002 -5324 29063 -5318
rect 29120 -5324 29180 -5298
rect 29238 -5324 29298 -5298
rect 28885 -5509 28943 -5324
rect 28885 -5535 28945 -5509
rect 29003 -5535 29063 -5324
rect 29356 -5330 29416 -5298
rect 29474 -5324 29534 -5298
rect 29592 -5324 29652 -5298
rect 29353 -5346 29419 -5330
rect 29353 -5380 29369 -5346
rect 29403 -5380 29419 -5346
rect 29353 -5396 29419 -5380
rect 29235 -5463 29301 -5447
rect 29235 -5497 29251 -5463
rect 29285 -5497 29301 -5463
rect 29235 -5513 29301 -5497
rect 29238 -5535 29298 -5513
rect 27484 -5708 27634 -5692
rect 27484 -5742 27500 -5708
rect 27534 -5742 27634 -5708
rect 27484 -5758 27634 -5742
rect 27574 -5796 27634 -5758
rect 23489 -5840 23505 -5806
rect 23539 -5840 23555 -5806
rect 23489 -5856 23555 -5840
rect 23371 -5923 23437 -5907
rect 23371 -5957 23387 -5923
rect 23421 -5957 23437 -5923
rect 23371 -5973 23437 -5957
rect 23374 -5995 23434 -5973
rect 20952 -6023 21012 -5997
rect 18176 -6223 18236 -6197
rect 18294 -6223 18354 -6197
rect 18412 -6223 18472 -6197
rect 18530 -6223 18590 -6197
rect 20074 -6223 20134 -6197
rect 20192 -6223 20252 -6197
rect 20310 -6223 20370 -6197
rect 20428 -6223 20488 -6197
rect 16399 -6418 16459 -6396
rect 16517 -6418 16577 -6396
rect 16396 -6434 16462 -6418
rect 9859 -6485 9925 -6469
rect 16396 -6468 16412 -6434
rect 16446 -6468 16462 -6434
rect 16396 -6484 16462 -6468
rect 16514 -6434 16580 -6418
rect 16514 -6468 16530 -6434
rect 16564 -6468 16580 -6434
rect 24378 -6022 24438 -5996
rect 23374 -6221 23434 -6195
rect 25676 -6022 25736 -5996
rect 26276 -6022 26336 -5996
rect 29238 -5761 29298 -5735
rect 28885 -5957 28945 -5935
rect 29003 -5957 29063 -5935
rect 28882 -5973 28948 -5957
rect 27574 -6022 27634 -5996
rect 28882 -6007 28898 -5973
rect 28932 -6007 28948 -5973
rect 28882 -6023 28948 -6007
rect 29000 -5973 29066 -5957
rect 29000 -6007 29016 -5973
rect 29050 -6007 29066 -5973
rect 29000 -6023 29066 -6007
rect 24798 -6222 24858 -6196
rect 24916 -6222 24976 -6196
rect 25034 -6222 25094 -6196
rect 25152 -6222 25212 -6196
rect 26696 -6222 26756 -6196
rect 26814 -6222 26874 -6196
rect 26932 -6222 26992 -6196
rect 27050 -6222 27110 -6196
rect 23021 -6417 23081 -6395
rect 23139 -6417 23199 -6395
rect 23018 -6433 23084 -6417
rect 16514 -6484 16580 -6468
rect 23018 -6467 23034 -6433
rect 23068 -6467 23084 -6433
rect 23018 -6483 23084 -6467
rect 23136 -6433 23202 -6417
rect 23136 -6467 23152 -6433
rect 23186 -6467 23202 -6433
rect 23136 -6483 23202 -6467
rect 30879 -6628 31175 -6577
rect 30879 -6643 30939 -6628
rect 30997 -6643 31057 -6628
rect 31115 -6643 31175 -6628
rect 31233 -6643 31293 -6617
rect 31351 -6643 31411 -6617
rect 31469 -6643 31529 -6617
rect 30395 -6843 30455 -6817
rect 30513 -6843 30573 -6817
rect 30631 -6843 30691 -6817
rect 31716 -6826 32012 -6775
rect 31716 -6843 31776 -6826
rect 31834 -6843 31894 -6826
rect 31952 -6843 32012 -6826
rect 32188 -6825 32484 -6789
rect 32188 -6846 32248 -6825
rect 32306 -6846 32366 -6825
rect 32424 -6846 32484 -6825
rect 32542 -6826 32838 -6790
rect 32542 -6846 32602 -6826
rect 32660 -6846 32720 -6826
rect 32778 -6846 32838 -6826
rect 32896 -6826 33192 -6790
rect 32896 -6846 32956 -6826
rect 33014 -6846 33074 -6826
rect 33132 -6846 33192 -6826
rect 30395 -7060 30455 -7043
rect 30513 -7060 30573 -7043
rect 30631 -7060 30691 -7043
rect 30879 -7060 30939 -7043
rect 30395 -7111 30939 -7060
rect 30997 -7069 31057 -7043
rect 31115 -7069 31175 -7043
rect 31233 -7062 31293 -7043
rect 31351 -7062 31411 -7043
rect 31469 -7062 31529 -7043
rect 31716 -7062 31776 -7043
rect 31834 -7062 31894 -7043
rect 30520 -7315 30580 -7111
rect 31233 -7113 31776 -7062
rect 31818 -7069 31894 -7062
rect 31952 -7069 32012 -7043
rect 31818 -7113 31893 -7069
rect 32188 -7072 32248 -7046
rect 32306 -7072 32366 -7046
rect 32424 -7072 32484 -7046
rect 32542 -7066 32602 -7046
rect 32542 -7072 32603 -7066
rect 32660 -7072 32720 -7046
rect 32778 -7072 32838 -7046
rect 31818 -7195 31878 -7113
rect 31818 -7213 32052 -7195
rect 31818 -7247 32001 -7213
rect 32035 -7247 32052 -7213
rect 30822 -7313 31118 -7253
rect 6998 -7352 7064 -7336
rect 6998 -7386 7014 -7352
rect 7048 -7386 7064 -7352
rect 6998 -7402 7064 -7386
rect 7116 -7352 7182 -7336
rect 7116 -7386 7132 -7352
rect 7166 -7386 7182 -7352
rect 7116 -7402 7182 -7386
rect 13552 -7347 13618 -7331
rect 13552 -7381 13568 -7347
rect 13602 -7381 13618 -7347
rect 13552 -7397 13618 -7381
rect 13670 -7347 13736 -7331
rect 30520 -7332 30651 -7315
rect 13670 -7381 13686 -7347
rect 13720 -7381 13736 -7347
rect 13670 -7397 13736 -7381
rect 20201 -7359 20267 -7343
rect 20201 -7393 20217 -7359
rect 20251 -7393 20267 -7359
rect 7001 -7424 7061 -7402
rect 7119 -7424 7179 -7402
rect 13555 -7419 13615 -7397
rect 13673 -7419 13733 -7397
rect 20201 -7409 20267 -7393
rect 20319 -7359 20385 -7343
rect 20319 -7393 20335 -7359
rect 20369 -7393 20385 -7359
rect 20319 -7409 20385 -7393
rect 30520 -7366 30601 -7332
rect 30635 -7366 30651 -7332
rect 30822 -7336 30882 -7313
rect 30940 -7336 31000 -7313
rect 31058 -7336 31118 -7313
rect 31176 -7312 31472 -7252
rect 31176 -7336 31236 -7312
rect 31294 -7336 31354 -7312
rect 31412 -7336 31472 -7312
rect 31818 -7263 32052 -7247
rect 32425 -7257 32483 -7072
rect 30520 -7383 30651 -7366
rect 7354 -7624 7414 -7598
rect 20204 -7431 20264 -7409
rect 20322 -7431 20382 -7409
rect 13908 -7619 13968 -7593
rect 7001 -7850 7061 -7824
rect 7001 -8035 7059 -7850
rect 7119 -8035 7179 -7824
rect 7354 -7846 7414 -7824
rect 13555 -7845 13615 -7819
rect 7351 -7862 7417 -7846
rect 7351 -7896 7367 -7862
rect 7401 -7896 7417 -7862
rect 7351 -7912 7417 -7896
rect 7469 -7979 7535 -7963
rect 7469 -8013 7485 -7979
rect 7519 -8013 7535 -7979
rect 7469 -8029 7535 -8013
rect 6764 -8061 6824 -8035
rect 6882 -8061 6942 -8035
rect 7000 -8061 7060 -8035
rect 7118 -8041 7179 -8035
rect 7118 -8061 7178 -8041
rect 7236 -8061 7296 -8035
rect 7354 -8061 7414 -8035
rect 7472 -8061 7532 -8029
rect 13555 -8030 13613 -7845
rect 13673 -8030 13733 -7819
rect 13908 -7841 13968 -7819
rect 20557 -7631 20617 -7605
rect 13905 -7857 13971 -7841
rect 13905 -7891 13921 -7857
rect 13955 -7891 13971 -7857
rect 13905 -7907 13971 -7891
rect 20204 -7857 20264 -7831
rect 14023 -7974 14089 -7958
rect 14023 -8008 14039 -7974
rect 14073 -8008 14089 -7974
rect 14023 -8024 14089 -8008
rect 7590 -8061 7650 -8035
rect 7708 -8061 7768 -8035
rect 13318 -8056 13378 -8030
rect 13436 -8056 13496 -8030
rect 13554 -8056 13614 -8030
rect 13672 -8036 13733 -8030
rect 13672 -8056 13732 -8036
rect 13790 -8056 13850 -8030
rect 13908 -8056 13968 -8030
rect 14026 -8056 14086 -8024
rect 14144 -8056 14204 -8030
rect 14262 -8056 14322 -8030
rect 20204 -8042 20262 -7857
rect 20322 -8042 20382 -7831
rect 20557 -7853 20617 -7831
rect 20554 -7869 20620 -7853
rect 20554 -7903 20570 -7869
rect 20604 -7903 20620 -7869
rect 20554 -7919 20620 -7903
rect 28655 -7922 28951 -7886
rect 28655 -7943 28715 -7922
rect 28773 -7943 28833 -7922
rect 28891 -7943 28951 -7922
rect 29009 -7923 29305 -7887
rect 29009 -7943 29069 -7923
rect 29127 -7943 29187 -7923
rect 29245 -7943 29305 -7923
rect 29363 -7923 29659 -7887
rect 29363 -7943 29423 -7923
rect 29481 -7943 29541 -7923
rect 29599 -7943 29659 -7923
rect 20672 -7986 20738 -7970
rect 20672 -8020 20688 -7986
rect 20722 -8020 20738 -7986
rect 20672 -8036 20738 -8020
rect 19967 -8068 20027 -8042
rect 20085 -8068 20145 -8042
rect 20203 -8068 20263 -8042
rect 20321 -8048 20382 -8042
rect 20321 -8068 20381 -8048
rect 20439 -8068 20499 -8042
rect 20557 -8068 20617 -8042
rect 20675 -8068 20735 -8036
rect 20793 -8068 20853 -8042
rect 20911 -8068 20971 -8042
rect 6764 -8282 6824 -8261
rect 6882 -8282 6942 -8261
rect 7000 -8282 7060 -8261
rect 6764 -8318 7060 -8282
rect 7118 -8281 7178 -8261
rect 7236 -8281 7296 -8261
rect 7354 -8281 7414 -8261
rect 7118 -8317 7414 -8281
rect 7472 -8281 7532 -8261
rect 7590 -8281 7650 -8261
rect 7708 -8281 7768 -8261
rect 7472 -8317 7768 -8281
rect 13318 -8277 13378 -8256
rect 13436 -8277 13496 -8256
rect 13554 -8277 13614 -8256
rect 13318 -8313 13614 -8277
rect 13672 -8276 13732 -8256
rect 13790 -8276 13850 -8256
rect 13908 -8276 13968 -8256
rect 13672 -8312 13968 -8276
rect 14026 -8276 14086 -8256
rect 14144 -8276 14204 -8256
rect 14262 -8276 14322 -8256
rect 30520 -7963 30580 -7383
rect 30822 -7762 30882 -7736
rect 30790 -7903 30857 -7896
rect 30940 -7903 31000 -7736
rect 31058 -7762 31118 -7736
rect 31176 -7762 31236 -7736
rect 30790 -7912 31000 -7903
rect 30790 -7946 30806 -7912
rect 30840 -7946 31000 -7912
rect 30790 -7962 31000 -7946
rect 30520 -7979 30671 -7963
rect 30520 -8013 30621 -7979
rect 30655 -8013 30671 -7979
rect 30520 -8029 30671 -8013
rect 30520 -8068 30580 -8029
rect 30940 -8068 31000 -7962
rect 31294 -7903 31354 -7736
rect 31412 -7762 31472 -7736
rect 31437 -7903 31504 -7896
rect 31294 -7912 31504 -7903
rect 31294 -7946 31454 -7912
rect 31488 -7946 31504 -7912
rect 31294 -7962 31504 -7946
rect 31056 -7996 31122 -7980
rect 31056 -8030 31072 -7996
rect 31106 -8030 31122 -7996
rect 31056 -8046 31122 -8030
rect 31174 -7995 31240 -7980
rect 31174 -8029 31190 -7995
rect 31224 -8029 31240 -7995
rect 31174 -8045 31240 -8029
rect 31058 -8068 31118 -8046
rect 31176 -8068 31236 -8045
rect 31294 -8068 31354 -7962
rect 31818 -7964 31878 -7263
rect 32425 -7283 32485 -7257
rect 32543 -7283 32603 -7072
rect 32896 -7078 32956 -7046
rect 33014 -7072 33074 -7046
rect 33132 -7072 33192 -7046
rect 32893 -7094 32959 -7078
rect 32893 -7128 32909 -7094
rect 32943 -7128 32959 -7094
rect 32893 -7144 32959 -7128
rect 32775 -7211 32841 -7195
rect 32775 -7245 32791 -7211
rect 32825 -7245 32841 -7211
rect 32775 -7261 32841 -7245
rect 32778 -7283 32838 -7261
rect 32778 -7509 32838 -7483
rect 32425 -7705 32485 -7683
rect 32543 -7705 32603 -7683
rect 32422 -7721 32488 -7705
rect 32422 -7755 32438 -7721
rect 32472 -7755 32488 -7721
rect 32422 -7771 32488 -7755
rect 32540 -7721 32606 -7705
rect 32540 -7755 32556 -7721
rect 32590 -7755 32606 -7721
rect 32540 -7771 32606 -7755
rect 31728 -7980 31878 -7964
rect 31728 -8014 31744 -7980
rect 31778 -8014 31878 -7980
rect 31728 -8030 31878 -8014
rect 31818 -8068 31878 -8030
rect 28655 -8169 28715 -8143
rect 28773 -8169 28833 -8143
rect 28891 -8169 28951 -8143
rect 29009 -8163 29069 -8143
rect 29009 -8169 29070 -8163
rect 29127 -8169 29187 -8143
rect 29245 -8169 29305 -8143
rect 14026 -8312 14322 -8276
rect 19967 -8289 20027 -8268
rect 20085 -8289 20145 -8268
rect 20203 -8289 20263 -8268
rect 19967 -8325 20263 -8289
rect 20321 -8288 20381 -8268
rect 20439 -8288 20499 -8268
rect 20557 -8288 20617 -8268
rect 20321 -8324 20617 -8288
rect 20675 -8288 20735 -8268
rect 20793 -8288 20853 -8268
rect 20911 -8288 20971 -8268
rect 20675 -8324 20971 -8288
rect 28892 -8354 28950 -8169
rect 28892 -8380 28952 -8354
rect 29010 -8380 29070 -8169
rect 29363 -8175 29423 -8143
rect 29481 -8169 29541 -8143
rect 29599 -8169 29659 -8143
rect 29360 -8191 29426 -8175
rect 29360 -8225 29376 -8191
rect 29410 -8225 29426 -8191
rect 29360 -8241 29426 -8225
rect 29242 -8308 29308 -8292
rect 30520 -8294 30580 -8268
rect 29242 -8342 29258 -8308
rect 29292 -8342 29308 -8308
rect 29242 -8358 29308 -8342
rect 29245 -8380 29305 -8358
rect 31818 -8294 31878 -8268
rect 30940 -8494 31000 -8468
rect 31058 -8494 31118 -8468
rect 31176 -8494 31236 -8468
rect 31294 -8494 31354 -8468
rect 29245 -8606 29305 -8580
rect 28892 -8802 28952 -8780
rect 29010 -8802 29070 -8780
rect 28889 -8818 28955 -8802
rect 28889 -8852 28905 -8818
rect 28939 -8852 28955 -8818
rect 28889 -8868 28955 -8852
rect 29007 -8818 29073 -8802
rect 29007 -8852 29023 -8818
rect 29057 -8852 29073 -8818
rect 29007 -8868 29073 -8852
<< polycont >>
rect 7450 5361 7484 5395
rect 7332 5244 7366 5278
rect 13999 5360 14033 5394
rect 13881 5243 13915 5277
rect 20653 5381 20687 5415
rect 20535 5264 20569 5298
rect 29306 5214 29340 5248
rect 29188 5097 29222 5131
rect 6979 4734 7013 4768
rect 7097 4734 7131 4768
rect 13528 4733 13562 4767
rect 13646 4733 13680 4767
rect 20182 4754 20216 4788
rect 20300 4754 20334 4788
rect 28835 4587 28869 4621
rect 28953 4587 28987 4621
rect 31999 4687 32033 4721
rect 30599 4568 30633 4602
rect 5119 3678 5153 3712
rect 6249 3684 6283 3718
rect 11668 3766 11702 3800
rect 12798 3772 12832 3806
rect 11668 3648 11702 3682
rect 12798 3652 12832 3686
rect 18322 3698 18356 3732
rect 19452 3704 19486 3738
rect 24947 3766 24981 3800
rect 26077 3772 26111 3806
rect 30804 3988 30838 4022
rect 30619 3921 30653 3955
rect 31452 3988 31486 4022
rect 31070 3904 31104 3938
rect 31188 3905 31222 3939
rect 32907 4806 32941 4840
rect 32789 4689 32823 4723
rect 32436 4179 32470 4213
rect 32554 4179 32588 4213
rect 31742 3920 31776 3954
rect 5119 3560 5153 3594
rect 6249 3564 6283 3598
rect 786 3461 820 3495
rect 668 3344 702 3378
rect 3676 3194 3710 3228
rect 3558 3077 3592 3111
rect 315 2834 349 2868
rect 433 2834 467 2868
rect 5439 2804 5473 2838
rect 10225 3282 10259 3316
rect 24947 3648 24981 3682
rect 18322 3580 18356 3614
rect 19452 3584 19486 3618
rect 26077 3652 26111 3686
rect 10107 3165 10141 3199
rect 6581 2808 6615 2842
rect 3205 2567 3239 2601
rect 3323 2567 3357 2601
rect 11988 2892 12022 2926
rect 16879 3214 16913 3248
rect 16761 3097 16795 3131
rect 13130 2896 13164 2930
rect 9754 2655 9788 2689
rect 9872 2655 9906 2689
rect 18642 2824 18676 2858
rect 23504 3282 23538 3316
rect 23386 3165 23420 3199
rect 19784 2828 19818 2862
rect 16408 2587 16442 2621
rect 16526 2587 16560 2621
rect 25267 2892 25301 2926
rect 26409 2896 26443 2930
rect 23033 2655 23067 2689
rect 23151 2655 23185 2689
rect 29301 2643 29335 2677
rect 29183 2526 29217 2560
rect 28830 2016 28864 2050
rect 28948 2016 28982 2050
rect 3690 1544 3724 1578
rect 10239 1632 10273 1666
rect 10121 1515 10155 1549
rect 3572 1427 3606 1461
rect 778 876 812 910
rect 3219 917 3253 951
rect 3337 917 3371 951
rect 660 759 694 793
rect 307 249 341 283
rect 425 249 459 283
rect 5851 749 5885 783
rect 4844 106 4878 140
rect 4659 39 4693 73
rect 5492 106 5526 140
rect 5110 22 5144 56
rect 5228 23 5262 57
rect 5782 38 5816 72
rect 9768 1005 9802 1039
rect 9886 1005 9920 1039
rect 16893 1564 16927 1598
rect 16775 1447 16809 1481
rect 23518 1632 23552 1666
rect 23400 1515 23434 1549
rect 7958 728 7992 762
rect 6472 233 6506 267
rect 6742 106 6776 140
rect 6557 39 6591 73
rect 7388 107 7422 141
rect 7008 22 7042 56
rect 7126 23 7160 57
rect 12400 837 12434 871
rect 11393 194 11427 228
rect 11208 127 11242 161
rect 7680 38 7714 72
rect 3685 -60 3719 -26
rect 3567 -177 3601 -143
rect 12041 194 12075 228
rect 11659 110 11693 144
rect 11777 111 11811 145
rect 12331 126 12365 160
rect 16422 937 16456 971
rect 16540 937 16574 971
rect 14507 816 14541 850
rect 13021 321 13055 355
rect 13291 194 13325 228
rect 13106 127 13140 161
rect 13937 195 13971 229
rect 13557 110 13591 144
rect 13675 111 13709 145
rect 14229 126 14263 160
rect 10234 28 10268 62
rect 10116 -89 10150 -55
rect 19054 769 19088 803
rect 18047 126 18081 160
rect 17862 59 17896 93
rect 18695 126 18729 160
rect 18313 42 18347 76
rect 18431 43 18465 77
rect 18985 58 19019 92
rect 23047 1005 23081 1039
rect 23165 1005 23199 1039
rect 21161 748 21195 782
rect 19675 253 19709 287
rect 19945 126 19979 160
rect 19760 59 19794 93
rect 20591 127 20625 161
rect 20211 42 20245 76
rect 20329 43 20363 77
rect 25679 837 25713 871
rect 24672 194 24706 228
rect 24487 127 24521 161
rect 20883 58 20917 92
rect 16888 -40 16922 -6
rect 16770 -157 16804 -123
rect 3214 -687 3248 -653
rect 3332 -687 3366 -653
rect 9763 -599 9797 -565
rect 9881 -599 9915 -565
rect 25320 194 25354 228
rect 24938 110 24972 144
rect 25056 111 25090 145
rect 25610 126 25644 160
rect 27786 816 27820 850
rect 26300 321 26334 355
rect 26570 194 26604 228
rect 26385 127 26419 161
rect 27216 195 27250 229
rect 26836 110 26870 144
rect 26954 111 26988 145
rect 27508 126 27542 160
rect 32001 596 32035 630
rect 30601 477 30635 511
rect 23513 28 23547 62
rect 23395 -89 23429 -55
rect 30806 -103 30840 -69
rect 30621 -170 30655 -136
rect 31454 -103 31488 -69
rect 31072 -187 31106 -153
rect 31190 -186 31224 -152
rect 32909 715 32943 749
rect 32791 598 32825 632
rect 32438 88 32472 122
rect 32556 88 32590 122
rect 31744 -171 31778 -137
rect 16417 -667 16451 -633
rect 16535 -667 16569 -633
rect 23042 -599 23076 -565
rect 23160 -599 23194 -565
rect 29301 -390 29335 -356
rect 29183 -507 29217 -473
rect 28830 -1017 28864 -983
rect 28948 -1017 28982 -983
rect 5111 -2102 5145 -2068
rect 6241 -2096 6275 -2062
rect 11662 -2104 11696 -2070
rect 12792 -2098 12826 -2064
rect 5111 -2220 5145 -2186
rect 6241 -2216 6275 -2182
rect 18317 -2103 18351 -2069
rect 19447 -2097 19481 -2063
rect 11662 -2222 11696 -2188
rect 759 -2402 793 -2368
rect 641 -2519 675 -2485
rect 3668 -2586 3702 -2552
rect 12792 -2218 12826 -2184
rect 24939 -2102 24973 -2068
rect 26069 -2096 26103 -2062
rect 18317 -2221 18351 -2187
rect 3550 -2703 3584 -2669
rect 288 -3029 322 -2995
rect 406 -3029 440 -2995
rect 5431 -2976 5465 -2942
rect 10219 -2588 10253 -2554
rect 19447 -2217 19481 -2183
rect 24939 -2220 24973 -2186
rect 10101 -2705 10135 -2671
rect 6573 -2972 6607 -2938
rect 3197 -3213 3231 -3179
rect 3315 -3213 3349 -3179
rect 11982 -2978 12016 -2944
rect 16874 -2587 16908 -2553
rect 26069 -2216 26103 -2182
rect 16756 -2704 16790 -2670
rect 13124 -2974 13158 -2940
rect 9748 -3215 9782 -3181
rect 9866 -3215 9900 -3181
rect 18637 -2977 18671 -2943
rect 23496 -2586 23530 -2552
rect 29372 -2310 29406 -2276
rect 29254 -2427 29288 -2393
rect 23378 -2703 23412 -2669
rect 19779 -2973 19813 -2939
rect 16403 -3214 16437 -3180
rect 16521 -3214 16555 -3180
rect 25259 -2976 25293 -2942
rect 26401 -2972 26435 -2938
rect 28901 -2937 28935 -2903
rect 29019 -2937 29053 -2903
rect 32001 -2899 32035 -2865
rect 23025 -3213 23059 -3179
rect 23143 -3213 23177 -3179
rect 30601 -3018 30635 -2984
rect 30806 -3598 30840 -3564
rect 30621 -3665 30655 -3631
rect 31454 -3598 31488 -3564
rect 31072 -3682 31106 -3648
rect 31190 -3681 31224 -3647
rect 32909 -2780 32943 -2746
rect 32791 -2897 32825 -2863
rect 32438 -3407 32472 -3373
rect 32556 -3407 32590 -3373
rect 31744 -3666 31778 -3632
rect 3682 -4236 3716 -4202
rect 3564 -4353 3598 -4319
rect 3211 -4863 3245 -4829
rect 3329 -4863 3363 -4829
rect 10233 -4238 10267 -4204
rect 10115 -4355 10149 -4321
rect 775 -5162 809 -5128
rect 657 -5279 691 -5245
rect 304 -5789 338 -5755
rect 422 -5789 456 -5755
rect 5843 -5031 5877 -4997
rect 4836 -5674 4870 -5640
rect 4651 -5741 4685 -5707
rect 5484 -5674 5518 -5640
rect 5102 -5758 5136 -5724
rect 5220 -5757 5254 -5723
rect 5774 -5742 5808 -5708
rect 9762 -4865 9796 -4831
rect 9880 -4865 9914 -4831
rect 16888 -4237 16922 -4203
rect 16770 -4354 16804 -4320
rect 7950 -5052 7984 -5018
rect 6464 -5547 6498 -5513
rect 6734 -5674 6768 -5640
rect 6549 -5741 6583 -5707
rect 7380 -5673 7414 -5639
rect 7000 -5758 7034 -5724
rect 7118 -5757 7152 -5723
rect 7672 -5742 7706 -5708
rect 12394 -5033 12428 -4999
rect 11387 -5676 11421 -5642
rect 11202 -5743 11236 -5709
rect 3677 -5840 3711 -5806
rect 3559 -5957 3593 -5923
rect 12035 -5676 12069 -5642
rect 11653 -5760 11687 -5726
rect 11771 -5759 11805 -5725
rect 12325 -5744 12359 -5710
rect 16417 -4864 16451 -4830
rect 16535 -4864 16569 -4830
rect 23510 -4236 23544 -4202
rect 23392 -4353 23426 -4319
rect 14501 -5054 14535 -5020
rect 13015 -5549 13049 -5515
rect 13285 -5676 13319 -5642
rect 13100 -5743 13134 -5709
rect 13931 -5675 13965 -5641
rect 13551 -5760 13585 -5726
rect 13669 -5759 13703 -5725
rect 14223 -5744 14257 -5710
rect 19049 -5032 19083 -4998
rect 18042 -5675 18076 -5641
rect 17857 -5742 17891 -5708
rect 10228 -5842 10262 -5808
rect 10110 -5959 10144 -5925
rect 3206 -6467 3240 -6433
rect 3324 -6467 3358 -6433
rect 18690 -5675 18724 -5641
rect 18308 -5759 18342 -5725
rect 18426 -5758 18460 -5724
rect 18980 -5743 19014 -5709
rect 23039 -4863 23073 -4829
rect 23157 -4863 23191 -4829
rect 21156 -5053 21190 -5019
rect 19670 -5548 19704 -5514
rect 19940 -5675 19974 -5641
rect 19755 -5742 19789 -5708
rect 20586 -5674 20620 -5640
rect 20206 -5759 20240 -5725
rect 20324 -5758 20358 -5724
rect 20878 -5743 20912 -5709
rect 25671 -5031 25705 -4997
rect 24664 -5674 24698 -5640
rect 24479 -5741 24513 -5707
rect 16883 -5841 16917 -5807
rect 16765 -5958 16799 -5924
rect 9757 -6469 9791 -6435
rect 9875 -6469 9909 -6435
rect 25312 -5674 25346 -5640
rect 24930 -5758 24964 -5724
rect 25048 -5757 25082 -5723
rect 25602 -5742 25636 -5708
rect 27778 -5052 27812 -5018
rect 26292 -5547 26326 -5513
rect 26562 -5674 26596 -5640
rect 26377 -5741 26411 -5707
rect 27208 -5673 27242 -5639
rect 26828 -5758 26862 -5724
rect 26946 -5757 26980 -5723
rect 29369 -5380 29403 -5346
rect 29251 -5497 29285 -5463
rect 27500 -5742 27534 -5708
rect 23505 -5840 23539 -5806
rect 23387 -5957 23421 -5923
rect 16412 -6468 16446 -6434
rect 16530 -6468 16564 -6434
rect 28898 -6007 28932 -5973
rect 29016 -6007 29050 -5973
rect 23034 -6467 23068 -6433
rect 23152 -6467 23186 -6433
rect 32001 -7247 32035 -7213
rect 7014 -7386 7048 -7352
rect 7132 -7386 7166 -7352
rect 13568 -7381 13602 -7347
rect 13686 -7381 13720 -7347
rect 20217 -7393 20251 -7359
rect 20335 -7393 20369 -7359
rect 30601 -7366 30635 -7332
rect 7367 -7896 7401 -7862
rect 7485 -8013 7519 -7979
rect 13921 -7891 13955 -7857
rect 14039 -8008 14073 -7974
rect 20570 -7903 20604 -7869
rect 20688 -8020 20722 -7986
rect 30806 -7946 30840 -7912
rect 30621 -8013 30655 -7979
rect 31454 -7946 31488 -7912
rect 31072 -8030 31106 -7996
rect 31190 -8029 31224 -7995
rect 32909 -7128 32943 -7094
rect 32791 -7245 32825 -7211
rect 32438 -7755 32472 -7721
rect 32556 -7755 32590 -7721
rect 31744 -8014 31778 -7980
rect 29376 -8225 29410 -8191
rect 29258 -8342 29292 -8308
rect 28905 -8852 28939 -8818
rect 29023 -8852 29057 -8818
<< locali >>
rect 20175 5891 20343 5907
rect 6972 5871 7140 5887
rect 6972 5801 6988 5871
rect 7124 5801 7140 5871
rect 6972 5785 7140 5801
rect 13521 5870 13689 5886
rect 13521 5800 13537 5870
rect 13673 5800 13689 5870
rect 20175 5821 20191 5891
rect 20327 5821 20343 5891
rect 20175 5805 20343 5821
rect 30970 5817 31414 5823
rect 13521 5784 13689 5800
rect 7509 5681 7779 5715
rect 6683 5631 6717 5647
rect 6683 5439 6717 5455
rect 6801 5631 6835 5647
rect 6801 5439 6835 5455
rect 6919 5631 6953 5647
rect 6919 5439 6953 5455
rect 7037 5631 7071 5647
rect 7037 5439 7071 5455
rect 7155 5631 7189 5647
rect 7155 5439 7189 5455
rect 7273 5631 7307 5647
rect 7273 5439 7307 5455
rect 7391 5631 7425 5647
rect 7391 5439 7425 5455
rect 7509 5631 7543 5681
rect 7509 5439 7543 5455
rect 7627 5631 7661 5647
rect 7627 5439 7661 5455
rect 7745 5631 7779 5681
rect 14058 5680 14328 5714
rect 7745 5439 7779 5455
rect 13232 5630 13266 5646
rect 13232 5438 13266 5454
rect 13350 5630 13384 5646
rect 13350 5438 13384 5454
rect 13468 5630 13502 5646
rect 13468 5438 13502 5454
rect 13586 5630 13620 5646
rect 13586 5438 13620 5454
rect 13704 5630 13738 5646
rect 13704 5438 13738 5454
rect 13822 5630 13856 5646
rect 13822 5438 13856 5454
rect 13940 5630 13974 5646
rect 13940 5438 13974 5454
rect 14058 5630 14092 5680
rect 14058 5438 14092 5454
rect 14176 5630 14210 5646
rect 14176 5438 14210 5454
rect 14294 5630 14328 5680
rect 20712 5701 20982 5735
rect 19886 5651 19920 5667
rect 19886 5459 19920 5475
rect 20004 5651 20038 5667
rect 20004 5459 20038 5475
rect 20122 5651 20156 5667
rect 20122 5459 20156 5475
rect 20240 5651 20274 5667
rect 20240 5459 20274 5475
rect 20358 5651 20392 5667
rect 20358 5459 20392 5475
rect 20476 5651 20510 5667
rect 20476 5459 20510 5475
rect 20594 5651 20628 5667
rect 20594 5459 20628 5475
rect 20712 5651 20746 5701
rect 20712 5459 20746 5475
rect 20830 5651 20864 5667
rect 20830 5459 20864 5475
rect 20948 5651 20982 5701
rect 28828 5724 28996 5740
rect 28828 5654 28844 5724
rect 28980 5654 28996 5724
rect 28828 5638 28996 5654
rect 30970 5617 30981 5817
rect 31402 5617 31414 5817
rect 30970 5611 31414 5617
rect 29365 5534 29635 5568
rect 20948 5459 20982 5475
rect 28539 5484 28573 5500
rect 14294 5438 14328 5454
rect 7434 5361 7450 5395
rect 7484 5361 7500 5395
rect 13983 5360 13999 5394
rect 14033 5360 14049 5394
rect 20637 5381 20653 5415
rect 20687 5381 20703 5415
rect 7316 5244 7332 5278
rect 7366 5244 7382 5278
rect 13865 5243 13881 5277
rect 13915 5243 13931 5277
rect 20519 5264 20535 5298
rect 20569 5264 20585 5298
rect 28539 5292 28573 5308
rect 28657 5484 28691 5500
rect 28657 5292 28691 5308
rect 28775 5484 28809 5500
rect 28775 5292 28809 5308
rect 28893 5484 28927 5500
rect 28893 5292 28927 5308
rect 29011 5484 29045 5500
rect 29011 5292 29045 5308
rect 29129 5484 29163 5500
rect 29129 5292 29163 5308
rect 29247 5484 29281 5500
rect 29247 5292 29281 5308
rect 29365 5484 29399 5534
rect 29365 5292 29399 5308
rect 29483 5484 29517 5500
rect 29483 5292 29517 5308
rect 29601 5484 29635 5534
rect 29601 5292 29635 5308
rect 31185 5332 31455 5367
rect 30831 5279 30865 5295
rect 20123 5214 20157 5230
rect 6920 5194 6954 5210
rect 6920 4802 6954 4818
rect 7038 5194 7072 5210
rect 7038 4802 7072 4818
rect 7156 5194 7190 5210
rect 7273 5194 7307 5210
rect 7273 5002 7307 5018
rect 7391 5194 7425 5210
rect 7391 5002 7425 5018
rect 13469 5193 13503 5209
rect 7156 4802 7190 4818
rect 13469 4801 13503 4817
rect 13587 5193 13621 5209
rect 13587 4801 13621 4817
rect 13705 5193 13739 5209
rect 13822 5193 13856 5209
rect 13822 5001 13856 5017
rect 13940 5193 13974 5209
rect 13940 5001 13974 5017
rect 20123 4822 20157 4838
rect 20241 5214 20275 5230
rect 20241 4822 20275 4838
rect 20359 5214 20393 5230
rect 20476 5214 20510 5230
rect 20476 5022 20510 5038
rect 20594 5214 20628 5230
rect 29290 5214 29306 5248
rect 29340 5214 29356 5248
rect 30347 5133 30617 5168
rect 29172 5097 29188 5131
rect 29222 5097 29238 5131
rect 30347 5079 30381 5133
rect 20594 5022 20628 5038
rect 28776 5047 28810 5063
rect 20359 4822 20393 4838
rect 13705 4801 13739 4817
rect 19985 4790 20056 4792
rect 13154 4768 13434 4773
rect 6963 4734 6979 4768
rect 7013 4734 7029 4768
rect 7081 4734 7097 4768
rect 7131 4734 7147 4768
rect 13154 4722 13382 4768
rect 13431 4722 13434 4768
rect 13512 4733 13528 4767
rect 13562 4733 13578 4767
rect 13630 4733 13646 4767
rect 13680 4733 13696 4767
rect 19985 4742 19989 4790
rect 20050 4742 20056 4790
rect 20166 4754 20182 4788
rect 20216 4754 20232 4788
rect 20284 4754 20300 4788
rect 20334 4754 20350 4788
rect 13154 4717 13434 4722
rect 19985 4729 20056 4742
rect 7196 4663 7364 4681
rect 7196 4607 7212 4663
rect 7346 4607 7364 4663
rect 7196 4591 7364 4607
rect -926 4516 -818 4519
rect -926 4466 -902 4516
rect -841 4466 -818 4516
rect -926 2824 -818 4466
rect 13154 4435 13207 4717
rect 13745 4662 13913 4680
rect 13745 4606 13761 4662
rect 13895 4606 13913 4662
rect 13745 4590 13913 4606
rect -767 4382 13207 4435
rect -767 3943 -676 4382
rect 19985 4347 20048 4729
rect -637 4343 20048 4347
rect -637 4289 6801 4343
rect 6850 4289 20048 4343
rect -637 4281 20048 4289
rect 20082 4700 20143 4705
rect 20082 4662 20091 4700
rect 20136 4662 20143 4700
rect -637 4117 -527 4281
rect 20082 4236 20143 4662
rect 20399 4683 20567 4701
rect 20399 4627 20415 4683
rect 20549 4627 20567 4683
rect 28776 4655 28810 4671
rect 28894 5047 28928 5063
rect 28894 4655 28928 4671
rect 29012 5047 29046 5063
rect 29129 5047 29163 5063
rect 29129 4855 29163 4871
rect 29247 5047 29281 5063
rect 30347 4887 30381 4903
rect 30465 5079 30499 5095
rect 30465 4887 30499 4903
rect 30583 5079 30617 5133
rect 30583 4887 30617 4903
rect 30701 5079 30735 5095
rect 30701 4887 30735 4903
rect 30831 4887 30865 4903
rect 30949 5279 30983 5295
rect 30949 4887 30983 4903
rect 31067 5279 31101 5295
rect 31067 4887 31101 4903
rect 31185 5279 31219 5332
rect 31185 4887 31219 4903
rect 31303 5279 31337 5295
rect 31303 4887 31337 4903
rect 31421 5279 31455 5332
rect 32429 5316 32597 5332
rect 31421 4887 31455 4903
rect 31539 5279 31573 5295
rect 32429 5246 32445 5316
rect 32581 5246 32597 5316
rect 32429 5230 32597 5246
rect 32966 5126 33236 5160
rect 31539 4887 31573 4903
rect 31668 5079 31702 5095
rect 31668 4887 31702 4903
rect 31786 5079 31820 5095
rect 31786 4887 31820 4903
rect 31904 5079 31938 5095
rect 31904 4887 31938 4903
rect 32022 5079 32056 5095
rect 32022 4887 32056 4903
rect 32140 5076 32174 5092
rect 32140 4884 32174 4900
rect 32258 5076 32292 5092
rect 32258 4884 32292 4900
rect 32376 5076 32410 5092
rect 32376 4884 32410 4900
rect 32494 5076 32528 5092
rect 32494 4884 32528 4900
rect 32612 5076 32646 5092
rect 32612 4884 32646 4900
rect 32730 5076 32764 5092
rect 32730 4884 32764 4900
rect 32848 5076 32882 5092
rect 32848 4884 32882 4900
rect 32966 5076 33000 5126
rect 32966 4884 33000 4900
rect 33084 5076 33118 5092
rect 33084 4884 33118 4900
rect 33202 5076 33236 5126
rect 33202 4884 33236 4900
rect 29247 4855 29281 4871
rect 32891 4806 32907 4840
rect 32941 4806 32957 4840
rect 31999 4721 32033 4737
rect 32773 4689 32789 4723
rect 32823 4689 32839 4723
rect 31999 4671 32033 4687
rect 29012 4655 29046 4671
rect 20399 4611 20567 4627
rect 32377 4639 32411 4655
rect 28819 4587 28835 4621
rect 28869 4587 28885 4621
rect 28937 4587 28953 4621
rect 28987 4587 29003 4621
rect 30076 4615 30418 4621
rect 30076 4547 30326 4615
rect 30406 4547 30418 4615
rect 30593 4602 30649 4619
rect 30593 4568 30599 4602
rect 30633 4568 30649 4602
rect 30593 4551 30649 4568
rect 30774 4586 30808 4602
rect 30076 4541 30418 4547
rect 29052 4516 29220 4534
rect 29052 4460 29068 4516
rect 29202 4460 29220 4516
rect 29052 4444 29220 4460
rect -767 3898 -749 3943
rect -692 3898 -676 3943
rect -767 3891 -676 3898
rect -926 2823 -798 2824
rect -937 2809 -798 2823
rect -937 2742 -922 2809
rect -936 2725 -922 2742
rect -809 2725 -798 2809
rect -936 -9100 -798 2725
rect -638 -5593 -527 4117
rect 1619 4170 20143 4236
rect 308 3971 476 3987
rect 308 3901 324 3971
rect 460 3901 476 3971
rect 308 3885 476 3901
rect 845 3781 1115 3815
rect 19 3731 53 3747
rect 19 3539 53 3555
rect 137 3731 171 3747
rect 137 3539 171 3555
rect 255 3731 289 3747
rect 255 3539 289 3555
rect 373 3731 407 3747
rect 373 3539 407 3555
rect 491 3731 525 3747
rect 491 3539 525 3555
rect 609 3731 643 3747
rect 609 3539 643 3555
rect 727 3731 761 3747
rect 727 3539 761 3555
rect 845 3731 879 3781
rect 845 3539 879 3555
rect 963 3731 997 3747
rect 963 3539 997 3555
rect 1081 3731 1115 3781
rect 1081 3539 1115 3555
rect 770 3461 786 3495
rect 820 3461 836 3495
rect 652 3344 668 3378
rect 702 3344 718 3378
rect 256 3294 290 3310
rect -638 -5674 -630 -5593
rect -528 -5674 -527 -5593
rect -638 -5685 -527 -5674
rect -492 2987 -389 2995
rect -492 2911 -484 2987
rect -395 2911 -389 2987
rect -492 -8951 -389 2911
rect 256 2902 290 2918
rect 374 3294 408 3310
rect 374 2902 408 2918
rect 492 3294 526 3310
rect 609 3294 643 3310
rect 609 3102 643 3118
rect 727 3294 761 3310
rect 727 3102 761 3118
rect 492 2902 526 2918
rect 299 2834 315 2868
rect 349 2834 365 2868
rect 417 2834 433 2868
rect 467 2834 483 2868
rect -246 2793 69 2798
rect -246 2749 10 2793
rect 66 2749 69 2793
rect -246 2745 69 2749
rect 532 2763 700 2781
rect -246 -3061 -164 2745
rect 532 2707 548 2763
rect 682 2707 700 2763
rect 532 2691 700 2707
rect 300 1386 468 1402
rect 300 1316 316 1386
rect 452 1316 468 1386
rect 300 1300 468 1316
rect 837 1196 1107 1230
rect 11 1146 45 1162
rect 11 954 45 970
rect 129 1146 163 1162
rect 129 954 163 970
rect 247 1146 281 1162
rect 247 954 281 970
rect 365 1146 399 1162
rect 365 954 399 970
rect 483 1146 517 1162
rect 483 954 517 970
rect 601 1146 635 1162
rect 601 954 635 970
rect 719 1146 753 1162
rect 719 954 753 970
rect 837 1146 871 1196
rect 837 954 871 970
rect 955 1146 989 1162
rect 955 954 989 970
rect 1073 1146 1107 1196
rect 1073 954 1107 970
rect 762 876 778 910
rect 812 876 828 910
rect 644 759 660 793
rect 694 759 710 793
rect 248 709 282 725
rect 248 317 282 333
rect 366 709 400 725
rect 366 317 400 333
rect 484 709 518 725
rect 601 709 635 725
rect 601 517 635 533
rect 719 709 753 725
rect 719 517 753 533
rect 484 317 518 333
rect 291 249 307 283
rect 341 249 357 283
rect 409 249 425 283
rect 459 249 475 283
rect 524 178 692 196
rect 524 122 540 178
rect 674 122 692 178
rect 524 106 692 122
rect 281 -1892 449 -1876
rect 281 -1962 297 -1892
rect 433 -1962 449 -1892
rect 281 -1978 449 -1962
rect 818 -2082 1088 -2048
rect -8 -2132 26 -2116
rect -8 -2324 26 -2308
rect 110 -2132 144 -2116
rect 110 -2324 144 -2308
rect 228 -2132 262 -2116
rect 228 -2324 262 -2308
rect 346 -2132 380 -2116
rect 346 -2324 380 -2308
rect 464 -2132 498 -2116
rect 464 -2324 498 -2308
rect 582 -2132 616 -2116
rect 582 -2324 616 -2308
rect 700 -2132 734 -2116
rect 700 -2324 734 -2308
rect 818 -2132 852 -2082
rect 818 -2324 852 -2308
rect 936 -2132 970 -2116
rect 936 -2324 970 -2308
rect 1054 -2132 1088 -2082
rect 1054 -2324 1088 -2308
rect 743 -2402 759 -2368
rect 793 -2402 809 -2368
rect 625 -2519 641 -2485
rect 675 -2519 691 -2485
rect 229 -2569 263 -2553
rect 229 -2961 263 -2945
rect 347 -2569 381 -2553
rect 347 -2961 381 -2945
rect 465 -2569 499 -2553
rect 582 -2569 616 -2553
rect 582 -2761 616 -2745
rect 700 -2569 734 -2553
rect 700 -2761 734 -2745
rect 465 -2961 499 -2945
rect 272 -3029 288 -2995
rect 322 -3029 338 -2995
rect 390 -3029 406 -2995
rect 440 -3029 456 -2995
rect -246 -3066 19 -3061
rect -246 -3119 -46 -3066
rect 14 -3119 19 -3066
rect -246 -3123 19 -3119
rect 505 -3100 673 -3082
rect 505 -3156 521 -3100
rect 655 -3156 673 -3100
rect 505 -3172 673 -3156
rect 297 -4652 465 -4636
rect 297 -4722 313 -4652
rect 449 -4722 465 -4652
rect 297 -4738 465 -4722
rect 834 -4842 1104 -4808
rect 8 -4892 42 -4876
rect 8 -5084 42 -5068
rect 126 -4892 160 -4876
rect 126 -5084 160 -5068
rect 244 -4892 278 -4876
rect 244 -5084 278 -5068
rect 362 -4892 396 -4876
rect 362 -5084 396 -5068
rect 480 -4892 514 -4876
rect 480 -5084 514 -5068
rect 598 -4892 632 -4876
rect 598 -5084 632 -5068
rect 716 -4892 750 -4876
rect 716 -5084 750 -5068
rect 834 -4892 868 -4842
rect 834 -5084 868 -5068
rect 952 -4892 986 -4876
rect 952 -5084 986 -5068
rect 1070 -4892 1104 -4842
rect 1070 -5084 1104 -5068
rect 759 -5162 775 -5128
rect 809 -5162 825 -5128
rect 641 -5279 657 -5245
rect 691 -5279 707 -5245
rect 245 -5329 279 -5313
rect 245 -5721 279 -5705
rect 363 -5329 397 -5313
rect 363 -5721 397 -5705
rect 481 -5329 515 -5313
rect 598 -5329 632 -5313
rect 598 -5521 632 -5505
rect 716 -5329 750 -5313
rect 716 -5521 750 -5505
rect 481 -5721 515 -5705
rect 288 -5789 304 -5755
rect 338 -5789 354 -5755
rect 406 -5789 422 -5755
rect 456 -5789 472 -5755
rect 521 -5860 689 -5842
rect 521 -5916 537 -5860
rect 671 -5916 689 -5860
rect 521 -5932 689 -5916
rect -535 -8960 -344 -8951
rect -535 -9026 -510 -8960
rect -366 -9026 -344 -8960
rect -535 -9034 -344 -9026
rect -936 -9171 -925 -9100
rect -811 -9171 -798 -9100
rect -936 -9188 -798 -9171
rect 1619 -9223 1746 4170
rect 3304 3879 3527 3954
rect 3304 3878 3384 3879
rect 3304 3729 3383 3878
rect 3451 3730 3527 3879
rect 3450 3729 3527 3730
rect 3304 3623 3527 3729
rect 5786 3932 6009 4008
rect 5786 3783 5865 3932
rect 5932 3929 6009 3932
rect 5786 3780 5866 3783
rect 5933 3780 6009 3929
rect 5119 3712 5153 3728
rect 5119 3662 5153 3678
rect 5786 3677 6009 3780
rect 6933 3932 7156 4008
rect 6933 3931 7012 3932
rect 6933 3782 7008 3931
rect 7079 3783 7156 3932
rect 7075 3782 7156 3783
rect 6249 3718 6283 3734
rect 6249 3668 6283 3684
rect 6933 3677 7156 3782
rect 9853 3967 10076 4042
rect 9853 3966 9933 3967
rect 9853 3817 9932 3966
rect 10000 3818 10076 3967
rect 9999 3817 10076 3818
rect 9853 3711 10076 3817
rect 12335 4020 12558 4096
rect 12335 3871 12414 4020
rect 12481 4018 12558 4020
rect 12335 3869 12416 3871
rect 12483 3869 12558 4018
rect 11668 3800 11702 3816
rect 11668 3750 11702 3766
rect 12335 3765 12558 3869
rect 13482 4020 13705 4096
rect 13482 3871 13560 4020
rect 13628 3871 13705 4020
rect 12798 3806 12832 3822
rect 12798 3756 12832 3772
rect 13482 3765 13705 3871
rect 16507 3898 16730 3974
rect 16507 3748 16586 3898
rect 16653 3748 16730 3898
rect 18989 3953 19212 4028
rect 18989 3804 19067 3953
rect 19134 3952 19212 3953
rect 18989 3803 19068 3804
rect 19135 3803 19212 3952
rect 11668 3682 11702 3698
rect 5119 3594 5153 3610
rect 3735 3514 4005 3548
rect 5119 3544 5153 3560
rect 6249 3598 6283 3614
rect 10284 3602 10554 3636
rect 11668 3632 11702 3648
rect 12798 3686 12832 3702
rect 2909 3464 2943 3480
rect 2909 3272 2943 3288
rect 3027 3464 3061 3480
rect 3027 3272 3061 3288
rect 3145 3464 3179 3480
rect 3145 3272 3179 3288
rect 3263 3464 3297 3480
rect 3263 3272 3297 3288
rect 3381 3464 3415 3480
rect 3381 3272 3415 3288
rect 3499 3464 3533 3480
rect 3499 3272 3533 3288
rect 3617 3464 3651 3480
rect 3617 3272 3651 3288
rect 3735 3464 3769 3514
rect 3735 3272 3769 3288
rect 3853 3464 3887 3480
rect 3853 3272 3887 3288
rect 3971 3464 4005 3514
rect 3971 3272 4005 3288
rect 5234 3536 5268 3552
rect 3660 3194 3676 3228
rect 3710 3194 3726 3228
rect 5234 3144 5268 3160
rect 5352 3536 5386 3552
rect 5352 3144 5386 3160
rect 5470 3536 5504 3552
rect 5470 3144 5504 3160
rect 5588 3536 5622 3552
rect 5588 3144 5622 3160
rect 5706 3536 5740 3552
rect 5706 3144 5740 3160
rect 5824 3536 5858 3552
rect 5824 3144 5858 3160
rect 5942 3536 5976 3552
rect 6249 3548 6283 3564
rect 5942 3144 5976 3160
rect 6376 3540 6410 3556
rect 6376 3148 6410 3164
rect 6494 3540 6528 3556
rect 6494 3148 6528 3164
rect 6612 3540 6646 3556
rect 6612 3148 6646 3164
rect 6730 3540 6764 3556
rect 6730 3148 6764 3164
rect 6848 3540 6882 3556
rect 6848 3148 6882 3164
rect 6966 3540 7000 3556
rect 6966 3148 7000 3164
rect 7084 3540 7118 3556
rect 9458 3552 9492 3568
rect 9458 3360 9492 3376
rect 9576 3552 9610 3568
rect 9576 3360 9610 3376
rect 9694 3552 9728 3568
rect 9694 3360 9728 3376
rect 9812 3552 9846 3568
rect 9812 3360 9846 3376
rect 9930 3552 9964 3568
rect 9930 3360 9964 3376
rect 10048 3552 10082 3568
rect 10048 3360 10082 3376
rect 10166 3552 10200 3568
rect 10166 3360 10200 3376
rect 10284 3552 10318 3602
rect 10284 3360 10318 3376
rect 10402 3552 10436 3568
rect 10402 3360 10436 3376
rect 10520 3552 10554 3602
rect 10520 3360 10554 3376
rect 11783 3624 11817 3640
rect 10209 3282 10225 3316
rect 10259 3282 10275 3316
rect 11783 3232 11817 3248
rect 11901 3624 11935 3640
rect 11901 3232 11935 3248
rect 12019 3624 12053 3640
rect 12019 3232 12053 3248
rect 12137 3624 12171 3640
rect 12137 3232 12171 3248
rect 12255 3624 12289 3640
rect 12255 3232 12289 3248
rect 12373 3624 12407 3640
rect 12373 3232 12407 3248
rect 12491 3624 12525 3640
rect 12798 3636 12832 3652
rect 12491 3232 12525 3248
rect 12925 3628 12959 3644
rect 12925 3236 12959 3252
rect 13043 3628 13077 3644
rect 13043 3236 13077 3252
rect 13161 3628 13195 3644
rect 13161 3236 13195 3252
rect 13279 3628 13313 3644
rect 13279 3236 13313 3252
rect 13397 3628 13431 3644
rect 13397 3236 13431 3252
rect 13515 3628 13549 3644
rect 13515 3236 13549 3252
rect 13633 3628 13667 3644
rect 16507 3643 16730 3748
rect 18322 3732 18356 3748
rect 18322 3682 18356 3698
rect 18989 3697 19212 3803
rect 20136 3952 20359 4028
rect 20136 3803 20214 3952
rect 20282 3803 20359 3952
rect 19452 3738 19486 3754
rect 19452 3688 19486 3704
rect 20136 3697 20359 3803
rect 23132 3966 23355 4042
rect 23132 3817 23206 3966
rect 23278 3817 23355 3966
rect 23132 3711 23355 3817
rect 25614 4020 25837 4096
rect 25614 4018 25693 4020
rect 25614 3869 25690 4018
rect 25760 3871 25837 4020
rect 25757 3869 25837 3871
rect 24947 3800 24981 3816
rect 24947 3750 24981 3766
rect 25614 3765 25837 3869
rect 26761 4024 26984 4096
rect 26761 3875 26839 4024
rect 26906 4020 26984 4024
rect 26761 3871 26840 3875
rect 26907 3871 26984 4020
rect 26077 3806 26111 3822
rect 26077 3756 26111 3772
rect 26761 3765 26984 3871
rect 24947 3682 24981 3698
rect 18322 3614 18356 3630
rect 16938 3534 17208 3568
rect 18322 3564 18356 3580
rect 19452 3618 19486 3634
rect 16112 3484 16146 3500
rect 16112 3292 16146 3308
rect 16230 3484 16264 3500
rect 16230 3292 16264 3308
rect 16348 3484 16382 3500
rect 16348 3292 16382 3308
rect 16466 3484 16500 3500
rect 16466 3292 16500 3308
rect 16584 3484 16618 3500
rect 16584 3292 16618 3308
rect 16702 3484 16736 3500
rect 16702 3292 16736 3308
rect 16820 3484 16854 3500
rect 16820 3292 16854 3308
rect 16938 3484 16972 3534
rect 16938 3292 16972 3308
rect 17056 3484 17090 3500
rect 17056 3292 17090 3308
rect 17174 3484 17208 3534
rect 17174 3292 17208 3308
rect 18437 3556 18471 3572
rect 13633 3236 13667 3252
rect 16863 3214 16879 3248
rect 16913 3214 16929 3248
rect 10091 3165 10107 3199
rect 10141 3165 10157 3199
rect 18437 3164 18471 3180
rect 18555 3556 18589 3572
rect 18555 3164 18589 3180
rect 18673 3556 18707 3572
rect 18673 3164 18707 3180
rect 18791 3556 18825 3572
rect 18791 3164 18825 3180
rect 18909 3556 18943 3572
rect 18909 3164 18943 3180
rect 19027 3556 19061 3572
rect 19027 3164 19061 3180
rect 19145 3556 19179 3572
rect 19452 3568 19486 3584
rect 23563 3602 23833 3636
rect 24947 3632 24981 3648
rect 26077 3686 26111 3702
rect 19145 3164 19179 3180
rect 19579 3560 19613 3576
rect 19579 3168 19613 3184
rect 19697 3560 19731 3576
rect 19697 3168 19731 3184
rect 19815 3560 19849 3576
rect 19815 3168 19849 3184
rect 19933 3560 19967 3576
rect 19933 3168 19967 3184
rect 20051 3560 20085 3576
rect 20051 3168 20085 3184
rect 20169 3560 20203 3576
rect 20169 3168 20203 3184
rect 20287 3560 20321 3576
rect 22737 3552 22771 3568
rect 22737 3360 22771 3376
rect 22855 3552 22889 3568
rect 22855 3360 22889 3376
rect 22973 3552 23007 3568
rect 22973 3360 23007 3376
rect 23091 3552 23125 3568
rect 23091 3360 23125 3376
rect 23209 3552 23243 3568
rect 23209 3360 23243 3376
rect 23327 3552 23361 3568
rect 23327 3360 23361 3376
rect 23445 3552 23479 3568
rect 23445 3360 23479 3376
rect 23563 3552 23597 3602
rect 23563 3360 23597 3376
rect 23681 3552 23715 3568
rect 23681 3360 23715 3376
rect 23799 3552 23833 3602
rect 23799 3360 23833 3376
rect 25062 3624 25096 3640
rect 23488 3282 23504 3316
rect 23538 3282 23554 3316
rect 25062 3232 25096 3248
rect 25180 3624 25214 3640
rect 25180 3232 25214 3248
rect 25298 3624 25332 3640
rect 25298 3232 25332 3248
rect 25416 3624 25450 3640
rect 25416 3232 25450 3248
rect 25534 3624 25568 3640
rect 25534 3232 25568 3248
rect 25652 3624 25686 3640
rect 25652 3232 25686 3248
rect 25770 3624 25804 3640
rect 26077 3636 26111 3652
rect 25770 3232 25804 3248
rect 26204 3628 26238 3644
rect 26204 3236 26238 3252
rect 26322 3628 26356 3644
rect 26322 3236 26356 3252
rect 26440 3628 26474 3644
rect 26440 3236 26474 3252
rect 26558 3628 26592 3644
rect 26558 3236 26592 3252
rect 26676 3628 26710 3644
rect 26676 3236 26710 3252
rect 26794 3628 26828 3644
rect 26794 3236 26828 3252
rect 26912 3628 26946 3644
rect 26912 3236 26946 3252
rect 20287 3168 20321 3184
rect 23370 3165 23386 3199
rect 23420 3165 23436 3199
rect 7084 3148 7118 3164
rect 28823 3153 28991 3169
rect 9695 3115 9729 3131
rect 3542 3077 3558 3111
rect 3592 3077 3608 3111
rect 3146 3027 3180 3043
rect 3146 2635 3180 2651
rect 3264 3027 3298 3043
rect 3264 2635 3298 2651
rect 3382 3027 3416 3043
rect 3499 3027 3533 3043
rect 3499 2835 3533 2851
rect 3617 3027 3651 3043
rect 3617 2835 3651 2851
rect 5423 2804 5439 2838
rect 5473 2804 5489 2838
rect 6565 2808 6581 2842
rect 6615 2808 6631 2842
rect 5144 2753 5178 2769
rect 3382 2635 3416 2651
rect 3669 2701 3918 2744
rect 3669 2611 3716 2701
rect 3879 2611 3918 2701
rect 3189 2567 3205 2601
rect 3239 2567 3255 2601
rect 3307 2567 3323 2601
rect 3357 2567 3373 2601
rect 3669 2572 3918 2611
rect 5144 2561 5178 2577
rect 5262 2753 5296 2769
rect 5262 2561 5296 2577
rect 5380 2753 5414 2769
rect 5380 2561 5414 2577
rect 5498 2753 5532 2769
rect 5498 2561 5532 2577
rect 5663 2753 5697 2769
rect 5663 2561 5697 2577
rect 5781 2753 5815 2769
rect 5781 2561 5815 2577
rect 5899 2753 5933 2769
rect 5899 2561 5933 2577
rect 6017 2753 6051 2769
rect 6017 2561 6051 2577
rect 6286 2757 6320 2773
rect 6286 2565 6320 2581
rect 6404 2757 6438 2773
rect 6404 2565 6438 2581
rect 6522 2757 6556 2773
rect 6522 2565 6556 2581
rect 6640 2757 6674 2773
rect 6640 2565 6674 2581
rect 6805 2757 6839 2773
rect 6805 2565 6839 2581
rect 6923 2757 6957 2773
rect 6923 2565 6957 2581
rect 7041 2757 7075 2773
rect 7041 2565 7075 2581
rect 7159 2757 7193 2773
rect 9695 2723 9729 2739
rect 9813 3115 9847 3131
rect 9813 2723 9847 2739
rect 9931 3115 9965 3131
rect 10048 3115 10082 3131
rect 10048 2923 10082 2939
rect 10166 3115 10200 3131
rect 16745 3097 16761 3131
rect 16795 3097 16811 3131
rect 22974 3115 23008 3131
rect 10166 2923 10200 2939
rect 16349 3047 16383 3063
rect 11972 2892 11988 2926
rect 12022 2892 12038 2926
rect 13114 2896 13130 2930
rect 13164 2896 13180 2930
rect 11693 2841 11727 2857
rect 9931 2723 9965 2739
rect 10218 2789 10467 2832
rect 10218 2699 10265 2789
rect 10428 2699 10467 2789
rect 9738 2655 9754 2689
rect 9788 2655 9804 2689
rect 9856 2655 9872 2689
rect 9906 2655 9922 2689
rect 10218 2660 10467 2699
rect 11693 2649 11727 2665
rect 11811 2841 11845 2857
rect 11811 2649 11845 2665
rect 11929 2841 11963 2857
rect 11929 2649 11963 2665
rect 12047 2841 12081 2857
rect 12047 2649 12081 2665
rect 12212 2841 12246 2857
rect 12212 2649 12246 2665
rect 12330 2841 12364 2857
rect 12330 2649 12364 2665
rect 12448 2841 12482 2857
rect 12448 2649 12482 2665
rect 12566 2841 12600 2857
rect 12566 2649 12600 2665
rect 12835 2845 12869 2861
rect 12835 2653 12869 2669
rect 12953 2845 12987 2861
rect 12953 2653 12987 2669
rect 13071 2845 13105 2861
rect 13071 2653 13105 2669
rect 13189 2845 13223 2861
rect 13189 2653 13223 2669
rect 13354 2845 13388 2861
rect 13354 2653 13388 2669
rect 13472 2845 13506 2861
rect 13472 2653 13506 2669
rect 13590 2845 13624 2861
rect 13590 2653 13624 2669
rect 13708 2845 13742 2861
rect 13708 2653 13742 2669
rect 16349 2655 16383 2671
rect 16467 3047 16501 3063
rect 16467 2655 16501 2671
rect 16585 3047 16619 3063
rect 16702 3047 16736 3063
rect 16702 2855 16736 2871
rect 16820 3047 16854 3063
rect 16820 2855 16854 2871
rect 18626 2824 18642 2858
rect 18676 2824 18692 2858
rect 19768 2828 19784 2862
rect 19818 2828 19834 2862
rect 18347 2773 18381 2789
rect 16585 2655 16619 2671
rect 16872 2721 17121 2764
rect 16872 2631 16919 2721
rect 17082 2631 17121 2721
rect 16392 2587 16408 2621
rect 16442 2587 16458 2621
rect 16510 2587 16526 2621
rect 16560 2587 16576 2621
rect 16872 2592 17121 2631
rect 18347 2581 18381 2597
rect 18465 2773 18499 2789
rect 18465 2581 18499 2597
rect 18583 2773 18617 2789
rect 18583 2581 18617 2597
rect 18701 2773 18735 2789
rect 18701 2581 18735 2597
rect 18866 2773 18900 2789
rect 18866 2581 18900 2597
rect 18984 2773 19018 2789
rect 18984 2581 19018 2597
rect 19102 2773 19136 2789
rect 19102 2581 19136 2597
rect 19220 2773 19254 2789
rect 19220 2581 19254 2597
rect 19489 2777 19523 2793
rect 19489 2585 19523 2601
rect 19607 2777 19641 2793
rect 19607 2585 19641 2601
rect 19725 2777 19759 2793
rect 19725 2585 19759 2601
rect 19843 2777 19877 2793
rect 19843 2585 19877 2601
rect 20008 2777 20042 2793
rect 20008 2585 20042 2601
rect 20126 2777 20160 2793
rect 20126 2585 20160 2601
rect 20244 2777 20278 2793
rect 20244 2585 20278 2601
rect 20362 2777 20396 2793
rect 22974 2723 23008 2739
rect 23092 3115 23126 3131
rect 23092 2723 23126 2739
rect 23210 3115 23244 3131
rect 23327 3115 23361 3131
rect 23327 2923 23361 2939
rect 23445 3115 23479 3131
rect 28823 3083 28839 3153
rect 28975 3083 28991 3153
rect 28823 3067 28991 3083
rect 23445 2923 23479 2939
rect 29360 2963 29630 2997
rect 25251 2892 25267 2926
rect 25301 2892 25317 2926
rect 26393 2896 26409 2930
rect 26443 2896 26459 2930
rect 28534 2913 28568 2929
rect 24972 2841 25006 2857
rect 23210 2723 23244 2739
rect 23497 2789 23746 2832
rect 23497 2699 23544 2789
rect 23707 2699 23746 2789
rect 23017 2655 23033 2689
rect 23067 2655 23083 2689
rect 23135 2655 23151 2689
rect 23185 2655 23201 2689
rect 23497 2660 23746 2699
rect 24972 2649 25006 2665
rect 25090 2841 25124 2857
rect 25090 2649 25124 2665
rect 25208 2841 25242 2857
rect 25208 2649 25242 2665
rect 25326 2841 25360 2857
rect 25326 2649 25360 2665
rect 25491 2841 25525 2857
rect 25491 2649 25525 2665
rect 25609 2841 25643 2857
rect 25609 2649 25643 2665
rect 25727 2841 25761 2857
rect 25727 2649 25761 2665
rect 25845 2841 25879 2857
rect 25845 2649 25879 2665
rect 26114 2845 26148 2861
rect 26114 2653 26148 2669
rect 26232 2845 26266 2861
rect 26232 2653 26266 2669
rect 26350 2845 26384 2861
rect 26350 2653 26384 2669
rect 26468 2845 26502 2861
rect 26468 2653 26502 2669
rect 26633 2845 26667 2861
rect 26633 2653 26667 2669
rect 26751 2845 26785 2861
rect 26751 2653 26785 2669
rect 26869 2845 26903 2861
rect 26869 2653 26903 2669
rect 26987 2845 27021 2861
rect 28534 2721 28568 2737
rect 28652 2913 28686 2929
rect 28652 2721 28686 2737
rect 28770 2913 28804 2929
rect 28770 2721 28804 2737
rect 28888 2913 28922 2929
rect 28888 2721 28922 2737
rect 29006 2913 29040 2929
rect 29006 2721 29040 2737
rect 29124 2913 29158 2929
rect 29124 2721 29158 2737
rect 29242 2913 29276 2929
rect 29242 2721 29276 2737
rect 29360 2913 29394 2963
rect 29360 2721 29394 2737
rect 29478 2913 29512 2929
rect 29478 2721 29512 2737
rect 29596 2913 29630 2963
rect 29596 2721 29630 2737
rect 26987 2653 27021 2669
rect 29285 2643 29301 2677
rect 29335 2643 29351 2677
rect 20362 2585 20396 2601
rect 7159 2565 7193 2581
rect 29167 2526 29183 2560
rect 29217 2526 29233 2560
rect 28771 2476 28805 2492
rect 11708 2418 11880 2465
rect 5159 2330 5331 2377
rect 3318 2228 3541 2304
rect 3318 2079 3396 2228
rect 3464 2079 3541 2228
rect 5159 2167 5198 2330
rect 5288 2167 5331 2330
rect 5159 2128 5331 2167
rect 6301 2328 6473 2375
rect 6301 2165 6340 2328
rect 6430 2165 6473 2328
rect 6301 2126 6473 2165
rect 9867 2316 10090 2392
rect 9867 2167 9946 2316
rect 10013 2315 10090 2316
rect 9867 2166 9947 2167
rect 10014 2166 10090 2315
rect 11708 2255 11747 2418
rect 11837 2255 11880 2418
rect 11708 2216 11880 2255
rect 12850 2416 13022 2463
rect 12850 2253 12889 2416
rect 12979 2253 13022 2416
rect 24987 2418 25159 2465
rect 18362 2350 18534 2397
rect 12850 2214 13022 2253
rect 16521 2249 16744 2324
rect 16521 2248 16601 2249
rect 3318 1973 3541 2079
rect 9867 2061 10090 2166
rect 16521 2099 16600 2248
rect 16668 2100 16744 2249
rect 18362 2187 18401 2350
rect 18491 2187 18534 2350
rect 18362 2148 18534 2187
rect 19504 2348 19676 2395
rect 19504 2185 19543 2348
rect 19633 2185 19676 2348
rect 19504 2146 19676 2185
rect 23146 2316 23369 2392
rect 23146 2167 23225 2316
rect 23292 2315 23369 2316
rect 23146 2166 23229 2167
rect 23296 2166 23369 2315
rect 24987 2255 25026 2418
rect 25116 2255 25159 2418
rect 24987 2253 25030 2255
rect 25097 2253 25159 2255
rect 24987 2216 25159 2253
rect 26129 2416 26301 2463
rect 26129 2253 26168 2416
rect 26258 2253 26301 2416
rect 26129 2214 26301 2253
rect 16667 2099 16744 2100
rect 3749 1864 4019 1898
rect 2923 1814 2957 1830
rect 2923 1622 2957 1638
rect 3041 1814 3075 1830
rect 3041 1622 3075 1638
rect 3159 1814 3193 1830
rect 3159 1622 3193 1638
rect 3277 1814 3311 1830
rect 3277 1622 3311 1638
rect 3395 1814 3429 1830
rect 3395 1622 3429 1638
rect 3513 1814 3547 1830
rect 3513 1622 3547 1638
rect 3631 1814 3665 1830
rect 3631 1622 3665 1638
rect 3749 1814 3783 1864
rect 3749 1622 3783 1638
rect 3867 1814 3901 1830
rect 3867 1622 3901 1638
rect 3985 1814 4019 1864
rect 3985 1622 4019 1638
rect 7029 1886 7254 1961
rect 10298 1952 10568 1986
rect 7029 1736 7108 1886
rect 7175 1736 7254 1886
rect 7029 1630 7254 1736
rect 9472 1902 9506 1918
rect 9472 1710 9506 1726
rect 9590 1902 9624 1918
rect 9590 1710 9624 1726
rect 9708 1902 9742 1918
rect 9708 1710 9742 1726
rect 9826 1902 9860 1918
rect 9826 1710 9860 1726
rect 9944 1902 9978 1918
rect 9944 1710 9978 1726
rect 10062 1902 10096 1918
rect 10062 1710 10096 1726
rect 10180 1902 10214 1918
rect 10180 1710 10214 1726
rect 10298 1902 10332 1952
rect 10298 1710 10332 1726
rect 10416 1902 10450 1918
rect 10416 1710 10450 1726
rect 10534 1902 10568 1952
rect 10534 1710 10568 1726
rect 13578 1973 13803 2049
rect 16521 1993 16744 2099
rect 23146 2061 23369 2166
rect 28771 2084 28805 2100
rect 28889 2476 28923 2492
rect 28889 2084 28923 2100
rect 29007 2476 29041 2492
rect 29124 2476 29158 2492
rect 29124 2284 29158 2300
rect 29242 2476 29276 2492
rect 29242 2284 29276 2300
rect 29007 2084 29041 2100
rect 13578 1824 13657 1973
rect 13729 1824 13803 1973
rect 16952 1884 17222 1918
rect 13578 1718 13803 1824
rect 16126 1834 16160 1850
rect 10223 1632 10239 1666
rect 10273 1632 10289 1666
rect 16126 1642 16160 1658
rect 16244 1834 16278 1850
rect 16244 1642 16278 1658
rect 16362 1834 16396 1850
rect 16362 1642 16396 1658
rect 16480 1834 16514 1850
rect 16480 1642 16514 1658
rect 16598 1834 16632 1850
rect 16598 1642 16632 1658
rect 16716 1834 16750 1850
rect 16716 1642 16750 1658
rect 16834 1834 16868 1850
rect 16834 1642 16868 1658
rect 16952 1834 16986 1884
rect 16952 1642 16986 1658
rect 17070 1834 17104 1850
rect 17070 1642 17104 1658
rect 17188 1834 17222 1884
rect 17188 1642 17222 1658
rect 20232 1905 20457 1981
rect 23577 1952 23847 1986
rect 20232 1901 20311 1905
rect 20232 1752 20308 1901
rect 20378 1756 20457 1905
rect 20375 1752 20457 1756
rect 20232 1650 20457 1752
rect 22751 1902 22785 1918
rect 22751 1710 22785 1726
rect 22869 1902 22903 1918
rect 22869 1710 22903 1726
rect 22987 1902 23021 1918
rect 22987 1710 23021 1726
rect 23105 1902 23139 1918
rect 23105 1710 23139 1726
rect 23223 1902 23257 1918
rect 23223 1710 23257 1726
rect 23341 1902 23375 1918
rect 23341 1710 23375 1726
rect 23459 1902 23493 1918
rect 23459 1710 23493 1726
rect 23577 1902 23611 1952
rect 23577 1710 23611 1726
rect 23695 1902 23729 1918
rect 23695 1710 23729 1726
rect 23813 1902 23847 1952
rect 23813 1710 23847 1726
rect 26857 1973 27082 2049
rect 28814 2016 28830 2050
rect 28864 2016 28880 2050
rect 28932 2016 28948 2050
rect 28982 2016 28998 2050
rect 26857 1821 26936 1973
rect 27003 1821 27082 1973
rect 29047 1945 29215 1963
rect 29047 1889 29063 1945
rect 29197 1889 29215 1945
rect 29047 1873 29215 1889
rect 26857 1718 27082 1821
rect 23502 1632 23518 1666
rect 23552 1632 23568 1666
rect 3674 1544 3690 1578
rect 3724 1544 3740 1578
rect 10105 1515 10121 1549
rect 10155 1515 10171 1549
rect 11774 1538 12044 1573
rect 11420 1485 11454 1501
rect 3556 1427 3572 1461
rect 3606 1427 3622 1461
rect 5225 1450 5495 1485
rect 4871 1397 4905 1413
rect 3160 1377 3194 1393
rect 2014 1037 2274 1039
rect 2012 1008 2274 1037
rect 2012 898 2121 1008
rect 2239 898 2274 1008
rect 3160 985 3194 1001
rect 3278 1377 3312 1393
rect 3278 985 3312 1001
rect 3396 1377 3430 1393
rect 3513 1377 3547 1393
rect 3513 1185 3547 1201
rect 3631 1377 3665 1393
rect 3631 1185 3665 1201
rect 4387 1251 4657 1286
rect 4387 1197 4421 1251
rect 3396 985 3430 1001
rect 3683 1051 3932 1094
rect 3683 961 3730 1051
rect 3893 961 3932 1051
rect 4387 1005 4421 1021
rect 4505 1197 4539 1213
rect 4505 1005 4539 1021
rect 4623 1197 4657 1251
rect 4623 1005 4657 1021
rect 4741 1197 4775 1213
rect 4741 1005 4775 1021
rect 4871 1005 4905 1021
rect 4989 1397 5023 1413
rect 4989 1005 5023 1021
rect 5107 1397 5141 1413
rect 5107 1005 5141 1021
rect 5225 1397 5259 1450
rect 5225 1005 5259 1021
rect 5343 1397 5377 1413
rect 5343 1005 5377 1021
rect 5461 1397 5495 1450
rect 7123 1450 7393 1485
rect 5461 1005 5495 1021
rect 5579 1397 5613 1413
rect 6769 1397 6803 1413
rect 6285 1251 6555 1286
rect 5579 1005 5613 1021
rect 5708 1197 5742 1213
rect 5708 1005 5742 1021
rect 5826 1197 5860 1213
rect 5826 1005 5860 1021
rect 5944 1197 5978 1213
rect 5944 1005 5978 1021
rect 6062 1197 6096 1213
rect 6062 1005 6096 1021
rect 6285 1197 6319 1251
rect 6285 1005 6319 1021
rect 6403 1197 6437 1213
rect 6403 1005 6437 1021
rect 6521 1197 6555 1251
rect 6521 1005 6555 1021
rect 6639 1197 6673 1213
rect 6639 1005 6673 1021
rect 6769 1005 6803 1021
rect 6887 1397 6921 1413
rect 6887 1005 6921 1021
rect 7005 1397 7039 1413
rect 7005 1005 7039 1021
rect 7123 1397 7157 1450
rect 7123 1005 7157 1021
rect 7241 1397 7275 1413
rect 7241 1005 7275 1021
rect 7359 1397 7393 1450
rect 9709 1465 9743 1481
rect 7359 1005 7393 1021
rect 7477 1397 7511 1413
rect 7477 1005 7511 1021
rect 7606 1197 7640 1213
rect 7606 1005 7640 1021
rect 7724 1197 7758 1213
rect 7724 1005 7758 1021
rect 7842 1197 7876 1213
rect 7842 1005 7876 1021
rect 7960 1197 7994 1213
rect 9709 1073 9743 1089
rect 9827 1465 9861 1481
rect 9827 1073 9861 1089
rect 9945 1465 9979 1481
rect 10062 1465 10096 1481
rect 10062 1273 10096 1289
rect 10180 1465 10214 1481
rect 10180 1273 10214 1289
rect 10936 1339 11206 1374
rect 10936 1285 10970 1339
rect 9945 1073 9979 1089
rect 10232 1139 10481 1182
rect 10232 1049 10279 1139
rect 10442 1049 10481 1139
rect 10936 1093 10970 1109
rect 11054 1285 11088 1301
rect 11054 1093 11088 1109
rect 11172 1285 11206 1339
rect 11172 1093 11206 1109
rect 11290 1285 11324 1301
rect 11290 1093 11324 1109
rect 11420 1093 11454 1109
rect 11538 1485 11572 1501
rect 11538 1093 11572 1109
rect 11656 1485 11690 1501
rect 11656 1093 11690 1109
rect 11774 1485 11808 1538
rect 11774 1093 11808 1109
rect 11892 1485 11926 1501
rect 11892 1093 11926 1109
rect 12010 1485 12044 1538
rect 13672 1538 13942 1573
rect 16877 1564 16893 1598
rect 16927 1564 16943 1598
rect 12010 1093 12044 1109
rect 12128 1485 12162 1501
rect 13318 1485 13352 1501
rect 12834 1339 13104 1374
rect 12128 1093 12162 1109
rect 12257 1285 12291 1301
rect 12257 1093 12291 1109
rect 12375 1285 12409 1301
rect 12375 1093 12409 1109
rect 12493 1285 12527 1301
rect 12493 1093 12527 1109
rect 12611 1285 12645 1301
rect 12611 1093 12645 1109
rect 12834 1285 12868 1339
rect 12834 1093 12868 1109
rect 12952 1285 12986 1301
rect 12952 1093 12986 1109
rect 13070 1285 13104 1339
rect 13070 1093 13104 1109
rect 13188 1285 13222 1301
rect 13188 1093 13222 1109
rect 13318 1093 13352 1109
rect 13436 1485 13470 1501
rect 13436 1093 13470 1109
rect 13554 1485 13588 1501
rect 13554 1093 13588 1109
rect 13672 1485 13706 1538
rect 13672 1093 13706 1109
rect 13790 1485 13824 1501
rect 13790 1093 13824 1109
rect 13908 1485 13942 1538
rect 23384 1515 23400 1549
rect 23434 1515 23450 1549
rect 25053 1538 25323 1573
rect 13908 1093 13942 1109
rect 14026 1485 14060 1501
rect 16759 1447 16775 1481
rect 16809 1447 16825 1481
rect 18428 1470 18698 1505
rect 18074 1417 18108 1433
rect 16363 1397 16397 1413
rect 14026 1093 14060 1109
rect 14155 1285 14189 1301
rect 14155 1093 14189 1109
rect 14273 1285 14307 1301
rect 14273 1093 14307 1109
rect 14391 1285 14425 1301
rect 14391 1093 14425 1109
rect 14509 1285 14543 1301
rect 14509 1093 14543 1109
rect 7960 1005 7994 1021
rect 9752 1005 9768 1039
rect 9802 1005 9818 1039
rect 9870 1005 9886 1039
rect 9920 1005 9936 1039
rect 10232 1010 10481 1049
rect 15257 1037 15483 1059
rect 3203 917 3219 951
rect 3253 917 3269 951
rect 3321 917 3337 951
rect 3371 917 3387 951
rect 3683 922 3932 961
rect 15257 920 15323 1037
rect 15462 920 15483 1037
rect 16363 1005 16397 1021
rect 16481 1397 16515 1413
rect 16481 1005 16515 1021
rect 16599 1397 16633 1413
rect 16716 1397 16750 1413
rect 16716 1205 16750 1221
rect 16834 1397 16868 1413
rect 16834 1205 16868 1221
rect 17590 1271 17860 1306
rect 17590 1217 17624 1271
rect 16599 1005 16633 1021
rect 16886 1071 17135 1114
rect 16886 981 16933 1071
rect 17096 981 17135 1071
rect 17590 1025 17624 1041
rect 17708 1217 17742 1233
rect 17708 1025 17742 1041
rect 17826 1217 17860 1271
rect 17826 1025 17860 1041
rect 17944 1217 17978 1233
rect 17944 1025 17978 1041
rect 18074 1025 18108 1041
rect 18192 1417 18226 1433
rect 18192 1025 18226 1041
rect 18310 1417 18344 1433
rect 18310 1025 18344 1041
rect 18428 1417 18462 1470
rect 18428 1025 18462 1041
rect 18546 1417 18580 1433
rect 18546 1025 18580 1041
rect 18664 1417 18698 1470
rect 20326 1470 20596 1505
rect 24699 1485 24733 1501
rect 18664 1025 18698 1041
rect 18782 1417 18816 1433
rect 19972 1417 20006 1433
rect 19488 1271 19758 1306
rect 18782 1025 18816 1041
rect 18911 1217 18945 1233
rect 18911 1025 18945 1041
rect 19029 1217 19063 1233
rect 19029 1025 19063 1041
rect 19147 1217 19181 1233
rect 19147 1025 19181 1041
rect 19265 1217 19299 1233
rect 19265 1025 19299 1041
rect 19488 1217 19522 1271
rect 19488 1025 19522 1041
rect 19606 1217 19640 1233
rect 19606 1025 19640 1041
rect 19724 1217 19758 1271
rect 19724 1025 19758 1041
rect 19842 1217 19876 1233
rect 19842 1025 19876 1041
rect 19972 1025 20006 1041
rect 20090 1417 20124 1433
rect 20090 1025 20124 1041
rect 20208 1417 20242 1433
rect 20208 1025 20242 1041
rect 20326 1417 20360 1470
rect 20326 1025 20360 1041
rect 20444 1417 20478 1433
rect 20444 1025 20478 1041
rect 20562 1417 20596 1470
rect 22988 1465 23022 1481
rect 20562 1025 20596 1041
rect 20680 1417 20714 1433
rect 20680 1025 20714 1041
rect 20809 1217 20843 1233
rect 20809 1025 20843 1041
rect 20927 1217 20961 1233
rect 20927 1025 20961 1041
rect 21045 1217 21079 1233
rect 21045 1025 21079 1041
rect 21163 1217 21197 1233
rect 22988 1073 23022 1089
rect 23106 1465 23140 1481
rect 23106 1073 23140 1089
rect 23224 1465 23258 1481
rect 23341 1465 23375 1481
rect 23341 1273 23375 1289
rect 23459 1465 23493 1481
rect 23459 1273 23493 1289
rect 24215 1339 24485 1374
rect 24215 1285 24249 1339
rect 23224 1073 23258 1089
rect 23511 1139 23760 1182
rect 21163 1025 21197 1041
rect 23511 1049 23558 1139
rect 23721 1049 23760 1139
rect 24215 1093 24249 1109
rect 24333 1285 24367 1301
rect 24333 1093 24367 1109
rect 24451 1285 24485 1339
rect 24451 1093 24485 1109
rect 24569 1285 24603 1301
rect 24569 1093 24603 1109
rect 24699 1093 24733 1109
rect 24817 1485 24851 1501
rect 24817 1093 24851 1109
rect 24935 1485 24969 1501
rect 24935 1093 24969 1109
rect 25053 1485 25087 1538
rect 25053 1093 25087 1109
rect 25171 1485 25205 1501
rect 25171 1093 25205 1109
rect 25289 1485 25323 1538
rect 26951 1538 27221 1573
rect 25289 1093 25323 1109
rect 25407 1485 25441 1501
rect 26597 1485 26631 1501
rect 26113 1339 26383 1374
rect 25407 1093 25441 1109
rect 25536 1285 25570 1301
rect 25536 1093 25570 1109
rect 25654 1285 25688 1301
rect 25654 1093 25688 1109
rect 25772 1285 25806 1301
rect 25772 1093 25806 1109
rect 25890 1285 25924 1301
rect 25890 1093 25924 1109
rect 26113 1285 26147 1339
rect 26113 1093 26147 1109
rect 26231 1285 26265 1301
rect 26231 1093 26265 1109
rect 26349 1285 26383 1339
rect 26349 1093 26383 1109
rect 26467 1285 26501 1301
rect 26467 1093 26501 1109
rect 26597 1093 26631 1109
rect 26715 1485 26749 1501
rect 26715 1093 26749 1109
rect 26833 1485 26867 1501
rect 26833 1093 26867 1109
rect 26951 1485 26985 1538
rect 26951 1093 26985 1109
rect 27069 1485 27103 1501
rect 27069 1093 27103 1109
rect 27187 1485 27221 1538
rect 27187 1093 27221 1109
rect 27305 1485 27339 1501
rect 27305 1093 27339 1109
rect 27434 1285 27468 1301
rect 27434 1093 27468 1109
rect 27552 1285 27586 1301
rect 27552 1093 27586 1109
rect 27670 1285 27704 1301
rect 27670 1093 27704 1109
rect 27788 1285 27822 1301
rect 27788 1093 27822 1109
rect 23031 1005 23047 1039
rect 23081 1005 23097 1039
rect 23149 1005 23165 1039
rect 23199 1005 23215 1039
rect 23511 1010 23760 1049
rect 16406 937 16422 971
rect 16456 937 16472 971
rect 16524 937 16540 971
rect 16574 937 16590 971
rect 16886 942 17135 981
rect 15257 908 15483 920
rect 2012 888 2274 898
rect 2012 -1510 2176 888
rect 12400 871 12434 887
rect 12400 821 12434 837
rect 14490 850 14557 866
rect 14490 816 14507 850
rect 14541 816 14557 850
rect 5851 783 5885 799
rect 11363 792 11397 808
rect 5851 733 5885 749
rect 7941 762 8008 778
rect 7941 728 7958 762
rect 7992 728 8008 762
rect 4814 704 4848 720
rect 3313 624 3536 700
rect 3313 475 3392 624
rect 3459 622 3536 624
rect 3313 473 3394 475
rect 3461 473 3536 622
rect 3313 369 3536 473
rect 4932 704 4966 720
rect 4814 312 4848 328
rect 4931 328 4932 375
rect 5050 704 5084 720
rect 4966 328 4967 375
rect 3744 260 4014 294
rect 2918 210 2952 226
rect 2918 18 2952 34
rect 3036 210 3070 226
rect 3036 18 3070 34
rect 3154 210 3188 226
rect 3154 18 3188 34
rect 3272 210 3306 226
rect 3272 18 3306 34
rect 3390 210 3424 226
rect 3390 18 3424 34
rect 3508 210 3542 226
rect 3508 18 3542 34
rect 3626 210 3660 226
rect 3626 18 3660 34
rect 3744 210 3778 260
rect 3744 18 3778 34
rect 3862 210 3896 226
rect 3862 18 3896 34
rect 3980 210 4014 260
rect 4931 270 4967 328
rect 5168 704 5202 720
rect 5050 312 5084 328
rect 5166 328 5168 375
rect 5166 270 5202 328
rect 5286 704 5320 720
rect 5286 312 5320 328
rect 5404 704 5438 720
rect 5522 704 5556 720
rect 5438 328 5440 374
rect 5404 270 5440 328
rect 5522 312 5556 328
rect 6712 704 6746 720
rect 6830 704 6864 720
rect 6712 312 6746 328
rect 6829 328 6830 375
rect 6948 704 6982 720
rect 6864 328 6865 375
rect 6027 270 6524 288
rect 4931 267 6524 270
rect 4931 233 6472 267
rect 6506 233 6524 267
rect 4931 230 6524 233
rect 6829 270 6865 328
rect 7066 704 7100 720
rect 6948 312 6982 328
rect 7064 328 7066 375
rect 7064 270 7100 328
rect 7184 704 7218 720
rect 7184 312 7218 328
rect 7302 704 7336 720
rect 7420 704 7454 720
rect 7941 712 8008 728
rect 9862 715 10085 788
rect 7336 328 7338 374
rect 7302 270 7338 328
rect 9862 566 9939 715
rect 10006 712 10085 715
rect 9862 563 9941 566
rect 10008 563 10085 712
rect 9862 457 10085 563
rect 11481 792 11515 808
rect 11363 400 11397 416
rect 11480 416 11481 463
rect 11599 792 11633 808
rect 11515 416 11516 463
rect 7420 312 7454 328
rect 10293 348 10563 382
rect 7925 270 8188 300
rect 6829 230 8188 270
rect 4950 229 6524 230
rect 6848 229 8188 230
rect 4828 140 4895 156
rect 4828 106 4844 140
rect 4878 106 4895 140
rect 4828 90 4895 106
rect 3980 18 4014 34
rect 4659 73 4693 89
rect 4659 23 4693 39
rect 5005 -12 5039 229
rect 6027 212 6524 229
rect 5475 140 5542 156
rect 5475 106 5492 140
rect 5526 106 5542 140
rect 5475 90 5542 106
rect 6726 140 6793 156
rect 6726 106 6742 140
rect 6776 106 6793 140
rect 6726 90 6793 106
rect 5782 72 5816 88
rect 5094 22 5110 56
rect 5144 22 5160 56
rect 5212 23 5228 57
rect 5262 23 5278 57
rect 5782 22 5816 38
rect 6557 73 6591 89
rect 6557 23 6591 39
rect 6903 -12 6937 229
rect 7925 200 8188 229
rect 7371 141 7438 157
rect 7371 107 7388 141
rect 7422 107 7438 141
rect 7371 91 7438 107
rect 7680 72 7714 88
rect 6992 22 7008 56
rect 7042 22 7058 56
rect 7110 23 7126 57
rect 7160 23 7176 57
rect 7680 22 7714 38
rect 3669 -60 3685 -26
rect 3719 -60 3735 -26
rect 4512 -28 4546 -12
rect 3551 -177 3567 -143
rect 3601 -177 3617 -143
rect 3155 -227 3189 -211
rect 3155 -619 3189 -603
rect 3273 -227 3307 -211
rect 3273 -619 3307 -603
rect 3391 -227 3425 -211
rect 3508 -227 3542 -211
rect 3508 -419 3542 -403
rect 3626 -227 3660 -211
rect 4512 -220 4546 -204
rect 4630 -28 4664 -12
rect 4630 -220 4664 -204
rect 4932 -28 4966 -12
rect 3626 -419 3660 -403
rect 5005 -28 5084 -12
rect 5005 -58 5050 -28
rect 4932 -471 4967 -404
rect 5050 -420 5084 -404
rect 5168 -28 5202 -12
rect 5168 -420 5202 -404
rect 5286 -28 5320 -12
rect 5404 -28 5438 -12
rect 5810 -28 5844 -12
rect 5810 -220 5844 -204
rect 5928 -28 5962 -12
rect 5928 -220 5962 -204
rect 6410 -28 6444 -12
rect 6410 -220 6444 -204
rect 6528 -28 6562 -12
rect 6528 -220 6562 -204
rect 6830 -28 6864 -12
rect 5286 -420 5320 -404
rect 5403 -471 5438 -404
rect 4932 -506 5438 -471
rect 6903 -28 6982 -12
rect 6903 -58 6948 -28
rect 6830 -471 6865 -404
rect 6948 -420 6982 -404
rect 7066 -28 7100 -12
rect 7066 -420 7100 -404
rect 7184 -28 7218 -12
rect 7302 -28 7336 -12
rect 7708 -28 7742 -12
rect 7708 -220 7742 -204
rect 7826 -28 7860 -12
rect 7826 -220 7860 -204
rect 7184 -420 7218 -404
rect 7301 -471 7336 -404
rect 6830 -506 7336 -471
rect 3391 -619 3425 -603
rect 3678 -553 3927 -510
rect 3678 -643 3725 -553
rect 3888 -643 3927 -553
rect 3198 -687 3214 -653
rect 3248 -687 3264 -653
rect 3316 -687 3332 -653
rect 3366 -687 3382 -653
rect 3678 -682 3927 -643
rect 5103 -713 5275 -666
rect 5103 -876 5142 -713
rect 5232 -876 5275 -713
rect 5103 -916 5275 -876
rect 8056 -1258 8188 200
rect 9467 298 9501 314
rect 9467 106 9501 122
rect 9585 298 9619 314
rect 9585 106 9619 122
rect 9703 298 9737 314
rect 9703 106 9737 122
rect 9821 298 9855 314
rect 9821 106 9855 122
rect 9939 298 9973 314
rect 9939 106 9973 122
rect 10057 298 10091 314
rect 10057 106 10091 122
rect 10175 298 10209 314
rect 10175 106 10209 122
rect 10293 298 10327 348
rect 10293 106 10327 122
rect 10411 298 10445 314
rect 10411 106 10445 122
rect 10529 298 10563 348
rect 11480 358 11516 416
rect 11717 792 11751 808
rect 11599 400 11633 416
rect 11715 416 11717 463
rect 11715 358 11751 416
rect 11835 792 11869 808
rect 11835 400 11869 416
rect 11953 792 11987 808
rect 12071 792 12105 808
rect 11987 416 11989 462
rect 11953 358 11989 416
rect 12071 400 12105 416
rect 13261 792 13295 808
rect 13379 792 13413 808
rect 13261 400 13295 416
rect 13378 416 13379 463
rect 13497 792 13531 808
rect 13413 416 13414 463
rect 12576 358 13073 376
rect 11480 355 13073 358
rect 11480 321 13021 355
rect 13055 321 13073 355
rect 11480 318 13073 321
rect 13378 358 13414 416
rect 13615 792 13649 808
rect 13497 400 13531 416
rect 13613 416 13615 463
rect 13613 358 13649 416
rect 13733 792 13767 808
rect 13733 400 13767 416
rect 13851 792 13885 808
rect 13969 792 14003 808
rect 14490 800 14557 816
rect 13885 416 13887 462
rect 13851 358 13887 416
rect 13969 400 14003 416
rect 14474 387 14574 388
rect 14474 358 14630 387
rect 13378 318 14630 358
rect 11499 317 13073 318
rect 13397 317 14630 318
rect 11377 228 11444 244
rect 11377 194 11393 228
rect 11427 194 11444 228
rect 11377 178 11444 194
rect 10529 106 10563 122
rect 11208 161 11242 177
rect 11208 111 11242 127
rect 11554 76 11588 317
rect 12576 300 13073 317
rect 12024 228 12091 244
rect 12024 194 12041 228
rect 12075 194 12091 228
rect 12024 178 12091 194
rect 13275 228 13342 244
rect 13275 194 13291 228
rect 13325 194 13342 228
rect 13275 178 13342 194
rect 12331 160 12365 176
rect 11643 110 11659 144
rect 11693 110 11709 144
rect 11761 111 11777 145
rect 11811 111 11827 145
rect 12331 110 12365 126
rect 13106 161 13140 177
rect 13106 111 13140 127
rect 13452 76 13486 317
rect 14474 289 14630 317
rect 14474 288 14574 289
rect 13920 229 13987 245
rect 13920 195 13937 229
rect 13971 195 13987 229
rect 13920 179 13987 195
rect 14229 160 14263 176
rect 13541 110 13557 144
rect 13591 110 13607 144
rect 13659 111 13675 145
rect 13709 111 13725 145
rect 14229 110 14263 126
rect 10218 28 10234 62
rect 10268 28 10284 62
rect 11061 60 11095 76
rect 10100 -89 10116 -55
rect 10150 -89 10166 -55
rect 9704 -139 9738 -123
rect 9704 -531 9738 -515
rect 9822 -139 9856 -123
rect 9822 -531 9856 -515
rect 9940 -139 9974 -123
rect 10057 -139 10091 -123
rect 10057 -331 10091 -315
rect 10175 -139 10209 -123
rect 11061 -132 11095 -116
rect 11179 60 11213 76
rect 11179 -132 11213 -116
rect 11481 60 11515 76
rect 10175 -331 10209 -315
rect 11554 60 11633 76
rect 11554 30 11599 60
rect 11481 -383 11516 -316
rect 11599 -332 11633 -316
rect 11717 60 11751 76
rect 11717 -332 11751 -316
rect 11835 60 11869 76
rect 11953 60 11987 76
rect 12359 60 12393 76
rect 12359 -132 12393 -116
rect 12477 60 12511 76
rect 12477 -132 12511 -116
rect 12959 60 12993 76
rect 12959 -132 12993 -116
rect 13077 60 13111 76
rect 13077 -132 13111 -116
rect 13379 60 13413 76
rect 11835 -332 11869 -316
rect 11952 -383 11987 -316
rect 11481 -418 11987 -383
rect 13452 60 13531 76
rect 13452 30 13497 60
rect 13379 -383 13414 -316
rect 13497 -332 13531 -316
rect 13615 60 13649 76
rect 13615 -332 13649 -316
rect 13733 60 13767 76
rect 13851 60 13885 76
rect 14257 60 14291 76
rect 14257 -132 14291 -116
rect 14375 60 14409 76
rect 14375 -132 14409 -116
rect 13733 -332 13767 -316
rect 13850 -383 13885 -316
rect 13379 -418 13885 -383
rect 9940 -531 9974 -515
rect 10227 -465 10476 -422
rect 10227 -555 10274 -465
rect 10437 -555 10476 -465
rect 9747 -599 9763 -565
rect 9797 -599 9813 -565
rect 9865 -599 9881 -565
rect 9915 -599 9931 -565
rect 10227 -594 10476 -555
rect 11652 -625 11824 -578
rect 11652 -788 11691 -625
rect 11781 -788 11824 -625
rect 11652 -828 11824 -788
rect 15258 -1028 15421 908
rect 25679 871 25713 887
rect 25679 821 25713 837
rect 27769 850 27836 866
rect 19054 803 19088 819
rect 27769 816 27786 850
rect 27820 816 27836 850
rect 19054 753 19088 769
rect 21144 782 21211 798
rect 24642 792 24676 808
rect 21144 748 21161 782
rect 21195 748 21211 782
rect 18017 724 18051 740
rect 16516 646 16739 720
rect 16516 644 16596 646
rect 16516 495 16595 644
rect 16663 497 16739 646
rect 16662 495 16739 497
rect 16516 389 16739 495
rect 18135 724 18169 740
rect 18017 332 18051 348
rect 18134 348 18135 395
rect 18253 724 18287 740
rect 18169 348 18170 395
rect 16947 280 17217 314
rect 16121 230 16155 246
rect 16121 38 16155 54
rect 16239 230 16273 246
rect 16239 38 16273 54
rect 16357 230 16391 246
rect 16357 38 16391 54
rect 16475 230 16509 246
rect 16475 38 16509 54
rect 16593 230 16627 246
rect 16593 38 16627 54
rect 16711 230 16745 246
rect 16711 38 16745 54
rect 16829 230 16863 246
rect 16829 38 16863 54
rect 16947 230 16981 280
rect 16947 38 16981 54
rect 17065 230 17099 246
rect 17065 38 17099 54
rect 17183 230 17217 280
rect 18134 290 18170 348
rect 18371 724 18405 740
rect 18253 332 18287 348
rect 18369 348 18371 395
rect 18369 290 18405 348
rect 18489 724 18523 740
rect 18489 332 18523 348
rect 18607 724 18641 740
rect 18725 724 18759 740
rect 18641 348 18643 394
rect 18607 290 18643 348
rect 18725 332 18759 348
rect 19915 724 19949 740
rect 20033 724 20067 740
rect 19915 332 19949 348
rect 20032 348 20033 395
rect 20151 724 20185 740
rect 20067 348 20068 395
rect 19230 290 19727 308
rect 18134 287 19727 290
rect 18134 253 19675 287
rect 19709 253 19727 287
rect 18134 250 19727 253
rect 20032 290 20068 348
rect 20269 724 20303 740
rect 20151 332 20185 348
rect 20267 348 20269 395
rect 20267 290 20303 348
rect 20387 724 20421 740
rect 20387 332 20421 348
rect 20505 724 20539 740
rect 20623 724 20657 740
rect 21144 732 21211 748
rect 20539 348 20541 394
rect 20505 290 20541 348
rect 23141 712 23364 788
rect 23141 563 23220 712
rect 23287 707 23364 712
rect 23141 558 23221 563
rect 23288 558 23364 707
rect 23141 457 23364 558
rect 24760 792 24794 808
rect 24642 400 24676 416
rect 24759 416 24760 463
rect 24878 792 24912 808
rect 24794 416 24795 463
rect 20623 332 20657 348
rect 23572 348 23842 382
rect 21738 321 21847 327
rect 21214 320 21847 321
rect 21128 318 21847 320
rect 21128 290 21745 318
rect 20032 250 21745 290
rect 18153 249 19727 250
rect 20051 249 21745 250
rect 18031 160 18098 176
rect 18031 126 18047 160
rect 18081 126 18098 160
rect 18031 110 18098 126
rect 17183 38 17217 54
rect 17862 93 17896 109
rect 17862 43 17896 59
rect 18208 8 18242 249
rect 19230 232 19727 249
rect 18678 160 18745 176
rect 18678 126 18695 160
rect 18729 126 18745 160
rect 18678 110 18745 126
rect 19929 160 19996 176
rect 19929 126 19945 160
rect 19979 126 19996 160
rect 19929 110 19996 126
rect 18985 92 19019 108
rect 18297 42 18313 76
rect 18347 42 18363 76
rect 18415 43 18431 77
rect 18465 43 18481 77
rect 18985 42 19019 58
rect 19760 93 19794 109
rect 19760 43 19794 59
rect 20106 8 20140 249
rect 21128 220 21745 249
rect 21214 219 21745 220
rect 21738 218 21745 219
rect 21841 218 21847 318
rect 21738 212 21847 218
rect 22746 298 22780 314
rect 20574 161 20641 177
rect 20574 127 20591 161
rect 20625 127 20641 161
rect 20574 111 20641 127
rect 20883 92 20917 108
rect 22746 106 22780 122
rect 22864 298 22898 314
rect 22864 106 22898 122
rect 22982 298 23016 314
rect 22982 106 23016 122
rect 23100 298 23134 314
rect 23100 106 23134 122
rect 23218 298 23252 314
rect 23218 106 23252 122
rect 23336 298 23370 314
rect 23336 106 23370 122
rect 23454 298 23488 314
rect 23454 106 23488 122
rect 23572 298 23606 348
rect 23572 106 23606 122
rect 23690 298 23724 314
rect 23690 106 23724 122
rect 23808 298 23842 348
rect 24759 358 24795 416
rect 24996 792 25030 808
rect 24878 400 24912 416
rect 24994 416 24996 463
rect 24994 358 25030 416
rect 25114 792 25148 808
rect 25114 400 25148 416
rect 25232 792 25266 808
rect 25350 792 25384 808
rect 25266 416 25268 462
rect 25232 358 25268 416
rect 25350 400 25384 416
rect 26540 792 26574 808
rect 26658 792 26692 808
rect 26540 400 26574 416
rect 26657 416 26658 463
rect 26776 792 26810 808
rect 26692 416 26693 463
rect 25855 358 26352 376
rect 24759 355 26352 358
rect 24759 321 26300 355
rect 26334 321 26352 355
rect 24759 318 26352 321
rect 26657 358 26693 416
rect 26894 792 26928 808
rect 26776 400 26810 416
rect 26892 416 26894 463
rect 26892 358 26928 416
rect 27012 792 27046 808
rect 27012 400 27046 416
rect 27130 792 27164 808
rect 27248 792 27282 808
rect 27769 800 27836 816
rect 27164 416 27166 462
rect 27130 358 27166 416
rect 27248 400 27282 416
rect 27753 387 27853 388
rect 27753 358 27909 387
rect 26657 318 27909 358
rect 24778 317 26352 318
rect 26676 317 27909 318
rect 24656 228 24723 244
rect 24656 194 24672 228
rect 24706 194 24723 228
rect 24656 178 24723 194
rect 23808 106 23842 122
rect 24487 161 24521 177
rect 24487 111 24521 127
rect 20195 42 20211 76
rect 20245 42 20261 76
rect 20313 43 20329 77
rect 20363 43 20379 77
rect 24833 76 24867 317
rect 25855 300 26352 317
rect 25303 228 25370 244
rect 25303 194 25320 228
rect 25354 194 25370 228
rect 25303 178 25370 194
rect 26554 228 26621 244
rect 26554 194 26570 228
rect 26604 194 26621 228
rect 26554 178 26621 194
rect 25610 160 25644 176
rect 24922 110 24938 144
rect 24972 110 24988 144
rect 25040 111 25056 145
rect 25090 111 25106 145
rect 25610 110 25644 126
rect 26385 161 26419 177
rect 26385 111 26419 127
rect 26731 76 26765 317
rect 27753 289 27909 317
rect 27753 288 27853 289
rect 27199 229 27266 245
rect 27199 195 27216 229
rect 27250 195 27266 229
rect 27199 179 27266 195
rect 27508 160 27542 176
rect 26820 110 26836 144
rect 26870 110 26886 144
rect 26938 111 26954 145
rect 26988 111 27004 145
rect 27508 110 27542 126
rect 28823 120 28991 136
rect 20883 42 20917 58
rect 23497 28 23513 62
rect 23547 28 23563 62
rect 24340 60 24374 76
rect 16872 -40 16888 -6
rect 16922 -40 16938 -6
rect 17715 -8 17749 8
rect 16754 -157 16770 -123
rect 16804 -157 16820 -123
rect 16358 -207 16392 -191
rect 16358 -599 16392 -583
rect 16476 -207 16510 -191
rect 16476 -599 16510 -583
rect 16594 -207 16628 -191
rect 16711 -207 16745 -191
rect 16711 -399 16745 -383
rect 16829 -207 16863 -191
rect 17715 -200 17749 -184
rect 17833 -8 17867 8
rect 17833 -200 17867 -184
rect 18135 -8 18169 8
rect 16829 -399 16863 -383
rect 18208 -8 18287 8
rect 18208 -38 18253 -8
rect 18135 -451 18170 -384
rect 18253 -400 18287 -384
rect 18371 -8 18405 8
rect 18371 -400 18405 -384
rect 18489 -8 18523 8
rect 18607 -8 18641 8
rect 19013 -8 19047 8
rect 19013 -200 19047 -184
rect 19131 -8 19165 8
rect 19131 -200 19165 -184
rect 19613 -8 19647 8
rect 19613 -200 19647 -184
rect 19731 -8 19765 8
rect 19731 -200 19765 -184
rect 20033 -8 20067 8
rect 18489 -400 18523 -384
rect 18606 -451 18641 -384
rect 18135 -486 18641 -451
rect 20106 -8 20185 8
rect 20106 -38 20151 -8
rect 20033 -451 20068 -384
rect 20151 -400 20185 -384
rect 20269 -8 20303 8
rect 20269 -400 20303 -384
rect 20387 -8 20421 8
rect 20505 -8 20539 8
rect 20911 -8 20945 8
rect 20911 -200 20945 -184
rect 21029 -8 21063 8
rect 23379 -89 23395 -55
rect 23429 -89 23445 -55
rect 21029 -200 21063 -184
rect 22983 -139 23017 -123
rect 20387 -400 20421 -384
rect 20504 -451 20539 -384
rect 20033 -486 20539 -451
rect 16594 -599 16628 -583
rect 16881 -533 17130 -490
rect 22983 -531 23017 -515
rect 23101 -139 23135 -123
rect 23101 -531 23135 -515
rect 23219 -139 23253 -123
rect 23336 -139 23370 -123
rect 23336 -331 23370 -315
rect 23454 -139 23488 -123
rect 24340 -132 24374 -116
rect 24458 60 24492 76
rect 24458 -132 24492 -116
rect 24760 60 24794 76
rect 23454 -331 23488 -315
rect 24833 60 24912 76
rect 24833 30 24878 60
rect 24760 -383 24795 -316
rect 24878 -332 24912 -316
rect 24996 60 25030 76
rect 24996 -332 25030 -316
rect 25114 60 25148 76
rect 25232 60 25266 76
rect 25638 60 25672 76
rect 25638 -132 25672 -116
rect 25756 60 25790 76
rect 25756 -132 25790 -116
rect 26238 60 26272 76
rect 26238 -132 26272 -116
rect 26356 60 26390 76
rect 26356 -132 26390 -116
rect 26658 60 26692 76
rect 25114 -332 25148 -316
rect 25231 -383 25266 -316
rect 24760 -418 25266 -383
rect 26731 60 26810 76
rect 26731 30 26776 60
rect 26658 -383 26693 -316
rect 26776 -332 26810 -316
rect 26894 60 26928 76
rect 26894 -332 26928 -316
rect 27012 60 27046 76
rect 27130 60 27164 76
rect 27536 60 27570 76
rect 27536 -132 27570 -116
rect 27654 60 27688 76
rect 28823 50 28839 120
rect 28975 50 28991 120
rect 28823 34 28991 50
rect 29360 -70 29630 -36
rect 27654 -132 27688 -116
rect 28534 -120 28568 -104
rect 28534 -312 28568 -296
rect 28652 -120 28686 -104
rect 28652 -312 28686 -296
rect 28770 -120 28804 -104
rect 28770 -312 28804 -296
rect 28888 -120 28922 -104
rect 28888 -312 28922 -296
rect 29006 -120 29040 -104
rect 29006 -312 29040 -296
rect 29124 -120 29158 -104
rect 29124 -312 29158 -296
rect 29242 -120 29276 -104
rect 29242 -312 29276 -296
rect 29360 -120 29394 -70
rect 29360 -312 29394 -296
rect 29478 -120 29512 -104
rect 29478 -312 29512 -296
rect 29596 -120 29630 -70
rect 29596 -312 29630 -296
rect 27012 -332 27046 -316
rect 27129 -383 27164 -316
rect 26658 -418 27164 -383
rect 29285 -390 29301 -356
rect 29335 -390 29351 -356
rect 23219 -531 23253 -515
rect 23506 -465 23755 -422
rect 16881 -623 16928 -533
rect 17091 -623 17130 -533
rect 23506 -555 23553 -465
rect 23716 -555 23755 -465
rect 29167 -507 29183 -473
rect 29217 -507 29233 -473
rect 23026 -599 23042 -565
rect 23076 -599 23092 -565
rect 23144 -599 23160 -565
rect 23194 -599 23210 -565
rect 23506 -594 23755 -555
rect 28771 -557 28805 -541
rect 16401 -667 16417 -633
rect 16451 -667 16467 -633
rect 16519 -667 16535 -633
rect 16569 -667 16585 -633
rect 16881 -662 17130 -623
rect 24931 -625 25103 -578
rect 18306 -693 18478 -646
rect 18306 -856 18345 -693
rect 18435 -856 18478 -693
rect 24931 -788 24970 -625
rect 25060 -788 25103 -625
rect 24931 -828 25103 -788
rect 18306 -896 18478 -856
rect 28771 -949 28805 -933
rect 28889 -557 28923 -541
rect 28889 -949 28923 -933
rect 29007 -557 29041 -541
rect 29124 -557 29158 -541
rect 29124 -749 29158 -733
rect 29242 -557 29276 -541
rect 29242 -749 29276 -733
rect 29007 -949 29041 -933
rect 15258 -1096 15302 -1028
rect 15372 -1096 15421 -1028
rect 15258 -1112 15421 -1096
rect 21254 -1003 22526 -976
rect 21254 -1102 21285 -1003
rect 21391 -1102 22394 -1003
rect 22500 -1102 22526 -1003
rect 28814 -1017 28830 -983
rect 28864 -1017 28880 -983
rect 28932 -1017 28948 -983
rect 28982 -1017 28998 -983
rect 21254 -1129 22526 -1102
rect 29047 -1088 29215 -1070
rect 29047 -1144 29063 -1088
rect 29197 -1144 29215 -1088
rect 29047 -1160 29215 -1144
rect 15276 -1256 27548 -1255
rect 30076 -1256 30195 4541
rect 30892 4586 30926 4602
rect 30774 4194 30808 4210
rect 30891 4210 30892 4257
rect 31010 4586 31044 4602
rect 30926 4210 30927 4257
rect 30891 4152 30927 4210
rect 31128 4586 31162 4602
rect 31010 4194 31044 4210
rect 31126 4210 31128 4257
rect 31126 4152 31162 4210
rect 31246 4586 31280 4602
rect 31246 4194 31280 4210
rect 31364 4586 31398 4602
rect 31482 4586 31516 4602
rect 31398 4210 31400 4256
rect 31364 4152 31400 4210
rect 31644 4381 31714 4385
rect 31644 4290 31648 4381
rect 31710 4290 31714 4381
rect 31644 4285 31714 4290
rect 31482 4194 31516 4210
rect 31659 4152 31700 4285
rect 32377 4247 32411 4263
rect 32495 4639 32529 4655
rect 32495 4247 32529 4263
rect 32613 4639 32647 4655
rect 32730 4639 32764 4655
rect 32730 4447 32764 4463
rect 32848 4639 32882 4655
rect 32848 4447 32882 4463
rect 32613 4247 32647 4263
rect 32420 4179 32436 4213
rect 32470 4179 32486 4213
rect 32538 4179 32554 4213
rect 32588 4179 32604 4213
rect 30891 4112 31700 4152
rect 30910 4111 31700 4112
rect 30788 4022 30855 4038
rect 30788 3988 30804 4022
rect 30838 3988 30855 4022
rect 30788 3972 30855 3988
rect 30619 3955 30653 3971
rect 30619 3905 30653 3921
rect 30965 3870 30999 4111
rect 32653 4108 32821 4126
rect 32653 4052 32669 4108
rect 32803 4052 32821 4108
rect 31435 4022 31502 4038
rect 32653 4036 32821 4052
rect 31435 3988 31452 4022
rect 31486 3988 31502 4022
rect 31435 3972 31502 3988
rect 31742 3954 31776 3970
rect 31054 3904 31070 3938
rect 31104 3904 31120 3938
rect 31172 3905 31188 3939
rect 31222 3905 31238 3939
rect 31742 3904 31776 3920
rect 30472 3854 30506 3870
rect 30472 3662 30506 3678
rect 30590 3854 30624 3870
rect 30590 3662 30624 3678
rect 30892 3854 30926 3870
rect 30965 3854 31044 3870
rect 30965 3824 31010 3854
rect 30892 3411 30927 3478
rect 31010 3462 31044 3478
rect 31128 3854 31162 3870
rect 31128 3462 31162 3478
rect 31246 3854 31280 3870
rect 31364 3854 31398 3870
rect 31770 3854 31804 3870
rect 31770 3662 31804 3678
rect 31888 3854 31922 3870
rect 31888 3662 31922 3678
rect 31246 3462 31280 3478
rect 31363 3411 31398 3478
rect 30892 3376 31398 3411
rect 31039 3307 31281 3319
rect 31039 3205 31086 3307
rect 31221 3205 31281 3307
rect 31039 3188 31281 3205
rect 30972 1726 31416 1732
rect 30972 1526 30983 1726
rect 31404 1526 31416 1726
rect 30972 1520 31416 1526
rect 31187 1241 31457 1276
rect 30833 1188 30867 1204
rect 30349 1042 30619 1077
rect 30349 988 30383 1042
rect 30349 796 30383 812
rect 30467 988 30501 1004
rect 30467 796 30501 812
rect 30585 988 30619 1042
rect 30585 796 30619 812
rect 30703 988 30737 1004
rect 30703 796 30737 812
rect 30833 796 30867 812
rect 30951 1188 30985 1204
rect 30951 796 30985 812
rect 31069 1188 31103 1204
rect 31069 796 31103 812
rect 31187 1188 31221 1241
rect 31187 796 31221 812
rect 31305 1188 31339 1204
rect 31305 796 31339 812
rect 31423 1188 31457 1241
rect 32431 1225 32599 1241
rect 31423 796 31457 812
rect 31541 1188 31575 1204
rect 32431 1155 32447 1225
rect 32583 1155 32599 1225
rect 32431 1139 32599 1155
rect 32968 1035 33238 1069
rect 31541 796 31575 812
rect 31670 988 31704 1004
rect 31670 796 31704 812
rect 31788 988 31822 1004
rect 31788 796 31822 812
rect 31906 988 31940 1004
rect 31906 796 31940 812
rect 32024 988 32058 1004
rect 32024 796 32058 812
rect 32142 985 32176 1001
rect 32142 793 32176 809
rect 32260 985 32294 1001
rect 32260 793 32294 809
rect 32378 985 32412 1001
rect 32378 793 32412 809
rect 32496 985 32530 1001
rect 32496 793 32530 809
rect 32614 985 32648 1001
rect 32614 793 32648 809
rect 32732 985 32766 1001
rect 32732 793 32766 809
rect 32850 985 32884 1001
rect 32850 793 32884 809
rect 32968 985 33002 1035
rect 32968 793 33002 809
rect 33086 985 33120 1001
rect 33086 793 33120 809
rect 33204 985 33238 1035
rect 33204 793 33238 809
rect 32893 715 32909 749
rect 32943 715 32959 749
rect 32001 630 32035 646
rect 32775 598 32791 632
rect 32825 598 32841 632
rect 32001 580 32035 596
rect 32379 548 32413 564
rect 30595 511 30651 528
rect 30595 477 30601 511
rect 30635 477 30651 511
rect 30595 460 30651 477
rect 30776 495 30810 511
rect 30894 495 30928 511
rect 30776 103 30810 119
rect 30893 119 30894 166
rect 31012 495 31046 511
rect 30928 119 30929 166
rect 30893 61 30929 119
rect 31130 495 31164 511
rect 31012 103 31046 119
rect 31128 119 31130 166
rect 31128 61 31164 119
rect 31248 495 31282 511
rect 31248 103 31282 119
rect 31366 495 31400 511
rect 31484 495 31518 511
rect 31400 119 31402 165
rect 31366 61 31402 119
rect 31646 290 31716 294
rect 31646 199 31650 290
rect 31712 199 31716 290
rect 31646 194 31716 199
rect 31484 103 31518 119
rect 31661 61 31702 194
rect 32379 156 32413 172
rect 32497 548 32531 564
rect 32497 156 32531 172
rect 32615 548 32649 564
rect 32732 548 32766 564
rect 32732 356 32766 372
rect 32850 548 32884 564
rect 33082 538 33238 544
rect 33082 467 33097 538
rect 33224 467 33238 538
rect 33082 457 33238 467
rect 32850 356 32884 372
rect 32615 156 32649 172
rect 32422 88 32438 122
rect 32472 88 32488 122
rect 32540 88 32556 122
rect 32590 88 32606 122
rect 30893 21 31702 61
rect 30912 20 31702 21
rect 30790 -69 30857 -53
rect 30790 -103 30806 -69
rect 30840 -103 30857 -69
rect 30790 -119 30857 -103
rect 30621 -136 30655 -120
rect 30621 -186 30655 -170
rect 30967 -221 31001 20
rect 32655 17 32823 35
rect 32655 -39 32671 17
rect 32805 -39 32823 17
rect 31437 -69 31504 -53
rect 32655 -55 32823 -39
rect 31437 -103 31454 -69
rect 31488 -103 31504 -69
rect 31437 -119 31504 -103
rect 31744 -137 31778 -121
rect 31056 -187 31072 -153
rect 31106 -187 31122 -153
rect 31174 -186 31190 -152
rect 31224 -186 31240 -152
rect 31744 -187 31778 -171
rect 30474 -237 30508 -221
rect 30474 -429 30508 -413
rect 30592 -237 30626 -221
rect 30592 -429 30626 -413
rect 30894 -237 30928 -221
rect 30967 -237 31046 -221
rect 30967 -267 31012 -237
rect 30894 -680 30929 -613
rect 31012 -629 31046 -613
rect 31130 -237 31164 -221
rect 31130 -629 31164 -613
rect 31248 -237 31282 -221
rect 31366 -237 31400 -221
rect 31772 -237 31806 -221
rect 31772 -429 31806 -413
rect 31890 -237 31924 -221
rect 31890 -429 31924 -413
rect 31248 -629 31282 -613
rect 31365 -680 31400 -613
rect 30894 -715 31400 -680
rect 31041 -784 31283 -772
rect 31041 -886 31088 -784
rect 31223 -886 31283 -784
rect 31041 -903 31283 -886
rect 15276 -1257 30195 -1256
rect 12811 -1258 30195 -1257
rect 8056 -1367 30195 -1258
rect 8056 -1369 18483 -1367
rect 27534 -1368 30195 -1367
rect 8056 -1370 15060 -1369
rect 2011 -1512 30036 -1510
rect 33145 -1512 33238 457
rect 2011 -1639 33238 -1512
rect 13402 -1641 33238 -1639
rect 30972 -1769 31416 -1763
rect 3296 -1901 3519 -1826
rect 3296 -2050 3372 -1901
rect 3439 -1902 3519 -1901
rect 3296 -2051 3375 -2050
rect 3442 -2051 3519 -1902
rect 3296 -2157 3519 -2051
rect 5778 -1846 6001 -1772
rect 5778 -1995 5852 -1846
rect 5919 -1848 6001 -1846
rect 5778 -1997 5857 -1995
rect 5924 -1997 6001 -1848
rect 5111 -2068 5145 -2052
rect 5111 -2118 5145 -2102
rect 5778 -2103 6001 -1997
rect 6925 -1848 7148 -1772
rect 6925 -1997 7004 -1848
rect 7071 -1849 7148 -1848
rect 6925 -1998 7008 -1997
rect 7075 -1998 7148 -1849
rect 6241 -2062 6275 -2046
rect 6241 -2112 6275 -2096
rect 6925 -2103 7148 -1998
rect 9847 -1903 10070 -1828
rect 9847 -1904 9927 -1903
rect 9847 -2053 9926 -1904
rect 9994 -2052 10070 -1903
rect 9993 -2053 10070 -2052
rect 9847 -2159 10070 -2053
rect 12329 -1850 12552 -1774
rect 12329 -1999 12408 -1850
rect 12475 -1999 12552 -1850
rect 11662 -2070 11696 -2054
rect 11662 -2120 11696 -2104
rect 12329 -2105 12552 -1999
rect 13476 -1850 13699 -1774
rect 13476 -1999 13555 -1850
rect 13623 -1999 13699 -1850
rect 12792 -2064 12826 -2048
rect 12792 -2114 12826 -2098
rect 13476 -2105 13699 -1999
rect 15258 -1845 15420 -1829
rect 15258 -1913 15301 -1845
rect 15371 -1913 15420 -1845
rect 5111 -2186 5145 -2170
rect 3727 -2266 3997 -2232
rect 5111 -2236 5145 -2220
rect 6241 -2182 6275 -2166
rect 2901 -2316 2935 -2300
rect 2901 -2508 2935 -2492
rect 3019 -2316 3053 -2300
rect 3019 -2508 3053 -2492
rect 3137 -2316 3171 -2300
rect 3137 -2508 3171 -2492
rect 3255 -2316 3289 -2300
rect 3255 -2508 3289 -2492
rect 3373 -2316 3407 -2300
rect 3373 -2508 3407 -2492
rect 3491 -2316 3525 -2300
rect 3491 -2508 3525 -2492
rect 3609 -2316 3643 -2300
rect 3609 -2508 3643 -2492
rect 3727 -2316 3761 -2266
rect 3727 -2508 3761 -2492
rect 3845 -2316 3879 -2300
rect 3845 -2508 3879 -2492
rect 3963 -2316 3997 -2266
rect 3963 -2508 3997 -2492
rect 5226 -2244 5260 -2228
rect 3652 -2586 3668 -2552
rect 3702 -2586 3718 -2552
rect 5226 -2636 5260 -2620
rect 5344 -2244 5378 -2228
rect 5344 -2636 5378 -2620
rect 5462 -2244 5496 -2228
rect 5462 -2636 5496 -2620
rect 5580 -2244 5614 -2228
rect 5580 -2636 5614 -2620
rect 5698 -2244 5732 -2228
rect 5698 -2636 5732 -2620
rect 5816 -2244 5850 -2228
rect 5816 -2636 5850 -2620
rect 5934 -2244 5968 -2228
rect 6241 -2232 6275 -2216
rect 11662 -2188 11696 -2172
rect 5934 -2636 5968 -2620
rect 6368 -2240 6402 -2224
rect 6368 -2632 6402 -2616
rect 6486 -2240 6520 -2224
rect 6486 -2632 6520 -2616
rect 6604 -2240 6638 -2224
rect 6604 -2632 6638 -2616
rect 6722 -2240 6756 -2224
rect 6722 -2632 6756 -2616
rect 6840 -2240 6874 -2224
rect 6840 -2632 6874 -2616
rect 6958 -2240 6992 -2224
rect 6958 -2632 6992 -2616
rect 7076 -2240 7110 -2224
rect 10278 -2268 10548 -2234
rect 11662 -2238 11696 -2222
rect 12792 -2184 12826 -2168
rect 9452 -2318 9486 -2302
rect 9452 -2510 9486 -2494
rect 9570 -2318 9604 -2302
rect 9570 -2510 9604 -2494
rect 9688 -2318 9722 -2302
rect 9688 -2510 9722 -2494
rect 9806 -2318 9840 -2302
rect 9806 -2510 9840 -2494
rect 9924 -2318 9958 -2302
rect 9924 -2510 9958 -2494
rect 10042 -2318 10076 -2302
rect 10042 -2510 10076 -2494
rect 10160 -2318 10194 -2302
rect 10160 -2510 10194 -2494
rect 10278 -2318 10312 -2268
rect 10278 -2510 10312 -2494
rect 10396 -2318 10430 -2302
rect 10396 -2510 10430 -2494
rect 10514 -2318 10548 -2268
rect 10514 -2510 10548 -2494
rect 11777 -2246 11811 -2230
rect 10203 -2588 10219 -2554
rect 10253 -2588 10269 -2554
rect 7076 -2632 7110 -2616
rect 11777 -2638 11811 -2622
rect 11895 -2246 11929 -2230
rect 11895 -2638 11929 -2622
rect 12013 -2246 12047 -2230
rect 12013 -2638 12047 -2622
rect 12131 -2246 12165 -2230
rect 12131 -2638 12165 -2622
rect 12249 -2246 12283 -2230
rect 12249 -2638 12283 -2622
rect 12367 -2246 12401 -2230
rect 12367 -2638 12401 -2622
rect 12485 -2246 12519 -2230
rect 12792 -2234 12826 -2218
rect 12485 -2638 12519 -2622
rect 12919 -2242 12953 -2226
rect 12919 -2634 12953 -2618
rect 13037 -2242 13071 -2226
rect 13037 -2634 13071 -2618
rect 13155 -2242 13189 -2226
rect 13155 -2634 13189 -2618
rect 13273 -2242 13307 -2226
rect 13273 -2634 13307 -2618
rect 13391 -2242 13425 -2226
rect 13391 -2634 13425 -2618
rect 13509 -2242 13543 -2226
rect 13509 -2634 13543 -2618
rect 13627 -2242 13661 -2226
rect 15258 -2431 15420 -1913
rect 16502 -1903 16725 -1827
rect 16502 -1906 16581 -1903
rect 16502 -2055 16578 -1906
rect 16648 -2052 16725 -1903
rect 16645 -2055 16725 -2052
rect 18984 -1846 19207 -1773
rect 18984 -1998 19063 -1846
rect 19130 -1998 19207 -1846
rect 16502 -2158 16725 -2055
rect 18317 -2069 18351 -2053
rect 18317 -2119 18351 -2103
rect 18984 -2104 19207 -1998
rect 20131 -1849 20354 -1773
rect 20131 -1998 20210 -1849
rect 20279 -1998 20354 -1849
rect 19447 -2063 19481 -2047
rect 19447 -2113 19481 -2097
rect 20131 -2104 20354 -1998
rect 23124 -1901 23347 -1826
rect 23124 -2050 23202 -1901
rect 23269 -1902 23347 -1901
rect 23124 -2051 23203 -2050
rect 23270 -2051 23347 -1902
rect 23124 -2157 23347 -2051
rect 25606 -1848 25829 -1772
rect 25606 -1853 25685 -1848
rect 25606 -2002 25681 -1853
rect 25752 -1997 25829 -1848
rect 25748 -2002 25829 -1997
rect 24939 -2068 24973 -2052
rect 24939 -2118 24973 -2102
rect 25606 -2103 25829 -2002
rect 26753 -1847 26976 -1772
rect 26753 -1996 26829 -1847
rect 26896 -1848 26976 -1847
rect 26753 -1997 26832 -1996
rect 26899 -1997 26976 -1848
rect 28894 -1800 29062 -1784
rect 28894 -1870 28910 -1800
rect 29046 -1870 29062 -1800
rect 28894 -1886 29062 -1870
rect 26069 -2062 26103 -2046
rect 26069 -2112 26103 -2096
rect 26753 -2103 26976 -1997
rect 29431 -1990 29701 -1956
rect 30972 -1969 30983 -1769
rect 31404 -1969 31416 -1769
rect 30972 -1975 31416 -1969
rect 28605 -2040 28639 -2024
rect 18317 -2187 18351 -2171
rect 16933 -2267 17203 -2233
rect 18317 -2237 18351 -2221
rect 19447 -2183 19481 -2167
rect 16107 -2317 16141 -2301
rect 13627 -2634 13661 -2618
rect 3534 -2703 3550 -2669
rect 3584 -2703 3600 -2669
rect 10085 -2705 10101 -2671
rect 10135 -2705 10151 -2671
rect 3138 -2753 3172 -2737
rect 3138 -3145 3172 -3129
rect 3256 -2753 3290 -2737
rect 3256 -3145 3290 -3129
rect 3374 -2753 3408 -2737
rect 3491 -2753 3525 -2737
rect 3491 -2945 3525 -2929
rect 3609 -2753 3643 -2737
rect 3609 -2945 3643 -2929
rect 9689 -2755 9723 -2739
rect 5415 -2976 5431 -2942
rect 5465 -2976 5481 -2942
rect 6557 -2972 6573 -2938
rect 6607 -2972 6623 -2938
rect 5136 -3027 5170 -3011
rect 3374 -3145 3408 -3129
rect 3661 -3079 3910 -3036
rect 3661 -3169 3708 -3079
rect 3871 -3169 3910 -3079
rect 3181 -3213 3197 -3179
rect 3231 -3213 3247 -3179
rect 3299 -3213 3315 -3179
rect 3349 -3213 3365 -3179
rect 3661 -3208 3910 -3169
rect 5136 -3219 5170 -3203
rect 5254 -3027 5288 -3011
rect 5254 -3219 5288 -3203
rect 5372 -3027 5406 -3011
rect 5372 -3219 5406 -3203
rect 5490 -3027 5524 -3011
rect 5490 -3219 5524 -3203
rect 5655 -3027 5689 -3011
rect 5655 -3219 5689 -3203
rect 5773 -3027 5807 -3011
rect 5773 -3219 5807 -3203
rect 5891 -3027 5925 -3011
rect 5891 -3219 5925 -3203
rect 6009 -3027 6043 -3011
rect 6009 -3219 6043 -3203
rect 6278 -3023 6312 -3007
rect 6278 -3215 6312 -3199
rect 6396 -3023 6430 -3007
rect 6396 -3215 6430 -3199
rect 6514 -3023 6548 -3007
rect 6514 -3215 6548 -3199
rect 6632 -3023 6666 -3007
rect 6632 -3215 6666 -3199
rect 6797 -3023 6831 -3007
rect 6797 -3215 6831 -3199
rect 6915 -3023 6949 -3007
rect 6915 -3215 6949 -3199
rect 7033 -3023 7067 -3007
rect 7033 -3215 7067 -3199
rect 7151 -3023 7185 -3007
rect 9689 -3147 9723 -3131
rect 9807 -2755 9841 -2739
rect 9807 -3147 9841 -3131
rect 9925 -2755 9959 -2739
rect 10042 -2755 10076 -2739
rect 10042 -2947 10076 -2931
rect 10160 -2755 10194 -2739
rect 10160 -2947 10194 -2931
rect 11966 -2978 11982 -2944
rect 12016 -2978 12032 -2944
rect 13108 -2974 13124 -2940
rect 13158 -2974 13174 -2940
rect 11687 -3029 11721 -3013
rect 9925 -3147 9959 -3131
rect 10212 -3081 10461 -3038
rect 10212 -3171 10259 -3081
rect 10422 -3171 10461 -3081
rect 7151 -3215 7185 -3199
rect 9732 -3215 9748 -3181
rect 9782 -3215 9798 -3181
rect 9850 -3215 9866 -3181
rect 9900 -3215 9916 -3181
rect 10212 -3210 10461 -3171
rect 11687 -3221 11721 -3205
rect 11805 -3029 11839 -3013
rect 11805 -3221 11839 -3205
rect 11923 -3029 11957 -3013
rect 11923 -3221 11957 -3205
rect 12041 -3029 12075 -3013
rect 12041 -3221 12075 -3205
rect 12206 -3029 12240 -3013
rect 12206 -3221 12240 -3205
rect 12324 -3029 12358 -3013
rect 12324 -3221 12358 -3205
rect 12442 -3029 12476 -3013
rect 12442 -3221 12476 -3205
rect 12560 -3029 12594 -3013
rect 12560 -3221 12594 -3205
rect 12829 -3025 12863 -3009
rect 12829 -3217 12863 -3201
rect 12947 -3025 12981 -3009
rect 12947 -3217 12981 -3201
rect 13065 -3025 13099 -3009
rect 13065 -3217 13099 -3201
rect 13183 -3025 13217 -3009
rect 13183 -3217 13217 -3201
rect 13348 -3025 13382 -3009
rect 13348 -3217 13382 -3201
rect 13466 -3025 13500 -3009
rect 13466 -3217 13500 -3201
rect 13584 -3025 13618 -3009
rect 13584 -3217 13618 -3201
rect 13702 -3025 13736 -3009
rect 13702 -3217 13736 -3201
rect 5151 -3450 5323 -3403
rect 3310 -3552 3533 -3476
rect 3310 -3701 3389 -3552
rect 3456 -3554 3533 -3552
rect 3310 -3703 3393 -3701
rect 3460 -3703 3533 -3554
rect 5151 -3613 5190 -3450
rect 5280 -3613 5323 -3450
rect 5151 -3652 5323 -3613
rect 6293 -3452 6465 -3405
rect 6293 -3615 6332 -3452
rect 6422 -3615 6465 -3452
rect 11702 -3452 11874 -3405
rect 6293 -3654 6465 -3615
rect 9861 -3547 10084 -3478
rect 3310 -3807 3533 -3703
rect 9861 -3696 9938 -3547
rect 10005 -3554 10084 -3547
rect 9861 -3703 9940 -3696
rect 10007 -3703 10084 -3554
rect 11702 -3615 11741 -3452
rect 11831 -3615 11874 -3452
rect 11702 -3654 11874 -3615
rect 12844 -3454 13016 -3407
rect 12844 -3617 12883 -3454
rect 12973 -3617 13016 -3454
rect 12844 -3621 12891 -3617
rect 12958 -3621 13016 -3617
rect 12844 -3656 13016 -3621
rect 9861 -3809 10084 -3703
rect 3741 -3916 4011 -3882
rect 2915 -3966 2949 -3950
rect 2915 -4158 2949 -4142
rect 3033 -3966 3067 -3950
rect 3033 -4158 3067 -4142
rect 3151 -3966 3185 -3950
rect 3151 -4158 3185 -4142
rect 3269 -3966 3303 -3950
rect 3269 -4158 3303 -4142
rect 3387 -3966 3421 -3950
rect 3387 -4158 3421 -4142
rect 3505 -3966 3539 -3950
rect 3505 -4158 3539 -4142
rect 3623 -3966 3657 -3950
rect 3623 -4158 3657 -4142
rect 3741 -3966 3775 -3916
rect 3741 -4158 3775 -4142
rect 3859 -3966 3893 -3950
rect 3859 -4158 3893 -4142
rect 3977 -3966 4011 -3916
rect 3977 -4158 4011 -4142
rect 7021 -3895 7246 -3819
rect 7021 -4044 7099 -3895
rect 7167 -4044 7246 -3895
rect 10292 -3918 10562 -3884
rect 7021 -4150 7246 -4044
rect 9466 -3968 9500 -3952
rect 9466 -4160 9500 -4144
rect 9584 -3968 9618 -3952
rect 9584 -4160 9618 -4144
rect 9702 -3968 9736 -3952
rect 9702 -4160 9736 -4144
rect 9820 -3968 9854 -3952
rect 9820 -4160 9854 -4144
rect 9938 -3968 9972 -3952
rect 9938 -4160 9972 -4144
rect 10056 -3968 10090 -3952
rect 10056 -4160 10090 -4144
rect 10174 -3968 10208 -3952
rect 10174 -4160 10208 -4144
rect 10292 -3968 10326 -3918
rect 10292 -4160 10326 -4144
rect 10410 -3968 10444 -3952
rect 10410 -4160 10444 -4144
rect 10528 -3968 10562 -3918
rect 10528 -4160 10562 -4144
rect 13572 -3896 13797 -3821
rect 13572 -3897 13655 -3896
rect 13572 -4046 13651 -3897
rect 13722 -4045 13797 -3896
rect 13718 -4046 13797 -4045
rect 13572 -4152 13797 -4046
rect 3666 -4236 3682 -4202
rect 3716 -4236 3732 -4202
rect 10217 -4238 10233 -4204
rect 10267 -4238 10283 -4204
rect 3548 -4353 3564 -4319
rect 3598 -4353 3614 -4319
rect 5217 -4330 5487 -4295
rect 4863 -4383 4897 -4367
rect 3152 -4403 3186 -4387
rect 3152 -4795 3186 -4779
rect 3270 -4403 3304 -4387
rect 3270 -4795 3304 -4779
rect 3388 -4403 3422 -4387
rect 3505 -4403 3539 -4387
rect 3505 -4595 3539 -4579
rect 3623 -4403 3657 -4387
rect 3623 -4595 3657 -4579
rect 4379 -4529 4649 -4494
rect 4379 -4583 4413 -4529
rect 3388 -4795 3422 -4779
rect 3675 -4729 3924 -4686
rect 3675 -4819 3722 -4729
rect 3885 -4819 3924 -4729
rect 4379 -4775 4413 -4759
rect 4497 -4583 4531 -4567
rect 4497 -4775 4531 -4759
rect 4615 -4583 4649 -4529
rect 4615 -4775 4649 -4759
rect 4733 -4583 4767 -4567
rect 4733 -4775 4767 -4759
rect 4863 -4775 4897 -4759
rect 4981 -4383 5015 -4367
rect 4981 -4775 5015 -4759
rect 5099 -4383 5133 -4367
rect 5099 -4775 5133 -4759
rect 5217 -4383 5251 -4330
rect 5217 -4775 5251 -4759
rect 5335 -4383 5369 -4367
rect 5335 -4775 5369 -4759
rect 5453 -4383 5487 -4330
rect 7115 -4330 7385 -4295
rect 5453 -4775 5487 -4759
rect 5571 -4383 5605 -4367
rect 6761 -4383 6795 -4367
rect 6277 -4529 6547 -4494
rect 5571 -4775 5605 -4759
rect 5700 -4583 5734 -4567
rect 5700 -4775 5734 -4759
rect 5818 -4583 5852 -4567
rect 5818 -4775 5852 -4759
rect 5936 -4583 5970 -4567
rect 5936 -4775 5970 -4759
rect 6054 -4583 6088 -4567
rect 6054 -4775 6088 -4759
rect 6277 -4583 6311 -4529
rect 6277 -4775 6311 -4759
rect 6395 -4583 6429 -4567
rect 6395 -4775 6429 -4759
rect 6513 -4583 6547 -4529
rect 6513 -4775 6547 -4759
rect 6631 -4583 6665 -4567
rect 6631 -4775 6665 -4759
rect 6761 -4775 6795 -4759
rect 6879 -4383 6913 -4367
rect 6879 -4775 6913 -4759
rect 6997 -4383 7031 -4367
rect 6997 -4775 7031 -4759
rect 7115 -4383 7149 -4330
rect 7115 -4775 7149 -4759
rect 7233 -4383 7267 -4367
rect 7233 -4775 7267 -4759
rect 7351 -4383 7385 -4330
rect 10099 -4355 10115 -4321
rect 10149 -4355 10165 -4321
rect 11768 -4332 12038 -4297
rect 7351 -4775 7385 -4759
rect 7469 -4383 7503 -4367
rect 11414 -4385 11448 -4369
rect 9703 -4405 9737 -4389
rect 7469 -4775 7503 -4759
rect 7598 -4583 7632 -4567
rect 7598 -4775 7632 -4759
rect 7716 -4583 7750 -4567
rect 7716 -4775 7750 -4759
rect 7834 -4583 7868 -4567
rect 7834 -4775 7868 -4759
rect 7952 -4583 7986 -4567
rect 7952 -4775 7986 -4759
rect 9703 -4797 9737 -4781
rect 9821 -4405 9855 -4389
rect 9821 -4797 9855 -4781
rect 9939 -4405 9973 -4389
rect 10056 -4405 10090 -4389
rect 10056 -4597 10090 -4581
rect 10174 -4405 10208 -4389
rect 10174 -4597 10208 -4581
rect 10930 -4531 11200 -4496
rect 10930 -4585 10964 -4531
rect 9939 -4797 9973 -4781
rect 10226 -4731 10475 -4688
rect 3195 -4863 3211 -4829
rect 3245 -4863 3261 -4829
rect 3313 -4863 3329 -4829
rect 3363 -4863 3379 -4829
rect 3675 -4858 3924 -4819
rect 10226 -4821 10273 -4731
rect 10436 -4821 10475 -4731
rect 10930 -4777 10964 -4761
rect 11048 -4585 11082 -4569
rect 11048 -4777 11082 -4761
rect 11166 -4585 11200 -4531
rect 11166 -4777 11200 -4761
rect 11284 -4585 11318 -4569
rect 11284 -4777 11318 -4761
rect 11414 -4777 11448 -4761
rect 11532 -4385 11566 -4369
rect 11532 -4777 11566 -4761
rect 11650 -4385 11684 -4369
rect 11650 -4777 11684 -4761
rect 11768 -4385 11802 -4332
rect 11768 -4777 11802 -4761
rect 11886 -4385 11920 -4369
rect 11886 -4777 11920 -4761
rect 12004 -4385 12038 -4332
rect 13666 -4332 13936 -4297
rect 12004 -4777 12038 -4761
rect 12122 -4385 12156 -4369
rect 13312 -4385 13346 -4369
rect 12828 -4531 13098 -4496
rect 12122 -4777 12156 -4761
rect 12251 -4585 12285 -4569
rect 12251 -4777 12285 -4761
rect 12369 -4585 12403 -4569
rect 12369 -4777 12403 -4761
rect 12487 -4585 12521 -4569
rect 12487 -4777 12521 -4761
rect 12605 -4585 12639 -4569
rect 12605 -4777 12639 -4761
rect 12828 -4585 12862 -4531
rect 12828 -4777 12862 -4761
rect 12946 -4585 12980 -4569
rect 12946 -4777 12980 -4761
rect 13064 -4585 13098 -4531
rect 13064 -4777 13098 -4761
rect 13182 -4585 13216 -4569
rect 13182 -4777 13216 -4761
rect 13312 -4777 13346 -4761
rect 13430 -4385 13464 -4369
rect 13430 -4777 13464 -4761
rect 13548 -4385 13582 -4369
rect 13548 -4777 13582 -4761
rect 13666 -4385 13700 -4332
rect 13666 -4777 13700 -4761
rect 13784 -4385 13818 -4369
rect 13784 -4777 13818 -4761
rect 13902 -4385 13936 -4332
rect 13902 -4777 13936 -4761
rect 14020 -4385 14054 -4369
rect 14020 -4777 14054 -4761
rect 14149 -4585 14183 -4569
rect 14149 -4777 14183 -4761
rect 14267 -4585 14301 -4569
rect 14267 -4777 14301 -4761
rect 14385 -4585 14419 -4569
rect 14385 -4777 14419 -4761
rect 14503 -4585 14537 -4569
rect 14503 -4777 14537 -4761
rect 9746 -4865 9762 -4831
rect 9796 -4865 9812 -4831
rect 9864 -4865 9880 -4831
rect 9914 -4865 9930 -4831
rect 10226 -4860 10475 -4821
rect 5843 -4997 5877 -4981
rect 12394 -4999 12428 -4983
rect 5843 -5047 5877 -5031
rect 7933 -5018 8000 -5002
rect 7933 -5052 7950 -5018
rect 7984 -5052 8000 -5018
rect 12394 -5049 12428 -5033
rect 14484 -5020 14551 -5004
rect 4806 -5076 4840 -5060
rect 3305 -5153 3528 -5080
rect 3305 -5302 3382 -5153
rect 3449 -5156 3528 -5153
rect 3305 -5305 3384 -5302
rect 3451 -5305 3528 -5156
rect 3305 -5411 3528 -5305
rect 4924 -5076 4958 -5060
rect 4806 -5468 4840 -5452
rect 4923 -5452 4924 -5405
rect 5042 -5076 5076 -5060
rect 4958 -5452 4959 -5405
rect 3736 -5520 4006 -5486
rect 2910 -5570 2944 -5554
rect 2910 -5762 2944 -5746
rect 3028 -5570 3062 -5554
rect 3028 -5762 3062 -5746
rect 3146 -5570 3180 -5554
rect 3146 -5762 3180 -5746
rect 3264 -5570 3298 -5554
rect 3264 -5762 3298 -5746
rect 3382 -5570 3416 -5554
rect 3382 -5762 3416 -5746
rect 3500 -5570 3534 -5554
rect 3500 -5762 3534 -5746
rect 3618 -5570 3652 -5554
rect 3618 -5762 3652 -5746
rect 3736 -5570 3770 -5520
rect 3736 -5762 3770 -5746
rect 3854 -5570 3888 -5554
rect 3854 -5762 3888 -5746
rect 3972 -5570 4006 -5520
rect 4923 -5510 4959 -5452
rect 5160 -5076 5194 -5060
rect 5042 -5468 5076 -5452
rect 5158 -5452 5160 -5405
rect 5158 -5510 5194 -5452
rect 5278 -5076 5312 -5060
rect 5278 -5468 5312 -5452
rect 5396 -5076 5430 -5060
rect 5514 -5076 5548 -5060
rect 5430 -5452 5432 -5406
rect 5396 -5510 5432 -5452
rect 5514 -5468 5548 -5452
rect 6704 -5076 6738 -5060
rect 6822 -5076 6856 -5060
rect 6704 -5468 6738 -5452
rect 6821 -5452 6822 -5405
rect 6940 -5076 6974 -5060
rect 6856 -5452 6857 -5405
rect 6019 -5510 6516 -5492
rect 4923 -5513 6516 -5510
rect 4923 -5547 6464 -5513
rect 6498 -5547 6516 -5513
rect 4923 -5550 6516 -5547
rect 6821 -5510 6857 -5452
rect 7058 -5076 7092 -5060
rect 6940 -5468 6974 -5452
rect 7056 -5452 7058 -5405
rect 7056 -5510 7092 -5452
rect 7176 -5076 7210 -5060
rect 7176 -5468 7210 -5452
rect 7294 -5076 7328 -5060
rect 7412 -5076 7446 -5060
rect 7933 -5068 8000 -5052
rect 14484 -5054 14501 -5020
rect 14535 -5054 14551 -5020
rect 7328 -5452 7330 -5406
rect 7294 -5510 7330 -5452
rect 11357 -5078 11391 -5062
rect 9856 -5158 10079 -5082
rect 9856 -5307 9935 -5158
rect 10005 -5307 10079 -5158
rect 9856 -5413 10079 -5307
rect 7412 -5468 7446 -5452
rect 11475 -5078 11509 -5062
rect 11357 -5470 11391 -5454
rect 11474 -5454 11475 -5407
rect 11593 -5078 11627 -5062
rect 11509 -5454 11510 -5407
rect 7917 -5481 8017 -5480
rect 7917 -5510 8073 -5481
rect 6821 -5550 8073 -5510
rect 4942 -5551 6516 -5550
rect 6840 -5551 8073 -5550
rect 4820 -5640 4887 -5624
rect 4820 -5674 4836 -5640
rect 4870 -5674 4887 -5640
rect 4820 -5690 4887 -5674
rect 3972 -5762 4006 -5746
rect 4651 -5707 4685 -5691
rect 4651 -5757 4685 -5741
rect 4997 -5792 5031 -5551
rect 6019 -5568 6516 -5551
rect 5467 -5640 5534 -5624
rect 5467 -5674 5484 -5640
rect 5518 -5674 5534 -5640
rect 5467 -5690 5534 -5674
rect 6718 -5640 6785 -5624
rect 6718 -5674 6734 -5640
rect 6768 -5674 6785 -5640
rect 6718 -5690 6785 -5674
rect 5774 -5708 5808 -5692
rect 5086 -5758 5102 -5724
rect 5136 -5758 5152 -5724
rect 5204 -5757 5220 -5723
rect 5254 -5757 5270 -5723
rect 5774 -5758 5808 -5742
rect 6549 -5707 6583 -5691
rect 6549 -5757 6583 -5741
rect 6895 -5792 6929 -5551
rect 7917 -5579 8073 -5551
rect 10287 -5522 10557 -5488
rect 9461 -5572 9495 -5556
rect 7917 -5580 8017 -5579
rect 7363 -5639 7430 -5623
rect 7363 -5673 7380 -5639
rect 7414 -5673 7430 -5639
rect 7363 -5689 7430 -5673
rect 7672 -5708 7706 -5692
rect 6984 -5758 7000 -5724
rect 7034 -5758 7050 -5724
rect 7102 -5757 7118 -5723
rect 7152 -5757 7168 -5723
rect 7672 -5758 7706 -5742
rect 9461 -5764 9495 -5748
rect 9579 -5572 9613 -5556
rect 9579 -5764 9613 -5748
rect 9697 -5572 9731 -5556
rect 9697 -5764 9731 -5748
rect 9815 -5572 9849 -5556
rect 9815 -5764 9849 -5748
rect 9933 -5572 9967 -5556
rect 9933 -5764 9967 -5748
rect 10051 -5572 10085 -5556
rect 10051 -5764 10085 -5748
rect 10169 -5572 10203 -5556
rect 10169 -5764 10203 -5748
rect 10287 -5572 10321 -5522
rect 10287 -5764 10321 -5748
rect 10405 -5572 10439 -5556
rect 10405 -5764 10439 -5748
rect 10523 -5572 10557 -5522
rect 11474 -5512 11510 -5454
rect 11711 -5078 11745 -5062
rect 11593 -5470 11627 -5454
rect 11709 -5454 11711 -5407
rect 11709 -5512 11745 -5454
rect 11829 -5078 11863 -5062
rect 11829 -5470 11863 -5454
rect 11947 -5078 11981 -5062
rect 12065 -5078 12099 -5062
rect 11981 -5454 11983 -5408
rect 11947 -5512 11983 -5454
rect 12065 -5470 12099 -5454
rect 13255 -5078 13289 -5062
rect 13373 -5078 13407 -5062
rect 13255 -5470 13289 -5454
rect 13372 -5454 13373 -5407
rect 13491 -5078 13525 -5062
rect 13407 -5454 13408 -5407
rect 12570 -5512 13067 -5494
rect 11474 -5515 13067 -5512
rect 11474 -5549 13015 -5515
rect 13049 -5549 13067 -5515
rect 11474 -5552 13067 -5549
rect 13372 -5512 13408 -5454
rect 13609 -5078 13643 -5062
rect 13491 -5470 13525 -5454
rect 13607 -5454 13609 -5407
rect 13607 -5512 13643 -5454
rect 13727 -5078 13761 -5062
rect 13727 -5470 13761 -5454
rect 13845 -5078 13879 -5062
rect 13963 -5078 13997 -5062
rect 14484 -5070 14551 -5054
rect 13879 -5454 13881 -5408
rect 13845 -5512 13881 -5454
rect 13963 -5470 13997 -5454
rect 14468 -5512 14775 -5482
rect 13372 -5552 14775 -5512
rect 11493 -5553 13067 -5552
rect 13391 -5553 14775 -5552
rect 11371 -5642 11438 -5626
rect 11371 -5676 11387 -5642
rect 11421 -5676 11438 -5642
rect 11371 -5692 11438 -5676
rect 10523 -5764 10557 -5748
rect 11202 -5709 11236 -5693
rect 11202 -5759 11236 -5743
rect 3661 -5840 3677 -5806
rect 3711 -5840 3727 -5806
rect 4504 -5808 4538 -5792
rect 3543 -5957 3559 -5923
rect 3593 -5957 3609 -5923
rect 3147 -6007 3181 -5991
rect 3147 -6399 3181 -6383
rect 3265 -6007 3299 -5991
rect 3265 -6399 3299 -6383
rect 3383 -6007 3417 -5991
rect 3500 -6007 3534 -5991
rect 3500 -6199 3534 -6183
rect 3618 -6007 3652 -5991
rect 4504 -6000 4538 -5984
rect 4622 -5808 4656 -5792
rect 4622 -6000 4656 -5984
rect 4924 -5808 4958 -5792
rect 3618 -6199 3652 -6183
rect 4997 -5808 5076 -5792
rect 4997 -5838 5042 -5808
rect 4924 -6251 4959 -6184
rect 5042 -6200 5076 -6184
rect 5160 -5808 5194 -5792
rect 5160 -6200 5194 -6184
rect 5278 -5808 5312 -5792
rect 5396 -5808 5430 -5792
rect 5802 -5808 5836 -5792
rect 5802 -6000 5836 -5984
rect 5920 -5808 5954 -5792
rect 5920 -6000 5954 -5984
rect 6402 -5808 6436 -5792
rect 6402 -6000 6436 -5984
rect 6520 -5808 6554 -5792
rect 6520 -6000 6554 -5984
rect 6822 -5808 6856 -5792
rect 5278 -6200 5312 -6184
rect 5395 -6251 5430 -6184
rect 4924 -6286 5430 -6251
rect 6895 -5808 6974 -5792
rect 6895 -5838 6940 -5808
rect 6822 -6251 6857 -6184
rect 6940 -6200 6974 -6184
rect 7058 -5808 7092 -5792
rect 7058 -6200 7092 -6184
rect 7176 -5808 7210 -5792
rect 7294 -5808 7328 -5792
rect 7700 -5808 7734 -5792
rect 7700 -6000 7734 -5984
rect 7818 -5808 7852 -5792
rect 11548 -5794 11582 -5553
rect 12570 -5570 13067 -5553
rect 12018 -5642 12085 -5626
rect 12018 -5676 12035 -5642
rect 12069 -5676 12085 -5642
rect 12018 -5692 12085 -5676
rect 13269 -5642 13336 -5626
rect 13269 -5676 13285 -5642
rect 13319 -5676 13336 -5642
rect 13269 -5692 13336 -5676
rect 12325 -5710 12359 -5694
rect 11637 -5760 11653 -5726
rect 11687 -5760 11703 -5726
rect 11755 -5759 11771 -5725
rect 11805 -5759 11821 -5725
rect 12325 -5760 12359 -5744
rect 13100 -5709 13134 -5693
rect 13100 -5759 13134 -5743
rect 13446 -5794 13480 -5553
rect 14468 -5582 14775 -5553
rect 14540 -5583 14775 -5582
rect 13914 -5641 13981 -5625
rect 13914 -5675 13931 -5641
rect 13965 -5675 13981 -5641
rect 13914 -5691 13981 -5675
rect 14223 -5710 14257 -5694
rect 13535 -5760 13551 -5726
rect 13585 -5760 13601 -5726
rect 13653 -5759 13669 -5725
rect 13703 -5759 13719 -5725
rect 14223 -5760 14257 -5744
rect 10212 -5842 10228 -5808
rect 10262 -5842 10278 -5808
rect 11055 -5810 11089 -5794
rect 10094 -5959 10110 -5925
rect 10144 -5959 10160 -5925
rect 7818 -6000 7852 -5984
rect 7176 -6200 7210 -6184
rect 7293 -6251 7328 -6184
rect 6822 -6286 7328 -6251
rect 9698 -6009 9732 -5993
rect 3383 -6399 3417 -6383
rect 3670 -6333 3919 -6290
rect 3670 -6423 3717 -6333
rect 3880 -6423 3919 -6333
rect 9698 -6401 9732 -6385
rect 9816 -6009 9850 -5993
rect 9816 -6401 9850 -6385
rect 9934 -6009 9968 -5993
rect 10051 -6009 10085 -5993
rect 10051 -6201 10085 -6185
rect 10169 -6009 10203 -5993
rect 11055 -6002 11089 -5986
rect 11173 -5810 11207 -5794
rect 11173 -6002 11207 -5986
rect 11475 -5810 11509 -5794
rect 10169 -6201 10203 -6185
rect 11548 -5810 11627 -5794
rect 11548 -5840 11593 -5810
rect 11475 -6253 11510 -6186
rect 11593 -6202 11627 -6186
rect 11711 -5810 11745 -5794
rect 11711 -6202 11745 -6186
rect 11829 -5810 11863 -5794
rect 11947 -5810 11981 -5794
rect 12353 -5810 12387 -5794
rect 12353 -6002 12387 -5986
rect 12471 -5810 12505 -5794
rect 12471 -6002 12505 -5986
rect 12953 -5810 12987 -5794
rect 12953 -6002 12987 -5986
rect 13071 -5810 13105 -5794
rect 13071 -6002 13105 -5986
rect 13373 -5810 13407 -5794
rect 11829 -6202 11863 -6186
rect 11946 -6253 11981 -6186
rect 11475 -6288 11981 -6253
rect 13446 -5810 13525 -5794
rect 13446 -5840 13491 -5810
rect 13373 -6253 13408 -6186
rect 13491 -6202 13525 -6186
rect 13609 -5810 13643 -5794
rect 13609 -6202 13643 -6186
rect 13727 -5810 13761 -5794
rect 13845 -5810 13879 -5794
rect 14251 -5810 14285 -5794
rect 14251 -6002 14285 -5986
rect 14369 -5810 14403 -5794
rect 14369 -6002 14403 -5986
rect 13727 -6202 13761 -6186
rect 13844 -6253 13879 -6186
rect 13373 -6288 13879 -6253
rect 9934 -6401 9968 -6385
rect 10221 -6335 10470 -6292
rect 3190 -6467 3206 -6433
rect 3240 -6467 3256 -6433
rect 3308 -6467 3324 -6433
rect 3358 -6467 3374 -6433
rect 3670 -6462 3919 -6423
rect 10221 -6425 10268 -6335
rect 10431 -6425 10470 -6335
rect 5095 -6493 5267 -6446
rect 9741 -6469 9757 -6435
rect 9791 -6469 9807 -6435
rect 9859 -6469 9875 -6435
rect 9909 -6469 9925 -6435
rect 10221 -6464 10470 -6425
rect 5095 -6656 5134 -6493
rect 5224 -6656 5267 -6493
rect 5095 -6696 5267 -6656
rect 11646 -6495 11818 -6448
rect 11646 -6658 11685 -6495
rect 11775 -6658 11818 -6495
rect 11646 -6698 11818 -6658
rect 14641 -6938 14775 -5583
rect 15255 -6603 15423 -2431
rect 16107 -2509 16141 -2493
rect 16225 -2317 16259 -2301
rect 16225 -2509 16259 -2493
rect 16343 -2317 16377 -2301
rect 16343 -2509 16377 -2493
rect 16461 -2317 16495 -2301
rect 16461 -2509 16495 -2493
rect 16579 -2317 16613 -2301
rect 16579 -2509 16613 -2493
rect 16697 -2317 16731 -2301
rect 16697 -2509 16731 -2493
rect 16815 -2317 16849 -2301
rect 16815 -2509 16849 -2493
rect 16933 -2317 16967 -2267
rect 16933 -2509 16967 -2493
rect 17051 -2317 17085 -2301
rect 17051 -2509 17085 -2493
rect 17169 -2317 17203 -2267
rect 17169 -2509 17203 -2493
rect 18432 -2245 18466 -2229
rect 16858 -2587 16874 -2553
rect 16908 -2587 16924 -2553
rect 18432 -2637 18466 -2621
rect 18550 -2245 18584 -2229
rect 18550 -2637 18584 -2621
rect 18668 -2245 18702 -2229
rect 18668 -2637 18702 -2621
rect 18786 -2245 18820 -2229
rect 18786 -2637 18820 -2621
rect 18904 -2245 18938 -2229
rect 18904 -2637 18938 -2621
rect 19022 -2245 19056 -2229
rect 19022 -2637 19056 -2621
rect 19140 -2245 19174 -2229
rect 19447 -2233 19481 -2217
rect 24939 -2186 24973 -2170
rect 19140 -2637 19174 -2621
rect 19574 -2241 19608 -2225
rect 19574 -2633 19608 -2617
rect 19692 -2241 19726 -2225
rect 19692 -2633 19726 -2617
rect 19810 -2241 19844 -2225
rect 19810 -2633 19844 -2617
rect 19928 -2241 19962 -2225
rect 19928 -2633 19962 -2617
rect 20046 -2241 20080 -2225
rect 20046 -2633 20080 -2617
rect 20164 -2241 20198 -2225
rect 20164 -2633 20198 -2617
rect 20282 -2241 20316 -2225
rect 23555 -2266 23825 -2232
rect 24939 -2236 24973 -2220
rect 26069 -2182 26103 -2166
rect 22729 -2316 22763 -2300
rect 22729 -2508 22763 -2492
rect 22847 -2316 22881 -2300
rect 22847 -2508 22881 -2492
rect 22965 -2316 22999 -2300
rect 22965 -2508 22999 -2492
rect 23083 -2316 23117 -2300
rect 23083 -2508 23117 -2492
rect 23201 -2316 23235 -2300
rect 23201 -2508 23235 -2492
rect 23319 -2316 23353 -2300
rect 23319 -2508 23353 -2492
rect 23437 -2316 23471 -2300
rect 23437 -2508 23471 -2492
rect 23555 -2316 23589 -2266
rect 23555 -2508 23589 -2492
rect 23673 -2316 23707 -2300
rect 23673 -2508 23707 -2492
rect 23791 -2316 23825 -2266
rect 23791 -2508 23825 -2492
rect 25054 -2244 25088 -2228
rect 23480 -2586 23496 -2552
rect 23530 -2586 23546 -2552
rect 20282 -2633 20316 -2617
rect 25054 -2636 25088 -2620
rect 25172 -2244 25206 -2228
rect 25172 -2636 25206 -2620
rect 25290 -2244 25324 -2228
rect 25290 -2636 25324 -2620
rect 25408 -2244 25442 -2228
rect 25408 -2636 25442 -2620
rect 25526 -2244 25560 -2228
rect 25526 -2636 25560 -2620
rect 25644 -2244 25678 -2228
rect 25644 -2636 25678 -2620
rect 25762 -2244 25796 -2228
rect 26069 -2232 26103 -2216
rect 25762 -2636 25796 -2620
rect 26196 -2240 26230 -2224
rect 26196 -2632 26230 -2616
rect 26314 -2240 26348 -2224
rect 26314 -2632 26348 -2616
rect 26432 -2240 26466 -2224
rect 26432 -2632 26466 -2616
rect 26550 -2240 26584 -2224
rect 26550 -2632 26584 -2616
rect 26668 -2240 26702 -2224
rect 26668 -2632 26702 -2616
rect 26786 -2240 26820 -2224
rect 26786 -2632 26820 -2616
rect 26904 -2240 26938 -2224
rect 28605 -2232 28639 -2216
rect 28723 -2040 28757 -2024
rect 28723 -2232 28757 -2216
rect 28841 -2040 28875 -2024
rect 28841 -2232 28875 -2216
rect 28959 -2040 28993 -2024
rect 28959 -2232 28993 -2216
rect 29077 -2040 29111 -2024
rect 29077 -2232 29111 -2216
rect 29195 -2040 29229 -2024
rect 29195 -2232 29229 -2216
rect 29313 -2040 29347 -2024
rect 29313 -2232 29347 -2216
rect 29431 -2040 29465 -1990
rect 29431 -2232 29465 -2216
rect 29549 -2040 29583 -2024
rect 29549 -2232 29583 -2216
rect 29667 -2040 29701 -1990
rect 29667 -2232 29701 -2216
rect 31187 -2254 31457 -2219
rect 29356 -2310 29372 -2276
rect 29406 -2310 29422 -2276
rect 30833 -2307 30867 -2291
rect 29238 -2427 29254 -2393
rect 29288 -2427 29304 -2393
rect 30349 -2453 30619 -2418
rect 26904 -2632 26938 -2616
rect 28842 -2477 28876 -2461
rect 16740 -2704 16756 -2670
rect 16790 -2704 16806 -2670
rect 23362 -2703 23378 -2669
rect 23412 -2703 23428 -2669
rect 16344 -2754 16378 -2738
rect 16344 -3146 16378 -3130
rect 16462 -2754 16496 -2738
rect 16462 -3146 16496 -3130
rect 16580 -2754 16614 -2738
rect 16697 -2754 16731 -2738
rect 16697 -2946 16731 -2930
rect 16815 -2754 16849 -2738
rect 16815 -2946 16849 -2930
rect 22966 -2753 23000 -2737
rect 18621 -2977 18637 -2943
rect 18671 -2977 18687 -2943
rect 19763 -2973 19779 -2939
rect 19813 -2973 19829 -2939
rect 18342 -3028 18376 -3012
rect 16580 -3146 16614 -3130
rect 16867 -3080 17116 -3037
rect 16867 -3170 16914 -3080
rect 17077 -3170 17116 -3080
rect 16387 -3214 16403 -3180
rect 16437 -3214 16453 -3180
rect 16505 -3214 16521 -3180
rect 16555 -3214 16571 -3180
rect 16867 -3209 17116 -3170
rect 18342 -3220 18376 -3204
rect 18460 -3028 18494 -3012
rect 18460 -3220 18494 -3204
rect 18578 -3028 18612 -3012
rect 18578 -3220 18612 -3204
rect 18696 -3028 18730 -3012
rect 18696 -3220 18730 -3204
rect 18861 -3028 18895 -3012
rect 18861 -3220 18895 -3204
rect 18979 -3028 19013 -3012
rect 18979 -3220 19013 -3204
rect 19097 -3028 19131 -3012
rect 19097 -3220 19131 -3204
rect 19215 -3028 19249 -3012
rect 19215 -3220 19249 -3204
rect 19484 -3024 19518 -3008
rect 19484 -3216 19518 -3200
rect 19602 -3024 19636 -3008
rect 19602 -3216 19636 -3200
rect 19720 -3024 19754 -3008
rect 19720 -3216 19754 -3200
rect 19838 -3024 19872 -3008
rect 19838 -3216 19872 -3200
rect 20003 -3024 20037 -3008
rect 20003 -3216 20037 -3200
rect 20121 -3024 20155 -3008
rect 20121 -3216 20155 -3200
rect 20239 -3024 20273 -3008
rect 20239 -3216 20273 -3200
rect 20357 -3024 20391 -3008
rect 22966 -3145 23000 -3129
rect 23084 -2753 23118 -2737
rect 23084 -3145 23118 -3129
rect 23202 -2753 23236 -2737
rect 23319 -2753 23353 -2737
rect 23319 -2945 23353 -2929
rect 23437 -2753 23471 -2737
rect 28842 -2869 28876 -2853
rect 28960 -2477 28994 -2461
rect 28960 -2869 28994 -2853
rect 29078 -2477 29112 -2461
rect 29195 -2477 29229 -2461
rect 29195 -2669 29229 -2653
rect 29313 -2477 29347 -2461
rect 29313 -2669 29347 -2653
rect 30349 -2507 30383 -2453
rect 30349 -2699 30383 -2683
rect 30467 -2507 30501 -2491
rect 30467 -2699 30501 -2683
rect 30585 -2507 30619 -2453
rect 30585 -2699 30619 -2683
rect 30703 -2507 30737 -2491
rect 30703 -2699 30737 -2683
rect 30833 -2699 30867 -2683
rect 30951 -2307 30985 -2291
rect 30951 -2699 30985 -2683
rect 31069 -2307 31103 -2291
rect 31069 -2699 31103 -2683
rect 31187 -2307 31221 -2254
rect 31187 -2699 31221 -2683
rect 31305 -2307 31339 -2291
rect 31305 -2699 31339 -2683
rect 31423 -2307 31457 -2254
rect 32431 -2270 32599 -2254
rect 31423 -2699 31457 -2683
rect 31541 -2307 31575 -2291
rect 32431 -2340 32447 -2270
rect 32583 -2340 32599 -2270
rect 32431 -2356 32599 -2340
rect 32968 -2460 33238 -2426
rect 31541 -2699 31575 -2683
rect 31670 -2507 31704 -2491
rect 31670 -2699 31704 -2683
rect 31788 -2507 31822 -2491
rect 31788 -2699 31822 -2683
rect 31906 -2507 31940 -2491
rect 31906 -2699 31940 -2683
rect 32024 -2507 32058 -2491
rect 32024 -2699 32058 -2683
rect 32142 -2510 32176 -2494
rect 32142 -2702 32176 -2686
rect 32260 -2510 32294 -2494
rect 32260 -2702 32294 -2686
rect 32378 -2510 32412 -2494
rect 32378 -2702 32412 -2686
rect 32496 -2510 32530 -2494
rect 32496 -2702 32530 -2686
rect 32614 -2510 32648 -2494
rect 32614 -2702 32648 -2686
rect 32732 -2510 32766 -2494
rect 32732 -2702 32766 -2686
rect 32850 -2510 32884 -2494
rect 32850 -2702 32884 -2686
rect 32968 -2510 33002 -2460
rect 32968 -2702 33002 -2686
rect 33086 -2510 33120 -2494
rect 33086 -2702 33120 -2686
rect 33204 -2510 33238 -2460
rect 33204 -2702 33238 -2686
rect 32893 -2780 32909 -2746
rect 32943 -2780 32959 -2746
rect 29078 -2869 29112 -2853
rect 32001 -2865 32035 -2849
rect 32775 -2897 32791 -2863
rect 32825 -2897 32841 -2863
rect 23437 -2945 23471 -2929
rect 28885 -2937 28901 -2903
rect 28935 -2937 28951 -2903
rect 29003 -2937 29019 -2903
rect 29053 -2937 29069 -2903
rect 32001 -2915 32035 -2899
rect 25243 -2976 25259 -2942
rect 25293 -2976 25309 -2942
rect 26385 -2972 26401 -2938
rect 26435 -2972 26451 -2938
rect 32379 -2947 32413 -2931
rect 30595 -2984 30651 -2967
rect 24964 -3027 24998 -3011
rect 23202 -3145 23236 -3129
rect 23489 -3079 23738 -3036
rect 23489 -3169 23536 -3079
rect 23699 -3169 23738 -3079
rect 20357 -3216 20391 -3200
rect 23009 -3213 23025 -3179
rect 23059 -3213 23075 -3179
rect 23127 -3213 23143 -3179
rect 23177 -3213 23193 -3179
rect 23489 -3208 23738 -3169
rect 24964 -3219 24998 -3203
rect 25082 -3027 25116 -3011
rect 25082 -3219 25116 -3203
rect 25200 -3027 25234 -3011
rect 25200 -3219 25234 -3203
rect 25318 -3027 25352 -3011
rect 25318 -3219 25352 -3203
rect 25483 -3027 25517 -3011
rect 25483 -3219 25517 -3203
rect 25601 -3027 25635 -3011
rect 25601 -3219 25635 -3203
rect 25719 -3027 25753 -3011
rect 25719 -3219 25753 -3203
rect 25837 -3027 25871 -3011
rect 25837 -3219 25871 -3203
rect 26106 -3023 26140 -3007
rect 26106 -3215 26140 -3199
rect 26224 -3023 26258 -3007
rect 26224 -3215 26258 -3199
rect 26342 -3023 26376 -3007
rect 26342 -3215 26376 -3199
rect 26460 -3023 26494 -3007
rect 26460 -3215 26494 -3199
rect 26625 -3023 26659 -3007
rect 26625 -3215 26659 -3199
rect 26743 -3023 26777 -3007
rect 26743 -3215 26777 -3199
rect 26861 -3023 26895 -3007
rect 26861 -3215 26895 -3199
rect 26979 -3023 27013 -3007
rect 29118 -3008 29286 -2990
rect 29118 -3064 29134 -3008
rect 29268 -3064 29286 -3008
rect 30595 -3018 30601 -2984
rect 30635 -3018 30651 -2984
rect 30595 -3035 30651 -3018
rect 30776 -3000 30810 -2984
rect 29118 -3080 29286 -3064
rect 26979 -3215 27013 -3199
rect 30894 -3000 30928 -2984
rect 30776 -3392 30810 -3376
rect 30893 -3376 30894 -3329
rect 31012 -3000 31046 -2984
rect 30928 -3376 30929 -3329
rect 18357 -3451 18529 -3404
rect 16516 -3552 16739 -3477
rect 16516 -3553 16598 -3552
rect 16516 -3702 16595 -3553
rect 16665 -3701 16739 -3552
rect 18357 -3614 18396 -3451
rect 18486 -3614 18529 -3451
rect 18357 -3653 18529 -3614
rect 19499 -3453 19671 -3406
rect 19499 -3616 19538 -3453
rect 19628 -3616 19671 -3453
rect 24979 -3450 25151 -3403
rect 19499 -3655 19671 -3616
rect 23138 -3551 23361 -3476
rect 16662 -3702 16739 -3701
rect 16516 -3808 16739 -3702
rect 23138 -3701 23217 -3551
rect 23284 -3701 23361 -3551
rect 24979 -3613 25018 -3450
rect 25108 -3613 25151 -3450
rect 24979 -3652 25151 -3613
rect 26121 -3452 26293 -3405
rect 26121 -3615 26160 -3452
rect 26250 -3615 26293 -3452
rect 30893 -3434 30929 -3376
rect 31130 -3000 31164 -2984
rect 31012 -3392 31046 -3376
rect 31128 -3376 31130 -3329
rect 31128 -3434 31164 -3376
rect 31248 -3000 31282 -2984
rect 31248 -3392 31282 -3376
rect 31366 -3000 31400 -2984
rect 31484 -3000 31518 -2984
rect 31400 -3376 31402 -3330
rect 31366 -3434 31402 -3376
rect 31646 -3205 31716 -3201
rect 31646 -3296 31650 -3205
rect 31712 -3296 31716 -3205
rect 31646 -3301 31716 -3296
rect 31484 -3392 31518 -3376
rect 31661 -3434 31702 -3301
rect 32379 -3339 32413 -3323
rect 32497 -2947 32531 -2931
rect 32497 -3339 32531 -3323
rect 32615 -2947 32649 -2931
rect 32732 -2947 32766 -2931
rect 32732 -3139 32766 -3123
rect 32850 -2947 32884 -2931
rect 32850 -3139 32884 -3123
rect 32615 -3339 32649 -3323
rect 32422 -3407 32438 -3373
rect 32472 -3407 32488 -3373
rect 32540 -3407 32556 -3373
rect 32590 -3407 32606 -3373
rect 30893 -3474 31702 -3434
rect 30912 -3475 31702 -3474
rect 30790 -3564 30857 -3548
rect 30790 -3598 30806 -3564
rect 30840 -3598 30857 -3564
rect 30790 -3614 30857 -3598
rect 26121 -3654 26293 -3615
rect 30621 -3631 30655 -3615
rect 30621 -3681 30655 -3665
rect 23138 -3807 23361 -3701
rect 30967 -3716 31001 -3475
rect 32655 -3478 32823 -3460
rect 32655 -3534 32671 -3478
rect 32805 -3534 32823 -3478
rect 31437 -3564 31504 -3548
rect 32655 -3550 32823 -3534
rect 31437 -3598 31454 -3564
rect 31488 -3598 31504 -3564
rect 31437 -3614 31504 -3598
rect 31744 -3632 31778 -3616
rect 31056 -3682 31072 -3648
rect 31106 -3682 31122 -3648
rect 31174 -3681 31190 -3647
rect 31224 -3681 31240 -3647
rect 31744 -3682 31778 -3666
rect 30474 -3732 30508 -3716
rect 16947 -3917 17217 -3883
rect 16121 -3967 16155 -3951
rect 16121 -4159 16155 -4143
rect 16239 -3967 16273 -3951
rect 16239 -4159 16273 -4143
rect 16357 -3967 16391 -3951
rect 16357 -4159 16391 -4143
rect 16475 -3967 16509 -3951
rect 16475 -4159 16509 -4143
rect 16593 -3967 16627 -3951
rect 16593 -4159 16627 -4143
rect 16711 -3967 16745 -3951
rect 16711 -4159 16745 -4143
rect 16829 -3967 16863 -3951
rect 16829 -4159 16863 -4143
rect 16947 -3967 16981 -3917
rect 16947 -4159 16981 -4143
rect 17065 -3967 17099 -3951
rect 17065 -4159 17099 -4143
rect 17183 -3967 17217 -3917
rect 17183 -4159 17217 -4143
rect 20227 -3894 20452 -3820
rect 20227 -3896 20309 -3894
rect 20227 -4045 20306 -3896
rect 20376 -4043 20452 -3894
rect 23569 -3916 23839 -3882
rect 20373 -4045 20452 -4043
rect 20227 -4151 20452 -4045
rect 22743 -3966 22777 -3950
rect 22743 -4158 22777 -4142
rect 22861 -3966 22895 -3950
rect 22861 -4158 22895 -4142
rect 22979 -3966 23013 -3950
rect 22979 -4158 23013 -4142
rect 23097 -3966 23131 -3950
rect 23097 -4158 23131 -4142
rect 23215 -3966 23249 -3950
rect 23215 -4158 23249 -4142
rect 23333 -3966 23367 -3950
rect 23333 -4158 23367 -4142
rect 23451 -3966 23485 -3950
rect 23451 -4158 23485 -4142
rect 23569 -3966 23603 -3916
rect 23569 -4158 23603 -4142
rect 23687 -3966 23721 -3950
rect 23687 -4158 23721 -4142
rect 23805 -3966 23839 -3916
rect 23805 -4158 23839 -4142
rect 26849 -3895 27074 -3819
rect 26849 -4044 26928 -3895
rect 26995 -3896 27074 -3895
rect 26849 -4045 26930 -4044
rect 26997 -4045 27074 -3896
rect 30474 -3924 30508 -3908
rect 30592 -3732 30626 -3716
rect 30592 -3924 30626 -3908
rect 30894 -3732 30928 -3716
rect 26849 -4150 27074 -4045
rect 30967 -3732 31046 -3716
rect 30967 -3762 31012 -3732
rect 30894 -4175 30929 -4108
rect 31012 -4124 31046 -4108
rect 31130 -3732 31164 -3716
rect 31130 -4124 31164 -4108
rect 31248 -3732 31282 -3716
rect 31366 -3732 31400 -3716
rect 31772 -3732 31806 -3716
rect 31772 -3924 31806 -3908
rect 31890 -3732 31924 -3716
rect 31890 -3924 31924 -3908
rect 31248 -4124 31282 -4108
rect 31365 -4175 31400 -4108
rect 16872 -4237 16888 -4203
rect 16922 -4237 16938 -4203
rect 23494 -4236 23510 -4202
rect 23544 -4236 23560 -4202
rect 30894 -4210 31400 -4175
rect 31041 -4279 31283 -4267
rect 16754 -4354 16770 -4320
rect 16804 -4354 16820 -4320
rect 18423 -4331 18693 -4296
rect 18069 -4384 18103 -4368
rect 16358 -4404 16392 -4388
rect 16358 -4796 16392 -4780
rect 16476 -4404 16510 -4388
rect 16476 -4796 16510 -4780
rect 16594 -4404 16628 -4388
rect 16711 -4404 16745 -4388
rect 16711 -4596 16745 -4580
rect 16829 -4404 16863 -4388
rect 16829 -4596 16863 -4580
rect 17585 -4530 17855 -4495
rect 17585 -4584 17619 -4530
rect 16594 -4796 16628 -4780
rect 16881 -4730 17130 -4687
rect 16881 -4820 16928 -4730
rect 17091 -4820 17130 -4730
rect 17585 -4776 17619 -4760
rect 17703 -4584 17737 -4568
rect 17703 -4776 17737 -4760
rect 17821 -4584 17855 -4530
rect 17821 -4776 17855 -4760
rect 17939 -4584 17973 -4568
rect 17939 -4776 17973 -4760
rect 18069 -4776 18103 -4760
rect 18187 -4384 18221 -4368
rect 18187 -4776 18221 -4760
rect 18305 -4384 18339 -4368
rect 18305 -4776 18339 -4760
rect 18423 -4384 18457 -4331
rect 18423 -4776 18457 -4760
rect 18541 -4384 18575 -4368
rect 18541 -4776 18575 -4760
rect 18659 -4384 18693 -4331
rect 20321 -4331 20591 -4296
rect 18659 -4776 18693 -4760
rect 18777 -4384 18811 -4368
rect 19967 -4384 20001 -4368
rect 19483 -4530 19753 -4495
rect 18777 -4776 18811 -4760
rect 18906 -4584 18940 -4568
rect 18906 -4776 18940 -4760
rect 19024 -4584 19058 -4568
rect 19024 -4776 19058 -4760
rect 19142 -4584 19176 -4568
rect 19142 -4776 19176 -4760
rect 19260 -4584 19294 -4568
rect 19260 -4776 19294 -4760
rect 19483 -4584 19517 -4530
rect 19483 -4776 19517 -4760
rect 19601 -4584 19635 -4568
rect 19601 -4776 19635 -4760
rect 19719 -4584 19753 -4530
rect 19719 -4776 19753 -4760
rect 19837 -4584 19871 -4568
rect 19837 -4776 19871 -4760
rect 19967 -4776 20001 -4760
rect 20085 -4384 20119 -4368
rect 20085 -4776 20119 -4760
rect 20203 -4384 20237 -4368
rect 20203 -4776 20237 -4760
rect 20321 -4384 20355 -4331
rect 20321 -4776 20355 -4760
rect 20439 -4384 20473 -4368
rect 20439 -4776 20473 -4760
rect 20557 -4384 20591 -4331
rect 23376 -4353 23392 -4319
rect 23426 -4353 23442 -4319
rect 25045 -4330 25315 -4295
rect 20557 -4776 20591 -4760
rect 20675 -4384 20709 -4368
rect 24691 -4383 24725 -4367
rect 22980 -4403 23014 -4387
rect 20675 -4776 20709 -4760
rect 20804 -4584 20838 -4568
rect 20804 -4776 20838 -4760
rect 20922 -4584 20956 -4568
rect 20922 -4776 20956 -4760
rect 21040 -4584 21074 -4568
rect 21040 -4776 21074 -4760
rect 21158 -4584 21192 -4568
rect 21158 -4776 21192 -4760
rect 22980 -4795 23014 -4779
rect 23098 -4403 23132 -4387
rect 23098 -4795 23132 -4779
rect 23216 -4403 23250 -4387
rect 23333 -4403 23367 -4387
rect 23333 -4595 23367 -4579
rect 23451 -4403 23485 -4387
rect 23451 -4595 23485 -4579
rect 24207 -4529 24477 -4494
rect 24207 -4583 24241 -4529
rect 23216 -4795 23250 -4779
rect 23503 -4729 23752 -4686
rect 16401 -4864 16417 -4830
rect 16451 -4864 16467 -4830
rect 16519 -4864 16535 -4830
rect 16569 -4864 16585 -4830
rect 16881 -4859 17130 -4820
rect 23503 -4819 23550 -4729
rect 23713 -4819 23752 -4729
rect 24207 -4775 24241 -4759
rect 24325 -4583 24359 -4567
rect 24325 -4775 24359 -4759
rect 24443 -4583 24477 -4529
rect 24443 -4775 24477 -4759
rect 24561 -4583 24595 -4567
rect 24561 -4775 24595 -4759
rect 24691 -4775 24725 -4759
rect 24809 -4383 24843 -4367
rect 24809 -4775 24843 -4759
rect 24927 -4383 24961 -4367
rect 24927 -4775 24961 -4759
rect 25045 -4383 25079 -4330
rect 25045 -4775 25079 -4759
rect 25163 -4383 25197 -4367
rect 25163 -4775 25197 -4759
rect 25281 -4383 25315 -4330
rect 26943 -4330 27213 -4295
rect 25281 -4775 25315 -4759
rect 25399 -4383 25433 -4367
rect 26589 -4383 26623 -4367
rect 26105 -4529 26375 -4494
rect 25399 -4775 25433 -4759
rect 25528 -4583 25562 -4567
rect 25528 -4775 25562 -4759
rect 25646 -4583 25680 -4567
rect 25646 -4775 25680 -4759
rect 25764 -4583 25798 -4567
rect 25764 -4775 25798 -4759
rect 25882 -4583 25916 -4567
rect 25882 -4775 25916 -4759
rect 26105 -4583 26139 -4529
rect 26105 -4775 26139 -4759
rect 26223 -4583 26257 -4567
rect 26223 -4775 26257 -4759
rect 26341 -4583 26375 -4529
rect 26341 -4775 26375 -4759
rect 26459 -4583 26493 -4567
rect 26459 -4775 26493 -4759
rect 26589 -4775 26623 -4759
rect 26707 -4383 26741 -4367
rect 26707 -4775 26741 -4759
rect 26825 -4383 26859 -4367
rect 26825 -4775 26859 -4759
rect 26943 -4383 26977 -4330
rect 26943 -4775 26977 -4759
rect 27061 -4383 27095 -4367
rect 27061 -4775 27095 -4759
rect 27179 -4383 27213 -4330
rect 27179 -4775 27213 -4759
rect 27297 -4383 27331 -4367
rect 31041 -4381 31088 -4279
rect 31223 -4381 31283 -4279
rect 31041 -4398 31283 -4381
rect 27297 -4775 27331 -4759
rect 27426 -4583 27460 -4567
rect 27426 -4775 27460 -4759
rect 27544 -4583 27578 -4567
rect 27544 -4775 27578 -4759
rect 27662 -4583 27696 -4567
rect 27662 -4775 27696 -4759
rect 27780 -4583 27814 -4567
rect 27780 -4775 27814 -4759
rect 23023 -4863 23039 -4829
rect 23073 -4863 23089 -4829
rect 23141 -4863 23157 -4829
rect 23191 -4863 23207 -4829
rect 23503 -4858 23752 -4819
rect 28891 -4870 29059 -4854
rect 28891 -4940 28907 -4870
rect 29043 -4940 29059 -4870
rect 28891 -4956 29059 -4940
rect 19049 -4998 19083 -4982
rect 25671 -4997 25705 -4981
rect 19049 -5048 19083 -5032
rect 21139 -5019 21206 -5003
rect 21139 -5053 21156 -5019
rect 21190 -5053 21206 -5019
rect 25671 -5047 25705 -5031
rect 27761 -5018 27828 -5002
rect 18012 -5077 18046 -5061
rect 16511 -5157 16734 -5081
rect 16511 -5306 16590 -5157
rect 16657 -5160 16734 -5157
rect 16511 -5309 16593 -5306
rect 16660 -5309 16734 -5160
rect 16511 -5412 16734 -5309
rect 18130 -5077 18164 -5061
rect 18012 -5469 18046 -5453
rect 18129 -5453 18130 -5406
rect 18248 -5077 18282 -5061
rect 18164 -5453 18165 -5406
rect 16942 -5521 17212 -5487
rect 16116 -5571 16150 -5555
rect 16116 -5763 16150 -5747
rect 16234 -5571 16268 -5555
rect 16234 -5763 16268 -5747
rect 16352 -5571 16386 -5555
rect 16352 -5763 16386 -5747
rect 16470 -5571 16504 -5555
rect 16470 -5763 16504 -5747
rect 16588 -5571 16622 -5555
rect 16588 -5763 16622 -5747
rect 16706 -5571 16740 -5555
rect 16706 -5763 16740 -5747
rect 16824 -5571 16858 -5555
rect 16824 -5763 16858 -5747
rect 16942 -5571 16976 -5521
rect 16942 -5763 16976 -5747
rect 17060 -5571 17094 -5555
rect 17060 -5763 17094 -5747
rect 17178 -5571 17212 -5521
rect 18129 -5511 18165 -5453
rect 18366 -5077 18400 -5061
rect 18248 -5469 18282 -5453
rect 18364 -5453 18366 -5406
rect 18364 -5511 18400 -5453
rect 18484 -5077 18518 -5061
rect 18484 -5469 18518 -5453
rect 18602 -5077 18636 -5061
rect 18720 -5077 18754 -5061
rect 18636 -5453 18638 -5407
rect 18602 -5511 18638 -5453
rect 18720 -5469 18754 -5453
rect 19910 -5077 19944 -5061
rect 20028 -5077 20062 -5061
rect 19910 -5469 19944 -5453
rect 20027 -5453 20028 -5406
rect 20146 -5077 20180 -5061
rect 20062 -5453 20063 -5406
rect 19225 -5511 19722 -5493
rect 18129 -5514 19722 -5511
rect 18129 -5548 19670 -5514
rect 19704 -5548 19722 -5514
rect 18129 -5551 19722 -5548
rect 20027 -5511 20063 -5453
rect 20264 -5077 20298 -5061
rect 20146 -5469 20180 -5453
rect 20262 -5453 20264 -5406
rect 20262 -5511 20298 -5453
rect 20382 -5077 20416 -5061
rect 20382 -5469 20416 -5453
rect 20500 -5077 20534 -5061
rect 20618 -5077 20652 -5061
rect 21139 -5069 21206 -5053
rect 27761 -5052 27778 -5018
rect 27812 -5052 27828 -5018
rect 20534 -5453 20536 -5407
rect 20500 -5511 20536 -5453
rect 24634 -5076 24668 -5060
rect 23133 -5156 23356 -5080
rect 23133 -5305 23212 -5156
rect 23279 -5160 23356 -5156
rect 23133 -5309 23214 -5305
rect 23281 -5309 23356 -5160
rect 23133 -5411 23356 -5309
rect 20618 -5469 20652 -5453
rect 24752 -5076 24786 -5060
rect 24634 -5468 24668 -5452
rect 24751 -5452 24752 -5405
rect 24870 -5076 24904 -5060
rect 24786 -5452 24787 -5405
rect 21123 -5482 21223 -5481
rect 21123 -5511 21279 -5482
rect 20027 -5551 21279 -5511
rect 18148 -5552 19722 -5551
rect 20046 -5552 21279 -5551
rect 18026 -5641 18093 -5625
rect 18026 -5675 18042 -5641
rect 18076 -5675 18093 -5641
rect 18026 -5691 18093 -5675
rect 17178 -5763 17212 -5747
rect 17857 -5708 17891 -5692
rect 17857 -5758 17891 -5742
rect 18203 -5793 18237 -5552
rect 19225 -5569 19722 -5552
rect 18673 -5641 18740 -5625
rect 18673 -5675 18690 -5641
rect 18724 -5675 18740 -5641
rect 18673 -5691 18740 -5675
rect 19924 -5641 19991 -5625
rect 19924 -5675 19940 -5641
rect 19974 -5675 19991 -5641
rect 19924 -5691 19991 -5675
rect 18980 -5709 19014 -5693
rect 18292 -5759 18308 -5725
rect 18342 -5759 18358 -5725
rect 18410 -5758 18426 -5724
rect 18460 -5758 18476 -5724
rect 18980 -5759 19014 -5743
rect 19755 -5708 19789 -5692
rect 19755 -5758 19789 -5742
rect 20101 -5793 20135 -5552
rect 21123 -5580 21279 -5552
rect 23564 -5520 23834 -5486
rect 22738 -5570 22772 -5554
rect 21123 -5581 21223 -5580
rect 20569 -5640 20636 -5624
rect 20569 -5674 20586 -5640
rect 20620 -5674 20636 -5640
rect 20569 -5690 20636 -5674
rect 20878 -5709 20912 -5693
rect 20190 -5759 20206 -5725
rect 20240 -5759 20256 -5725
rect 20308 -5758 20324 -5724
rect 20358 -5758 20374 -5724
rect 20878 -5759 20912 -5743
rect 22738 -5762 22772 -5746
rect 22856 -5570 22890 -5554
rect 22856 -5762 22890 -5746
rect 22974 -5570 23008 -5554
rect 22974 -5762 23008 -5746
rect 23092 -5570 23126 -5554
rect 23092 -5762 23126 -5746
rect 23210 -5570 23244 -5554
rect 23210 -5762 23244 -5746
rect 23328 -5570 23362 -5554
rect 23328 -5762 23362 -5746
rect 23446 -5570 23480 -5554
rect 23446 -5762 23480 -5746
rect 23564 -5570 23598 -5520
rect 23564 -5762 23598 -5746
rect 23682 -5570 23716 -5554
rect 23682 -5762 23716 -5746
rect 23800 -5570 23834 -5520
rect 24751 -5510 24787 -5452
rect 24988 -5076 25022 -5060
rect 24870 -5468 24904 -5452
rect 24986 -5452 24988 -5405
rect 24986 -5510 25022 -5452
rect 25106 -5076 25140 -5060
rect 25106 -5468 25140 -5452
rect 25224 -5076 25258 -5060
rect 25342 -5076 25376 -5060
rect 25258 -5452 25260 -5406
rect 25224 -5510 25260 -5452
rect 25342 -5468 25376 -5452
rect 26532 -5076 26566 -5060
rect 26650 -5076 26684 -5060
rect 26532 -5468 26566 -5452
rect 26649 -5452 26650 -5405
rect 26768 -5076 26802 -5060
rect 26684 -5452 26685 -5405
rect 25847 -5510 26344 -5492
rect 24751 -5513 26344 -5510
rect 24751 -5547 26292 -5513
rect 26326 -5547 26344 -5513
rect 24751 -5550 26344 -5547
rect 26649 -5510 26685 -5452
rect 26886 -5076 26920 -5060
rect 26768 -5468 26802 -5452
rect 26884 -5452 26886 -5405
rect 26884 -5510 26920 -5452
rect 27004 -5076 27038 -5060
rect 27004 -5468 27038 -5452
rect 27122 -5076 27156 -5060
rect 27240 -5076 27274 -5060
rect 27761 -5068 27828 -5052
rect 29428 -5060 29698 -5026
rect 27156 -5452 27158 -5406
rect 27122 -5510 27158 -5452
rect 28602 -5110 28636 -5094
rect 28602 -5302 28636 -5286
rect 28720 -5110 28754 -5094
rect 28720 -5302 28754 -5286
rect 28838 -5110 28872 -5094
rect 28838 -5302 28872 -5286
rect 28956 -5110 28990 -5094
rect 28956 -5302 28990 -5286
rect 29074 -5110 29108 -5094
rect 29074 -5302 29108 -5286
rect 29192 -5110 29226 -5094
rect 29192 -5302 29226 -5286
rect 29310 -5110 29344 -5094
rect 29310 -5302 29344 -5286
rect 29428 -5110 29462 -5060
rect 29428 -5302 29462 -5286
rect 29546 -5110 29580 -5094
rect 29546 -5302 29580 -5286
rect 29664 -5110 29698 -5060
rect 29664 -5302 29698 -5286
rect 29353 -5380 29369 -5346
rect 29403 -5380 29419 -5346
rect 27240 -5468 27274 -5452
rect 27745 -5481 27845 -5480
rect 27745 -5510 27901 -5481
rect 26649 -5550 27901 -5510
rect 24770 -5551 26344 -5550
rect 26668 -5551 27901 -5550
rect 24648 -5640 24715 -5624
rect 24648 -5674 24664 -5640
rect 24698 -5674 24715 -5640
rect 24648 -5690 24715 -5674
rect 23800 -5762 23834 -5746
rect 24479 -5707 24513 -5691
rect 24479 -5757 24513 -5741
rect 24825 -5792 24859 -5551
rect 25847 -5568 26344 -5551
rect 25295 -5640 25362 -5624
rect 25295 -5674 25312 -5640
rect 25346 -5674 25362 -5640
rect 25295 -5690 25362 -5674
rect 26546 -5640 26613 -5624
rect 26546 -5674 26562 -5640
rect 26596 -5674 26613 -5640
rect 26546 -5690 26613 -5674
rect 25602 -5708 25636 -5692
rect 24914 -5758 24930 -5724
rect 24964 -5758 24980 -5724
rect 25032 -5757 25048 -5723
rect 25082 -5757 25098 -5723
rect 25602 -5758 25636 -5742
rect 26377 -5707 26411 -5691
rect 26377 -5757 26411 -5741
rect 26723 -5792 26757 -5551
rect 27745 -5579 27901 -5551
rect 29235 -5497 29251 -5463
rect 29285 -5497 29301 -5463
rect 28839 -5547 28873 -5531
rect 27745 -5580 27845 -5579
rect 27191 -5639 27258 -5623
rect 27191 -5673 27208 -5639
rect 27242 -5673 27258 -5639
rect 27191 -5689 27258 -5673
rect 27500 -5708 27534 -5692
rect 26812 -5758 26828 -5724
rect 26862 -5758 26878 -5724
rect 26930 -5757 26946 -5723
rect 26980 -5757 26996 -5723
rect 27500 -5758 27534 -5742
rect 16867 -5841 16883 -5807
rect 16917 -5841 16933 -5807
rect 17710 -5809 17744 -5793
rect 16749 -5958 16765 -5924
rect 16799 -5958 16815 -5924
rect 16353 -6008 16387 -5992
rect 16353 -6400 16387 -6384
rect 16471 -6008 16505 -5992
rect 16471 -6400 16505 -6384
rect 16589 -6008 16623 -5992
rect 16706 -6008 16740 -5992
rect 16706 -6200 16740 -6184
rect 16824 -6008 16858 -5992
rect 17710 -6001 17744 -5985
rect 17828 -5809 17862 -5793
rect 17828 -6001 17862 -5985
rect 18130 -5809 18164 -5793
rect 16824 -6200 16858 -6184
rect 18203 -5809 18282 -5793
rect 18203 -5839 18248 -5809
rect 18130 -6252 18165 -6185
rect 18248 -6201 18282 -6185
rect 18366 -5809 18400 -5793
rect 18366 -6201 18400 -6185
rect 18484 -5809 18518 -5793
rect 18602 -5809 18636 -5793
rect 19008 -5809 19042 -5793
rect 19008 -6001 19042 -5985
rect 19126 -5809 19160 -5793
rect 19126 -6001 19160 -5985
rect 19608 -5809 19642 -5793
rect 19608 -6001 19642 -5985
rect 19726 -5809 19760 -5793
rect 19726 -6001 19760 -5985
rect 20028 -5809 20062 -5793
rect 18484 -6201 18518 -6185
rect 18601 -6252 18636 -6185
rect 18130 -6287 18636 -6252
rect 20101 -5809 20180 -5793
rect 20101 -5839 20146 -5809
rect 20028 -6252 20063 -6185
rect 20146 -6201 20180 -6185
rect 20264 -5809 20298 -5793
rect 20264 -6201 20298 -6185
rect 20382 -5809 20416 -5793
rect 20500 -5809 20534 -5793
rect 20906 -5809 20940 -5793
rect 20906 -6001 20940 -5985
rect 21024 -5809 21058 -5793
rect 23489 -5840 23505 -5806
rect 23539 -5840 23555 -5806
rect 24332 -5808 24366 -5792
rect 23371 -5957 23387 -5923
rect 23421 -5957 23437 -5923
rect 21024 -6001 21058 -5985
rect 20382 -6201 20416 -6185
rect 20499 -6252 20534 -6185
rect 20028 -6287 20534 -6252
rect 22975 -6007 23009 -5991
rect 16589 -6400 16623 -6384
rect 16876 -6334 17125 -6291
rect 16876 -6424 16923 -6334
rect 17086 -6354 17125 -6334
rect 17089 -6421 17125 -6354
rect 22975 -6399 23009 -6383
rect 23093 -6007 23127 -5991
rect 23093 -6399 23127 -6383
rect 23211 -6007 23245 -5991
rect 23328 -6007 23362 -5991
rect 23328 -6199 23362 -6183
rect 23446 -6007 23480 -5991
rect 24332 -6000 24366 -5984
rect 24450 -5808 24484 -5792
rect 24450 -6000 24484 -5984
rect 24752 -5808 24786 -5792
rect 23446 -6199 23480 -6183
rect 24825 -5808 24904 -5792
rect 24825 -5838 24870 -5808
rect 24752 -6251 24787 -6184
rect 24870 -6200 24904 -6184
rect 24988 -5808 25022 -5792
rect 24988 -6200 25022 -6184
rect 25106 -5808 25140 -5792
rect 25224 -5808 25258 -5792
rect 25630 -5808 25664 -5792
rect 25630 -6000 25664 -5984
rect 25748 -5808 25782 -5792
rect 25748 -6000 25782 -5984
rect 26230 -5808 26264 -5792
rect 26230 -6000 26264 -5984
rect 26348 -5808 26382 -5792
rect 26348 -6000 26382 -5984
rect 26650 -5808 26684 -5792
rect 25106 -6200 25140 -6184
rect 25223 -6251 25258 -6184
rect 24752 -6286 25258 -6251
rect 26723 -5808 26802 -5792
rect 26723 -5838 26768 -5808
rect 26650 -6251 26685 -6184
rect 26768 -6200 26802 -6184
rect 26886 -5808 26920 -5792
rect 26886 -6200 26920 -6184
rect 27004 -5808 27038 -5792
rect 27122 -5808 27156 -5792
rect 27528 -5808 27562 -5792
rect 27528 -6000 27562 -5984
rect 27646 -5808 27680 -5792
rect 28839 -5939 28873 -5923
rect 28957 -5547 28991 -5531
rect 28957 -5939 28991 -5923
rect 29075 -5547 29109 -5531
rect 29192 -5547 29226 -5531
rect 29192 -5739 29226 -5723
rect 29310 -5547 29344 -5531
rect 29310 -5739 29344 -5723
rect 29075 -5939 29109 -5923
rect 27646 -6000 27680 -5984
rect 28882 -6007 28898 -5973
rect 28932 -6007 28948 -5973
rect 29000 -6007 29016 -5973
rect 29050 -6007 29066 -5973
rect 29115 -6078 29283 -6060
rect 29115 -6134 29131 -6078
rect 29265 -6134 29283 -6078
rect 29115 -6150 29283 -6134
rect 30972 -6117 31416 -6111
rect 27004 -6200 27038 -6184
rect 27121 -6251 27156 -6184
rect 26650 -6286 27156 -6251
rect 23211 -6399 23245 -6383
rect 23498 -6333 23747 -6290
rect 30972 -6317 30983 -6117
rect 31404 -6317 31416 -6117
rect 30972 -6323 31416 -6317
rect 17086 -6424 17125 -6421
rect 16396 -6468 16412 -6434
rect 16446 -6468 16462 -6434
rect 16514 -6468 16530 -6434
rect 16564 -6468 16580 -6434
rect 16876 -6463 17125 -6424
rect 23498 -6423 23545 -6333
rect 23708 -6423 23747 -6333
rect 15255 -6671 15301 -6603
rect 15371 -6671 15423 -6603
rect 15255 -6684 15423 -6671
rect 18301 -6494 18473 -6447
rect 23018 -6467 23034 -6433
rect 23068 -6467 23084 -6433
rect 23136 -6467 23152 -6433
rect 23186 -6467 23202 -6433
rect 23498 -6462 23747 -6423
rect 18301 -6657 18340 -6494
rect 18430 -6657 18473 -6494
rect 18301 -6697 18473 -6657
rect 24923 -6493 25095 -6446
rect 24923 -6656 24962 -6493
rect 25052 -6656 25095 -6493
rect 31187 -6602 31457 -6567
rect 24923 -6696 25095 -6656
rect 30833 -6655 30867 -6639
rect 30349 -6801 30619 -6766
rect 30349 -6855 30383 -6801
rect 14641 -7090 29987 -6938
rect 30349 -7047 30383 -7031
rect 30467 -6855 30501 -6839
rect 30467 -7047 30501 -7031
rect 30585 -6855 30619 -6801
rect 30585 -7047 30619 -7031
rect 30703 -6855 30737 -6839
rect 30703 -7047 30737 -7031
rect 30833 -7047 30867 -7031
rect 30951 -6655 30985 -6639
rect 30951 -7047 30985 -7031
rect 31069 -6655 31103 -6639
rect 31069 -7047 31103 -7031
rect 31187 -6655 31221 -6602
rect 31187 -7047 31221 -7031
rect 31305 -6655 31339 -6639
rect 31305 -7047 31339 -7031
rect 31423 -6655 31457 -6602
rect 32431 -6618 32599 -6602
rect 31423 -7047 31457 -7031
rect 31541 -6655 31575 -6639
rect 32431 -6688 32447 -6618
rect 32583 -6688 32599 -6618
rect 32431 -6704 32599 -6688
rect 32968 -6808 33238 -6774
rect 31541 -7047 31575 -7031
rect 31670 -6855 31704 -6839
rect 31670 -7047 31704 -7031
rect 31788 -6855 31822 -6839
rect 31788 -7047 31822 -7031
rect 31906 -6855 31940 -6839
rect 31906 -7047 31940 -7031
rect 32024 -6855 32058 -6839
rect 32024 -7047 32058 -7031
rect 32142 -6858 32176 -6842
rect 32142 -7050 32176 -7034
rect 32260 -6858 32294 -6842
rect 32260 -7050 32294 -7034
rect 32378 -6858 32412 -6842
rect 32378 -7050 32412 -7034
rect 32496 -6858 32530 -6842
rect 32496 -7050 32530 -7034
rect 32614 -6858 32648 -6842
rect 32614 -7050 32648 -7034
rect 32732 -6858 32766 -6842
rect 32732 -7050 32766 -7034
rect 32850 -6858 32884 -6842
rect 32850 -7050 32884 -7034
rect 32968 -6858 33002 -6808
rect 32968 -7050 33002 -7034
rect 33086 -6858 33120 -6842
rect 33086 -7050 33120 -7034
rect 33204 -6858 33238 -6808
rect 33204 -7050 33238 -7034
rect 29895 -7187 29987 -7090
rect 32893 -7128 32909 -7094
rect 32943 -7128 32959 -7094
rect 29895 -7193 30415 -7187
rect 7231 -7225 7399 -7209
rect 7231 -7281 7247 -7225
rect 7381 -7281 7399 -7225
rect 7231 -7299 7399 -7281
rect 13785 -7220 13953 -7204
rect 13785 -7276 13801 -7220
rect 13935 -7276 13953 -7220
rect 13785 -7294 13953 -7276
rect 20434 -7232 20602 -7216
rect 20434 -7288 20450 -7232
rect 20584 -7288 20602 -7232
rect 29895 -7263 30329 -7193
rect 29896 -7264 30329 -7263
rect 30402 -7264 30415 -7193
rect 32001 -7213 32035 -7197
rect 32775 -7245 32791 -7211
rect 32825 -7245 32841 -7211
rect 32001 -7263 32035 -7247
rect 29896 -7271 30415 -7264
rect 20434 -7306 20602 -7288
rect 32379 -7295 32413 -7279
rect 30595 -7332 30651 -7315
rect 6998 -7386 7014 -7352
rect 7048 -7386 7064 -7352
rect 7116 -7386 7132 -7352
rect 7166 -7386 7182 -7352
rect 13552 -7381 13568 -7347
rect 13602 -7381 13618 -7347
rect 13670 -7381 13686 -7347
rect 13720 -7381 13736 -7347
rect 20201 -7393 20217 -7359
rect 20251 -7393 20267 -7359
rect 20319 -7393 20335 -7359
rect 20369 -7393 20385 -7359
rect 30595 -7366 30601 -7332
rect 30635 -7366 30651 -7332
rect 30595 -7383 30651 -7366
rect 30776 -7348 30810 -7332
rect 6955 -7436 6989 -7420
rect 6955 -7828 6989 -7812
rect 7073 -7436 7107 -7420
rect 7073 -7828 7107 -7812
rect 7191 -7436 7225 -7420
rect 13509 -7431 13543 -7415
rect 7191 -7828 7225 -7812
rect 7308 -7636 7342 -7620
rect 7308 -7828 7342 -7812
rect 7426 -7636 7460 -7620
rect 7426 -7828 7460 -7812
rect 13509 -7823 13543 -7807
rect 13627 -7431 13661 -7415
rect 13627 -7823 13661 -7807
rect 13745 -7431 13779 -7415
rect 20158 -7443 20192 -7427
rect 13745 -7823 13779 -7807
rect 13862 -7631 13896 -7615
rect 13862 -7823 13896 -7807
rect 13980 -7631 14014 -7615
rect 13980 -7823 14014 -7807
rect 20158 -7835 20192 -7819
rect 20276 -7443 20310 -7427
rect 20276 -7835 20310 -7819
rect 20394 -7443 20428 -7427
rect 20394 -7835 20428 -7819
rect 20511 -7643 20545 -7627
rect 20511 -7835 20545 -7819
rect 20629 -7643 20663 -7627
rect 28898 -7715 29066 -7699
rect 28898 -7785 28914 -7715
rect 29050 -7785 29066 -7715
rect 30894 -7348 30928 -7332
rect 30776 -7740 30810 -7724
rect 30893 -7724 30894 -7677
rect 31012 -7348 31046 -7332
rect 30928 -7724 30929 -7677
rect 28898 -7801 29066 -7785
rect 30893 -7782 30929 -7724
rect 31130 -7348 31164 -7332
rect 31012 -7740 31046 -7724
rect 31128 -7724 31130 -7677
rect 31128 -7782 31164 -7724
rect 31248 -7348 31282 -7332
rect 31248 -7740 31282 -7724
rect 31366 -7348 31400 -7332
rect 31484 -7348 31518 -7332
rect 31400 -7724 31402 -7678
rect 31366 -7782 31402 -7724
rect 31646 -7553 31716 -7549
rect 31646 -7644 31650 -7553
rect 31712 -7644 31716 -7553
rect 31646 -7649 31716 -7644
rect 31484 -7740 31518 -7724
rect 31661 -7782 31702 -7649
rect 32379 -7687 32413 -7671
rect 32497 -7295 32531 -7279
rect 32497 -7687 32531 -7671
rect 32615 -7295 32649 -7279
rect 32732 -7295 32766 -7279
rect 32732 -7487 32766 -7471
rect 32850 -7295 32884 -7279
rect 32850 -7487 32884 -7471
rect 32615 -7687 32649 -7671
rect 32422 -7755 32438 -7721
rect 32472 -7755 32488 -7721
rect 32540 -7755 32556 -7721
rect 32590 -7755 32606 -7721
rect 20629 -7835 20663 -7819
rect 30893 -7822 31702 -7782
rect 30912 -7823 31702 -7822
rect 7351 -7896 7367 -7862
rect 7401 -7896 7417 -7862
rect 13905 -7891 13921 -7857
rect 13955 -7891 13971 -7857
rect 20554 -7903 20570 -7869
rect 20604 -7903 20620 -7869
rect 29435 -7905 29705 -7871
rect 28609 -7955 28643 -7939
rect 7469 -8013 7485 -7979
rect 7519 -8013 7535 -7979
rect 14023 -8008 14039 -7974
rect 14073 -8008 14089 -7974
rect 20672 -8020 20688 -7986
rect 20722 -8020 20738 -7986
rect 6718 -8073 6752 -8057
rect 6718 -8265 6752 -8249
rect 6836 -8073 6870 -8057
rect 6836 -8265 6870 -8249
rect 6954 -8073 6988 -8057
rect 6954 -8265 6988 -8249
rect 7072 -8073 7106 -8057
rect 7072 -8265 7106 -8249
rect 7190 -8073 7224 -8057
rect 7190 -8265 7224 -8249
rect 7308 -8073 7342 -8057
rect 7308 -8265 7342 -8249
rect 7426 -8073 7460 -8057
rect 7426 -8265 7460 -8249
rect 7544 -8073 7578 -8057
rect 7544 -8299 7578 -8249
rect 7662 -8073 7696 -8057
rect 7662 -8265 7696 -8249
rect 7780 -8073 7814 -8057
rect 7780 -8299 7814 -8249
rect 13272 -8068 13306 -8052
rect 13272 -8260 13306 -8244
rect 13390 -8068 13424 -8052
rect 13390 -8260 13424 -8244
rect 13508 -8068 13542 -8052
rect 13508 -8260 13542 -8244
rect 13626 -8068 13660 -8052
rect 13626 -8260 13660 -8244
rect 13744 -8068 13778 -8052
rect 13744 -8260 13778 -8244
rect 13862 -8068 13896 -8052
rect 13862 -8260 13896 -8244
rect 13980 -8068 14014 -8052
rect 13980 -8260 14014 -8244
rect 14098 -8068 14132 -8052
rect 7544 -8333 7814 -8299
rect 14098 -8294 14132 -8244
rect 14216 -8068 14250 -8052
rect 14216 -8260 14250 -8244
rect 14334 -8068 14368 -8052
rect 14334 -8294 14368 -8244
rect 19921 -8080 19955 -8064
rect 19921 -8272 19955 -8256
rect 20039 -8080 20073 -8064
rect 20039 -8272 20073 -8256
rect 20157 -8080 20191 -8064
rect 20157 -8272 20191 -8256
rect 20275 -8080 20309 -8064
rect 20275 -8272 20309 -8256
rect 20393 -8080 20427 -8064
rect 20393 -8272 20427 -8256
rect 20511 -8080 20545 -8064
rect 20511 -8272 20545 -8256
rect 20629 -8080 20663 -8064
rect 20629 -8272 20663 -8256
rect 20747 -8080 20781 -8064
rect 14098 -8328 14368 -8294
rect 20747 -8306 20781 -8256
rect 20865 -8080 20899 -8064
rect 20865 -8272 20899 -8256
rect 20983 -8080 21017 -8064
rect 28609 -8147 28643 -8131
rect 28727 -7955 28761 -7939
rect 28727 -8147 28761 -8131
rect 28845 -7955 28879 -7939
rect 28845 -8147 28879 -8131
rect 28963 -7955 28997 -7939
rect 28963 -8147 28997 -8131
rect 29081 -7955 29115 -7939
rect 29081 -8147 29115 -8131
rect 29199 -7955 29233 -7939
rect 29199 -8147 29233 -8131
rect 29317 -7955 29351 -7939
rect 29317 -8147 29351 -8131
rect 29435 -7955 29469 -7905
rect 29435 -8147 29469 -8131
rect 29553 -7955 29587 -7939
rect 29553 -8147 29587 -8131
rect 29671 -7955 29705 -7905
rect 30790 -7912 30857 -7896
rect 30790 -7946 30806 -7912
rect 30840 -7946 30857 -7912
rect 30790 -7962 30857 -7946
rect 30621 -7979 30655 -7963
rect 30621 -8029 30655 -8013
rect 30967 -8064 31001 -7823
rect 32655 -7826 32823 -7808
rect 32655 -7882 32671 -7826
rect 32805 -7882 32823 -7826
rect 31437 -7912 31504 -7896
rect 32655 -7898 32823 -7882
rect 31437 -7946 31454 -7912
rect 31488 -7946 31504 -7912
rect 31437 -7962 31504 -7946
rect 31744 -7980 31778 -7964
rect 31056 -8030 31072 -7996
rect 31106 -8030 31122 -7996
rect 31174 -8029 31190 -7995
rect 31224 -8029 31240 -7995
rect 31744 -8030 31778 -8014
rect 29671 -8147 29705 -8131
rect 30474 -8080 30508 -8064
rect 29360 -8225 29376 -8191
rect 29410 -8225 29426 -8191
rect 20983 -8306 21017 -8256
rect 30474 -8272 30508 -8256
rect 30592 -8080 30626 -8064
rect 30592 -8272 30626 -8256
rect 30894 -8080 30928 -8064
rect 20747 -8340 21017 -8306
rect 29242 -8342 29258 -8308
rect 29292 -8342 29308 -8308
rect 28846 -8392 28880 -8376
rect 7007 -8419 7175 -8403
rect 7007 -8489 7023 -8419
rect 7159 -8489 7175 -8419
rect 7007 -8505 7175 -8489
rect 13561 -8414 13729 -8398
rect 13561 -8484 13577 -8414
rect 13713 -8484 13729 -8414
rect 13561 -8500 13729 -8484
rect 20210 -8426 20378 -8410
rect 20210 -8496 20226 -8426
rect 20362 -8496 20378 -8426
rect 20210 -8512 20378 -8496
rect 28846 -8784 28880 -8768
rect 28964 -8392 28998 -8376
rect 28964 -8784 28998 -8768
rect 29082 -8392 29116 -8376
rect 29199 -8392 29233 -8376
rect 29199 -8584 29233 -8568
rect 29317 -8392 29351 -8376
rect 30967 -8080 31046 -8064
rect 30967 -8110 31012 -8080
rect 30894 -8523 30929 -8456
rect 31012 -8472 31046 -8456
rect 31130 -8080 31164 -8064
rect 31130 -8472 31164 -8456
rect 31248 -8080 31282 -8064
rect 31366 -8080 31400 -8064
rect 31772 -8080 31806 -8064
rect 31772 -8272 31806 -8256
rect 31890 -8080 31924 -8064
rect 31890 -8272 31924 -8256
rect 31248 -8472 31282 -8456
rect 31365 -8523 31400 -8456
rect 30894 -8558 31400 -8523
rect 29317 -8584 29351 -8568
rect 31041 -8627 31283 -8615
rect 31041 -8729 31088 -8627
rect 31223 -8729 31283 -8627
rect 31041 -8746 31283 -8729
rect 29082 -8784 29116 -8768
rect 28889 -8852 28905 -8818
rect 28939 -8852 28955 -8818
rect 29007 -8852 29023 -8818
rect 29057 -8852 29073 -8818
rect 29122 -8923 29290 -8905
rect 29122 -8979 29138 -8923
rect 29272 -8979 29290 -8923
rect 29122 -8995 29290 -8979
rect 1594 -9238 1785 -9223
rect 1594 -9304 1619 -9238
rect 1763 -9304 1785 -9238
rect 1594 -9325 1785 -9304
<< viali >>
rect 7024 5807 7084 5869
rect 13573 5806 13633 5868
rect 20227 5827 20287 5889
rect 6683 5455 6717 5631
rect 6801 5455 6835 5631
rect 6919 5455 6953 5631
rect 7037 5455 7071 5631
rect 7155 5455 7189 5631
rect 7273 5455 7307 5631
rect 7391 5455 7425 5631
rect 7509 5455 7543 5631
rect 7627 5455 7661 5631
rect 7745 5455 7779 5631
rect 13232 5454 13266 5630
rect 13350 5454 13384 5630
rect 13468 5454 13502 5630
rect 13586 5454 13620 5630
rect 13704 5454 13738 5630
rect 13822 5454 13856 5630
rect 13940 5454 13974 5630
rect 14058 5454 14092 5630
rect 14176 5454 14210 5630
rect 14294 5454 14328 5630
rect 19886 5475 19920 5651
rect 20004 5475 20038 5651
rect 20122 5475 20156 5651
rect 20240 5475 20274 5651
rect 20358 5475 20392 5651
rect 20476 5475 20510 5651
rect 20594 5475 20628 5651
rect 20712 5475 20746 5651
rect 20830 5475 20864 5651
rect 20948 5475 20982 5651
rect 28880 5660 28940 5722
rect 30981 5783 31402 5817
rect 30981 5638 31044 5783
rect 31044 5638 31353 5783
rect 31353 5638 31402 5783
rect 30981 5617 31402 5638
rect 7450 5361 7484 5395
rect 13999 5360 14033 5394
rect 20653 5381 20687 5415
rect 28539 5308 28573 5484
rect 7332 5244 7366 5278
rect 13881 5243 13915 5277
rect 20535 5264 20569 5298
rect 28657 5308 28691 5484
rect 28775 5308 28809 5484
rect 28893 5308 28927 5484
rect 29011 5308 29045 5484
rect 29129 5308 29163 5484
rect 29247 5308 29281 5484
rect 29365 5308 29399 5484
rect 29483 5308 29517 5484
rect 29601 5308 29635 5484
rect 6920 4818 6954 5194
rect 7038 4818 7072 5194
rect 7156 4818 7190 5194
rect 7273 5018 7307 5194
rect 7391 5018 7425 5194
rect 13469 4817 13503 5193
rect 13587 4817 13621 5193
rect 13705 4817 13739 5193
rect 13822 5017 13856 5193
rect 13940 5017 13974 5193
rect 20123 4838 20157 5214
rect 20241 4838 20275 5214
rect 20359 4838 20393 5214
rect 20476 5038 20510 5214
rect 29306 5214 29340 5248
rect 20594 5038 20628 5214
rect 29188 5097 29222 5131
rect 6979 4734 7013 4768
rect 7097 4734 7131 4768
rect 13382 4722 13431 4768
rect 13528 4733 13562 4767
rect 13646 4733 13680 4767
rect 19989 4742 20050 4790
rect 20182 4754 20216 4788
rect 20300 4754 20334 4788
rect 7252 4611 7304 4657
rect -902 4466 -841 4516
rect 13801 4610 13853 4656
rect 6801 4289 6850 4343
rect 20091 4662 20136 4700
rect 20455 4631 20507 4677
rect 28776 4671 28810 5047
rect 28894 4671 28928 5047
rect 29012 4671 29046 5047
rect 29129 4871 29163 5047
rect 29247 4871 29281 5047
rect 30347 4903 30381 5079
rect 30465 4903 30499 5079
rect 30583 4903 30617 5079
rect 30701 4903 30735 5079
rect 30831 4903 30865 5279
rect 30949 4903 30983 5279
rect 31067 4903 31101 5279
rect 31185 4903 31219 5279
rect 31303 4903 31337 5279
rect 31421 4903 31455 5279
rect 31539 4903 31573 5279
rect 32481 5252 32541 5314
rect 31668 4903 31702 5079
rect 31786 4903 31820 5079
rect 31904 4903 31938 5079
rect 32022 4903 32056 5079
rect 32140 4900 32174 5076
rect 32258 4900 32292 5076
rect 32376 4900 32410 5076
rect 32494 4900 32528 5076
rect 32612 4900 32646 5076
rect 32730 4900 32764 5076
rect 32848 4900 32882 5076
rect 32966 4900 33000 5076
rect 33084 4900 33118 5076
rect 33202 4900 33236 5076
rect 32907 4806 32941 4840
rect 31999 4687 32033 4721
rect 32789 4689 32823 4723
rect 28835 4587 28869 4621
rect 28953 4587 28987 4621
rect 30326 4547 30406 4615
rect 30599 4568 30633 4602
rect 29108 4464 29160 4510
rect -749 3898 -692 3943
rect -922 2725 -809 2809
rect 360 3907 420 3969
rect 19 3555 53 3731
rect 137 3555 171 3731
rect 255 3555 289 3731
rect 373 3555 407 3731
rect 491 3555 525 3731
rect 609 3555 643 3731
rect 727 3555 761 3731
rect 845 3555 879 3731
rect 963 3555 997 3731
rect 1081 3555 1115 3731
rect 786 3461 820 3495
rect 668 3344 702 3378
rect -630 -5674 -528 -5593
rect -484 2911 -395 2987
rect 256 2918 290 3294
rect 374 2918 408 3294
rect 492 2918 526 3294
rect 609 3118 643 3294
rect 727 3118 761 3294
rect 315 2834 349 2868
rect 433 2834 467 2868
rect 10 2749 66 2793
rect 588 2711 640 2757
rect 352 1322 412 1384
rect 11 970 45 1146
rect 129 970 163 1146
rect 247 970 281 1146
rect 365 970 399 1146
rect 483 970 517 1146
rect 601 970 635 1146
rect 719 970 753 1146
rect 837 970 871 1146
rect 955 970 989 1146
rect 1073 970 1107 1146
rect 778 876 812 910
rect 660 759 694 793
rect 248 333 282 709
rect 366 333 400 709
rect 484 333 518 709
rect 601 533 635 709
rect 719 533 753 709
rect 307 249 341 283
rect 425 249 459 283
rect 580 126 632 172
rect 333 -1956 393 -1894
rect -8 -2308 26 -2132
rect 110 -2308 144 -2132
rect 228 -2308 262 -2132
rect 346 -2308 380 -2132
rect 464 -2308 498 -2132
rect 582 -2308 616 -2132
rect 700 -2308 734 -2132
rect 818 -2308 852 -2132
rect 936 -2308 970 -2132
rect 1054 -2308 1088 -2132
rect 759 -2402 793 -2368
rect 641 -2519 675 -2485
rect 229 -2945 263 -2569
rect 347 -2945 381 -2569
rect 465 -2945 499 -2569
rect 582 -2745 616 -2569
rect 700 -2745 734 -2569
rect 288 -3029 322 -2995
rect 406 -3029 440 -2995
rect -46 -3119 14 -3066
rect 561 -3152 613 -3106
rect 349 -4716 409 -4654
rect 8 -5068 42 -4892
rect 126 -5068 160 -4892
rect 244 -5068 278 -4892
rect 362 -5068 396 -4892
rect 480 -5068 514 -4892
rect 598 -5068 632 -4892
rect 716 -5068 750 -4892
rect 834 -5068 868 -4892
rect 952 -5068 986 -4892
rect 1070 -5068 1104 -4892
rect 775 -5162 809 -5128
rect 657 -5279 691 -5245
rect 245 -5705 279 -5329
rect 363 -5705 397 -5329
rect 481 -5705 515 -5329
rect 598 -5505 632 -5329
rect 716 -5505 750 -5329
rect 304 -5789 338 -5755
rect 422 -5789 456 -5755
rect 577 -5912 629 -5866
rect -510 -9026 -366 -8960
rect -925 -9171 -811 -9100
rect 3384 3878 3451 3879
rect 3384 3730 3450 3878
rect 3450 3730 3451 3878
rect 5866 3783 5932 3929
rect 5932 3783 5933 3929
rect 5866 3780 5933 3783
rect 5119 3678 5153 3712
rect 7008 3783 7012 3931
rect 7012 3783 7075 3931
rect 7008 3782 7075 3783
rect 6249 3684 6283 3718
rect 9933 3966 10000 3967
rect 9933 3818 9999 3966
rect 9999 3818 10000 3966
rect 12416 3871 12481 4018
rect 12481 3871 12483 4018
rect 12416 3869 12483 3871
rect 11668 3766 11702 3800
rect 13560 3871 13561 4020
rect 13561 3871 13627 4020
rect 12798 3772 12832 3806
rect 16586 3749 16653 3897
rect 16586 3748 16653 3749
rect 19067 3952 19134 3953
rect 19067 3804 19068 3952
rect 19068 3804 19134 3952
rect 11668 3648 11702 3682
rect 5119 3560 5153 3594
rect 6249 3564 6283 3598
rect 12798 3652 12832 3686
rect 2909 3288 2943 3464
rect 3027 3288 3061 3464
rect 3145 3288 3179 3464
rect 3263 3288 3297 3464
rect 3381 3288 3415 3464
rect 3499 3288 3533 3464
rect 3617 3288 3651 3464
rect 3735 3288 3769 3464
rect 3853 3288 3887 3464
rect 3971 3288 4005 3464
rect 3676 3194 3710 3228
rect 5234 3160 5268 3536
rect 5352 3160 5386 3536
rect 5470 3160 5504 3536
rect 5588 3160 5622 3536
rect 5706 3160 5740 3536
rect 5824 3160 5858 3536
rect 5942 3160 5976 3536
rect 6376 3164 6410 3540
rect 6494 3164 6528 3540
rect 6612 3164 6646 3540
rect 6730 3164 6764 3540
rect 6848 3164 6882 3540
rect 6966 3164 7000 3540
rect 7084 3164 7118 3540
rect 9458 3376 9492 3552
rect 9576 3376 9610 3552
rect 9694 3376 9728 3552
rect 9812 3376 9846 3552
rect 9930 3376 9964 3552
rect 10048 3376 10082 3552
rect 10166 3376 10200 3552
rect 10284 3376 10318 3552
rect 10402 3376 10436 3552
rect 10520 3376 10554 3552
rect 10225 3282 10259 3316
rect 11783 3248 11817 3624
rect 11901 3248 11935 3624
rect 12019 3248 12053 3624
rect 12137 3248 12171 3624
rect 12255 3248 12289 3624
rect 12373 3248 12407 3624
rect 12491 3248 12525 3624
rect 12925 3252 12959 3628
rect 13043 3252 13077 3628
rect 13161 3252 13195 3628
rect 13279 3252 13313 3628
rect 13397 3252 13431 3628
rect 13515 3252 13549 3628
rect 18322 3698 18356 3732
rect 20214 3803 20215 3952
rect 20215 3803 20281 3952
rect 19452 3704 19486 3738
rect 23206 3817 23211 3966
rect 23211 3817 23273 3966
rect 25690 3871 25693 4018
rect 25693 3871 25757 4018
rect 25690 3869 25757 3871
rect 24947 3766 24981 3800
rect 26839 4020 26906 4024
rect 26839 3875 26840 4020
rect 26840 3875 26906 4020
rect 26077 3772 26111 3806
rect 24947 3648 24981 3682
rect 13633 3252 13667 3628
rect 18322 3580 18356 3614
rect 19452 3584 19486 3618
rect 16112 3308 16146 3484
rect 16230 3308 16264 3484
rect 16348 3308 16382 3484
rect 16466 3308 16500 3484
rect 16584 3308 16618 3484
rect 16702 3308 16736 3484
rect 16820 3308 16854 3484
rect 16938 3308 16972 3484
rect 17056 3308 17090 3484
rect 17174 3308 17208 3484
rect 16879 3214 16913 3248
rect 10107 3165 10141 3199
rect 18437 3180 18471 3556
rect 18555 3180 18589 3556
rect 18673 3180 18707 3556
rect 18791 3180 18825 3556
rect 18909 3180 18943 3556
rect 19027 3180 19061 3556
rect 26077 3652 26111 3686
rect 19145 3180 19179 3556
rect 19579 3184 19613 3560
rect 19697 3184 19731 3560
rect 19815 3184 19849 3560
rect 19933 3184 19967 3560
rect 20051 3184 20085 3560
rect 20169 3184 20203 3560
rect 20287 3184 20321 3560
rect 22737 3376 22771 3552
rect 22855 3376 22889 3552
rect 22973 3376 23007 3552
rect 23091 3376 23125 3552
rect 23209 3376 23243 3552
rect 23327 3376 23361 3552
rect 23445 3376 23479 3552
rect 23563 3376 23597 3552
rect 23681 3376 23715 3552
rect 23799 3376 23833 3552
rect 23504 3282 23538 3316
rect 25062 3248 25096 3624
rect 25180 3248 25214 3624
rect 25298 3248 25332 3624
rect 25416 3248 25450 3624
rect 25534 3248 25568 3624
rect 25652 3248 25686 3624
rect 25770 3248 25804 3624
rect 26204 3252 26238 3628
rect 26322 3252 26356 3628
rect 26440 3252 26474 3628
rect 26558 3252 26592 3628
rect 26676 3252 26710 3628
rect 26794 3252 26828 3628
rect 26912 3252 26946 3628
rect 23386 3165 23420 3199
rect 3558 3077 3592 3111
rect 3146 2651 3180 3027
rect 3264 2651 3298 3027
rect 3382 2651 3416 3027
rect 3499 2851 3533 3027
rect 3617 2851 3651 3027
rect 5439 2804 5473 2838
rect 6581 2808 6615 2842
rect 3725 2623 3874 2690
rect 3205 2567 3239 2601
rect 3323 2567 3357 2601
rect 5144 2577 5178 2753
rect 5262 2577 5296 2753
rect 5380 2577 5414 2753
rect 5498 2577 5532 2753
rect 5663 2577 5697 2753
rect 5781 2577 5815 2753
rect 5899 2577 5933 2753
rect 6017 2577 6051 2753
rect 6286 2581 6320 2757
rect 6404 2581 6438 2757
rect 6522 2581 6556 2757
rect 6640 2581 6674 2757
rect 6805 2581 6839 2757
rect 6923 2581 6957 2757
rect 7041 2581 7075 2757
rect 7159 2581 7193 2757
rect 9695 2739 9729 3115
rect 9813 2739 9847 3115
rect 9931 2739 9965 3115
rect 10048 2939 10082 3115
rect 10166 2939 10200 3115
rect 16761 3097 16795 3131
rect 11988 2892 12022 2926
rect 13130 2896 13164 2930
rect 10271 2705 10420 2772
rect 9754 2655 9788 2689
rect 9872 2655 9906 2689
rect 11693 2665 11727 2841
rect 11811 2665 11845 2841
rect 11929 2665 11963 2841
rect 12047 2665 12081 2841
rect 12212 2665 12246 2841
rect 12330 2665 12364 2841
rect 12448 2665 12482 2841
rect 12566 2665 12600 2841
rect 12835 2669 12869 2845
rect 12953 2669 12987 2845
rect 13071 2669 13105 2845
rect 13189 2669 13223 2845
rect 13354 2669 13388 2845
rect 13472 2669 13506 2845
rect 13590 2669 13624 2845
rect 13708 2669 13742 2845
rect 16349 2671 16383 3047
rect 16467 2671 16501 3047
rect 16585 2671 16619 3047
rect 16702 2871 16736 3047
rect 16820 2871 16854 3047
rect 18642 2824 18676 2858
rect 19784 2828 19818 2862
rect 16921 2639 17070 2706
rect 16408 2587 16442 2621
rect 16526 2587 16560 2621
rect 18347 2597 18381 2773
rect 18465 2597 18499 2773
rect 18583 2597 18617 2773
rect 18701 2597 18735 2773
rect 18866 2597 18900 2773
rect 18984 2597 19018 2773
rect 19102 2597 19136 2773
rect 19220 2597 19254 2773
rect 19489 2601 19523 2777
rect 19607 2601 19641 2777
rect 19725 2601 19759 2777
rect 19843 2601 19877 2777
rect 20008 2601 20042 2777
rect 20126 2601 20160 2777
rect 20244 2601 20278 2777
rect 20362 2601 20396 2777
rect 22974 2739 23008 3115
rect 23092 2739 23126 3115
rect 23210 2739 23244 3115
rect 23327 2939 23361 3115
rect 23445 2939 23479 3115
rect 28875 3089 28935 3151
rect 25267 2892 25301 2926
rect 26409 2896 26443 2930
rect 23553 2715 23702 2782
rect 23033 2655 23067 2689
rect 23151 2655 23185 2689
rect 24972 2665 25006 2841
rect 25090 2665 25124 2841
rect 25208 2665 25242 2841
rect 25326 2665 25360 2841
rect 25491 2665 25525 2841
rect 25609 2665 25643 2841
rect 25727 2665 25761 2841
rect 25845 2665 25879 2841
rect 26114 2669 26148 2845
rect 26232 2669 26266 2845
rect 26350 2669 26384 2845
rect 26468 2669 26502 2845
rect 26633 2669 26667 2845
rect 26751 2669 26785 2845
rect 26869 2669 26903 2845
rect 26987 2669 27021 2845
rect 28534 2737 28568 2913
rect 28652 2737 28686 2913
rect 28770 2737 28804 2913
rect 28888 2737 28922 2913
rect 29006 2737 29040 2913
rect 29124 2737 29158 2913
rect 29242 2737 29276 2913
rect 29360 2737 29394 2913
rect 29478 2737 29512 2913
rect 29596 2737 29630 2913
rect 29301 2643 29335 2677
rect 29183 2526 29217 2560
rect 3396 2079 3397 2228
rect 3397 2079 3463 2228
rect 5211 2170 5278 2319
rect 6349 2172 6416 2321
rect 9947 2167 10013 2315
rect 10013 2167 10014 2315
rect 9947 2166 10014 2167
rect 11756 2266 11823 2415
rect 12895 2258 12962 2407
rect 16601 2248 16668 2249
rect 16601 2100 16667 2248
rect 16667 2100 16668 2248
rect 18409 2194 18476 2343
rect 19555 2197 19622 2346
rect 23229 2167 23292 2315
rect 23292 2167 23296 2315
rect 23229 2166 23296 2167
rect 25030 2255 25097 2402
rect 25030 2253 25097 2255
rect 26173 2255 26240 2404
rect 2923 1638 2957 1814
rect 3041 1638 3075 1814
rect 3159 1638 3193 1814
rect 3277 1638 3311 1814
rect 3395 1638 3429 1814
rect 3513 1638 3547 1814
rect 3631 1638 3665 1814
rect 3749 1638 3783 1814
rect 3867 1638 3901 1814
rect 3985 1638 4019 1814
rect 7108 1885 7175 1886
rect 7108 1737 7175 1885
rect 9472 1726 9506 1902
rect 9590 1726 9624 1902
rect 9708 1726 9742 1902
rect 9826 1726 9860 1902
rect 9944 1726 9978 1902
rect 10062 1726 10096 1902
rect 10180 1726 10214 1902
rect 10298 1726 10332 1902
rect 10416 1726 10450 1902
rect 10534 1726 10568 1902
rect 28771 2100 28805 2476
rect 28889 2100 28923 2476
rect 29007 2100 29041 2476
rect 29124 2300 29158 2476
rect 29242 2300 29276 2476
rect 13662 1824 13724 1973
rect 13724 1824 13729 1973
rect 10239 1632 10273 1666
rect 16126 1658 16160 1834
rect 16244 1658 16278 1834
rect 16362 1658 16396 1834
rect 16480 1658 16514 1834
rect 16598 1658 16632 1834
rect 16716 1658 16750 1834
rect 16834 1658 16868 1834
rect 16952 1658 16986 1834
rect 17070 1658 17104 1834
rect 17188 1658 17222 1834
rect 20308 1756 20311 1901
rect 20311 1756 20375 1901
rect 20308 1752 20375 1756
rect 22751 1726 22785 1902
rect 22869 1726 22903 1902
rect 22987 1726 23021 1902
rect 23105 1726 23139 1902
rect 23223 1726 23257 1902
rect 23341 1726 23375 1902
rect 23459 1726 23493 1902
rect 23577 1726 23611 1902
rect 23695 1726 23729 1902
rect 23813 1726 23847 1902
rect 28830 2016 28864 2050
rect 28948 2016 28982 2050
rect 26936 1824 27003 1970
rect 26936 1821 27003 1824
rect 29103 1893 29155 1939
rect 23518 1632 23552 1666
rect 3690 1544 3724 1578
rect 10121 1515 10155 1549
rect 3572 1427 3606 1461
rect 2121 898 2239 1008
rect 3160 1001 3194 1377
rect 3278 1001 3312 1377
rect 3396 1001 3430 1377
rect 3513 1201 3547 1377
rect 3631 1201 3665 1377
rect 3740 973 3889 1040
rect 4387 1021 4421 1197
rect 4505 1021 4539 1197
rect 4623 1021 4657 1197
rect 4741 1021 4775 1197
rect 4871 1021 4905 1397
rect 4989 1021 5023 1397
rect 5107 1021 5141 1397
rect 5225 1021 5259 1397
rect 5343 1021 5377 1397
rect 5461 1021 5495 1397
rect 5579 1021 5613 1397
rect 5708 1021 5742 1197
rect 5826 1021 5860 1197
rect 5944 1021 5978 1197
rect 6062 1021 6096 1197
rect 6285 1021 6319 1197
rect 6403 1021 6437 1197
rect 6521 1021 6555 1197
rect 6639 1021 6673 1197
rect 6769 1021 6803 1397
rect 6887 1021 6921 1397
rect 7005 1021 7039 1397
rect 7123 1021 7157 1397
rect 7241 1021 7275 1397
rect 7359 1021 7393 1397
rect 7477 1021 7511 1397
rect 7606 1021 7640 1197
rect 7724 1021 7758 1197
rect 7842 1021 7876 1197
rect 7960 1021 7994 1197
rect 9709 1089 9743 1465
rect 9827 1089 9861 1465
rect 9945 1089 9979 1465
rect 10062 1289 10096 1465
rect 10180 1289 10214 1465
rect 10289 1055 10438 1122
rect 10936 1109 10970 1285
rect 11054 1109 11088 1285
rect 11172 1109 11206 1285
rect 11290 1109 11324 1285
rect 11420 1109 11454 1485
rect 11538 1109 11572 1485
rect 11656 1109 11690 1485
rect 11774 1109 11808 1485
rect 11892 1109 11926 1485
rect 16893 1564 16927 1598
rect 12010 1109 12044 1485
rect 12128 1109 12162 1485
rect 12257 1109 12291 1285
rect 12375 1109 12409 1285
rect 12493 1109 12527 1285
rect 12611 1109 12645 1285
rect 12834 1109 12868 1285
rect 12952 1109 12986 1285
rect 13070 1109 13104 1285
rect 13188 1109 13222 1285
rect 13318 1109 13352 1485
rect 13436 1109 13470 1485
rect 13554 1109 13588 1485
rect 13672 1109 13706 1485
rect 13790 1109 13824 1485
rect 23400 1515 23434 1549
rect 13908 1109 13942 1485
rect 14026 1109 14060 1485
rect 16775 1447 16809 1481
rect 14155 1109 14189 1285
rect 14273 1109 14307 1285
rect 14391 1109 14425 1285
rect 14509 1109 14543 1285
rect 9768 1005 9802 1039
rect 9886 1005 9920 1039
rect 3219 917 3253 951
rect 3337 917 3371 951
rect 15323 920 15462 1037
rect 16363 1021 16397 1397
rect 16481 1021 16515 1397
rect 16599 1021 16633 1397
rect 16716 1221 16750 1397
rect 16834 1221 16868 1397
rect 16938 988 17087 1055
rect 17590 1041 17624 1217
rect 17708 1041 17742 1217
rect 17826 1041 17860 1217
rect 17944 1041 17978 1217
rect 18074 1041 18108 1417
rect 18192 1041 18226 1417
rect 18310 1041 18344 1417
rect 18428 1041 18462 1417
rect 18546 1041 18580 1417
rect 18664 1041 18698 1417
rect 18782 1041 18816 1417
rect 18911 1041 18945 1217
rect 19029 1041 19063 1217
rect 19147 1041 19181 1217
rect 19265 1041 19299 1217
rect 19488 1041 19522 1217
rect 19606 1041 19640 1217
rect 19724 1041 19758 1217
rect 19842 1041 19876 1217
rect 19972 1041 20006 1417
rect 20090 1041 20124 1417
rect 20208 1041 20242 1417
rect 20326 1041 20360 1417
rect 20444 1041 20478 1417
rect 20562 1041 20596 1417
rect 20680 1041 20714 1417
rect 20809 1041 20843 1217
rect 20927 1041 20961 1217
rect 21045 1041 21079 1217
rect 21163 1041 21197 1217
rect 22988 1089 23022 1465
rect 23106 1089 23140 1465
rect 23224 1089 23258 1465
rect 23341 1289 23375 1465
rect 23459 1289 23493 1465
rect 23558 1054 23707 1121
rect 24215 1109 24249 1285
rect 24333 1109 24367 1285
rect 24451 1109 24485 1285
rect 24569 1109 24603 1285
rect 24699 1109 24733 1485
rect 24817 1109 24851 1485
rect 24935 1109 24969 1485
rect 25053 1109 25087 1485
rect 25171 1109 25205 1485
rect 25289 1109 25323 1485
rect 25407 1109 25441 1485
rect 25536 1109 25570 1285
rect 25654 1109 25688 1285
rect 25772 1109 25806 1285
rect 25890 1109 25924 1285
rect 26113 1109 26147 1285
rect 26231 1109 26265 1285
rect 26349 1109 26383 1285
rect 26467 1109 26501 1285
rect 26597 1109 26631 1485
rect 26715 1109 26749 1485
rect 26833 1109 26867 1485
rect 26951 1109 26985 1485
rect 27069 1109 27103 1485
rect 27187 1109 27221 1485
rect 27305 1109 27339 1485
rect 27434 1109 27468 1285
rect 27552 1109 27586 1285
rect 27670 1109 27704 1285
rect 27788 1109 27822 1285
rect 23047 1005 23081 1039
rect 23165 1005 23199 1039
rect 16422 937 16456 971
rect 16540 937 16574 971
rect 12400 837 12434 871
rect 14507 816 14541 850
rect 5851 749 5885 783
rect 7958 728 7992 762
rect 3394 475 3459 622
rect 3459 475 3461 622
rect 3394 473 3461 475
rect 4814 328 4848 704
rect 4932 328 4966 704
rect 2918 34 2952 210
rect 3036 34 3070 210
rect 3154 34 3188 210
rect 3272 34 3306 210
rect 3390 34 3424 210
rect 3508 34 3542 210
rect 3626 34 3660 210
rect 3744 34 3778 210
rect 3862 34 3896 210
rect 5050 328 5084 704
rect 5168 328 5202 704
rect 5286 328 5320 704
rect 5404 328 5438 704
rect 5522 328 5556 704
rect 6712 328 6746 704
rect 6830 328 6864 704
rect 6948 328 6982 704
rect 7066 328 7100 704
rect 7184 328 7218 704
rect 7302 328 7336 704
rect 7420 328 7454 704
rect 9939 712 10006 715
rect 9939 566 9941 712
rect 9941 566 10006 712
rect 11363 416 11397 792
rect 11481 416 11515 792
rect 3980 34 4014 210
rect 4844 106 4878 140
rect 4659 39 4693 73
rect 5492 106 5526 140
rect 6742 106 6776 140
rect 5110 22 5144 56
rect 5228 23 5262 57
rect 5782 38 5816 72
rect 6557 39 6591 73
rect 7388 107 7422 141
rect 7008 22 7042 56
rect 7126 23 7160 57
rect 7680 38 7714 72
rect 3685 -60 3719 -26
rect 3567 -177 3601 -143
rect 4512 -204 4546 -28
rect 3155 -603 3189 -227
rect 3273 -603 3307 -227
rect 3391 -603 3425 -227
rect 3508 -403 3542 -227
rect 4630 -204 4664 -28
rect 3626 -403 3660 -227
rect 4932 -404 4966 -28
rect 5050 -404 5084 -28
rect 5168 -404 5202 -28
rect 5286 -404 5320 -28
rect 5404 -404 5438 -28
rect 5810 -204 5844 -28
rect 5928 -204 5962 -28
rect 6410 -204 6444 -28
rect 6528 -204 6562 -28
rect 6830 -404 6864 -28
rect 6948 -404 6982 -28
rect 7066 -404 7100 -28
rect 7184 -404 7218 -28
rect 7302 -404 7336 -28
rect 7708 -204 7742 -28
rect 7826 -204 7860 -28
rect 3738 -635 3887 -568
rect 3214 -687 3248 -653
rect 3332 -687 3366 -653
rect 5151 -870 5218 -721
rect 9467 122 9501 298
rect 9585 122 9619 298
rect 9703 122 9737 298
rect 9821 122 9855 298
rect 9939 122 9973 298
rect 10057 122 10091 298
rect 10175 122 10209 298
rect 10293 122 10327 298
rect 10411 122 10445 298
rect 11599 416 11633 792
rect 11717 416 11751 792
rect 11835 416 11869 792
rect 11953 416 11987 792
rect 12071 416 12105 792
rect 13261 416 13295 792
rect 13379 416 13413 792
rect 13497 416 13531 792
rect 13615 416 13649 792
rect 13733 416 13767 792
rect 13851 416 13885 792
rect 13969 416 14003 792
rect 10529 122 10563 298
rect 11393 194 11427 228
rect 11208 127 11242 161
rect 12041 194 12075 228
rect 13291 194 13325 228
rect 11659 110 11693 144
rect 11777 111 11811 145
rect 12331 126 12365 160
rect 13106 127 13140 161
rect 14630 289 14762 387
rect 13937 195 13971 229
rect 13557 110 13591 144
rect 13675 111 13709 145
rect 14229 126 14263 160
rect 10234 28 10268 62
rect 10116 -89 10150 -55
rect 11061 -116 11095 60
rect 9704 -515 9738 -139
rect 9822 -515 9856 -139
rect 9940 -515 9974 -139
rect 10057 -315 10091 -139
rect 11179 -116 11213 60
rect 10175 -315 10209 -139
rect 11481 -316 11515 60
rect 11599 -316 11633 60
rect 11717 -316 11751 60
rect 11835 -316 11869 60
rect 11953 -316 11987 60
rect 12359 -116 12393 60
rect 12477 -116 12511 60
rect 12959 -116 12993 60
rect 13077 -116 13111 60
rect 13379 -316 13413 60
rect 13497 -316 13531 60
rect 13615 -316 13649 60
rect 13733 -316 13767 60
rect 13851 -316 13885 60
rect 14257 -116 14291 60
rect 14375 -116 14409 60
rect 10286 -546 10435 -479
rect 9763 -599 9797 -565
rect 9881 -599 9915 -565
rect 11700 -785 11767 -636
rect 25679 837 25713 871
rect 27786 816 27820 850
rect 19054 769 19088 803
rect 21161 748 21195 782
rect 16596 644 16663 646
rect 16596 497 16662 644
rect 16662 497 16663 644
rect 18017 348 18051 724
rect 18135 348 18169 724
rect 16121 54 16155 230
rect 16239 54 16273 230
rect 16357 54 16391 230
rect 16475 54 16509 230
rect 16593 54 16627 230
rect 16711 54 16745 230
rect 16829 54 16863 230
rect 16947 54 16981 230
rect 17065 54 17099 230
rect 18253 348 18287 724
rect 18371 348 18405 724
rect 18489 348 18523 724
rect 18607 348 18641 724
rect 18725 348 18759 724
rect 19915 348 19949 724
rect 20033 348 20067 724
rect 20151 348 20185 724
rect 20269 348 20303 724
rect 20387 348 20421 724
rect 20505 348 20539 724
rect 20623 348 20657 724
rect 23221 563 23287 707
rect 23287 563 23288 707
rect 23221 558 23288 563
rect 24642 416 24676 792
rect 24760 416 24794 792
rect 17183 54 17217 230
rect 18047 126 18081 160
rect 17862 59 17896 93
rect 18695 126 18729 160
rect 19945 126 19979 160
rect 18313 42 18347 76
rect 18431 43 18465 77
rect 18985 58 19019 92
rect 19760 59 19794 93
rect 21745 218 21841 318
rect 20591 127 20625 161
rect 22746 122 22780 298
rect 22864 122 22898 298
rect 22982 122 23016 298
rect 23100 122 23134 298
rect 23218 122 23252 298
rect 23336 122 23370 298
rect 23454 122 23488 298
rect 23572 122 23606 298
rect 23690 122 23724 298
rect 24878 416 24912 792
rect 24996 416 25030 792
rect 25114 416 25148 792
rect 25232 416 25266 792
rect 25350 416 25384 792
rect 26540 416 26574 792
rect 26658 416 26692 792
rect 26776 416 26810 792
rect 26894 416 26928 792
rect 27012 416 27046 792
rect 27130 416 27164 792
rect 27248 416 27282 792
rect 23808 122 23842 298
rect 24672 194 24706 228
rect 24487 127 24521 161
rect 20211 42 20245 76
rect 20329 43 20363 77
rect 20883 58 20917 92
rect 25320 194 25354 228
rect 26570 194 26604 228
rect 24938 110 24972 144
rect 25056 111 25090 145
rect 25610 126 25644 160
rect 26385 127 26419 161
rect 27909 289 28041 387
rect 27216 195 27250 229
rect 26836 110 26870 144
rect 26954 111 26988 145
rect 27508 126 27542 160
rect 23513 28 23547 62
rect 16888 -40 16922 -6
rect 16770 -157 16804 -123
rect 17715 -184 17749 -8
rect 16358 -583 16392 -207
rect 16476 -583 16510 -207
rect 16594 -583 16628 -207
rect 16711 -383 16745 -207
rect 17833 -184 17867 -8
rect 16829 -383 16863 -207
rect 18135 -384 18169 -8
rect 18253 -384 18287 -8
rect 18371 -384 18405 -8
rect 18489 -384 18523 -8
rect 18607 -384 18641 -8
rect 19013 -184 19047 -8
rect 19131 -184 19165 -8
rect 19613 -184 19647 -8
rect 19731 -184 19765 -8
rect 20033 -384 20067 -8
rect 20151 -384 20185 -8
rect 20269 -384 20303 -8
rect 20387 -384 20421 -8
rect 20505 -384 20539 -8
rect 20911 -184 20945 -8
rect 21029 -184 21063 -8
rect 23395 -89 23429 -55
rect 24340 -116 24374 60
rect 22983 -515 23017 -139
rect 23101 -515 23135 -139
rect 23219 -515 23253 -139
rect 23336 -315 23370 -139
rect 24458 -116 24492 60
rect 23454 -315 23488 -139
rect 24760 -316 24794 60
rect 24878 -316 24912 60
rect 24996 -316 25030 60
rect 25114 -316 25148 60
rect 25232 -316 25266 60
rect 25638 -116 25672 60
rect 25756 -116 25790 60
rect 26238 -116 26272 60
rect 26356 -116 26390 60
rect 26658 -316 26692 60
rect 26776 -316 26810 60
rect 26894 -316 26928 60
rect 27012 -316 27046 60
rect 27130 -316 27164 60
rect 27536 -116 27570 60
rect 27654 -116 27688 60
rect 28875 56 28935 118
rect 28534 -296 28568 -120
rect 28652 -296 28686 -120
rect 28770 -296 28804 -120
rect 28888 -296 28922 -120
rect 29006 -296 29040 -120
rect 29124 -296 29158 -120
rect 29242 -296 29276 -120
rect 29360 -296 29394 -120
rect 29478 -296 29512 -120
rect 29596 -296 29630 -120
rect 29301 -390 29335 -356
rect 16940 -617 17089 -550
rect 23564 -551 23713 -484
rect 29183 -507 29217 -473
rect 23042 -599 23076 -565
rect 23160 -599 23194 -565
rect 16417 -667 16451 -633
rect 16535 -667 16569 -633
rect 18349 -851 18416 -702
rect 24980 -785 25047 -636
rect 28771 -933 28805 -557
rect 28889 -933 28923 -557
rect 29007 -933 29041 -557
rect 29124 -733 29158 -557
rect 29242 -733 29276 -557
rect 15302 -1096 15372 -1028
rect 21285 -1102 21391 -1003
rect 22394 -1102 22500 -1003
rect 28830 -1017 28864 -983
rect 28948 -1017 28982 -983
rect 29103 -1140 29155 -1094
rect 30774 4210 30808 4586
rect 30892 4210 30926 4586
rect 31010 4210 31044 4586
rect 31128 4210 31162 4586
rect 31246 4210 31280 4586
rect 31364 4210 31398 4586
rect 31482 4210 31516 4586
rect 31648 4290 31710 4381
rect 32377 4263 32411 4639
rect 32495 4263 32529 4639
rect 32613 4263 32647 4639
rect 32730 4463 32764 4639
rect 32848 4463 32882 4639
rect 32436 4179 32470 4213
rect 32554 4179 32588 4213
rect 30804 3988 30838 4022
rect 30619 3921 30653 3955
rect 32709 4056 32761 4102
rect 31452 3988 31486 4022
rect 31070 3904 31104 3938
rect 31188 3905 31222 3939
rect 31742 3920 31776 3954
rect 30472 3678 30506 3854
rect 30590 3678 30624 3854
rect 30892 3478 30926 3854
rect 31010 3478 31044 3854
rect 31128 3478 31162 3854
rect 31246 3478 31280 3854
rect 31364 3478 31398 3854
rect 31770 3678 31804 3854
rect 31888 3678 31922 3854
rect 31086 3205 31221 3307
rect 30983 1692 31404 1726
rect 30983 1547 31046 1692
rect 31046 1547 31355 1692
rect 31355 1547 31404 1692
rect 30983 1526 31404 1547
rect 30349 812 30383 988
rect 30467 812 30501 988
rect 30585 812 30619 988
rect 30703 812 30737 988
rect 30833 812 30867 1188
rect 30951 812 30985 1188
rect 31069 812 31103 1188
rect 31187 812 31221 1188
rect 31305 812 31339 1188
rect 31423 812 31457 1188
rect 31541 812 31575 1188
rect 32483 1161 32543 1223
rect 31670 812 31704 988
rect 31788 812 31822 988
rect 31906 812 31940 988
rect 32024 812 32058 988
rect 32142 809 32176 985
rect 32260 809 32294 985
rect 32378 809 32412 985
rect 32496 809 32530 985
rect 32614 809 32648 985
rect 32732 809 32766 985
rect 32850 809 32884 985
rect 32968 809 33002 985
rect 33086 809 33120 985
rect 33204 809 33238 985
rect 32909 715 32943 749
rect 32001 596 32035 630
rect 32791 598 32825 632
rect 30601 477 30635 511
rect 30776 119 30810 495
rect 30894 119 30928 495
rect 31012 119 31046 495
rect 31130 119 31164 495
rect 31248 119 31282 495
rect 31366 119 31400 495
rect 31484 119 31518 495
rect 31650 199 31712 290
rect 32379 172 32413 548
rect 32497 172 32531 548
rect 32615 172 32649 548
rect 32732 372 32766 548
rect 32850 372 32884 548
rect 33097 467 33224 538
rect 32438 88 32472 122
rect 32556 88 32590 122
rect 30806 -103 30840 -69
rect 30621 -170 30655 -136
rect 32711 -35 32763 11
rect 31454 -103 31488 -69
rect 31072 -187 31106 -153
rect 31190 -186 31224 -152
rect 31744 -171 31778 -137
rect 30474 -413 30508 -237
rect 30592 -413 30626 -237
rect 30894 -613 30928 -237
rect 31012 -613 31046 -237
rect 31130 -613 31164 -237
rect 31248 -613 31282 -237
rect 31366 -613 31400 -237
rect 31772 -413 31806 -237
rect 31890 -413 31924 -237
rect 31088 -886 31223 -784
rect 3372 -1902 3439 -1901
rect 3372 -2050 3375 -1902
rect 3375 -2050 3439 -1902
rect 5852 -1848 5919 -1846
rect 5852 -1995 5857 -1848
rect 5857 -1995 5919 -1848
rect 5111 -2102 5145 -2068
rect 7008 -1997 7071 -1849
rect 7071 -1997 7075 -1849
rect 7008 -1998 7075 -1997
rect 6241 -2096 6275 -2062
rect 9927 -1904 9994 -1903
rect 9927 -2052 9993 -1904
rect 9993 -2052 9994 -1904
rect 12408 -1999 12475 -1850
rect 11662 -2104 11696 -2070
rect 13556 -1999 13622 -1850
rect 13622 -1999 13623 -1850
rect 12792 -2098 12826 -2064
rect 15301 -1913 15371 -1845
rect 5111 -2220 5145 -2186
rect 6241 -2216 6275 -2182
rect 2901 -2492 2935 -2316
rect 3019 -2492 3053 -2316
rect 3137 -2492 3171 -2316
rect 3255 -2492 3289 -2316
rect 3373 -2492 3407 -2316
rect 3491 -2492 3525 -2316
rect 3609 -2492 3643 -2316
rect 3727 -2492 3761 -2316
rect 3845 -2492 3879 -2316
rect 3963 -2492 3997 -2316
rect 3668 -2586 3702 -2552
rect 5226 -2620 5260 -2244
rect 5344 -2620 5378 -2244
rect 5462 -2620 5496 -2244
rect 5580 -2620 5614 -2244
rect 5698 -2620 5732 -2244
rect 5816 -2620 5850 -2244
rect 11662 -2222 11696 -2188
rect 5934 -2620 5968 -2244
rect 6368 -2616 6402 -2240
rect 6486 -2616 6520 -2240
rect 6604 -2616 6638 -2240
rect 6722 -2616 6756 -2240
rect 6840 -2616 6874 -2240
rect 6958 -2616 6992 -2240
rect 7076 -2616 7110 -2240
rect 12792 -2218 12826 -2184
rect 9452 -2494 9486 -2318
rect 9570 -2494 9604 -2318
rect 9688 -2494 9722 -2318
rect 9806 -2494 9840 -2318
rect 9924 -2494 9958 -2318
rect 10042 -2494 10076 -2318
rect 10160 -2494 10194 -2318
rect 10278 -2494 10312 -2318
rect 10396 -2494 10430 -2318
rect 10514 -2494 10548 -2318
rect 10219 -2588 10253 -2554
rect 11777 -2622 11811 -2246
rect 11895 -2622 11929 -2246
rect 12013 -2622 12047 -2246
rect 12131 -2622 12165 -2246
rect 12249 -2622 12283 -2246
rect 12367 -2622 12401 -2246
rect 12485 -2622 12519 -2246
rect 12919 -2618 12953 -2242
rect 13037 -2618 13071 -2242
rect 13155 -2618 13189 -2242
rect 13273 -2618 13307 -2242
rect 13391 -2618 13425 -2242
rect 13509 -2618 13543 -2242
rect 13627 -2618 13661 -2242
rect 16578 -2052 16581 -1906
rect 16581 -2052 16645 -1906
rect 16578 -2055 16645 -2052
rect 19063 -1849 19130 -1846
rect 19063 -1995 19130 -1849
rect 18317 -2103 18351 -2069
rect 20212 -1998 20277 -1849
rect 20277 -1998 20279 -1849
rect 19447 -2097 19481 -2063
rect 23202 -1902 23269 -1901
rect 23202 -2050 23203 -1902
rect 23203 -2050 23269 -1902
rect 25681 -1997 25685 -1853
rect 25685 -1997 25748 -1853
rect 25681 -2002 25748 -1997
rect 24939 -2102 24973 -2068
rect 26829 -1848 26896 -1847
rect 26829 -1996 26832 -1848
rect 26832 -1996 26896 -1848
rect 28946 -1864 29006 -1802
rect 26069 -2096 26103 -2062
rect 30983 -1803 31404 -1769
rect 30983 -1948 31046 -1803
rect 31046 -1948 31355 -1803
rect 31355 -1948 31404 -1803
rect 30983 -1969 31404 -1948
rect 18317 -2221 18351 -2187
rect 19447 -2217 19481 -2183
rect 3550 -2703 3584 -2669
rect 10101 -2705 10135 -2671
rect 3138 -3129 3172 -2753
rect 3256 -3129 3290 -2753
rect 3374 -3129 3408 -2753
rect 3491 -2929 3525 -2753
rect 3609 -2929 3643 -2753
rect 5431 -2976 5465 -2942
rect 6573 -2972 6607 -2938
rect 3715 -3164 3864 -3097
rect 3197 -3213 3231 -3179
rect 3315 -3213 3349 -3179
rect 5136 -3203 5170 -3027
rect 5254 -3203 5288 -3027
rect 5372 -3203 5406 -3027
rect 5490 -3203 5524 -3027
rect 5655 -3203 5689 -3027
rect 5773 -3203 5807 -3027
rect 5891 -3203 5925 -3027
rect 6009 -3203 6043 -3027
rect 6278 -3199 6312 -3023
rect 6396 -3199 6430 -3023
rect 6514 -3199 6548 -3023
rect 6632 -3199 6666 -3023
rect 6797 -3199 6831 -3023
rect 6915 -3199 6949 -3023
rect 7033 -3199 7067 -3023
rect 7151 -3199 7185 -3023
rect 9689 -3131 9723 -2755
rect 9807 -3131 9841 -2755
rect 9925 -3131 9959 -2755
rect 10042 -2931 10076 -2755
rect 10160 -2931 10194 -2755
rect 11982 -2978 12016 -2944
rect 13124 -2974 13158 -2940
rect 10265 -3170 10414 -3103
rect 9748 -3215 9782 -3181
rect 9866 -3215 9900 -3181
rect 11687 -3205 11721 -3029
rect 11805 -3205 11839 -3029
rect 11923 -3205 11957 -3029
rect 12041 -3205 12075 -3029
rect 12206 -3205 12240 -3029
rect 12324 -3205 12358 -3029
rect 12442 -3205 12476 -3029
rect 12560 -3205 12594 -3029
rect 12829 -3201 12863 -3025
rect 12947 -3201 12981 -3025
rect 13065 -3201 13099 -3025
rect 13183 -3201 13217 -3025
rect 13348 -3201 13382 -3025
rect 13466 -3201 13500 -3025
rect 13584 -3201 13618 -3025
rect 13702 -3201 13736 -3025
rect 3393 -3701 3456 -3554
rect 3456 -3701 3460 -3554
rect 3393 -3703 3460 -3701
rect 5192 -3607 5259 -3458
rect 6345 -3612 6412 -3463
rect 9938 -3554 10005 -3547
rect 9938 -3696 9940 -3554
rect 9940 -3696 10005 -3554
rect 11750 -3610 11817 -3461
rect 12891 -3617 12958 -3472
rect 12891 -3621 12958 -3617
rect 2915 -4142 2949 -3966
rect 3033 -4142 3067 -3966
rect 3151 -4142 3185 -3966
rect 3269 -4142 3303 -3966
rect 3387 -4142 3421 -3966
rect 3505 -4142 3539 -3966
rect 3623 -4142 3657 -3966
rect 3741 -4142 3775 -3966
rect 3859 -4142 3893 -3966
rect 3977 -4142 4011 -3966
rect 7099 -4044 7100 -3895
rect 7100 -4044 7166 -3895
rect 9466 -4144 9500 -3968
rect 9584 -4144 9618 -3968
rect 9702 -4144 9736 -3968
rect 9820 -4144 9854 -3968
rect 9938 -4144 9972 -3968
rect 10056 -4144 10090 -3968
rect 10174 -4144 10208 -3968
rect 10292 -4144 10326 -3968
rect 10410 -4144 10444 -3968
rect 10528 -4144 10562 -3968
rect 13655 -3897 13722 -3896
rect 13655 -4045 13718 -3897
rect 13718 -4045 13722 -3897
rect 3682 -4236 3716 -4202
rect 10233 -4238 10267 -4204
rect 3564 -4353 3598 -4319
rect 3152 -4779 3186 -4403
rect 3270 -4779 3304 -4403
rect 3388 -4779 3422 -4403
rect 3505 -4579 3539 -4403
rect 3623 -4579 3657 -4403
rect 3723 -4814 3872 -4747
rect 4379 -4759 4413 -4583
rect 4497 -4759 4531 -4583
rect 4615 -4759 4649 -4583
rect 4733 -4759 4767 -4583
rect 4863 -4759 4897 -4383
rect 4981 -4759 5015 -4383
rect 5099 -4759 5133 -4383
rect 5217 -4759 5251 -4383
rect 5335 -4759 5369 -4383
rect 5453 -4759 5487 -4383
rect 5571 -4759 5605 -4383
rect 5700 -4759 5734 -4583
rect 5818 -4759 5852 -4583
rect 5936 -4759 5970 -4583
rect 6054 -4759 6088 -4583
rect 6277 -4759 6311 -4583
rect 6395 -4759 6429 -4583
rect 6513 -4759 6547 -4583
rect 6631 -4759 6665 -4583
rect 6761 -4759 6795 -4383
rect 6879 -4759 6913 -4383
rect 6997 -4759 7031 -4383
rect 7115 -4759 7149 -4383
rect 7233 -4759 7267 -4383
rect 10115 -4355 10149 -4321
rect 7351 -4759 7385 -4383
rect 7469 -4759 7503 -4383
rect 7598 -4759 7632 -4583
rect 7716 -4759 7750 -4583
rect 7834 -4759 7868 -4583
rect 7952 -4759 7986 -4583
rect 9703 -4781 9737 -4405
rect 9821 -4781 9855 -4405
rect 9939 -4781 9973 -4405
rect 10056 -4581 10090 -4405
rect 10174 -4581 10208 -4405
rect 3211 -4863 3245 -4829
rect 3329 -4863 3363 -4829
rect 10281 -4815 10430 -4748
rect 10930 -4761 10964 -4585
rect 11048 -4761 11082 -4585
rect 11166 -4761 11200 -4585
rect 11284 -4761 11318 -4585
rect 11414 -4761 11448 -4385
rect 11532 -4761 11566 -4385
rect 11650 -4761 11684 -4385
rect 11768 -4761 11802 -4385
rect 11886 -4761 11920 -4385
rect 12004 -4761 12038 -4385
rect 12122 -4761 12156 -4385
rect 12251 -4761 12285 -4585
rect 12369 -4761 12403 -4585
rect 12487 -4761 12521 -4585
rect 12605 -4761 12639 -4585
rect 12828 -4761 12862 -4585
rect 12946 -4761 12980 -4585
rect 13064 -4761 13098 -4585
rect 13182 -4761 13216 -4585
rect 13312 -4761 13346 -4385
rect 13430 -4761 13464 -4385
rect 13548 -4761 13582 -4385
rect 13666 -4761 13700 -4385
rect 13784 -4761 13818 -4385
rect 13902 -4761 13936 -4385
rect 14020 -4761 14054 -4385
rect 14149 -4761 14183 -4585
rect 14267 -4761 14301 -4585
rect 14385 -4761 14419 -4585
rect 14503 -4761 14537 -4585
rect 9762 -4865 9796 -4831
rect 9880 -4865 9914 -4831
rect 5843 -5031 5877 -4997
rect 7950 -5052 7984 -5018
rect 12394 -5033 12428 -4999
rect 3382 -5156 3449 -5153
rect 3382 -5302 3384 -5156
rect 3384 -5302 3449 -5156
rect 4806 -5452 4840 -5076
rect 4924 -5452 4958 -5076
rect 2910 -5746 2944 -5570
rect 3028 -5746 3062 -5570
rect 3146 -5746 3180 -5570
rect 3264 -5746 3298 -5570
rect 3382 -5746 3416 -5570
rect 3500 -5746 3534 -5570
rect 3618 -5746 3652 -5570
rect 3736 -5746 3770 -5570
rect 3854 -5746 3888 -5570
rect 5042 -5452 5076 -5076
rect 5160 -5452 5194 -5076
rect 5278 -5452 5312 -5076
rect 5396 -5452 5430 -5076
rect 5514 -5452 5548 -5076
rect 6704 -5452 6738 -5076
rect 6822 -5452 6856 -5076
rect 6940 -5452 6974 -5076
rect 7058 -5452 7092 -5076
rect 7176 -5452 7210 -5076
rect 7294 -5452 7328 -5076
rect 14501 -5054 14535 -5020
rect 7412 -5452 7446 -5076
rect 9938 -5307 10002 -5158
rect 10002 -5307 10005 -5158
rect 11357 -5454 11391 -5078
rect 11475 -5454 11509 -5078
rect 3972 -5746 4006 -5570
rect 4836 -5674 4870 -5640
rect 4651 -5741 4685 -5707
rect 5484 -5674 5518 -5640
rect 6734 -5674 6768 -5640
rect 5102 -5758 5136 -5724
rect 5220 -5757 5254 -5723
rect 5774 -5742 5808 -5708
rect 6549 -5741 6583 -5707
rect 8073 -5579 8205 -5481
rect 7380 -5673 7414 -5639
rect 7000 -5758 7034 -5724
rect 7118 -5757 7152 -5723
rect 7672 -5742 7706 -5708
rect 9461 -5748 9495 -5572
rect 9579 -5748 9613 -5572
rect 9697 -5748 9731 -5572
rect 9815 -5748 9849 -5572
rect 9933 -5748 9967 -5572
rect 10051 -5748 10085 -5572
rect 10169 -5748 10203 -5572
rect 10287 -5748 10321 -5572
rect 10405 -5748 10439 -5572
rect 11593 -5454 11627 -5078
rect 11711 -5454 11745 -5078
rect 11829 -5454 11863 -5078
rect 11947 -5454 11981 -5078
rect 12065 -5454 12099 -5078
rect 13255 -5454 13289 -5078
rect 13373 -5454 13407 -5078
rect 13491 -5454 13525 -5078
rect 13609 -5454 13643 -5078
rect 13727 -5454 13761 -5078
rect 13845 -5454 13879 -5078
rect 13963 -5454 13997 -5078
rect 10523 -5748 10557 -5572
rect 11387 -5676 11421 -5642
rect 11202 -5743 11236 -5709
rect 3677 -5840 3711 -5806
rect 3559 -5957 3593 -5923
rect 4504 -5984 4538 -5808
rect 3147 -6383 3181 -6007
rect 3265 -6383 3299 -6007
rect 3383 -6383 3417 -6007
rect 3500 -6183 3534 -6007
rect 4622 -5984 4656 -5808
rect 3618 -6183 3652 -6007
rect 4924 -6184 4958 -5808
rect 5042 -6184 5076 -5808
rect 5160 -6184 5194 -5808
rect 5278 -6184 5312 -5808
rect 5396 -6184 5430 -5808
rect 5802 -5984 5836 -5808
rect 5920 -5984 5954 -5808
rect 6402 -5984 6436 -5808
rect 6520 -5984 6554 -5808
rect 6822 -6184 6856 -5808
rect 6940 -6184 6974 -5808
rect 7058 -6184 7092 -5808
rect 7176 -6184 7210 -5808
rect 7294 -6184 7328 -5808
rect 7700 -5984 7734 -5808
rect 12035 -5676 12069 -5642
rect 13285 -5676 13319 -5642
rect 11653 -5760 11687 -5726
rect 11771 -5759 11805 -5725
rect 12325 -5744 12359 -5710
rect 13100 -5743 13134 -5709
rect 13931 -5675 13965 -5641
rect 13551 -5760 13585 -5726
rect 13669 -5759 13703 -5725
rect 14223 -5744 14257 -5710
rect 7818 -5984 7852 -5808
rect 10228 -5842 10262 -5808
rect 10110 -5959 10144 -5925
rect 11055 -5986 11089 -5810
rect 3723 -6406 3872 -6339
rect 9698 -6385 9732 -6009
rect 9816 -6385 9850 -6009
rect 9934 -6385 9968 -6009
rect 10051 -6185 10085 -6009
rect 11173 -5986 11207 -5810
rect 10169 -6185 10203 -6009
rect 11475 -6186 11509 -5810
rect 11593 -6186 11627 -5810
rect 11711 -6186 11745 -5810
rect 11829 -6186 11863 -5810
rect 11947 -6186 11981 -5810
rect 12353 -5986 12387 -5810
rect 12471 -5986 12505 -5810
rect 12953 -5986 12987 -5810
rect 13071 -5986 13105 -5810
rect 13373 -6186 13407 -5810
rect 13491 -6186 13525 -5810
rect 13609 -6186 13643 -5810
rect 13727 -6186 13761 -5810
rect 13845 -6186 13879 -5810
rect 14251 -5986 14285 -5810
rect 14369 -5986 14403 -5810
rect 3206 -6467 3240 -6433
rect 3324 -6467 3358 -6433
rect 10270 -6415 10419 -6348
rect 9757 -6469 9791 -6435
rect 9875 -6469 9909 -6435
rect 5144 -6656 5211 -6507
rect 11692 -6657 11759 -6508
rect 16107 -2493 16141 -2317
rect 16225 -2493 16259 -2317
rect 16343 -2493 16377 -2317
rect 16461 -2493 16495 -2317
rect 16579 -2493 16613 -2317
rect 16697 -2493 16731 -2317
rect 16815 -2493 16849 -2317
rect 16933 -2493 16967 -2317
rect 17051 -2493 17085 -2317
rect 17169 -2493 17203 -2317
rect 16874 -2587 16908 -2553
rect 18432 -2621 18466 -2245
rect 18550 -2621 18584 -2245
rect 18668 -2621 18702 -2245
rect 18786 -2621 18820 -2245
rect 18904 -2621 18938 -2245
rect 19022 -2621 19056 -2245
rect 24939 -2220 24973 -2186
rect 19140 -2621 19174 -2245
rect 19574 -2617 19608 -2241
rect 19692 -2617 19726 -2241
rect 19810 -2617 19844 -2241
rect 19928 -2617 19962 -2241
rect 20046 -2617 20080 -2241
rect 20164 -2617 20198 -2241
rect 20282 -2617 20316 -2241
rect 26069 -2216 26103 -2182
rect 22729 -2492 22763 -2316
rect 22847 -2492 22881 -2316
rect 22965 -2492 22999 -2316
rect 23083 -2492 23117 -2316
rect 23201 -2492 23235 -2316
rect 23319 -2492 23353 -2316
rect 23437 -2492 23471 -2316
rect 23555 -2492 23589 -2316
rect 23673 -2492 23707 -2316
rect 23791 -2492 23825 -2316
rect 23496 -2586 23530 -2552
rect 25054 -2620 25088 -2244
rect 25172 -2620 25206 -2244
rect 25290 -2620 25324 -2244
rect 25408 -2620 25442 -2244
rect 25526 -2620 25560 -2244
rect 25644 -2620 25678 -2244
rect 28605 -2216 28639 -2040
rect 25762 -2620 25796 -2244
rect 26196 -2616 26230 -2240
rect 26314 -2616 26348 -2240
rect 26432 -2616 26466 -2240
rect 26550 -2616 26584 -2240
rect 26668 -2616 26702 -2240
rect 26786 -2616 26820 -2240
rect 28723 -2216 28757 -2040
rect 28841 -2216 28875 -2040
rect 28959 -2216 28993 -2040
rect 29077 -2216 29111 -2040
rect 29195 -2216 29229 -2040
rect 29313 -2216 29347 -2040
rect 29431 -2216 29465 -2040
rect 29549 -2216 29583 -2040
rect 29667 -2216 29701 -2040
rect 26904 -2616 26938 -2240
rect 29372 -2310 29406 -2276
rect 29254 -2427 29288 -2393
rect 16756 -2704 16790 -2670
rect 23378 -2703 23412 -2669
rect 16344 -3130 16378 -2754
rect 16462 -3130 16496 -2754
rect 16580 -3130 16614 -2754
rect 16697 -2930 16731 -2754
rect 16815 -2930 16849 -2754
rect 18637 -2977 18671 -2943
rect 19779 -2973 19813 -2939
rect 16926 -3161 17075 -3094
rect 16403 -3214 16437 -3180
rect 16521 -3214 16555 -3180
rect 18342 -3204 18376 -3028
rect 18460 -3204 18494 -3028
rect 18578 -3204 18612 -3028
rect 18696 -3204 18730 -3028
rect 18861 -3204 18895 -3028
rect 18979 -3204 19013 -3028
rect 19097 -3204 19131 -3028
rect 19215 -3204 19249 -3028
rect 19484 -3200 19518 -3024
rect 19602 -3200 19636 -3024
rect 19720 -3200 19754 -3024
rect 19838 -3200 19872 -3024
rect 20003 -3200 20037 -3024
rect 20121 -3200 20155 -3024
rect 20239 -3200 20273 -3024
rect 20357 -3200 20391 -3024
rect 22966 -3129 23000 -2753
rect 23084 -3129 23118 -2753
rect 23202 -3129 23236 -2753
rect 23319 -2929 23353 -2753
rect 23437 -2929 23471 -2753
rect 28842 -2853 28876 -2477
rect 28960 -2853 28994 -2477
rect 29078 -2853 29112 -2477
rect 29195 -2653 29229 -2477
rect 29313 -2653 29347 -2477
rect 30349 -2683 30383 -2507
rect 30467 -2683 30501 -2507
rect 30585 -2683 30619 -2507
rect 30703 -2683 30737 -2507
rect 30833 -2683 30867 -2307
rect 30951 -2683 30985 -2307
rect 31069 -2683 31103 -2307
rect 31187 -2683 31221 -2307
rect 31305 -2683 31339 -2307
rect 31423 -2683 31457 -2307
rect 31541 -2683 31575 -2307
rect 32483 -2334 32543 -2272
rect 31670 -2683 31704 -2507
rect 31788 -2683 31822 -2507
rect 31906 -2683 31940 -2507
rect 32024 -2683 32058 -2507
rect 32142 -2686 32176 -2510
rect 32260 -2686 32294 -2510
rect 32378 -2686 32412 -2510
rect 32496 -2686 32530 -2510
rect 32614 -2686 32648 -2510
rect 32732 -2686 32766 -2510
rect 32850 -2686 32884 -2510
rect 32968 -2686 33002 -2510
rect 33086 -2686 33120 -2510
rect 33204 -2686 33238 -2510
rect 32909 -2780 32943 -2746
rect 32001 -2899 32035 -2865
rect 32791 -2897 32825 -2863
rect 28901 -2937 28935 -2903
rect 29019 -2937 29053 -2903
rect 25259 -2976 25293 -2942
rect 26401 -2972 26435 -2938
rect 23542 -3156 23691 -3089
rect 23025 -3213 23059 -3179
rect 23143 -3213 23177 -3179
rect 24964 -3203 24998 -3027
rect 25082 -3203 25116 -3027
rect 25200 -3203 25234 -3027
rect 25318 -3203 25352 -3027
rect 25483 -3203 25517 -3027
rect 25601 -3203 25635 -3027
rect 25719 -3203 25753 -3027
rect 25837 -3203 25871 -3027
rect 26106 -3199 26140 -3023
rect 26224 -3199 26258 -3023
rect 26342 -3199 26376 -3023
rect 26460 -3199 26494 -3023
rect 26625 -3199 26659 -3023
rect 26743 -3199 26777 -3023
rect 26861 -3199 26895 -3023
rect 26979 -3199 27013 -3023
rect 29174 -3060 29226 -3014
rect 30601 -3018 30635 -2984
rect 30776 -3376 30810 -3000
rect 30894 -3376 30928 -3000
rect 16598 -3553 16665 -3552
rect 16598 -3701 16662 -3553
rect 16662 -3701 16665 -3553
rect 18402 -3606 18469 -3457
rect 19548 -3603 19615 -3454
rect 23217 -3552 23284 -3551
rect 23217 -3700 23284 -3552
rect 25033 -3602 25100 -3453
rect 26167 -3611 26234 -3462
rect 31012 -3376 31046 -3000
rect 31130 -3376 31164 -3000
rect 31248 -3376 31282 -3000
rect 31366 -3376 31400 -3000
rect 31484 -3376 31518 -3000
rect 31650 -3296 31712 -3205
rect 32379 -3323 32413 -2947
rect 32497 -3323 32531 -2947
rect 32615 -3323 32649 -2947
rect 32732 -3123 32766 -2947
rect 32850 -3123 32884 -2947
rect 32438 -3407 32472 -3373
rect 32556 -3407 32590 -3373
rect 30806 -3598 30840 -3564
rect 30621 -3665 30655 -3631
rect 32711 -3530 32763 -3484
rect 31454 -3598 31488 -3564
rect 31072 -3682 31106 -3648
rect 31190 -3681 31224 -3647
rect 31744 -3666 31778 -3632
rect 16121 -4143 16155 -3967
rect 16239 -4143 16273 -3967
rect 16357 -4143 16391 -3967
rect 16475 -4143 16509 -3967
rect 16593 -4143 16627 -3967
rect 16711 -4143 16745 -3967
rect 16829 -4143 16863 -3967
rect 16947 -4143 16981 -3967
rect 17065 -4143 17099 -3967
rect 17183 -4143 17217 -3967
rect 20309 -3896 20376 -3894
rect 20309 -4043 20373 -3896
rect 20373 -4043 20376 -3896
rect 22743 -4142 22777 -3966
rect 22861 -4142 22895 -3966
rect 22979 -4142 23013 -3966
rect 23097 -4142 23131 -3966
rect 23215 -4142 23249 -3966
rect 23333 -4142 23367 -3966
rect 23451 -4142 23485 -3966
rect 23569 -4142 23603 -3966
rect 23687 -4142 23721 -3966
rect 23805 -4142 23839 -3966
rect 26930 -4044 26995 -3896
rect 26995 -4044 26997 -3896
rect 26930 -4045 26997 -4044
rect 30474 -3908 30508 -3732
rect 30592 -3908 30626 -3732
rect 30894 -4108 30928 -3732
rect 31012 -4108 31046 -3732
rect 31130 -4108 31164 -3732
rect 31248 -4108 31282 -3732
rect 31366 -4108 31400 -3732
rect 31772 -3908 31806 -3732
rect 31890 -3908 31924 -3732
rect 16888 -4237 16922 -4203
rect 23510 -4236 23544 -4202
rect 16770 -4354 16804 -4320
rect 16358 -4780 16392 -4404
rect 16476 -4780 16510 -4404
rect 16594 -4780 16628 -4404
rect 16711 -4580 16745 -4404
rect 16829 -4580 16863 -4404
rect 16937 -4812 17086 -4745
rect 17585 -4760 17619 -4584
rect 17703 -4760 17737 -4584
rect 17821 -4760 17855 -4584
rect 17939 -4760 17973 -4584
rect 18069 -4760 18103 -4384
rect 18187 -4760 18221 -4384
rect 18305 -4760 18339 -4384
rect 18423 -4760 18457 -4384
rect 18541 -4760 18575 -4384
rect 18659 -4760 18693 -4384
rect 18777 -4760 18811 -4384
rect 18906 -4760 18940 -4584
rect 19024 -4760 19058 -4584
rect 19142 -4760 19176 -4584
rect 19260 -4760 19294 -4584
rect 19483 -4760 19517 -4584
rect 19601 -4760 19635 -4584
rect 19719 -4760 19753 -4584
rect 19837 -4760 19871 -4584
rect 19967 -4760 20001 -4384
rect 20085 -4760 20119 -4384
rect 20203 -4760 20237 -4384
rect 20321 -4760 20355 -4384
rect 20439 -4760 20473 -4384
rect 23392 -4353 23426 -4319
rect 20557 -4760 20591 -4384
rect 20675 -4760 20709 -4384
rect 20804 -4760 20838 -4584
rect 20922 -4760 20956 -4584
rect 21040 -4760 21074 -4584
rect 21158 -4760 21192 -4584
rect 22980 -4779 23014 -4403
rect 23098 -4779 23132 -4403
rect 23216 -4779 23250 -4403
rect 23333 -4579 23367 -4403
rect 23451 -4579 23485 -4403
rect 16417 -4864 16451 -4830
rect 16535 -4864 16569 -4830
rect 23560 -4805 23709 -4738
rect 24207 -4759 24241 -4583
rect 24325 -4759 24359 -4583
rect 24443 -4759 24477 -4583
rect 24561 -4759 24595 -4583
rect 24691 -4759 24725 -4383
rect 24809 -4759 24843 -4383
rect 24927 -4759 24961 -4383
rect 25045 -4759 25079 -4383
rect 25163 -4759 25197 -4383
rect 25281 -4759 25315 -4383
rect 25399 -4759 25433 -4383
rect 25528 -4759 25562 -4583
rect 25646 -4759 25680 -4583
rect 25764 -4759 25798 -4583
rect 25882 -4759 25916 -4583
rect 26105 -4759 26139 -4583
rect 26223 -4759 26257 -4583
rect 26341 -4759 26375 -4583
rect 26459 -4759 26493 -4583
rect 26589 -4759 26623 -4383
rect 26707 -4759 26741 -4383
rect 26825 -4759 26859 -4383
rect 26943 -4759 26977 -4383
rect 27061 -4759 27095 -4383
rect 27179 -4759 27213 -4383
rect 27297 -4759 27331 -4383
rect 31088 -4381 31223 -4279
rect 27426 -4759 27460 -4583
rect 27544 -4759 27578 -4583
rect 27662 -4759 27696 -4583
rect 27780 -4759 27814 -4583
rect 23039 -4863 23073 -4829
rect 23157 -4863 23191 -4829
rect 28943 -4934 29003 -4872
rect 19049 -5032 19083 -4998
rect 21156 -5053 21190 -5019
rect 25671 -5031 25705 -4997
rect 16593 -5306 16657 -5160
rect 16657 -5306 16660 -5160
rect 16593 -5309 16660 -5306
rect 18012 -5453 18046 -5077
rect 18130 -5453 18164 -5077
rect 16116 -5747 16150 -5571
rect 16234 -5747 16268 -5571
rect 16352 -5747 16386 -5571
rect 16470 -5747 16504 -5571
rect 16588 -5747 16622 -5571
rect 16706 -5747 16740 -5571
rect 16824 -5747 16858 -5571
rect 16942 -5747 16976 -5571
rect 17060 -5747 17094 -5571
rect 18248 -5453 18282 -5077
rect 18366 -5453 18400 -5077
rect 18484 -5453 18518 -5077
rect 18602 -5453 18636 -5077
rect 18720 -5453 18754 -5077
rect 19910 -5453 19944 -5077
rect 20028 -5453 20062 -5077
rect 20146 -5453 20180 -5077
rect 20264 -5453 20298 -5077
rect 20382 -5453 20416 -5077
rect 20500 -5453 20534 -5077
rect 27778 -5052 27812 -5018
rect 20618 -5453 20652 -5077
rect 23214 -5305 23279 -5160
rect 23279 -5305 23281 -5160
rect 23214 -5309 23281 -5305
rect 24634 -5452 24668 -5076
rect 24752 -5452 24786 -5076
rect 17178 -5747 17212 -5571
rect 18042 -5675 18076 -5641
rect 17857 -5742 17891 -5708
rect 18690 -5675 18724 -5641
rect 19940 -5675 19974 -5641
rect 18308 -5759 18342 -5725
rect 18426 -5758 18460 -5724
rect 18980 -5743 19014 -5709
rect 19755 -5742 19789 -5708
rect 21279 -5580 21411 -5482
rect 20586 -5674 20620 -5640
rect 20206 -5759 20240 -5725
rect 20324 -5758 20358 -5724
rect 20878 -5743 20912 -5709
rect 22738 -5746 22772 -5570
rect 22856 -5746 22890 -5570
rect 22974 -5746 23008 -5570
rect 23092 -5746 23126 -5570
rect 23210 -5746 23244 -5570
rect 23328 -5746 23362 -5570
rect 23446 -5746 23480 -5570
rect 23564 -5746 23598 -5570
rect 23682 -5746 23716 -5570
rect 24870 -5452 24904 -5076
rect 24988 -5452 25022 -5076
rect 25106 -5452 25140 -5076
rect 25224 -5452 25258 -5076
rect 25342 -5452 25376 -5076
rect 26532 -5452 26566 -5076
rect 26650 -5452 26684 -5076
rect 26768 -5452 26802 -5076
rect 26886 -5452 26920 -5076
rect 27004 -5452 27038 -5076
rect 27122 -5452 27156 -5076
rect 27240 -5452 27274 -5076
rect 28602 -5286 28636 -5110
rect 28720 -5286 28754 -5110
rect 28838 -5286 28872 -5110
rect 28956 -5286 28990 -5110
rect 29074 -5286 29108 -5110
rect 29192 -5286 29226 -5110
rect 29310 -5286 29344 -5110
rect 29428 -5286 29462 -5110
rect 29546 -5286 29580 -5110
rect 29664 -5286 29698 -5110
rect 29369 -5380 29403 -5346
rect 23800 -5746 23834 -5570
rect 24664 -5674 24698 -5640
rect 24479 -5741 24513 -5707
rect 25312 -5674 25346 -5640
rect 26562 -5674 26596 -5640
rect 24930 -5758 24964 -5724
rect 25048 -5757 25082 -5723
rect 25602 -5742 25636 -5708
rect 26377 -5741 26411 -5707
rect 27901 -5579 28033 -5481
rect 29251 -5497 29285 -5463
rect 27208 -5673 27242 -5639
rect 26828 -5758 26862 -5724
rect 26946 -5757 26980 -5723
rect 27500 -5742 27534 -5708
rect 16883 -5841 16917 -5807
rect 16765 -5958 16799 -5924
rect 17710 -5985 17744 -5809
rect 16353 -6384 16387 -6008
rect 16471 -6384 16505 -6008
rect 16589 -6384 16623 -6008
rect 16706 -6184 16740 -6008
rect 17828 -5985 17862 -5809
rect 16824 -6184 16858 -6008
rect 18130 -6185 18164 -5809
rect 18248 -6185 18282 -5809
rect 18366 -6185 18400 -5809
rect 18484 -6185 18518 -5809
rect 18602 -6185 18636 -5809
rect 19008 -5985 19042 -5809
rect 19126 -5985 19160 -5809
rect 19608 -5985 19642 -5809
rect 19726 -5985 19760 -5809
rect 20028 -6185 20062 -5809
rect 20146 -6185 20180 -5809
rect 20264 -6185 20298 -5809
rect 20382 -6185 20416 -5809
rect 20500 -6185 20534 -5809
rect 20906 -5985 20940 -5809
rect 21024 -5985 21058 -5809
rect 23505 -5840 23539 -5806
rect 23387 -5957 23421 -5923
rect 24332 -5984 24366 -5808
rect 16940 -6421 17086 -6354
rect 17086 -6421 17089 -6354
rect 22975 -6383 23009 -6007
rect 23093 -6383 23127 -6007
rect 23211 -6383 23245 -6007
rect 23328 -6183 23362 -6007
rect 24450 -5984 24484 -5808
rect 23446 -6183 23480 -6007
rect 24752 -6184 24786 -5808
rect 24870 -6184 24904 -5808
rect 24988 -6184 25022 -5808
rect 25106 -6184 25140 -5808
rect 25224 -6184 25258 -5808
rect 25630 -5984 25664 -5808
rect 25748 -5984 25782 -5808
rect 26230 -5984 26264 -5808
rect 26348 -5984 26382 -5808
rect 26650 -6184 26684 -5808
rect 26768 -6184 26802 -5808
rect 26886 -6184 26920 -5808
rect 27004 -6184 27038 -5808
rect 27122 -6184 27156 -5808
rect 27528 -5984 27562 -5808
rect 27646 -5984 27680 -5808
rect 28839 -5923 28873 -5547
rect 28957 -5923 28991 -5547
rect 29075 -5923 29109 -5547
rect 29192 -5723 29226 -5547
rect 29310 -5723 29344 -5547
rect 28898 -6007 28932 -5973
rect 29016 -6007 29050 -5973
rect 29171 -6130 29223 -6084
rect 30983 -6151 31404 -6117
rect 30983 -6296 31046 -6151
rect 31046 -6296 31355 -6151
rect 31355 -6296 31404 -6151
rect 30983 -6317 31404 -6296
rect 16412 -6468 16446 -6434
rect 16530 -6468 16564 -6434
rect 23551 -6422 23700 -6355
rect 15301 -6671 15371 -6603
rect 23034 -6467 23068 -6433
rect 23152 -6467 23186 -6433
rect 18342 -6656 18409 -6507
rect 24970 -6650 25037 -6501
rect 30349 -7031 30383 -6855
rect 30467 -7031 30501 -6855
rect 30585 -7031 30619 -6855
rect 30703 -7031 30737 -6855
rect 30833 -7031 30867 -6655
rect 30951 -7031 30985 -6655
rect 31069 -7031 31103 -6655
rect 31187 -7031 31221 -6655
rect 31305 -7031 31339 -6655
rect 31423 -7031 31457 -6655
rect 31541 -7031 31575 -6655
rect 32483 -6682 32543 -6620
rect 31670 -7031 31704 -6855
rect 31788 -7031 31822 -6855
rect 31906 -7031 31940 -6855
rect 32024 -7031 32058 -6855
rect 32142 -7034 32176 -6858
rect 32260 -7034 32294 -6858
rect 32378 -7034 32412 -6858
rect 32496 -7034 32530 -6858
rect 32614 -7034 32648 -6858
rect 32732 -7034 32766 -6858
rect 32850 -7034 32884 -6858
rect 32968 -7034 33002 -6858
rect 33086 -7034 33120 -6858
rect 33204 -7034 33238 -6858
rect 32909 -7128 32943 -7094
rect 7287 -7275 7339 -7229
rect 13841 -7270 13893 -7224
rect 20490 -7282 20542 -7236
rect 30329 -7264 30402 -7193
rect 32001 -7247 32035 -7213
rect 32791 -7245 32825 -7211
rect 7014 -7386 7048 -7352
rect 7132 -7386 7166 -7352
rect 13568 -7381 13602 -7347
rect 13686 -7381 13720 -7347
rect 20217 -7393 20251 -7359
rect 20335 -7393 20369 -7359
rect 30601 -7366 30635 -7332
rect 6955 -7812 6989 -7436
rect 7073 -7812 7107 -7436
rect 7191 -7812 7225 -7436
rect 7308 -7812 7342 -7636
rect 7426 -7812 7460 -7636
rect 13509 -7807 13543 -7431
rect 13627 -7807 13661 -7431
rect 13745 -7807 13779 -7431
rect 13862 -7807 13896 -7631
rect 13980 -7807 14014 -7631
rect 20158 -7819 20192 -7443
rect 20276 -7819 20310 -7443
rect 20394 -7819 20428 -7443
rect 20511 -7819 20545 -7643
rect 20629 -7819 20663 -7643
rect 28950 -7779 29010 -7717
rect 30776 -7724 30810 -7348
rect 30894 -7724 30928 -7348
rect 31012 -7724 31046 -7348
rect 31130 -7724 31164 -7348
rect 31248 -7724 31282 -7348
rect 31366 -7724 31400 -7348
rect 31484 -7724 31518 -7348
rect 31650 -7644 31712 -7553
rect 32379 -7671 32413 -7295
rect 32497 -7671 32531 -7295
rect 32615 -7671 32649 -7295
rect 32732 -7471 32766 -7295
rect 32850 -7471 32884 -7295
rect 32438 -7755 32472 -7721
rect 32556 -7755 32590 -7721
rect 7367 -7896 7401 -7862
rect 13921 -7891 13955 -7857
rect 20570 -7903 20604 -7869
rect 7485 -8013 7519 -7979
rect 14039 -8008 14073 -7974
rect 20688 -8020 20722 -7986
rect 6718 -8249 6752 -8073
rect 6836 -8249 6870 -8073
rect 6954 -8249 6988 -8073
rect 7072 -8249 7106 -8073
rect 7190 -8249 7224 -8073
rect 7308 -8249 7342 -8073
rect 7426 -8249 7460 -8073
rect 7544 -8249 7578 -8073
rect 7662 -8249 7696 -8073
rect 7780 -8249 7814 -8073
rect 13272 -8244 13306 -8068
rect 13390 -8244 13424 -8068
rect 13508 -8244 13542 -8068
rect 13626 -8244 13660 -8068
rect 13744 -8244 13778 -8068
rect 13862 -8244 13896 -8068
rect 13980 -8244 14014 -8068
rect 14098 -8244 14132 -8068
rect 14216 -8244 14250 -8068
rect 14334 -8244 14368 -8068
rect 19921 -8256 19955 -8080
rect 20039 -8256 20073 -8080
rect 20157 -8256 20191 -8080
rect 20275 -8256 20309 -8080
rect 20393 -8256 20427 -8080
rect 20511 -8256 20545 -8080
rect 20629 -8256 20663 -8080
rect 20747 -8256 20781 -8080
rect 20865 -8256 20899 -8080
rect 20983 -8256 21017 -8080
rect 28609 -8131 28643 -7955
rect 28727 -8131 28761 -7955
rect 28845 -8131 28879 -7955
rect 28963 -8131 28997 -7955
rect 29081 -8131 29115 -7955
rect 29199 -8131 29233 -7955
rect 29317 -8131 29351 -7955
rect 29435 -8131 29469 -7955
rect 29553 -8131 29587 -7955
rect 29671 -8131 29705 -7955
rect 30806 -7946 30840 -7912
rect 30621 -8013 30655 -7979
rect 32711 -7878 32763 -7832
rect 31454 -7946 31488 -7912
rect 31072 -8030 31106 -7996
rect 31190 -8029 31224 -7995
rect 31744 -8014 31778 -7980
rect 29376 -8225 29410 -8191
rect 30474 -8256 30508 -8080
rect 30592 -8256 30626 -8080
rect 29258 -8342 29292 -8308
rect 7059 -8487 7119 -8425
rect 13613 -8482 13673 -8420
rect 20262 -8494 20322 -8432
rect 28846 -8768 28880 -8392
rect 28964 -8768 28998 -8392
rect 29082 -8768 29116 -8392
rect 29199 -8568 29233 -8392
rect 29317 -8568 29351 -8392
rect 30894 -8456 30928 -8080
rect 31012 -8456 31046 -8080
rect 31130 -8456 31164 -8080
rect 31248 -8456 31282 -8080
rect 31366 -8456 31400 -8080
rect 31772 -8256 31806 -8080
rect 31890 -8256 31924 -8080
rect 31088 -8729 31223 -8627
rect 28905 -8852 28939 -8818
rect 29023 -8852 29057 -8818
rect 29178 -8975 29230 -8929
rect 1619 -9304 1763 -9238
<< metal1 >>
rect 27799 5939 27912 6232
rect 20191 5889 20327 5909
rect 6988 5869 7124 5889
rect 6988 5807 7024 5869
rect 7084 5807 7124 5869
rect 6988 5779 7124 5807
rect 13537 5868 13673 5888
rect 13537 5806 13573 5868
rect 13633 5806 13673 5868
rect 6684 5749 7661 5779
rect 13537 5778 13673 5806
rect 20191 5827 20227 5889
rect 20287 5827 20327 5889
rect 20191 5799 20327 5827
rect 6684 5643 6716 5749
rect 6920 5643 6952 5749
rect 7156 5643 7188 5749
rect 7392 5643 7424 5749
rect 7627 5643 7661 5749
rect 13233 5748 14210 5778
rect 6677 5631 6723 5643
rect 6677 5455 6683 5631
rect 6717 5455 6723 5631
rect 6677 5443 6723 5455
rect 6795 5631 6841 5643
rect 6795 5455 6801 5631
rect 6835 5455 6841 5631
rect 6795 5443 6841 5455
rect 6913 5631 6959 5643
rect 6913 5455 6919 5631
rect 6953 5455 6959 5631
rect 6913 5443 6959 5455
rect 7031 5631 7077 5643
rect 7031 5455 7037 5631
rect 7071 5455 7077 5631
rect 7031 5443 7077 5455
rect 7149 5631 7195 5643
rect 7149 5455 7155 5631
rect 7189 5455 7195 5631
rect 7149 5443 7195 5455
rect 7267 5631 7313 5643
rect 7267 5455 7273 5631
rect 7307 5455 7313 5631
rect 7267 5443 7313 5455
rect 7385 5631 7431 5643
rect 7385 5455 7391 5631
rect 7425 5455 7431 5631
rect 7385 5443 7431 5455
rect 7503 5631 7549 5643
rect 7503 5455 7509 5631
rect 7543 5455 7549 5631
rect 7503 5443 7549 5455
rect 7621 5631 7667 5643
rect 7621 5455 7627 5631
rect 7661 5455 7667 5631
rect 7621 5443 7667 5455
rect 7739 5631 7785 5643
rect 13233 5642 13265 5748
rect 13469 5642 13501 5748
rect 13705 5642 13737 5748
rect 13941 5642 13973 5748
rect 14176 5642 14210 5748
rect 19887 5769 20864 5799
rect 19887 5663 19919 5769
rect 20123 5663 20155 5769
rect 20359 5663 20391 5769
rect 20595 5663 20627 5769
rect 20830 5663 20864 5769
rect 19880 5651 19926 5663
rect 7739 5455 7745 5631
rect 7779 5455 7785 5631
rect 7739 5443 7785 5455
rect 13226 5630 13272 5642
rect 13226 5454 13232 5630
rect 13266 5454 13272 5630
rect 6800 5349 6836 5443
rect 7036 5349 7072 5443
rect 7272 5350 7308 5443
rect 7434 5395 7500 5402
rect 7434 5361 7450 5395
rect 7484 5361 7500 5395
rect 7434 5350 7500 5361
rect 7272 5349 7500 5350
rect 6800 5320 7500 5349
rect 6800 5319 7382 5320
rect 6920 5206 6954 5319
rect 7316 5278 7382 5319
rect 7316 5244 7332 5278
rect 7366 5244 7382 5278
rect 7316 5237 7382 5244
rect 7744 5212 7779 5443
rect 13226 5442 13272 5454
rect 13344 5630 13390 5642
rect 13344 5454 13350 5630
rect 13384 5454 13390 5630
rect 13344 5442 13390 5454
rect 13462 5630 13508 5642
rect 13462 5454 13468 5630
rect 13502 5454 13508 5630
rect 13462 5442 13508 5454
rect 13580 5630 13626 5642
rect 13580 5454 13586 5630
rect 13620 5454 13626 5630
rect 13580 5442 13626 5454
rect 13698 5630 13744 5642
rect 13698 5454 13704 5630
rect 13738 5454 13744 5630
rect 13698 5442 13744 5454
rect 13816 5630 13862 5642
rect 13816 5454 13822 5630
rect 13856 5454 13862 5630
rect 13816 5442 13862 5454
rect 13934 5630 13980 5642
rect 13934 5454 13940 5630
rect 13974 5454 13980 5630
rect 13934 5442 13980 5454
rect 14052 5630 14098 5642
rect 14052 5454 14058 5630
rect 14092 5454 14098 5630
rect 14052 5442 14098 5454
rect 14170 5630 14216 5642
rect 14170 5454 14176 5630
rect 14210 5454 14216 5630
rect 14170 5442 14216 5454
rect 14288 5630 14334 5642
rect 14288 5454 14294 5630
rect 14328 5454 14334 5630
rect 19880 5475 19886 5651
rect 19920 5475 19926 5651
rect 19880 5463 19926 5475
rect 19998 5651 20044 5663
rect 19998 5475 20004 5651
rect 20038 5475 20044 5651
rect 19998 5463 20044 5475
rect 20116 5651 20162 5663
rect 20116 5475 20122 5651
rect 20156 5475 20162 5651
rect 20116 5463 20162 5475
rect 20234 5651 20280 5663
rect 20234 5475 20240 5651
rect 20274 5475 20280 5651
rect 20234 5463 20280 5475
rect 20352 5651 20398 5663
rect 20352 5475 20358 5651
rect 20392 5475 20398 5651
rect 20352 5463 20398 5475
rect 20470 5651 20516 5663
rect 20470 5475 20476 5651
rect 20510 5475 20516 5651
rect 20470 5463 20516 5475
rect 20588 5651 20634 5663
rect 20588 5475 20594 5651
rect 20628 5475 20634 5651
rect 20588 5463 20634 5475
rect 20706 5651 20752 5663
rect 20706 5475 20712 5651
rect 20746 5475 20752 5651
rect 20706 5463 20752 5475
rect 20824 5651 20870 5663
rect 20824 5475 20830 5651
rect 20864 5475 20870 5651
rect 20824 5463 20870 5475
rect 20942 5651 20988 5663
rect 20942 5475 20948 5651
rect 20982 5475 20988 5651
rect 20942 5463 20988 5475
rect 14288 5442 14334 5454
rect 13349 5348 13385 5442
rect 13585 5348 13621 5442
rect 13821 5349 13857 5442
rect 13983 5394 14049 5401
rect 13983 5360 13999 5394
rect 14033 5360 14049 5394
rect 13983 5349 14049 5360
rect 13821 5348 14049 5349
rect 13349 5319 14049 5348
rect 13349 5318 13931 5319
rect 7674 5210 8991 5212
rect 7390 5206 8991 5210
rect 6914 5194 6960 5206
rect 6914 4818 6920 5194
rect 6954 4818 6960 5194
rect 6914 4806 6960 4818
rect 7032 5194 7078 5206
rect 7032 4818 7038 5194
rect 7072 4818 7078 5194
rect 7032 4806 7078 4818
rect 7150 5194 7196 5206
rect 7150 4818 7156 5194
rect 7190 4845 7196 5194
rect 7267 5194 7313 5206
rect 7267 5018 7273 5194
rect 7307 5018 7313 5194
rect 7267 5011 7313 5018
rect 7385 5194 8991 5206
rect 13469 5205 13503 5318
rect 13865 5277 13931 5318
rect 13865 5243 13881 5277
rect 13915 5243 13931 5277
rect 13865 5236 13931 5243
rect 14293 5244 14328 5442
rect 20003 5369 20039 5463
rect 20239 5369 20275 5463
rect 20475 5370 20511 5463
rect 20637 5415 20703 5422
rect 20637 5381 20653 5415
rect 20687 5381 20703 5415
rect 20637 5370 20703 5381
rect 20475 5369 20703 5370
rect 20003 5340 20703 5369
rect 20003 5339 20585 5340
rect 14293 5209 14329 5244
rect 20123 5226 20157 5339
rect 20519 5298 20585 5339
rect 20519 5264 20535 5298
rect 20569 5264 20585 5298
rect 20519 5257 20585 5264
rect 20947 5230 20982 5463
rect 20593 5226 22267 5230
rect 20117 5214 20163 5226
rect 13939 5205 15641 5209
rect 7385 5018 7391 5194
rect 7425 5181 8991 5194
rect 7425 5018 7431 5181
rect 7674 5100 8991 5181
rect 7267 5006 7316 5011
rect 7385 5006 7431 5018
rect 7273 4845 7316 5006
rect 7190 4818 7316 4845
rect 7150 4806 7316 4818
rect 7156 4802 7316 4806
rect 6661 4768 7029 4774
rect 6661 4734 6979 4768
rect 7013 4734 7029 4768
rect 6661 4718 7029 4734
rect 7081 4768 7147 4774
rect 7081 4734 7097 4768
rect 7131 4734 7147 4768
rect 6661 4526 6740 4718
rect 7081 4689 7147 4734
rect -926 4516 6740 4526
rect -926 4466 -902 4516
rect -841 4466 6740 4516
rect -926 4456 6740 4466
rect 6798 4681 7147 4689
rect 6798 4649 7148 4681
rect 7240 4665 7316 4802
rect 6798 4355 6852 4649
rect 7236 4605 7246 4665
rect 7308 4605 7318 4665
rect 6795 4343 6856 4355
rect -1129 4331 -900 4340
rect -1129 4273 -994 4331
rect -910 4273 -900 4331
rect 6795 4289 6801 4343
rect 6850 4289 6856 4343
rect 6795 4277 6856 4289
rect -1129 4272 -900 4273
rect 324 3969 460 3989
rect -761 3946 -680 3949
rect -766 3894 -756 3946
rect -688 3894 -678 3946
rect 324 3907 360 3969
rect 420 3907 460 3969
rect -761 3892 -680 3894
rect 324 3879 460 3907
rect 5860 3929 5939 3941
rect 3378 3879 3457 3891
rect 20 3849 997 3879
rect 20 3743 52 3849
rect 256 3743 288 3849
rect 492 3743 524 3849
rect 728 3743 760 3849
rect 963 3743 997 3849
rect 3378 3782 3384 3879
rect 3306 3762 3384 3782
rect 3451 3782 3457 3879
rect 5860 3816 5866 3929
rect 5933 3816 5939 3929
rect 7002 3931 7081 3943
rect 7002 3816 7008 3931
rect 7075 3816 7081 3931
rect 3451 3762 3526 3782
rect 13 3731 59 3743
rect 13 3555 19 3731
rect 53 3555 59 3731
rect 13 3543 59 3555
rect 131 3731 177 3743
rect 131 3555 137 3731
rect 171 3555 177 3731
rect 131 3543 177 3555
rect 249 3731 295 3743
rect 249 3555 255 3731
rect 289 3555 295 3731
rect 249 3543 295 3555
rect 367 3731 413 3743
rect 367 3555 373 3731
rect 407 3555 413 3731
rect 367 3543 413 3555
rect 485 3731 531 3743
rect 485 3555 491 3731
rect 525 3555 531 3731
rect 485 3543 531 3555
rect 603 3731 649 3743
rect 603 3555 609 3731
rect 643 3555 649 3731
rect 603 3543 649 3555
rect 721 3731 767 3743
rect 721 3555 727 3731
rect 761 3555 767 3731
rect 721 3543 767 3555
rect 839 3731 885 3743
rect 839 3555 845 3731
rect 879 3555 885 3731
rect 839 3543 885 3555
rect 957 3731 1003 3743
rect 957 3555 963 3731
rect 997 3555 1003 3731
rect 957 3543 1003 3555
rect 1075 3731 1121 3743
rect 1075 3555 1081 3731
rect 1115 3555 1121 3731
rect 3306 3654 3350 3762
rect 3482 3654 3526 3762
rect 5103 3720 5159 3728
rect 3306 3612 3526 3654
rect 4177 3712 5159 3720
rect 4177 3678 5119 3712
rect 5153 3678 5159 3712
rect 5822 3708 5832 3816
rect 5964 3753 5974 3816
rect 5964 3742 5976 3753
rect 5964 3708 5977 3742
rect 6233 3732 6289 3734
rect 4177 3662 5159 3678
rect 5832 3670 5977 3708
rect 4177 3661 5156 3662
rect 1075 3543 1121 3555
rect 2910 3582 3887 3612
rect 136 3449 172 3543
rect 372 3449 408 3543
rect 608 3450 644 3543
rect 770 3495 836 3502
rect 770 3461 786 3495
rect 820 3461 836 3495
rect 770 3450 836 3461
rect 608 3449 836 3450
rect 136 3420 836 3449
rect 136 3419 718 3420
rect 256 3306 290 3419
rect 652 3378 718 3419
rect 652 3344 668 3378
rect 702 3344 718 3378
rect 652 3337 718 3344
rect 1080 3310 1115 3543
rect 2910 3476 2942 3582
rect 3146 3476 3178 3582
rect 3382 3476 3414 3582
rect 3618 3476 3650 3582
rect 3853 3476 3887 3582
rect 726 3306 1115 3310
rect 250 3294 296 3306
rect -1124 2987 210 3004
rect -1124 2911 -484 2987
rect -395 2911 210 2987
rect -1124 2904 210 2911
rect 250 2918 256 3294
rect 290 2918 296 3294
rect 250 2906 296 2918
rect 368 3294 414 3306
rect 368 2918 374 3294
rect 408 2918 414 3294
rect 368 2906 414 2918
rect 486 3294 532 3306
rect 486 2918 492 3294
rect 526 2945 532 3294
rect 603 3294 649 3306
rect 603 3118 609 3294
rect 643 3118 649 3294
rect 603 3111 649 3118
rect 721 3294 1115 3306
rect 721 3118 727 3294
rect 761 3281 1115 3294
rect 761 3118 767 3281
rect 603 3106 652 3111
rect 721 3106 767 3118
rect 609 2945 652 3106
rect 526 2918 652 2945
rect 486 2906 652 2918
rect 134 2874 188 2904
rect 492 2902 652 2906
rect 134 2868 365 2874
rect 134 2834 315 2868
rect 349 2834 365 2868
rect -1125 2809 78 2824
rect 134 2818 365 2834
rect 417 2868 483 2874
rect 417 2834 433 2868
rect 467 2834 483 2868
rect -1125 2733 -922 2809
rect -1124 2725 -922 2733
rect -809 2793 78 2809
rect -809 2749 10 2793
rect 66 2789 78 2793
rect 417 2789 483 2834
rect 66 2781 483 2789
rect 66 2749 484 2781
rect 576 2765 652 2902
rect -809 2725 79 2749
rect -1124 2713 79 2725
rect 572 2705 582 2765
rect 644 2705 654 2765
rect 1011 2637 1115 3281
rect 2903 3464 2949 3476
rect 2903 3288 2909 3464
rect 2943 3288 2949 3464
rect 2903 3276 2949 3288
rect 3021 3464 3067 3476
rect 3021 3288 3027 3464
rect 3061 3288 3067 3464
rect 3021 3276 3067 3288
rect 3139 3464 3185 3476
rect 3139 3288 3145 3464
rect 3179 3288 3185 3464
rect 3139 3276 3185 3288
rect 3257 3464 3303 3476
rect 3257 3288 3263 3464
rect 3297 3288 3303 3464
rect 3257 3276 3303 3288
rect 3375 3464 3421 3476
rect 3375 3288 3381 3464
rect 3415 3288 3421 3464
rect 3375 3276 3421 3288
rect 3493 3464 3539 3476
rect 3493 3288 3499 3464
rect 3533 3288 3539 3464
rect 3493 3276 3539 3288
rect 3611 3464 3657 3476
rect 3611 3288 3617 3464
rect 3651 3288 3657 3464
rect 3611 3276 3657 3288
rect 3729 3464 3775 3476
rect 3729 3288 3735 3464
rect 3769 3288 3775 3464
rect 3729 3276 3775 3288
rect 3847 3464 3893 3476
rect 3847 3288 3853 3464
rect 3887 3288 3893 3464
rect 3847 3276 3893 3288
rect 3965 3464 4011 3476
rect 3965 3288 3971 3464
rect 4005 3288 4011 3464
rect 3965 3276 4011 3288
rect 3026 3182 3062 3276
rect 3262 3182 3298 3276
rect 3498 3183 3534 3276
rect 3660 3228 3726 3235
rect 3660 3194 3676 3228
rect 3710 3194 3726 3228
rect 3660 3183 3726 3194
rect 3498 3182 3726 3183
rect 3026 3153 3726 3182
rect 3026 3152 3608 3153
rect 3146 3039 3180 3152
rect 3542 3111 3608 3152
rect 3542 3077 3558 3111
rect 3592 3077 3608 3111
rect 3542 3070 3608 3077
rect 3970 3071 4005 3276
rect 4177 3071 4244 3661
rect 5936 3638 5977 3670
rect 6223 3666 6233 3732
rect 6289 3666 6299 3732
rect 6969 3708 6979 3816
rect 7111 3753 7121 3816
rect 7111 3742 7123 3753
rect 7111 3708 7124 3742
rect 6979 3670 7124 3708
rect 7083 3642 7124 3670
rect 5352 3610 5622 3638
rect 5093 3544 5103 3610
rect 5169 3544 5179 3610
rect 5352 3548 5386 3610
rect 5588 3548 5622 3610
rect 5706 3610 5977 3638
rect 6494 3614 6764 3642
rect 5706 3548 5740 3610
rect 5942 3548 5977 3610
rect 6118 3598 6289 3614
rect 6118 3564 6249 3598
rect 6283 3564 6289 3598
rect 6118 3548 6289 3564
rect 6494 3552 6528 3614
rect 6730 3552 6764 3614
rect 6848 3614 7124 3642
rect 6848 3552 6882 3614
rect 7084 3552 7124 3614
rect 5228 3536 5274 3548
rect 5228 3160 5234 3536
rect 5268 3160 5274 3536
rect 5228 3148 5274 3160
rect 5346 3536 5392 3548
rect 5346 3160 5352 3536
rect 5386 3160 5392 3536
rect 5346 3148 5392 3160
rect 5464 3536 5510 3548
rect 5464 3160 5470 3536
rect 5504 3160 5510 3536
rect 5464 3148 5510 3160
rect 5582 3536 5628 3548
rect 5582 3160 5588 3536
rect 5622 3160 5628 3536
rect 5582 3148 5628 3160
rect 5700 3536 5746 3548
rect 5700 3160 5706 3536
rect 5740 3160 5746 3536
rect 5700 3148 5746 3160
rect 5818 3536 5864 3548
rect 5818 3160 5824 3536
rect 5858 3160 5864 3536
rect 5818 3148 5864 3160
rect 5936 3536 5982 3548
rect 5936 3160 5942 3536
rect 5976 3160 5982 3536
rect 5936 3148 5982 3160
rect 3970 3043 4244 3071
rect 3616 3039 4244 3043
rect 3140 3027 3186 3039
rect 3140 2651 3146 3027
rect 3180 2651 3186 3027
rect 3140 2639 3186 2651
rect 3258 3027 3304 3039
rect 3258 2651 3264 3027
rect 3298 2651 3304 3027
rect 3258 2639 3304 2651
rect 3376 3027 3422 3039
rect 3376 2651 3382 3027
rect 3416 2675 3422 3027
rect 3493 3027 3539 3039
rect 3493 2851 3499 3027
rect 3533 2851 3539 3027
rect 3493 2839 3539 2851
rect 3611 3027 4244 3039
rect 3611 2851 3617 3027
rect 3651 3014 4244 3027
rect 5234 3106 5268 3148
rect 5470 3106 5504 3148
rect 5234 3078 5504 3106
rect 5588 3107 5622 3148
rect 5824 3107 5858 3148
rect 5588 3078 5858 3107
rect 5234 3030 5268 3078
rect 3651 2851 3657 3014
rect 5234 3000 5297 3030
rect 3611 2839 3657 2851
rect 5262 2908 5297 3000
rect 5262 2872 5489 2908
rect 5759 2897 5769 2994
rect 5868 2897 5878 2994
rect 5942 2965 5976 3148
rect 5942 2911 6051 2965
rect 3499 2723 3534 2839
rect 5262 2765 5297 2872
rect 5423 2838 5489 2872
rect 5423 2804 5439 2838
rect 5473 2804 5489 2838
rect 5770 2896 5867 2897
rect 5770 2829 5827 2896
rect 5423 2798 5489 2804
rect 5664 2793 5933 2829
rect 5664 2765 5697 2793
rect 5900 2765 5933 2793
rect 6017 2765 6051 2911
rect 5138 2753 5184 2765
rect 3630 2723 3738 2733
rect 3499 2675 3630 2723
rect 3738 2690 3886 2696
rect 3416 2651 3630 2675
rect 3376 2639 3630 2651
rect 1011 2636 1118 2637
rect 1011 2635 1707 2636
rect 3382 2635 3630 2639
rect 1011 2634 2257 2635
rect 1011 2607 3018 2634
rect 1011 2601 3255 2607
rect 1011 2567 3205 2601
rect 3239 2567 3255 2601
rect 1011 2551 3255 2567
rect 3307 2601 3373 2607
rect 3307 2567 3323 2601
rect 3357 2567 3373 2601
rect 3556 2591 3630 2635
rect 3874 2623 3886 2690
rect 3738 2617 3886 2623
rect 3630 2581 3738 2591
rect 1011 2535 3018 2551
rect 1011 2534 2955 2535
rect 1011 2530 2490 2534
rect 1011 2529 2257 2530
rect 1011 2527 2098 2529
rect 1300 2119 2274 2148
rect 1300 2013 2122 2119
rect 2234 2106 2274 2119
rect 2234 2013 2276 2106
rect 1300 2002 2276 2013
rect 1300 2001 2274 2002
rect 316 1384 452 1404
rect 316 1322 352 1384
rect 412 1322 452 1384
rect 316 1294 452 1322
rect 12 1264 989 1294
rect 12 1158 44 1264
rect 248 1158 280 1264
rect 484 1158 516 1264
rect 720 1158 752 1264
rect 955 1158 989 1264
rect 5 1146 51 1158
rect 5 970 11 1146
rect 45 970 51 1146
rect 5 958 51 970
rect 123 1146 169 1158
rect 123 970 129 1146
rect 163 970 169 1146
rect 123 958 169 970
rect 241 1146 287 1158
rect 241 970 247 1146
rect 281 970 287 1146
rect 241 958 287 970
rect 359 1146 405 1158
rect 359 970 365 1146
rect 399 970 405 1146
rect 359 958 405 970
rect 477 1146 523 1158
rect 477 970 483 1146
rect 517 970 523 1146
rect 477 958 523 970
rect 595 1146 641 1158
rect 595 970 601 1146
rect 635 970 641 1146
rect 595 958 641 970
rect 713 1146 759 1158
rect 713 970 719 1146
rect 753 970 759 1146
rect 713 958 759 970
rect 831 1146 877 1158
rect 831 970 837 1146
rect 871 970 877 1146
rect 831 958 877 970
rect 949 1146 995 1158
rect 949 970 955 1146
rect 989 970 995 1146
rect 949 958 995 970
rect 1067 1146 1113 1158
rect 1067 970 1073 1146
rect 1107 970 1113 1146
rect 1067 958 1113 970
rect 128 864 164 958
rect 364 864 400 958
rect 600 865 636 958
rect 762 910 828 917
rect 762 876 778 910
rect 812 876 828 910
rect 762 865 828 876
rect 600 864 828 865
rect 128 835 828 864
rect 128 834 710 835
rect 248 721 282 834
rect 644 793 710 834
rect 644 759 660 793
rect 694 759 710 793
rect 644 752 710 759
rect 1072 725 1107 958
rect 1300 725 1420 2001
rect 2092 1008 2273 1038
rect 2092 898 2121 1008
rect 2239 994 2273 1008
rect 2239 898 2274 994
rect 2092 890 2274 898
rect 2092 888 2273 890
rect 718 721 1420 725
rect 242 709 288 721
rect 242 333 248 709
rect 282 333 288 709
rect 242 321 288 333
rect 360 709 406 721
rect 360 333 366 709
rect 400 333 406 709
rect 360 321 406 333
rect 478 709 524 721
rect 478 333 484 709
rect 518 360 524 709
rect 595 709 641 721
rect 595 533 601 709
rect 635 533 641 709
rect 595 526 641 533
rect 713 709 1420 721
rect 713 533 719 709
rect 753 696 1420 709
rect 753 533 759 696
rect 1003 617 1420 696
rect 2397 636 2490 2530
rect 2553 2471 3019 2493
rect 3307 2471 3373 2567
rect 5138 2577 5144 2753
rect 5178 2577 5184 2753
rect 5138 2565 5184 2577
rect 5256 2753 5302 2765
rect 5256 2577 5262 2753
rect 5296 2577 5302 2753
rect 5256 2565 5302 2577
rect 5374 2753 5420 2765
rect 5374 2577 5380 2753
rect 5414 2577 5420 2753
rect 5374 2565 5420 2577
rect 5492 2753 5538 2765
rect 5492 2577 5498 2753
rect 5532 2698 5538 2753
rect 5657 2753 5703 2765
rect 5657 2698 5663 2753
rect 5532 2610 5663 2698
rect 5532 2577 5538 2610
rect 5492 2565 5538 2577
rect 5657 2577 5663 2610
rect 5697 2577 5703 2753
rect 5657 2565 5703 2577
rect 5775 2753 5821 2765
rect 5775 2577 5781 2753
rect 5815 2577 5821 2753
rect 5775 2565 5821 2577
rect 5893 2753 5939 2765
rect 5893 2577 5899 2753
rect 5933 2577 5939 2753
rect 5893 2565 5939 2577
rect 6011 2753 6057 2765
rect 6011 2577 6017 2753
rect 6051 2577 6057 2753
rect 6011 2565 6057 2577
rect 5144 2526 5178 2565
rect 5380 2526 5414 2565
rect 5144 2491 5414 2526
rect 5781 2527 5814 2565
rect 6017 2527 6050 2565
rect 5781 2491 6050 2527
rect 2553 2423 3373 2471
rect 5178 2490 5414 2491
rect 2553 2392 3019 2423
rect 5178 2416 5310 2490
rect 2553 2136 2658 2392
rect 5168 2308 5178 2416
rect 5310 2308 5320 2416
rect 3390 2228 3469 2240
rect 2553 2030 2616 2136
rect 2728 2030 2738 2136
rect 3390 2132 3396 2228
rect 3320 2112 3396 2132
rect 3463 2132 3469 2228
rect 5205 2170 5211 2308
rect 5278 2170 5284 2308
rect 5205 2158 5284 2170
rect 3463 2112 3540 2132
rect 2553 2019 2702 2030
rect 2553 842 2658 2019
rect 3320 2004 3364 2112
rect 3496 2004 3540 2112
rect 3320 1962 3540 2004
rect 6118 1977 6180 3548
rect 6370 3540 6416 3552
rect 6370 3164 6376 3540
rect 6410 3164 6416 3540
rect 6370 3152 6416 3164
rect 6488 3540 6534 3552
rect 6488 3164 6494 3540
rect 6528 3164 6534 3540
rect 6488 3152 6534 3164
rect 6606 3540 6652 3552
rect 6606 3164 6612 3540
rect 6646 3164 6652 3540
rect 6606 3152 6652 3164
rect 6724 3540 6770 3552
rect 6724 3164 6730 3540
rect 6764 3164 6770 3540
rect 6724 3152 6770 3164
rect 6842 3540 6888 3552
rect 6842 3164 6848 3540
rect 6882 3164 6888 3540
rect 6842 3152 6888 3164
rect 6960 3540 7006 3552
rect 6960 3164 6966 3540
rect 7000 3164 7006 3540
rect 6960 3152 7006 3164
rect 7078 3540 7124 3552
rect 7078 3164 7084 3540
rect 7118 3164 7124 3540
rect 7078 3152 7124 3164
rect 6376 3110 6410 3152
rect 6612 3110 6646 3152
rect 6376 3082 6646 3110
rect 6730 3111 6764 3152
rect 6966 3111 7000 3152
rect 6730 3082 7000 3111
rect 6376 3034 6410 3082
rect 6376 3004 6439 3034
rect 6404 2912 6439 3004
rect 6911 2974 7011 2995
rect 6911 2920 6925 2974
rect 6990 2920 7011 2974
rect 6911 2915 7011 2920
rect 7084 2969 7118 3152
rect 7084 2915 7193 2969
rect 8810 2930 8991 5100
rect 13463 5193 13509 5205
rect 13463 4817 13469 5193
rect 13503 4817 13509 5193
rect 13463 4805 13509 4817
rect 13581 5193 13627 5205
rect 13581 4817 13587 5193
rect 13621 4817 13627 5193
rect 13581 4805 13627 4817
rect 13699 5193 13745 5205
rect 13699 4817 13705 5193
rect 13739 4844 13745 5193
rect 13816 5193 13862 5205
rect 13816 5017 13822 5193
rect 13856 5017 13862 5193
rect 13816 5010 13862 5017
rect 13934 5193 15641 5205
rect 13934 5017 13940 5193
rect 13974 5180 15641 5193
rect 13974 5017 13980 5180
rect 14224 5100 15641 5180
rect 14228 5099 15641 5100
rect 13816 5005 13865 5010
rect 13934 5005 13980 5017
rect 13822 4844 13865 5005
rect 13739 4817 13865 4844
rect 13699 4805 13865 4817
rect 13705 4801 13865 4805
rect 13370 4773 13443 4774
rect 13370 4768 13578 4773
rect 13370 4722 13382 4768
rect 13431 4767 13578 4768
rect 13431 4733 13528 4767
rect 13562 4733 13578 4767
rect 13431 4722 13578 4733
rect 13370 4717 13578 4722
rect 13630 4767 13696 4773
rect 13630 4733 13646 4767
rect 13680 4733 13696 4767
rect 13370 4716 13443 4717
rect 13630 4688 13696 4733
rect 13233 4680 13696 4688
rect 13233 4648 13697 4680
rect 13789 4664 13865 4801
rect 13233 4229 13279 4648
rect 13785 4604 13795 4664
rect 13857 4604 13867 4664
rect 13219 4175 13229 4229
rect 13286 4175 13296 4229
rect 15460 4191 15641 5099
rect 20117 4838 20123 5214
rect 20157 4838 20163 5214
rect 20117 4826 20163 4838
rect 20235 5214 20281 5226
rect 20235 4838 20241 5214
rect 20275 4838 20281 5214
rect 20235 4826 20281 4838
rect 20353 5214 20399 5226
rect 20353 4838 20359 5214
rect 20393 4865 20399 5214
rect 20470 5214 20516 5226
rect 20470 5038 20476 5214
rect 20510 5038 20516 5214
rect 20470 5031 20516 5038
rect 20588 5214 22267 5226
rect 20588 5038 20594 5214
rect 20628 5201 22267 5214
rect 20628 5038 20634 5201
rect 20878 5120 22267 5201
rect 20470 5026 20519 5031
rect 20588 5026 20634 5038
rect 20476 4865 20519 5026
rect 20393 4838 20519 4865
rect 20353 4826 20519 4838
rect 20359 4822 20519 4826
rect 19977 4794 20062 4796
rect 19977 4790 20232 4794
rect 19977 4742 19989 4790
rect 20050 4788 20232 4790
rect 20050 4754 20182 4788
rect 20216 4754 20232 4788
rect 20050 4742 20232 4754
rect 19977 4738 20232 4742
rect 20284 4788 20350 4794
rect 20284 4754 20300 4788
rect 20334 4754 20350 4788
rect 19977 4736 20062 4738
rect 20284 4708 20350 4754
rect 20078 4701 20350 4708
rect 20078 4700 20351 4701
rect 20078 4662 20091 4700
rect 20136 4669 20351 4700
rect 20443 4685 20519 4822
rect 20136 4662 20150 4669
rect 20078 4653 20150 4662
rect 20439 4625 20449 4685
rect 20511 4625 20521 4685
rect 22086 4259 22267 5120
rect 12410 4018 12489 4030
rect 9927 3967 10006 3979
rect 9927 3870 9933 3967
rect 9855 3850 9933 3870
rect 10000 3870 10006 3967
rect 12410 3904 12416 4018
rect 12483 3904 12489 4018
rect 13554 4020 13633 4032
rect 13554 3904 13560 4020
rect 13627 3904 13633 4020
rect 10000 3850 10075 3870
rect 9855 3742 9899 3850
rect 10031 3742 10075 3850
rect 11652 3808 11708 3816
rect 9855 3700 10075 3742
rect 10726 3800 11708 3808
rect 10726 3766 11668 3800
rect 11702 3766 11708 3800
rect 12371 3796 12381 3904
rect 12513 3841 12523 3904
rect 12513 3830 12525 3841
rect 12513 3796 12526 3830
rect 12782 3820 12838 3822
rect 10726 3750 11708 3766
rect 12381 3758 12526 3796
rect 10726 3749 11705 3750
rect 9459 3670 10436 3700
rect 9459 3564 9491 3670
rect 9695 3564 9727 3670
rect 9931 3564 9963 3670
rect 10167 3564 10199 3670
rect 10402 3564 10436 3670
rect 9452 3552 9498 3564
rect 9452 3376 9458 3552
rect 9492 3376 9498 3552
rect 9452 3364 9498 3376
rect 9570 3552 9616 3564
rect 9570 3376 9576 3552
rect 9610 3376 9616 3552
rect 9570 3364 9616 3376
rect 9688 3552 9734 3564
rect 9688 3376 9694 3552
rect 9728 3376 9734 3552
rect 9688 3364 9734 3376
rect 9806 3552 9852 3564
rect 9806 3376 9812 3552
rect 9846 3376 9852 3552
rect 9806 3364 9852 3376
rect 9924 3552 9970 3564
rect 9924 3376 9930 3552
rect 9964 3376 9970 3552
rect 9924 3364 9970 3376
rect 10042 3552 10088 3564
rect 10042 3376 10048 3552
rect 10082 3376 10088 3552
rect 10042 3364 10088 3376
rect 10160 3552 10206 3564
rect 10160 3376 10166 3552
rect 10200 3376 10206 3552
rect 10160 3364 10206 3376
rect 10278 3552 10324 3564
rect 10278 3376 10284 3552
rect 10318 3376 10324 3552
rect 10278 3364 10324 3376
rect 10396 3552 10442 3564
rect 10396 3376 10402 3552
rect 10436 3376 10442 3552
rect 10396 3364 10442 3376
rect 10514 3552 10560 3564
rect 10514 3376 10520 3552
rect 10554 3376 10560 3552
rect 10514 3364 10560 3376
rect 9575 3270 9611 3364
rect 9811 3270 9847 3364
rect 10047 3271 10083 3364
rect 10209 3316 10275 3323
rect 10209 3282 10225 3316
rect 10259 3282 10275 3316
rect 10209 3271 10275 3282
rect 10047 3270 10275 3271
rect 9575 3241 10275 3270
rect 9575 3240 10157 3241
rect 9695 3127 9729 3240
rect 10091 3199 10157 3240
rect 10091 3165 10107 3199
rect 10141 3165 10157 3199
rect 10091 3158 10157 3165
rect 10519 3159 10554 3364
rect 10726 3159 10793 3749
rect 12485 3726 12526 3758
rect 12772 3754 12782 3820
rect 12838 3754 12848 3820
rect 13518 3796 13528 3904
rect 13660 3841 13670 3904
rect 13660 3830 13672 3841
rect 13660 3796 13673 3830
rect 13528 3758 13673 3796
rect 13632 3730 13673 3758
rect 11901 3698 12171 3726
rect 11642 3632 11652 3698
rect 11718 3632 11728 3698
rect 11901 3636 11935 3698
rect 12137 3636 12171 3698
rect 12255 3698 12526 3726
rect 13043 3702 13313 3730
rect 12255 3636 12289 3698
rect 12491 3636 12526 3698
rect 12667 3686 12838 3702
rect 12667 3652 12798 3686
rect 12832 3652 12838 3686
rect 12667 3636 12838 3652
rect 13043 3640 13077 3702
rect 13279 3640 13313 3702
rect 13397 3702 13673 3730
rect 13397 3640 13431 3702
rect 13633 3640 13673 3702
rect 11777 3624 11823 3636
rect 11777 3248 11783 3624
rect 11817 3248 11823 3624
rect 11777 3236 11823 3248
rect 11895 3624 11941 3636
rect 11895 3248 11901 3624
rect 11935 3248 11941 3624
rect 11895 3236 11941 3248
rect 12013 3624 12059 3636
rect 12013 3248 12019 3624
rect 12053 3248 12059 3624
rect 12013 3236 12059 3248
rect 12131 3624 12177 3636
rect 12131 3248 12137 3624
rect 12171 3248 12177 3624
rect 12131 3236 12177 3248
rect 12249 3624 12295 3636
rect 12249 3248 12255 3624
rect 12289 3248 12295 3624
rect 12249 3236 12295 3248
rect 12367 3624 12413 3636
rect 12367 3248 12373 3624
rect 12407 3248 12413 3624
rect 12367 3236 12413 3248
rect 12485 3624 12531 3636
rect 12485 3248 12491 3624
rect 12525 3248 12531 3624
rect 12485 3236 12531 3248
rect 10519 3131 10793 3159
rect 10165 3127 10793 3131
rect 6404 2876 6631 2912
rect 6404 2769 6439 2876
rect 6565 2842 6631 2876
rect 6565 2808 6581 2842
rect 6615 2808 6631 2842
rect 6912 2900 7009 2915
rect 6912 2833 6969 2900
rect 6565 2802 6631 2808
rect 6806 2797 7075 2833
rect 6806 2769 6839 2797
rect 7042 2769 7075 2797
rect 7159 2769 7193 2915
rect 6280 2757 6326 2769
rect 6280 2581 6286 2757
rect 6320 2581 6326 2757
rect 6280 2569 6326 2581
rect 6398 2757 6444 2769
rect 6398 2581 6404 2757
rect 6438 2581 6444 2757
rect 6398 2569 6444 2581
rect 6516 2757 6562 2769
rect 6516 2581 6522 2757
rect 6556 2581 6562 2757
rect 6516 2569 6562 2581
rect 6634 2757 6680 2769
rect 6634 2581 6640 2757
rect 6674 2702 6680 2757
rect 6799 2757 6845 2769
rect 6799 2702 6805 2757
rect 6674 2614 6805 2702
rect 6674 2581 6680 2614
rect 6634 2569 6680 2581
rect 6799 2581 6805 2614
rect 6839 2581 6845 2757
rect 6799 2569 6845 2581
rect 6917 2757 6963 2769
rect 6917 2581 6923 2757
rect 6957 2581 6963 2757
rect 6917 2569 6963 2581
rect 7035 2757 7081 2769
rect 7035 2581 7041 2757
rect 7075 2581 7081 2757
rect 7035 2569 7081 2581
rect 7153 2757 7199 2769
rect 7153 2581 7159 2757
rect 7193 2581 7199 2757
rect 8811 2722 8991 2930
rect 9689 3115 9735 3127
rect 9689 2739 9695 3115
rect 9729 2739 9735 3115
rect 9689 2727 9735 2739
rect 9807 3115 9853 3127
rect 9807 2739 9813 3115
rect 9847 2739 9853 3115
rect 9807 2727 9853 2739
rect 9925 3115 9971 3127
rect 9925 2739 9931 3115
rect 9965 2763 9971 3115
rect 10042 3115 10088 3127
rect 10042 2939 10048 3115
rect 10082 2939 10088 3115
rect 10042 2927 10088 2939
rect 10160 3115 10793 3127
rect 10160 2939 10166 3115
rect 10200 3102 10793 3115
rect 11783 3194 11817 3236
rect 12019 3194 12053 3236
rect 11783 3166 12053 3194
rect 12137 3195 12171 3236
rect 12373 3195 12407 3236
rect 12137 3166 12407 3195
rect 11783 3118 11817 3166
rect 10200 2939 10206 3102
rect 11783 3088 11846 3118
rect 10160 2927 10206 2939
rect 11811 2996 11846 3088
rect 11811 2960 12038 2996
rect 12308 2985 12318 3082
rect 12417 2985 12427 3082
rect 12491 3053 12525 3236
rect 12491 2999 12600 3053
rect 10048 2811 10083 2927
rect 11811 2853 11846 2960
rect 11972 2926 12038 2960
rect 11972 2892 11988 2926
rect 12022 2892 12038 2926
rect 12319 2984 12416 2985
rect 12319 2917 12376 2984
rect 11972 2886 12038 2892
rect 12213 2881 12482 2917
rect 12213 2853 12246 2881
rect 12449 2853 12482 2881
rect 12566 2853 12600 2999
rect 11687 2841 11733 2853
rect 10179 2811 10287 2821
rect 10048 2763 10179 2811
rect 10287 2772 10432 2778
rect 9965 2739 10179 2763
rect 9925 2727 10179 2739
rect 9931 2723 10179 2727
rect 8811 2695 9567 2722
rect 8811 2689 9804 2695
rect 8811 2655 9754 2689
rect 9788 2655 9804 2689
rect 8811 2639 9804 2655
rect 9856 2689 9922 2695
rect 9856 2655 9872 2689
rect 9906 2655 9922 2689
rect 10105 2679 10179 2723
rect 10420 2705 10432 2772
rect 10287 2699 10432 2705
rect 10179 2669 10287 2679
rect 8811 2623 9567 2639
rect 8811 2622 9504 2623
rect 8811 2618 9039 2622
rect 7153 2569 7199 2581
rect 6286 2530 6320 2569
rect 6522 2530 6556 2569
rect 6286 2494 6556 2530
rect 6923 2531 6956 2569
rect 7159 2531 7192 2569
rect 6923 2495 7192 2531
rect 6286 2493 6452 2494
rect 6320 2414 6452 2493
rect 6310 2306 6320 2414
rect 6452 2306 6462 2414
rect 6343 2172 6349 2306
rect 6416 2172 6422 2306
rect 6343 2160 6422 2172
rect 8310 2207 8823 2239
rect 8310 2101 8671 2207
rect 8783 2194 8823 2207
rect 8783 2101 8825 2194
rect 8310 2090 8825 2101
rect 8310 2089 8823 2090
rect 2924 1932 3901 1962
rect 6118 1960 6181 1977
rect 6043 1956 6181 1960
rect 2924 1826 2956 1932
rect 3160 1826 3192 1932
rect 3396 1826 3428 1932
rect 3632 1826 3664 1932
rect 3867 1826 3901 1932
rect 4211 1922 6181 1956
rect 4209 1893 6181 1922
rect 4209 1877 4255 1893
rect 6043 1891 6181 1893
rect 2917 1814 2963 1826
rect 2917 1638 2923 1814
rect 2957 1638 2963 1814
rect 2917 1626 2963 1638
rect 3035 1814 3081 1826
rect 3035 1638 3041 1814
rect 3075 1638 3081 1814
rect 3035 1626 3081 1638
rect 3153 1814 3199 1826
rect 3153 1638 3159 1814
rect 3193 1638 3199 1814
rect 3153 1626 3199 1638
rect 3271 1814 3317 1826
rect 3271 1638 3277 1814
rect 3311 1638 3317 1814
rect 3271 1626 3317 1638
rect 3389 1814 3435 1826
rect 3389 1638 3395 1814
rect 3429 1638 3435 1814
rect 3389 1626 3435 1638
rect 3507 1814 3553 1826
rect 3507 1638 3513 1814
rect 3547 1638 3553 1814
rect 3507 1626 3553 1638
rect 3625 1814 3671 1826
rect 3625 1638 3631 1814
rect 3665 1638 3671 1814
rect 3625 1626 3671 1638
rect 3743 1814 3789 1826
rect 3743 1638 3749 1814
rect 3783 1638 3789 1814
rect 3743 1626 3789 1638
rect 3861 1814 3907 1826
rect 3861 1638 3867 1814
rect 3901 1638 3907 1814
rect 3861 1626 3907 1638
rect 3979 1814 4025 1826
rect 3979 1638 3985 1814
rect 4019 1638 4025 1814
rect 3979 1626 4025 1638
rect 3040 1532 3076 1626
rect 3276 1532 3312 1626
rect 3512 1533 3548 1626
rect 3674 1578 3740 1585
rect 3674 1544 3690 1578
rect 3724 1544 3740 1578
rect 3674 1533 3740 1544
rect 3512 1532 3740 1533
rect 3040 1503 3740 1532
rect 3040 1502 3622 1503
rect 3160 1389 3194 1502
rect 3556 1461 3622 1502
rect 3556 1427 3572 1461
rect 3606 1427 3622 1461
rect 3556 1420 3622 1427
rect 3984 1408 4019 1626
rect 4208 1425 4255 1877
rect 7102 1886 7181 1898
rect 7102 1769 7108 1886
rect 7175 1769 7181 1886
rect 5167 1661 5177 1769
rect 5309 1661 5319 1769
rect 7065 1661 7075 1769
rect 7207 1661 7217 1769
rect 5177 1621 5309 1661
rect 7075 1621 7207 1661
rect 5176 1555 5309 1621
rect 7074 1555 7207 1621
rect 4505 1512 5978 1555
rect 4208 1409 4254 1425
rect 4173 1408 4254 1409
rect 3984 1393 4254 1408
rect 3630 1389 4254 1393
rect 3154 1377 3200 1389
rect 2889 899 2899 1017
rect 3017 985 3027 1017
rect 3154 1001 3160 1377
rect 3194 1001 3200 1377
rect 3154 989 3200 1001
rect 3272 1377 3318 1389
rect 3272 1001 3278 1377
rect 3312 1001 3318 1377
rect 3272 989 3318 1001
rect 3390 1377 3436 1389
rect 3390 1001 3396 1377
rect 3430 1025 3436 1377
rect 3507 1377 3553 1389
rect 3507 1201 3513 1377
rect 3547 1201 3553 1377
rect 3507 1189 3553 1201
rect 3625 1377 4254 1389
rect 3625 1201 3631 1377
rect 3665 1365 4254 1377
rect 3665 1364 3907 1365
rect 3665 1201 3671 1364
rect 4173 1363 4254 1365
rect 4505 1209 4539 1512
rect 4871 1409 4905 1512
rect 5107 1409 5141 1512
rect 5343 1409 5377 1512
rect 5579 1409 5613 1512
rect 4865 1397 4911 1409
rect 3625 1189 3671 1201
rect 4381 1197 4427 1209
rect 3513 1073 3548 1189
rect 3644 1073 3752 1083
rect 3513 1025 3644 1073
rect 3752 1040 3901 1046
rect 3430 1001 3644 1025
rect 3390 989 3644 1001
rect 3396 985 3644 989
rect 3017 957 3032 985
rect 3017 951 3269 957
rect 3017 917 3219 951
rect 3253 917 3269 951
rect 3017 901 3269 917
rect 3321 951 3387 957
rect 3321 917 3337 951
rect 3371 917 3387 951
rect 3570 941 3644 985
rect 3889 973 3901 1040
rect 4381 1021 4387 1197
rect 4421 1021 4427 1197
rect 4381 1009 4427 1021
rect 4499 1197 4545 1209
rect 4499 1021 4505 1197
rect 4539 1021 4545 1197
rect 4499 1009 4545 1021
rect 4617 1197 4663 1209
rect 4617 1021 4623 1197
rect 4657 1021 4663 1197
rect 4617 1009 4663 1021
rect 4735 1197 4781 1209
rect 4865 1197 4871 1397
rect 4735 1021 4741 1197
rect 4775 1021 4871 1197
rect 4905 1021 4911 1397
rect 4735 1009 4781 1021
rect 4865 1009 4911 1021
rect 4983 1397 5029 1409
rect 4983 1021 4989 1397
rect 5023 1021 5029 1397
rect 4983 1009 5029 1021
rect 5101 1397 5147 1409
rect 5101 1021 5107 1397
rect 5141 1021 5147 1397
rect 5101 1009 5147 1021
rect 5219 1397 5265 1409
rect 5219 1021 5225 1397
rect 5259 1021 5265 1397
rect 5219 1009 5265 1021
rect 5337 1397 5383 1409
rect 5337 1021 5343 1397
rect 5377 1021 5383 1397
rect 5337 1009 5383 1021
rect 5455 1397 5501 1409
rect 5455 1021 5461 1397
rect 5495 1021 5501 1397
rect 5455 1009 5501 1021
rect 5573 1397 5619 1409
rect 5573 1021 5579 1397
rect 5613 1197 5619 1397
rect 5944 1209 5978 1512
rect 6403 1512 7876 1555
rect 6403 1209 6437 1512
rect 6769 1409 6803 1512
rect 7005 1409 7039 1512
rect 7241 1409 7275 1512
rect 7477 1409 7511 1512
rect 6763 1397 6809 1409
rect 5702 1197 5748 1209
rect 5613 1021 5708 1197
rect 5742 1021 5748 1197
rect 5573 1009 5619 1021
rect 5702 1009 5748 1021
rect 5820 1197 5866 1209
rect 5820 1021 5826 1197
rect 5860 1021 5866 1197
rect 5820 1009 5866 1021
rect 5938 1197 5984 1209
rect 5938 1021 5944 1197
rect 5978 1021 5984 1197
rect 5938 1009 5984 1021
rect 6056 1197 6102 1209
rect 6056 1021 6062 1197
rect 6096 1021 6102 1197
rect 6056 1009 6102 1021
rect 6279 1197 6325 1209
rect 6279 1021 6285 1197
rect 6319 1021 6325 1197
rect 6279 1009 6325 1021
rect 6397 1197 6443 1209
rect 6397 1021 6403 1197
rect 6437 1021 6443 1197
rect 6397 1009 6443 1021
rect 6515 1197 6561 1209
rect 6515 1021 6521 1197
rect 6555 1021 6561 1197
rect 6515 1009 6561 1021
rect 6633 1197 6679 1209
rect 6763 1197 6769 1397
rect 6633 1021 6639 1197
rect 6673 1021 6769 1197
rect 6803 1021 6809 1397
rect 6633 1009 6679 1021
rect 6763 1009 6809 1021
rect 6881 1397 6927 1409
rect 6881 1021 6887 1397
rect 6921 1021 6927 1397
rect 6881 1009 6927 1021
rect 6999 1397 7045 1409
rect 6999 1021 7005 1397
rect 7039 1021 7045 1397
rect 6999 1009 7045 1021
rect 7117 1397 7163 1409
rect 7117 1021 7123 1397
rect 7157 1021 7163 1397
rect 7117 1009 7163 1021
rect 7235 1397 7281 1409
rect 7235 1021 7241 1397
rect 7275 1021 7281 1397
rect 7235 1009 7281 1021
rect 7353 1397 7399 1409
rect 7353 1021 7359 1397
rect 7393 1021 7399 1397
rect 7353 1009 7399 1021
rect 7471 1397 7517 1409
rect 7471 1021 7477 1397
rect 7511 1197 7517 1397
rect 7842 1209 7876 1512
rect 7600 1197 7646 1209
rect 7511 1021 7606 1197
rect 7640 1021 7646 1197
rect 7471 1009 7517 1021
rect 7600 1009 7646 1021
rect 7718 1197 7764 1209
rect 7718 1021 7724 1197
rect 7758 1021 7764 1197
rect 7718 1009 7764 1021
rect 7836 1197 7882 1209
rect 7836 1021 7842 1197
rect 7876 1021 7882 1197
rect 7836 1009 7882 1021
rect 7954 1197 8000 1209
rect 7954 1021 7960 1197
rect 7994 1021 8000 1197
rect 7954 1009 8000 1021
rect 3752 967 3901 973
rect 4387 975 4421 1009
rect 4989 975 5023 1009
rect 5225 975 5259 1009
rect 3644 931 3752 941
rect 4387 940 4546 975
rect 4989 940 5259 975
rect 5826 975 5860 1009
rect 6062 975 6096 1009
rect 5826 940 6096 975
rect 6285 975 6319 1009
rect 6887 975 6921 1009
rect 7123 975 7157 1009
rect 6285 940 6444 975
rect 6887 940 7157 975
rect 7724 975 7758 1009
rect 7960 975 7994 1009
rect 7724 940 7994 975
rect 3017 899 3032 901
rect 2932 885 3032 899
rect 2932 842 3032 843
rect 2553 821 3032 842
rect 3321 821 3387 917
rect 2553 773 3387 821
rect 2553 744 3032 773
rect 2553 742 2658 744
rect 2932 743 3032 744
rect 2386 557 2396 636
rect 2489 557 2499 636
rect 3388 622 3467 634
rect 595 521 644 526
rect 713 521 759 533
rect 601 360 644 521
rect 518 333 644 360
rect 478 321 644 333
rect 484 317 644 321
rect -352 283 357 289
rect -352 249 307 283
rect 341 249 357 283
rect -352 233 357 249
rect 409 283 475 289
rect 409 249 425 283
rect 459 249 475 283
rect -1124 195 -857 200
rect -1124 91 -955 195
rect -868 91 -857 195
rect -1124 85 -857 91
rect -352 -5457 -247 233
rect 409 204 475 249
rect -189 196 475 204
rect -189 190 476 196
rect -189 94 -158 190
rect -81 164 476 190
rect 568 180 644 317
rect -81 94 -71 164
rect 564 120 574 180
rect 636 120 646 180
rect -189 -2697 -71 94
rect 2397 -617 2490 557
rect 3388 528 3394 622
rect 3315 508 3394 528
rect 3461 528 3467 622
rect 3461 508 3535 528
rect 3315 400 3359 508
rect 3491 400 3535 508
rect 3315 358 3535 400
rect 2919 328 3896 358
rect 2919 222 2951 328
rect 3155 222 3187 328
rect 3391 222 3423 328
rect 3627 222 3659 328
rect 3862 222 3896 328
rect 2912 210 2958 222
rect 2912 34 2918 210
rect 2952 34 2958 210
rect 2912 22 2958 34
rect 3030 210 3076 222
rect 3030 34 3036 210
rect 3070 34 3076 210
rect 3030 22 3076 34
rect 3148 210 3194 222
rect 3148 34 3154 210
rect 3188 34 3194 210
rect 3148 22 3194 34
rect 3266 210 3312 222
rect 3266 34 3272 210
rect 3306 34 3312 210
rect 3266 22 3312 34
rect 3384 210 3430 222
rect 3384 34 3390 210
rect 3424 34 3430 210
rect 3384 22 3430 34
rect 3502 210 3548 222
rect 3502 34 3508 210
rect 3542 34 3548 210
rect 3502 22 3548 34
rect 3620 210 3666 222
rect 3620 34 3626 210
rect 3660 34 3666 210
rect 3620 22 3666 34
rect 3738 210 3784 222
rect 3738 34 3744 210
rect 3778 34 3784 210
rect 3738 22 3784 34
rect 3856 210 3902 222
rect 3856 34 3862 210
rect 3896 34 3902 210
rect 3856 22 3902 34
rect 3974 210 4020 222
rect 3974 34 3980 210
rect 4014 34 4020 210
rect 3974 22 4020 34
rect 4512 156 4546 940
rect 5225 878 5259 940
rect 4814 840 5556 878
rect 4814 716 4848 840
rect 5050 716 5084 840
rect 5286 716 5320 840
rect 5522 716 5556 840
rect 5812 733 5822 799
rect 5885 733 5895 799
rect 4808 704 4854 716
rect 4808 328 4814 704
rect 4848 328 4854 704
rect 4808 316 4854 328
rect 4926 704 4972 716
rect 4926 328 4932 704
rect 4966 328 4972 704
rect 4926 316 4972 328
rect 5044 704 5090 716
rect 5044 328 5050 704
rect 5084 328 5090 704
rect 5044 316 5090 328
rect 5162 704 5208 716
rect 5162 328 5168 704
rect 5202 328 5208 704
rect 5162 316 5208 328
rect 5280 704 5326 716
rect 5280 328 5286 704
rect 5320 328 5326 704
rect 5280 316 5326 328
rect 5398 704 5444 716
rect 5398 328 5404 704
rect 5438 328 5444 704
rect 5398 316 5444 328
rect 5516 704 5562 716
rect 5516 328 5522 704
rect 5556 328 5562 704
rect 5516 316 5562 328
rect 5928 157 5962 940
rect 5655 156 5962 157
rect 4512 151 4828 156
rect 5542 151 5962 156
rect 4512 140 4895 151
rect 4512 113 4844 140
rect 3035 -72 3071 22
rect 3271 -72 3307 22
rect 3507 -71 3543 22
rect 3669 -26 3735 -19
rect 3669 -60 3685 -26
rect 3719 -60 3735 -26
rect 3669 -71 3735 -60
rect 3507 -72 3735 -71
rect 3035 -101 3735 -72
rect 3035 -102 3617 -101
rect 3155 -215 3189 -102
rect 3551 -143 3617 -102
rect 3551 -177 3567 -143
rect 3601 -177 3617 -143
rect 3551 -184 3617 -177
rect 3979 -211 4014 22
rect 4512 -16 4546 113
rect 4828 106 4844 113
rect 4878 106 4895 140
rect 4828 100 4895 106
rect 5475 140 5962 151
rect 5475 106 5492 140
rect 5526 113 5962 140
rect 5526 106 5542 113
rect 5655 112 5962 113
rect 5475 100 5542 106
rect 4653 73 4709 85
rect 4653 39 4659 73
rect 4693 72 4709 73
rect 5766 72 5822 84
rect 4693 56 5160 72
rect 4693 39 5110 56
rect 4653 23 5110 39
rect 5094 22 5110 23
rect 5144 22 5160 56
rect 5094 15 5160 22
rect 5212 57 5782 72
rect 5212 23 5228 57
rect 5262 38 5782 57
rect 5816 38 5822 72
rect 5262 23 5822 38
rect 5212 13 5279 23
rect 5766 22 5822 23
rect 5928 -16 5962 112
rect 6410 156 6444 940
rect 7123 878 7157 940
rect 6712 840 7454 878
rect 6712 716 6746 840
rect 6948 716 6982 840
rect 7184 716 7218 840
rect 7420 716 7454 840
rect 6706 704 6752 716
rect 6706 328 6712 704
rect 6746 328 6752 704
rect 6706 316 6752 328
rect 6824 704 6870 716
rect 6824 328 6830 704
rect 6864 328 6870 704
rect 6824 316 6870 328
rect 6942 704 6988 716
rect 6942 328 6948 704
rect 6982 328 6988 704
rect 6942 316 6988 328
rect 7060 704 7106 716
rect 7060 328 7066 704
rect 7100 328 7106 704
rect 7060 316 7106 328
rect 7178 704 7224 716
rect 7178 328 7184 704
rect 7218 328 7224 704
rect 7178 316 7224 328
rect 7296 704 7342 716
rect 7296 328 7302 704
rect 7336 328 7342 704
rect 7296 316 7342 328
rect 7414 704 7460 716
rect 7414 328 7420 704
rect 7454 328 7460 704
rect 7414 316 7460 328
rect 7826 157 7860 940
rect 7438 156 7507 157
rect 7553 156 7860 157
rect 6410 151 6726 156
rect 7438 152 7860 156
rect 6410 140 6793 151
rect 6410 113 6742 140
rect 6410 -16 6444 113
rect 6726 106 6742 113
rect 6776 106 6793 140
rect 6726 100 6793 106
rect 7371 141 7860 152
rect 7371 107 7388 141
rect 7422 113 7860 141
rect 7422 107 7438 113
rect 7553 112 7860 113
rect 7371 101 7438 107
rect 6551 73 6607 85
rect 6551 39 6557 73
rect 6591 72 6607 73
rect 7664 72 7720 84
rect 6591 56 7058 72
rect 6591 39 7008 56
rect 6551 23 7008 39
rect 6992 22 7008 23
rect 7042 22 7058 56
rect 6992 15 7058 22
rect 7110 57 7680 72
rect 7110 23 7126 57
rect 7160 38 7680 57
rect 7714 38 7720 72
rect 7160 23 7720 38
rect 7110 13 7177 23
rect 7664 22 7720 23
rect 7826 -16 7860 112
rect 7941 762 8008 786
rect 7941 728 7958 762
rect 7992 728 8008 762
rect 3625 -215 4014 -211
rect 3149 -227 3195 -215
rect 3149 -603 3155 -227
rect 3189 -603 3195 -227
rect 3149 -615 3195 -603
rect 3267 -227 3313 -215
rect 3267 -603 3273 -227
rect 3307 -603 3313 -227
rect 3267 -615 3313 -603
rect 3385 -227 3431 -215
rect 3385 -603 3391 -227
rect 3425 -579 3431 -227
rect 3502 -227 3548 -215
rect 3502 -403 3508 -227
rect 3542 -403 3548 -227
rect 3502 -415 3548 -403
rect 3620 -227 4014 -215
rect 4506 -28 4552 -16
rect 4506 -204 4512 -28
rect 4546 -204 4552 -28
rect 4506 -216 4552 -204
rect 4624 -28 4670 -16
rect 4624 -204 4630 -28
rect 4664 -204 4670 -28
rect 4624 -216 4670 -204
rect 4926 -28 4972 -16
rect 3620 -403 3626 -227
rect 3660 -240 4014 -227
rect 3660 -403 3666 -240
rect 3936 -243 4014 -240
rect 3936 -295 3946 -243
rect 4009 -295 4019 -243
rect 3941 -301 4014 -295
rect 3620 -415 3666 -403
rect 3508 -531 3543 -415
rect 4629 -510 4663 -216
rect 4926 -404 4932 -28
rect 4966 -404 4972 -28
rect 4926 -416 4972 -404
rect 5044 -28 5090 -16
rect 5044 -404 5050 -28
rect 5084 -404 5090 -28
rect 5044 -416 5090 -404
rect 5162 -28 5208 -16
rect 5162 -404 5168 -28
rect 5202 -404 5208 -28
rect 5162 -416 5208 -404
rect 5280 -28 5326 -16
rect 5280 -404 5286 -28
rect 5320 -404 5326 -28
rect 5280 -416 5326 -404
rect 5398 -28 5444 -16
rect 5398 -404 5404 -28
rect 5438 -404 5444 -28
rect 5804 -28 5850 -16
rect 5804 -204 5810 -28
rect 5844 -204 5850 -28
rect 5804 -216 5850 -204
rect 5922 -28 5968 -16
rect 5922 -204 5928 -28
rect 5962 -204 5968 -28
rect 5922 -216 5968 -204
rect 6404 -28 6450 -16
rect 6404 -204 6410 -28
rect 6444 -204 6450 -28
rect 6404 -216 6450 -204
rect 6522 -28 6568 -16
rect 6522 -204 6528 -28
rect 6562 -204 6568 -28
rect 6522 -216 6568 -204
rect 6824 -28 6870 -16
rect 5398 -416 5444 -404
rect 5286 -510 5320 -416
rect 5810 -510 5843 -216
rect 3639 -531 3747 -521
rect 3508 -579 3639 -531
rect 4629 -542 5843 -510
rect 6527 -510 6561 -216
rect 6824 -404 6830 -28
rect 6864 -404 6870 -28
rect 6824 -416 6870 -404
rect 6942 -28 6988 -16
rect 6942 -404 6948 -28
rect 6982 -404 6988 -28
rect 6942 -416 6988 -404
rect 7060 -28 7106 -16
rect 7060 -404 7066 -28
rect 7100 -404 7106 -28
rect 7060 -416 7106 -404
rect 7178 -28 7224 -16
rect 7178 -404 7184 -28
rect 7218 -404 7224 -28
rect 7178 -416 7224 -404
rect 7296 -28 7342 -16
rect 7296 -404 7302 -28
rect 7336 -404 7342 -28
rect 7702 -28 7748 -16
rect 7702 -204 7708 -28
rect 7742 -204 7748 -28
rect 7702 -216 7748 -204
rect 7820 -28 7866 -16
rect 7820 -204 7826 -28
rect 7860 -204 7866 -28
rect 7820 -216 7866 -204
rect 7296 -416 7342 -404
rect 7184 -510 7218 -416
rect 7708 -510 7741 -216
rect 6527 -542 7741 -510
rect 3747 -568 3899 -562
rect 3425 -603 3639 -579
rect 3385 -615 3639 -603
rect 2397 -619 2982 -617
rect 3391 -619 3639 -615
rect 2397 -647 3027 -619
rect 2397 -653 3264 -647
rect 2397 -687 3214 -653
rect 3248 -687 3264 -653
rect 2397 -703 3264 -687
rect 3316 -653 3382 -647
rect 3316 -687 3332 -653
rect 3366 -687 3382 -653
rect 3565 -663 3639 -619
rect 3887 -635 3899 -568
rect 5122 -627 5254 -542
rect 7020 -627 7152 -542
rect 3747 -641 3899 -635
rect 3639 -673 3747 -663
rect 2397 -719 3027 -703
rect 2397 -723 2982 -719
rect 2397 -724 2498 -723
rect 2927 -772 3027 -761
rect 2891 -878 2901 -772
rect 3013 -783 3027 -772
rect 3316 -783 3382 -687
rect 5112 -735 5122 -627
rect 5254 -735 5264 -627
rect 7010 -735 7020 -627
rect 7152 -735 7162 -627
rect 7941 -655 8008 728
rect 3013 -831 3382 -783
rect 3013 -861 3027 -831
rect 3013 -878 3023 -861
rect 3315 -934 3381 -831
rect 5145 -870 5151 -735
rect 5218 -870 5224 -735
rect 5145 -882 5224 -870
rect 7941 -934 8007 -655
rect 3313 -1014 8007 -934
rect 5846 -1846 5925 -1834
rect 297 -1894 433 -1874
rect 297 -1956 333 -1894
rect 393 -1956 433 -1894
rect 297 -1984 433 -1956
rect 3366 -1901 3445 -1889
rect -7 -2014 970 -1984
rect 3366 -1998 3372 -1901
rect -7 -2120 25 -2014
rect 229 -2120 261 -2014
rect 465 -2120 497 -2014
rect 701 -2120 733 -2014
rect 936 -2120 970 -2014
rect 3298 -2018 3372 -1998
rect 3439 -1998 3445 -1901
rect 5846 -1964 5852 -1846
rect 5919 -1964 5925 -1846
rect 7002 -1849 7081 -1837
rect 7002 -1964 7008 -1849
rect 7075 -1964 7081 -1849
rect 3439 -2018 3518 -1998
rect -14 -2132 32 -2120
rect -14 -2308 -8 -2132
rect 26 -2308 32 -2132
rect -14 -2320 32 -2308
rect 104 -2132 150 -2120
rect 104 -2308 110 -2132
rect 144 -2308 150 -2132
rect 104 -2320 150 -2308
rect 222 -2132 268 -2120
rect 222 -2308 228 -2132
rect 262 -2308 268 -2132
rect 222 -2320 268 -2308
rect 340 -2132 386 -2120
rect 340 -2308 346 -2132
rect 380 -2308 386 -2132
rect 340 -2320 386 -2308
rect 458 -2132 504 -2120
rect 458 -2308 464 -2132
rect 498 -2308 504 -2132
rect 458 -2320 504 -2308
rect 576 -2132 622 -2120
rect 576 -2308 582 -2132
rect 616 -2308 622 -2132
rect 576 -2320 622 -2308
rect 694 -2132 740 -2120
rect 694 -2308 700 -2132
rect 734 -2308 740 -2132
rect 694 -2320 740 -2308
rect 812 -2132 858 -2120
rect 812 -2308 818 -2132
rect 852 -2308 858 -2132
rect 812 -2320 858 -2308
rect 930 -2132 976 -2120
rect 930 -2308 936 -2132
rect 970 -2308 976 -2132
rect 930 -2320 976 -2308
rect 1048 -2132 1094 -2120
rect 1048 -2308 1054 -2132
rect 1088 -2308 1094 -2132
rect 3298 -2126 3342 -2018
rect 3474 -2126 3518 -2018
rect 5095 -2060 5151 -2052
rect 3298 -2168 3518 -2126
rect 4169 -2068 5151 -2060
rect 4169 -2102 5111 -2068
rect 5145 -2102 5151 -2068
rect 5814 -2072 5824 -1964
rect 5956 -2027 5966 -1964
rect 5956 -2038 5968 -2027
rect 5956 -2072 5969 -2038
rect 6225 -2048 6281 -2046
rect 4169 -2118 5151 -2102
rect 5824 -2110 5969 -2072
rect 4169 -2119 5148 -2118
rect 2902 -2198 3879 -2168
rect 2902 -2304 2934 -2198
rect 3138 -2304 3170 -2198
rect 3374 -2304 3406 -2198
rect 3610 -2304 3642 -2198
rect 3845 -2304 3879 -2198
rect 1048 -2320 1094 -2308
rect 2895 -2316 2941 -2304
rect 109 -2414 145 -2320
rect 345 -2414 381 -2320
rect 581 -2413 617 -2320
rect 743 -2368 809 -2361
rect 743 -2402 759 -2368
rect 793 -2402 809 -2368
rect 743 -2413 809 -2402
rect 581 -2414 809 -2413
rect 109 -2443 809 -2414
rect 109 -2444 691 -2443
rect 229 -2557 263 -2444
rect 625 -2485 691 -2444
rect 625 -2519 641 -2485
rect 675 -2519 691 -2485
rect 625 -2526 691 -2519
rect 1053 -2553 1088 -2320
rect 2895 -2492 2901 -2316
rect 2935 -2492 2941 -2316
rect 2895 -2504 2941 -2492
rect 3013 -2316 3059 -2304
rect 3013 -2492 3019 -2316
rect 3053 -2492 3059 -2316
rect 3013 -2504 3059 -2492
rect 3131 -2316 3177 -2304
rect 3131 -2492 3137 -2316
rect 3171 -2492 3177 -2316
rect 3131 -2504 3177 -2492
rect 3249 -2316 3295 -2304
rect 3249 -2492 3255 -2316
rect 3289 -2492 3295 -2316
rect 3249 -2504 3295 -2492
rect 3367 -2316 3413 -2304
rect 3367 -2492 3373 -2316
rect 3407 -2492 3413 -2316
rect 3367 -2504 3413 -2492
rect 3485 -2316 3531 -2304
rect 3485 -2492 3491 -2316
rect 3525 -2492 3531 -2316
rect 3485 -2504 3531 -2492
rect 3603 -2316 3649 -2304
rect 3603 -2492 3609 -2316
rect 3643 -2492 3649 -2316
rect 3603 -2504 3649 -2492
rect 3721 -2316 3767 -2304
rect 3721 -2492 3727 -2316
rect 3761 -2492 3767 -2316
rect 3721 -2504 3767 -2492
rect 3839 -2316 3885 -2304
rect 3839 -2492 3845 -2316
rect 3879 -2492 3885 -2316
rect 3839 -2504 3885 -2492
rect 3957 -2316 4003 -2304
rect 3957 -2492 3963 -2316
rect 3997 -2492 4003 -2316
rect 3957 -2504 4003 -2492
rect 699 -2557 1088 -2553
rect 223 -2569 269 -2557
rect -189 -2797 183 -2697
rect 107 -2989 161 -2797
rect 223 -2945 229 -2569
rect 263 -2945 269 -2569
rect 223 -2957 269 -2945
rect 341 -2569 387 -2557
rect 341 -2945 347 -2569
rect 381 -2945 387 -2569
rect 341 -2957 387 -2945
rect 459 -2569 505 -2557
rect 459 -2945 465 -2569
rect 499 -2918 505 -2569
rect 576 -2569 622 -2557
rect 576 -2745 582 -2569
rect 616 -2745 622 -2569
rect 576 -2752 622 -2745
rect 694 -2569 1088 -2557
rect 694 -2745 700 -2569
rect 734 -2578 1088 -2569
rect 734 -2582 1090 -2578
rect 734 -2745 740 -2582
rect 576 -2757 625 -2752
rect 694 -2757 740 -2745
rect 582 -2918 625 -2757
rect 499 -2945 625 -2918
rect 459 -2957 625 -2945
rect 465 -2961 625 -2957
rect 107 -2995 338 -2989
rect 107 -3029 288 -2995
rect 322 -3029 338 -2995
rect 107 -3045 338 -3029
rect 390 -2995 456 -2989
rect 390 -3029 406 -2995
rect 440 -3029 456 -2995
rect -58 -3066 26 -3060
rect -58 -3119 -46 -3066
rect 14 -3074 26 -3066
rect 390 -3074 456 -3029
rect 14 -3082 456 -3074
rect 14 -3114 457 -3082
rect 549 -3098 625 -2961
rect 983 -3058 1090 -2582
rect 3018 -2598 3054 -2504
rect 3254 -2598 3290 -2504
rect 3490 -2597 3526 -2504
rect 3652 -2552 3718 -2545
rect 3652 -2586 3668 -2552
rect 3702 -2586 3718 -2552
rect 3652 -2597 3718 -2586
rect 3490 -2598 3718 -2597
rect 3018 -2627 3718 -2598
rect 3018 -2628 3600 -2627
rect 3138 -2741 3172 -2628
rect 3534 -2669 3600 -2628
rect 3534 -2703 3550 -2669
rect 3584 -2703 3600 -2669
rect 3534 -2710 3600 -2703
rect 3962 -2709 3997 -2504
rect 4169 -2709 4236 -2119
rect 5928 -2142 5969 -2110
rect 6215 -2114 6225 -2048
rect 6281 -2114 6291 -2048
rect 6961 -2072 6971 -1964
rect 7103 -2027 7113 -1964
rect 7103 -2038 7115 -2027
rect 7103 -2072 7116 -2038
rect 6971 -2110 7116 -2072
rect 7075 -2138 7116 -2110
rect 5344 -2170 5614 -2142
rect 5085 -2236 5095 -2170
rect 5161 -2236 5171 -2170
rect 5344 -2232 5378 -2170
rect 5580 -2232 5614 -2170
rect 5698 -2170 5969 -2142
rect 6486 -2166 6756 -2138
rect 5698 -2232 5732 -2170
rect 5934 -2232 5969 -2170
rect 6110 -2182 6281 -2166
rect 6110 -2216 6241 -2182
rect 6275 -2216 6281 -2182
rect 6110 -2232 6281 -2216
rect 6486 -2228 6520 -2166
rect 6722 -2228 6756 -2166
rect 6840 -2166 7116 -2138
rect 6840 -2228 6874 -2166
rect 7076 -2228 7116 -2166
rect 5220 -2244 5266 -2232
rect 5220 -2620 5226 -2244
rect 5260 -2620 5266 -2244
rect 5220 -2632 5266 -2620
rect 5338 -2244 5384 -2232
rect 5338 -2620 5344 -2244
rect 5378 -2620 5384 -2244
rect 5338 -2632 5384 -2620
rect 5456 -2244 5502 -2232
rect 5456 -2620 5462 -2244
rect 5496 -2620 5502 -2244
rect 5456 -2632 5502 -2620
rect 5574 -2244 5620 -2232
rect 5574 -2620 5580 -2244
rect 5614 -2620 5620 -2244
rect 5574 -2632 5620 -2620
rect 5692 -2244 5738 -2232
rect 5692 -2620 5698 -2244
rect 5732 -2620 5738 -2244
rect 5692 -2632 5738 -2620
rect 5810 -2244 5856 -2232
rect 5810 -2620 5816 -2244
rect 5850 -2620 5856 -2244
rect 5810 -2632 5856 -2620
rect 5928 -2244 5974 -2232
rect 5928 -2620 5934 -2244
rect 5968 -2620 5974 -2244
rect 5928 -2632 5974 -2620
rect 3962 -2737 4236 -2709
rect 3608 -2741 4236 -2737
rect 14 -3119 26 -3114
rect -58 -3125 26 -3119
rect 545 -3158 555 -3098
rect 617 -3158 627 -3098
rect 982 -3146 1090 -3058
rect 3132 -2753 3178 -2741
rect 3132 -3129 3138 -2753
rect 3172 -3129 3178 -2753
rect 3132 -3141 3178 -3129
rect 3250 -2753 3296 -2741
rect 3250 -3129 3256 -2753
rect 3290 -3129 3296 -2753
rect 3250 -3141 3296 -3129
rect 3368 -2753 3414 -2741
rect 3368 -3129 3374 -2753
rect 3408 -3105 3414 -2753
rect 3485 -2753 3531 -2741
rect 3485 -2929 3491 -2753
rect 3525 -2929 3531 -2753
rect 3485 -2941 3531 -2929
rect 3603 -2753 4236 -2741
rect 3603 -2929 3609 -2753
rect 3643 -2766 4236 -2753
rect 5226 -2674 5260 -2632
rect 5462 -2674 5496 -2632
rect 5226 -2702 5496 -2674
rect 5580 -2673 5614 -2632
rect 5816 -2673 5850 -2632
rect 5580 -2702 5850 -2673
rect 5226 -2750 5260 -2702
rect 3643 -2929 3649 -2766
rect 5226 -2780 5289 -2750
rect 3603 -2941 3649 -2929
rect 5254 -2872 5289 -2780
rect 5254 -2908 5481 -2872
rect 5751 -2883 5761 -2786
rect 5860 -2883 5870 -2786
rect 5934 -2815 5968 -2632
rect 5934 -2869 6043 -2815
rect 3491 -3057 3526 -2941
rect 5254 -3015 5289 -2908
rect 5415 -2942 5481 -2908
rect 5415 -2976 5431 -2942
rect 5465 -2976 5481 -2942
rect 5762 -2884 5859 -2883
rect 5762 -2951 5819 -2884
rect 5415 -2982 5481 -2976
rect 5656 -2987 5925 -2951
rect 5656 -3015 5689 -2987
rect 5892 -3015 5925 -2987
rect 6009 -3015 6043 -2869
rect 5130 -3027 5176 -3015
rect 3622 -3057 3730 -3047
rect 3491 -3105 3622 -3057
rect 3730 -3097 3876 -3091
rect 3408 -3129 3622 -3105
rect 3368 -3141 3622 -3129
rect 3374 -3145 3622 -3141
rect 982 -3173 3010 -3146
rect 982 -3179 3247 -3173
rect 982 -3213 3197 -3179
rect 3231 -3213 3247 -3179
rect 982 -3229 3247 -3213
rect 3299 -3179 3365 -3173
rect 3299 -3213 3315 -3179
rect 3349 -3213 3365 -3179
rect 3548 -3189 3622 -3145
rect 3864 -3164 3876 -3097
rect 3730 -3170 3876 -3164
rect 3622 -3199 3730 -3189
rect 982 -3245 3010 -3229
rect 982 -3246 2947 -3245
rect 982 -3247 2482 -3246
rect 1977 -3634 2266 -3633
rect 1481 -3635 2266 -3634
rect 1298 -3661 2266 -3635
rect 1298 -3767 2114 -3661
rect 2226 -3674 2266 -3661
rect 2226 -3767 2268 -3674
rect 1298 -3778 2268 -3767
rect 1298 -3779 2266 -3778
rect 313 -4654 449 -4634
rect 313 -4716 349 -4654
rect 409 -4716 449 -4654
rect 313 -4744 449 -4716
rect 9 -4774 986 -4744
rect 9 -4880 41 -4774
rect 245 -4880 277 -4774
rect 481 -4880 513 -4774
rect 717 -4880 749 -4774
rect 952 -4880 986 -4774
rect 2 -4892 48 -4880
rect 2 -5068 8 -4892
rect 42 -5068 48 -4892
rect 2 -5080 48 -5068
rect 120 -4892 166 -4880
rect 120 -5068 126 -4892
rect 160 -5068 166 -4892
rect 120 -5080 166 -5068
rect 238 -4892 284 -4880
rect 238 -5068 244 -4892
rect 278 -5068 284 -4892
rect 238 -5080 284 -5068
rect 356 -4892 402 -4880
rect 356 -5068 362 -4892
rect 396 -5068 402 -4892
rect 356 -5080 402 -5068
rect 474 -4892 520 -4880
rect 474 -5068 480 -4892
rect 514 -5068 520 -4892
rect 474 -5080 520 -5068
rect 592 -4892 638 -4880
rect 592 -5068 598 -4892
rect 632 -5068 638 -4892
rect 592 -5080 638 -5068
rect 710 -4892 756 -4880
rect 710 -5068 716 -4892
rect 750 -5068 756 -4892
rect 710 -5080 756 -5068
rect 828 -4892 874 -4880
rect 828 -5068 834 -4892
rect 868 -5068 874 -4892
rect 828 -5080 874 -5068
rect 946 -4892 992 -4880
rect 946 -5068 952 -4892
rect 986 -5068 992 -4892
rect 946 -5080 992 -5068
rect 1064 -4892 1110 -4880
rect 1064 -5068 1070 -4892
rect 1104 -5068 1110 -4892
rect 1064 -5080 1110 -5068
rect 125 -5174 161 -5080
rect 361 -5174 397 -5080
rect 597 -5173 633 -5080
rect 759 -5128 825 -5121
rect 759 -5162 775 -5128
rect 809 -5162 825 -5128
rect 759 -5173 825 -5162
rect 597 -5174 825 -5173
rect 125 -5203 825 -5174
rect 125 -5204 707 -5203
rect 245 -5317 279 -5204
rect 641 -5245 707 -5204
rect 641 -5279 657 -5245
rect 691 -5279 707 -5245
rect 641 -5286 707 -5279
rect 1069 -5313 1104 -5080
rect 1298 -5313 1421 -3779
rect 2389 -5144 2482 -3247
rect 2545 -3309 3011 -3287
rect 3299 -3309 3365 -3213
rect 5130 -3203 5136 -3027
rect 5170 -3203 5176 -3027
rect 5130 -3215 5176 -3203
rect 5248 -3027 5294 -3015
rect 5248 -3203 5254 -3027
rect 5288 -3203 5294 -3027
rect 5248 -3215 5294 -3203
rect 5366 -3027 5412 -3015
rect 5366 -3203 5372 -3027
rect 5406 -3203 5412 -3027
rect 5366 -3215 5412 -3203
rect 5484 -3027 5530 -3015
rect 5484 -3203 5490 -3027
rect 5524 -3082 5530 -3027
rect 5649 -3027 5695 -3015
rect 5649 -3082 5655 -3027
rect 5524 -3170 5655 -3082
rect 5524 -3203 5530 -3170
rect 5484 -3215 5530 -3203
rect 5649 -3203 5655 -3170
rect 5689 -3203 5695 -3027
rect 5649 -3215 5695 -3203
rect 5767 -3027 5813 -3015
rect 5767 -3203 5773 -3027
rect 5807 -3203 5813 -3027
rect 5767 -3215 5813 -3203
rect 5885 -3027 5931 -3015
rect 5885 -3203 5891 -3027
rect 5925 -3203 5931 -3027
rect 5885 -3215 5931 -3203
rect 6003 -3027 6049 -3015
rect 6003 -3203 6009 -3027
rect 6043 -3203 6049 -3027
rect 6003 -3215 6049 -3203
rect 5136 -3254 5170 -3215
rect 5372 -3254 5406 -3215
rect 5136 -3289 5406 -3254
rect 5773 -3253 5806 -3215
rect 6009 -3253 6042 -3215
rect 5773 -3289 6042 -3253
rect 2545 -3357 3365 -3309
rect 5170 -3290 5406 -3289
rect 2545 -3388 3011 -3357
rect 5170 -3364 5302 -3290
rect 2545 -3644 2650 -3388
rect 5160 -3472 5170 -3364
rect 5302 -3472 5312 -3364
rect 3387 -3554 3466 -3542
rect 2545 -3750 2608 -3644
rect 2720 -3750 2730 -3644
rect 3387 -3648 3393 -3554
rect 3312 -3668 3393 -3648
rect 3460 -3648 3466 -3554
rect 5186 -3607 5192 -3472
rect 5259 -3607 5265 -3472
rect 5186 -3619 5265 -3607
rect 3460 -3668 3532 -3648
rect 2545 -3761 2694 -3750
rect 2545 -4938 2650 -3761
rect 3312 -3776 3356 -3668
rect 3488 -3776 3532 -3668
rect 3312 -3818 3532 -3776
rect 6110 -3803 6172 -2232
rect 6362 -2240 6408 -2228
rect 6362 -2616 6368 -2240
rect 6402 -2616 6408 -2240
rect 6362 -2628 6408 -2616
rect 6480 -2240 6526 -2228
rect 6480 -2616 6486 -2240
rect 6520 -2616 6526 -2240
rect 6480 -2628 6526 -2616
rect 6598 -2240 6644 -2228
rect 6598 -2616 6604 -2240
rect 6638 -2616 6644 -2240
rect 6598 -2628 6644 -2616
rect 6716 -2240 6762 -2228
rect 6716 -2616 6722 -2240
rect 6756 -2616 6762 -2240
rect 6716 -2628 6762 -2616
rect 6834 -2240 6880 -2228
rect 6834 -2616 6840 -2240
rect 6874 -2616 6880 -2240
rect 6834 -2628 6880 -2616
rect 6952 -2240 6998 -2228
rect 6952 -2616 6958 -2240
rect 6992 -2616 6998 -2240
rect 6952 -2628 6998 -2616
rect 7070 -2240 7116 -2228
rect 7070 -2616 7076 -2240
rect 7110 -2616 7116 -2240
rect 7070 -2628 7116 -2616
rect 6368 -2670 6402 -2628
rect 6604 -2670 6638 -2628
rect 6368 -2698 6638 -2670
rect 6722 -2669 6756 -2628
rect 6958 -2669 6992 -2628
rect 6722 -2698 6992 -2669
rect 6368 -2746 6402 -2698
rect 6368 -2776 6431 -2746
rect 6396 -2868 6431 -2776
rect 6903 -2806 7003 -2785
rect 6903 -2860 6917 -2806
rect 6982 -2860 7003 -2806
rect 6903 -2865 7003 -2860
rect 7076 -2811 7110 -2628
rect 8310 -2796 8422 2089
rect 8946 724 9039 2618
rect 9102 2559 9568 2581
rect 9856 2559 9922 2655
rect 11687 2665 11693 2841
rect 11727 2665 11733 2841
rect 11687 2653 11733 2665
rect 11805 2841 11851 2853
rect 11805 2665 11811 2841
rect 11845 2665 11851 2841
rect 11805 2653 11851 2665
rect 11923 2841 11969 2853
rect 11923 2665 11929 2841
rect 11963 2665 11969 2841
rect 11923 2653 11969 2665
rect 12041 2841 12087 2853
rect 12041 2665 12047 2841
rect 12081 2786 12087 2841
rect 12206 2841 12252 2853
rect 12206 2786 12212 2841
rect 12081 2698 12212 2786
rect 12081 2665 12087 2698
rect 12041 2653 12087 2665
rect 12206 2665 12212 2698
rect 12246 2665 12252 2841
rect 12206 2653 12252 2665
rect 12324 2841 12370 2853
rect 12324 2665 12330 2841
rect 12364 2665 12370 2841
rect 12324 2653 12370 2665
rect 12442 2841 12488 2853
rect 12442 2665 12448 2841
rect 12482 2665 12488 2841
rect 12442 2653 12488 2665
rect 12560 2841 12606 2853
rect 12560 2665 12566 2841
rect 12600 2665 12606 2841
rect 12560 2653 12606 2665
rect 11693 2614 11727 2653
rect 11929 2614 11963 2653
rect 11693 2579 11963 2614
rect 12330 2615 12363 2653
rect 12566 2615 12599 2653
rect 12330 2579 12599 2615
rect 9102 2511 9922 2559
rect 11727 2578 11963 2579
rect 9102 2480 9568 2511
rect 11727 2504 11859 2578
rect 9102 2224 9207 2480
rect 11717 2396 11727 2504
rect 11859 2396 11869 2504
rect 9941 2315 10020 2327
rect 9102 2118 9165 2224
rect 9277 2118 9287 2224
rect 9941 2220 9947 2315
rect 9869 2200 9947 2220
rect 10014 2220 10020 2315
rect 11750 2266 11756 2396
rect 11823 2266 11829 2396
rect 11750 2254 11829 2266
rect 10014 2200 10089 2220
rect 9102 2107 9251 2118
rect 9102 930 9207 2107
rect 9869 2092 9913 2200
rect 10045 2092 10089 2200
rect 9869 2050 10089 2092
rect 12667 2065 12729 3636
rect 12919 3628 12965 3640
rect 12919 3252 12925 3628
rect 12959 3252 12965 3628
rect 12919 3240 12965 3252
rect 13037 3628 13083 3640
rect 13037 3252 13043 3628
rect 13077 3252 13083 3628
rect 13037 3240 13083 3252
rect 13155 3628 13201 3640
rect 13155 3252 13161 3628
rect 13195 3252 13201 3628
rect 13155 3240 13201 3252
rect 13273 3628 13319 3640
rect 13273 3252 13279 3628
rect 13313 3252 13319 3628
rect 13273 3240 13319 3252
rect 13391 3628 13437 3640
rect 13391 3252 13397 3628
rect 13431 3252 13437 3628
rect 13391 3240 13437 3252
rect 13509 3628 13555 3640
rect 13509 3252 13515 3628
rect 13549 3252 13555 3628
rect 13509 3240 13555 3252
rect 13627 3628 13673 3640
rect 13627 3252 13633 3628
rect 13667 3252 13673 3628
rect 13627 3240 13673 3252
rect 12925 3198 12959 3240
rect 13161 3198 13195 3240
rect 12925 3170 13195 3198
rect 13279 3199 13313 3240
rect 13515 3199 13549 3240
rect 13279 3170 13549 3199
rect 12925 3122 12959 3170
rect 12925 3092 12988 3122
rect 12953 3000 12988 3092
rect 13460 3062 13560 3083
rect 13460 3008 13474 3062
rect 13539 3008 13560 3062
rect 13460 3003 13560 3008
rect 13633 3057 13667 3240
rect 13633 3003 13742 3057
rect 12953 2964 13180 3000
rect 12953 2857 12988 2964
rect 13114 2930 13180 2964
rect 13114 2896 13130 2930
rect 13164 2896 13180 2930
rect 13461 2988 13558 3003
rect 13461 2921 13518 2988
rect 13114 2890 13180 2896
rect 13355 2885 13624 2921
rect 13355 2857 13388 2885
rect 13591 2857 13624 2885
rect 13708 2857 13742 3003
rect 14559 2996 14569 3071
rect 14637 2996 15031 3071
rect 14586 2995 15031 2996
rect 12829 2845 12875 2857
rect 12829 2669 12835 2845
rect 12869 2669 12875 2845
rect 12829 2657 12875 2669
rect 12947 2845 12993 2857
rect 12947 2669 12953 2845
rect 12987 2669 12993 2845
rect 12947 2657 12993 2669
rect 13065 2845 13111 2857
rect 13065 2669 13071 2845
rect 13105 2669 13111 2845
rect 13065 2657 13111 2669
rect 13183 2845 13229 2857
rect 13183 2669 13189 2845
rect 13223 2790 13229 2845
rect 13348 2845 13394 2857
rect 13348 2790 13354 2845
rect 13223 2702 13354 2790
rect 13223 2669 13229 2702
rect 13183 2657 13229 2669
rect 13348 2669 13354 2702
rect 13388 2669 13394 2845
rect 13348 2657 13394 2669
rect 13466 2845 13512 2857
rect 13466 2669 13472 2845
rect 13506 2669 13512 2845
rect 13466 2657 13512 2669
rect 13584 2845 13630 2857
rect 13584 2669 13590 2845
rect 13624 2669 13630 2845
rect 13584 2657 13630 2669
rect 13702 2845 13748 2857
rect 13702 2669 13708 2845
rect 13742 2669 13748 2845
rect 13702 2657 13748 2669
rect 12835 2618 12869 2657
rect 13071 2618 13105 2657
rect 12835 2582 13105 2618
rect 13472 2619 13505 2657
rect 13708 2619 13741 2657
rect 13472 2583 13741 2619
rect 12835 2581 13001 2582
rect 12869 2502 13001 2581
rect 12859 2394 12869 2502
rect 13001 2394 13011 2502
rect 12889 2258 12895 2394
rect 12962 2258 12968 2394
rect 12889 2246 12968 2258
rect 9473 2020 10450 2050
rect 12667 2048 12730 2065
rect 12592 2044 12730 2048
rect 9473 1914 9505 2020
rect 9709 1914 9741 2020
rect 9945 1914 9977 2020
rect 10181 1914 10213 2020
rect 10416 1914 10450 2020
rect 10760 2010 12730 2044
rect 10758 1981 12730 2010
rect 10758 1965 10804 1981
rect 12592 1979 12730 1981
rect 9466 1902 9512 1914
rect 9466 1726 9472 1902
rect 9506 1726 9512 1902
rect 9466 1714 9512 1726
rect 9584 1902 9630 1914
rect 9584 1726 9590 1902
rect 9624 1726 9630 1902
rect 9584 1714 9630 1726
rect 9702 1902 9748 1914
rect 9702 1726 9708 1902
rect 9742 1726 9748 1902
rect 9702 1714 9748 1726
rect 9820 1902 9866 1914
rect 9820 1726 9826 1902
rect 9860 1726 9866 1902
rect 9820 1714 9866 1726
rect 9938 1902 9984 1914
rect 9938 1726 9944 1902
rect 9978 1726 9984 1902
rect 9938 1714 9984 1726
rect 10056 1902 10102 1914
rect 10056 1726 10062 1902
rect 10096 1726 10102 1902
rect 10056 1714 10102 1726
rect 10174 1902 10220 1914
rect 10174 1726 10180 1902
rect 10214 1726 10220 1902
rect 10174 1714 10220 1726
rect 10292 1902 10338 1914
rect 10292 1726 10298 1902
rect 10332 1726 10338 1902
rect 10292 1714 10338 1726
rect 10410 1902 10456 1914
rect 10410 1726 10416 1902
rect 10450 1726 10456 1902
rect 10410 1714 10456 1726
rect 10528 1902 10574 1914
rect 10528 1726 10534 1902
rect 10568 1726 10574 1902
rect 10528 1714 10574 1726
rect 9589 1620 9625 1714
rect 9825 1620 9861 1714
rect 10061 1621 10097 1714
rect 10223 1666 10289 1673
rect 10223 1632 10239 1666
rect 10273 1632 10289 1666
rect 10223 1621 10289 1632
rect 10061 1620 10289 1621
rect 9589 1591 10289 1620
rect 9589 1590 10171 1591
rect 9709 1477 9743 1590
rect 10105 1549 10171 1590
rect 10105 1515 10121 1549
rect 10155 1515 10171 1549
rect 10105 1508 10171 1515
rect 10533 1496 10568 1714
rect 10757 1513 10804 1965
rect 13656 1973 13735 1985
rect 13656 1857 13662 1973
rect 13729 1857 13735 1973
rect 11716 1749 11726 1857
rect 11858 1749 11868 1857
rect 13614 1749 13624 1857
rect 13756 1749 13766 1857
rect 11726 1709 11858 1749
rect 13624 1709 13756 1749
rect 11725 1643 11858 1709
rect 13623 1643 13756 1709
rect 11054 1600 12527 1643
rect 10757 1497 10803 1513
rect 10722 1496 10803 1497
rect 10533 1481 10803 1496
rect 10179 1477 10803 1481
rect 9703 1465 9749 1477
rect 9438 987 9448 1105
rect 9566 1073 9576 1105
rect 9703 1089 9709 1465
rect 9743 1089 9749 1465
rect 9703 1077 9749 1089
rect 9821 1465 9867 1477
rect 9821 1089 9827 1465
rect 9861 1089 9867 1465
rect 9821 1077 9867 1089
rect 9939 1465 9985 1477
rect 9939 1089 9945 1465
rect 9979 1113 9985 1465
rect 10056 1465 10102 1477
rect 10056 1289 10062 1465
rect 10096 1289 10102 1465
rect 10056 1277 10102 1289
rect 10174 1465 10803 1477
rect 10174 1289 10180 1465
rect 10214 1453 10803 1465
rect 10214 1452 10456 1453
rect 10214 1289 10220 1452
rect 10722 1451 10803 1453
rect 11054 1297 11088 1600
rect 11420 1497 11454 1600
rect 11656 1497 11690 1600
rect 11892 1497 11926 1600
rect 12128 1497 12162 1600
rect 11414 1485 11460 1497
rect 10174 1277 10220 1289
rect 10930 1285 10976 1297
rect 10062 1161 10097 1277
rect 10193 1161 10301 1171
rect 10062 1113 10193 1161
rect 10301 1122 10450 1128
rect 9979 1089 10193 1113
rect 9939 1077 10193 1089
rect 9945 1073 10193 1077
rect 9566 1045 9581 1073
rect 9566 1039 9818 1045
rect 9566 1005 9768 1039
rect 9802 1005 9818 1039
rect 9566 989 9818 1005
rect 9870 1039 9936 1045
rect 9870 1005 9886 1039
rect 9920 1005 9936 1039
rect 10119 1029 10193 1073
rect 10438 1055 10450 1122
rect 10930 1109 10936 1285
rect 10970 1109 10976 1285
rect 10930 1097 10976 1109
rect 11048 1285 11094 1297
rect 11048 1109 11054 1285
rect 11088 1109 11094 1285
rect 11048 1097 11094 1109
rect 11166 1285 11212 1297
rect 11166 1109 11172 1285
rect 11206 1109 11212 1285
rect 11166 1097 11212 1109
rect 11284 1285 11330 1297
rect 11414 1285 11420 1485
rect 11284 1109 11290 1285
rect 11324 1109 11420 1285
rect 11454 1109 11460 1485
rect 11284 1097 11330 1109
rect 11414 1097 11460 1109
rect 11532 1485 11578 1497
rect 11532 1109 11538 1485
rect 11572 1109 11578 1485
rect 11532 1097 11578 1109
rect 11650 1485 11696 1497
rect 11650 1109 11656 1485
rect 11690 1109 11696 1485
rect 11650 1097 11696 1109
rect 11768 1485 11814 1497
rect 11768 1109 11774 1485
rect 11808 1109 11814 1485
rect 11768 1097 11814 1109
rect 11886 1485 11932 1497
rect 11886 1109 11892 1485
rect 11926 1109 11932 1485
rect 11886 1097 11932 1109
rect 12004 1485 12050 1497
rect 12004 1109 12010 1485
rect 12044 1109 12050 1485
rect 12004 1097 12050 1109
rect 12122 1485 12168 1497
rect 12122 1109 12128 1485
rect 12162 1285 12168 1485
rect 12493 1297 12527 1600
rect 12952 1600 14425 1643
rect 12952 1297 12986 1600
rect 13318 1497 13352 1600
rect 13554 1497 13588 1600
rect 13790 1497 13824 1600
rect 14026 1497 14060 1600
rect 13312 1485 13358 1497
rect 12251 1285 12297 1297
rect 12162 1109 12257 1285
rect 12291 1109 12297 1285
rect 12122 1097 12168 1109
rect 12251 1097 12297 1109
rect 12369 1285 12415 1297
rect 12369 1109 12375 1285
rect 12409 1109 12415 1285
rect 12369 1097 12415 1109
rect 12487 1285 12533 1297
rect 12487 1109 12493 1285
rect 12527 1109 12533 1285
rect 12487 1097 12533 1109
rect 12605 1285 12651 1297
rect 12605 1109 12611 1285
rect 12645 1109 12651 1285
rect 12605 1097 12651 1109
rect 12828 1285 12874 1297
rect 12828 1109 12834 1285
rect 12868 1109 12874 1285
rect 12828 1097 12874 1109
rect 12946 1285 12992 1297
rect 12946 1109 12952 1285
rect 12986 1109 12992 1285
rect 12946 1097 12992 1109
rect 13064 1285 13110 1297
rect 13064 1109 13070 1285
rect 13104 1109 13110 1285
rect 13064 1097 13110 1109
rect 13182 1285 13228 1297
rect 13312 1285 13318 1485
rect 13182 1109 13188 1285
rect 13222 1109 13318 1285
rect 13352 1109 13358 1485
rect 13182 1097 13228 1109
rect 13312 1097 13358 1109
rect 13430 1485 13476 1497
rect 13430 1109 13436 1485
rect 13470 1109 13476 1485
rect 13430 1097 13476 1109
rect 13548 1485 13594 1497
rect 13548 1109 13554 1485
rect 13588 1109 13594 1485
rect 13548 1097 13594 1109
rect 13666 1485 13712 1497
rect 13666 1109 13672 1485
rect 13706 1109 13712 1485
rect 13666 1097 13712 1109
rect 13784 1485 13830 1497
rect 13784 1109 13790 1485
rect 13824 1109 13830 1485
rect 13784 1097 13830 1109
rect 13902 1485 13948 1497
rect 13902 1109 13908 1485
rect 13942 1109 13948 1485
rect 13902 1097 13948 1109
rect 14020 1485 14066 1497
rect 14020 1109 14026 1485
rect 14060 1285 14066 1485
rect 14391 1297 14425 1600
rect 14149 1285 14195 1297
rect 14060 1109 14155 1285
rect 14189 1109 14195 1285
rect 14020 1097 14066 1109
rect 14149 1097 14195 1109
rect 14267 1285 14313 1297
rect 14267 1109 14273 1285
rect 14307 1109 14313 1285
rect 14267 1097 14313 1109
rect 14385 1285 14431 1297
rect 14385 1109 14391 1285
rect 14425 1109 14431 1285
rect 14385 1097 14431 1109
rect 14503 1285 14549 1297
rect 14503 1109 14509 1285
rect 14543 1109 14549 1285
rect 14503 1097 14549 1109
rect 10301 1049 10450 1055
rect 10936 1063 10970 1097
rect 11538 1063 11572 1097
rect 11774 1063 11808 1097
rect 10193 1019 10301 1029
rect 10936 1028 11095 1063
rect 11538 1028 11808 1063
rect 12375 1063 12409 1097
rect 12611 1063 12645 1097
rect 12375 1028 12645 1063
rect 12834 1063 12868 1097
rect 13436 1063 13470 1097
rect 13672 1063 13706 1097
rect 12834 1028 12993 1063
rect 13436 1028 13706 1063
rect 14273 1063 14307 1097
rect 14509 1063 14543 1097
rect 14273 1028 14543 1063
rect 9566 987 9581 989
rect 9481 973 9581 987
rect 9481 930 9581 931
rect 9102 909 9581 930
rect 9870 909 9936 1005
rect 9102 861 9936 909
rect 9102 832 9581 861
rect 9102 830 9207 832
rect 9481 831 9581 832
rect 8935 645 8945 724
rect 9038 645 9048 724
rect 9933 715 10012 727
rect 8946 -529 9039 645
rect 9933 616 9939 715
rect 9864 596 9939 616
rect 10006 616 10012 715
rect 10006 596 10084 616
rect 9864 488 9908 596
rect 10040 488 10084 596
rect 9864 446 10084 488
rect 9468 416 10445 446
rect 9468 310 9500 416
rect 9704 310 9736 416
rect 9940 310 9972 416
rect 10176 310 10208 416
rect 10411 310 10445 416
rect 9461 298 9507 310
rect 9461 122 9467 298
rect 9501 122 9507 298
rect 9461 110 9507 122
rect 9579 298 9625 310
rect 9579 122 9585 298
rect 9619 122 9625 298
rect 9579 110 9625 122
rect 9697 298 9743 310
rect 9697 122 9703 298
rect 9737 122 9743 298
rect 9697 110 9743 122
rect 9815 298 9861 310
rect 9815 122 9821 298
rect 9855 122 9861 298
rect 9815 110 9861 122
rect 9933 298 9979 310
rect 9933 122 9939 298
rect 9973 122 9979 298
rect 9933 110 9979 122
rect 10051 298 10097 310
rect 10051 122 10057 298
rect 10091 122 10097 298
rect 10051 110 10097 122
rect 10169 298 10215 310
rect 10169 122 10175 298
rect 10209 122 10215 298
rect 10169 110 10215 122
rect 10287 298 10333 310
rect 10287 122 10293 298
rect 10327 122 10333 298
rect 10287 110 10333 122
rect 10405 298 10451 310
rect 10405 122 10411 298
rect 10445 122 10451 298
rect 10405 110 10451 122
rect 10523 298 10569 310
rect 10523 122 10529 298
rect 10563 122 10569 298
rect 10523 110 10569 122
rect 11061 244 11095 1028
rect 11774 966 11808 1028
rect 11363 928 12105 966
rect 11363 804 11397 928
rect 11599 804 11633 928
rect 11835 804 11869 928
rect 12071 804 12105 928
rect 12361 821 12371 887
rect 12434 821 12444 887
rect 11357 792 11403 804
rect 11357 416 11363 792
rect 11397 416 11403 792
rect 11357 404 11403 416
rect 11475 792 11521 804
rect 11475 416 11481 792
rect 11515 416 11521 792
rect 11475 404 11521 416
rect 11593 792 11639 804
rect 11593 416 11599 792
rect 11633 416 11639 792
rect 11593 404 11639 416
rect 11711 792 11757 804
rect 11711 416 11717 792
rect 11751 416 11757 792
rect 11711 404 11757 416
rect 11829 792 11875 804
rect 11829 416 11835 792
rect 11869 416 11875 792
rect 11829 404 11875 416
rect 11947 792 11993 804
rect 11947 416 11953 792
rect 11987 416 11993 792
rect 11947 404 11993 416
rect 12065 792 12111 804
rect 12065 416 12071 792
rect 12105 416 12111 792
rect 12065 404 12111 416
rect 12477 245 12511 1028
rect 12204 244 12511 245
rect 11061 239 11377 244
rect 12091 239 12511 244
rect 11061 228 11444 239
rect 11061 201 11393 228
rect 9584 16 9620 110
rect 9820 16 9856 110
rect 10056 17 10092 110
rect 10218 62 10284 69
rect 10218 28 10234 62
rect 10268 28 10284 62
rect 10218 17 10284 28
rect 10056 16 10284 17
rect 9584 -13 10284 16
rect 9584 -14 10166 -13
rect 9704 -127 9738 -14
rect 10100 -55 10166 -14
rect 10100 -89 10116 -55
rect 10150 -89 10166 -55
rect 10100 -96 10166 -89
rect 10528 -123 10563 110
rect 11061 72 11095 201
rect 11377 194 11393 201
rect 11427 194 11444 228
rect 11377 188 11444 194
rect 12024 228 12511 239
rect 12024 194 12041 228
rect 12075 201 12511 228
rect 12075 194 12091 201
rect 12204 200 12511 201
rect 12024 188 12091 194
rect 11202 161 11258 173
rect 11202 127 11208 161
rect 11242 160 11258 161
rect 12315 160 12371 172
rect 11242 144 11709 160
rect 11242 127 11659 144
rect 11202 111 11659 127
rect 11643 110 11659 111
rect 11693 110 11709 144
rect 11643 103 11709 110
rect 11761 145 12331 160
rect 11761 111 11777 145
rect 11811 126 12331 145
rect 12365 126 12371 160
rect 11811 111 12371 126
rect 11761 101 11828 111
rect 12315 110 12371 111
rect 12477 72 12511 200
rect 12959 244 12993 1028
rect 13672 966 13706 1028
rect 13261 928 14003 966
rect 13261 804 13295 928
rect 13497 804 13531 928
rect 13733 804 13767 928
rect 13969 804 14003 928
rect 13255 792 13301 804
rect 13255 416 13261 792
rect 13295 416 13301 792
rect 13255 404 13301 416
rect 13373 792 13419 804
rect 13373 416 13379 792
rect 13413 416 13419 792
rect 13373 404 13419 416
rect 13491 792 13537 804
rect 13491 416 13497 792
rect 13531 416 13537 792
rect 13491 404 13537 416
rect 13609 792 13655 804
rect 13609 416 13615 792
rect 13649 416 13655 792
rect 13609 404 13655 416
rect 13727 792 13773 804
rect 13727 416 13733 792
rect 13767 416 13773 792
rect 13727 404 13773 416
rect 13845 792 13891 804
rect 13845 416 13851 792
rect 13885 416 13891 792
rect 13845 404 13891 416
rect 13963 792 14009 804
rect 13963 416 13969 792
rect 14003 416 14009 792
rect 13963 404 14009 416
rect 14375 245 14409 1028
rect 13987 244 14056 245
rect 14102 244 14409 245
rect 12959 239 13275 244
rect 13987 240 14409 244
rect 12959 228 13342 239
rect 12959 201 13291 228
rect 12959 72 12993 201
rect 13275 194 13291 201
rect 13325 194 13342 228
rect 13275 188 13342 194
rect 13920 229 14409 240
rect 13920 195 13937 229
rect 13971 201 14409 229
rect 13971 195 13987 201
rect 14102 200 14409 201
rect 13920 189 13987 195
rect 13100 161 13156 173
rect 13100 127 13106 161
rect 13140 160 13156 161
rect 14213 160 14269 172
rect 13140 144 13607 160
rect 13140 127 13557 144
rect 13100 111 13557 127
rect 13541 110 13557 111
rect 13591 110 13607 144
rect 13541 103 13607 110
rect 13659 145 14229 160
rect 13659 111 13675 145
rect 13709 126 14229 145
rect 14263 126 14269 160
rect 13709 111 14269 126
rect 13659 101 13726 111
rect 14213 110 14269 111
rect 14375 72 14409 200
rect 14490 850 14557 874
rect 14490 816 14507 850
rect 14541 816 14557 850
rect 10174 -127 10563 -123
rect 9698 -139 9744 -127
rect 9698 -515 9704 -139
rect 9738 -515 9744 -139
rect 9698 -527 9744 -515
rect 9816 -139 9862 -127
rect 9816 -515 9822 -139
rect 9856 -515 9862 -139
rect 9816 -527 9862 -515
rect 9934 -139 9980 -127
rect 9934 -515 9940 -139
rect 9974 -491 9980 -139
rect 10051 -139 10097 -127
rect 10051 -315 10057 -139
rect 10091 -315 10097 -139
rect 10051 -327 10097 -315
rect 10169 -139 10563 -127
rect 11055 60 11101 72
rect 11055 -116 11061 60
rect 11095 -116 11101 60
rect 11055 -128 11101 -116
rect 11173 60 11219 72
rect 11173 -116 11179 60
rect 11213 -116 11219 60
rect 11173 -128 11219 -116
rect 11475 60 11521 72
rect 10169 -315 10175 -139
rect 10209 -152 10563 -139
rect 10209 -315 10215 -152
rect 10485 -155 10563 -152
rect 10485 -207 10495 -155
rect 10558 -207 10568 -155
rect 10490 -213 10563 -207
rect 10169 -327 10215 -315
rect 10057 -443 10092 -327
rect 11178 -422 11212 -128
rect 11475 -316 11481 60
rect 11515 -316 11521 60
rect 11475 -328 11521 -316
rect 11593 60 11639 72
rect 11593 -316 11599 60
rect 11633 -316 11639 60
rect 11593 -328 11639 -316
rect 11711 60 11757 72
rect 11711 -316 11717 60
rect 11751 -316 11757 60
rect 11711 -328 11757 -316
rect 11829 60 11875 72
rect 11829 -316 11835 60
rect 11869 -316 11875 60
rect 11829 -328 11875 -316
rect 11947 60 11993 72
rect 11947 -316 11953 60
rect 11987 -316 11993 60
rect 12353 60 12399 72
rect 12353 -116 12359 60
rect 12393 -116 12399 60
rect 12353 -128 12399 -116
rect 12471 60 12517 72
rect 12471 -116 12477 60
rect 12511 -116 12517 60
rect 12471 -128 12517 -116
rect 12953 60 12999 72
rect 12953 -116 12959 60
rect 12993 -116 12999 60
rect 12953 -128 12999 -116
rect 13071 60 13117 72
rect 13071 -116 13077 60
rect 13111 -116 13117 60
rect 13071 -128 13117 -116
rect 13373 60 13419 72
rect 11947 -328 11993 -316
rect 11835 -422 11869 -328
rect 12359 -422 12392 -128
rect 10188 -443 10296 -433
rect 10057 -491 10188 -443
rect 11178 -454 12392 -422
rect 13076 -422 13110 -128
rect 13373 -316 13379 60
rect 13413 -316 13419 60
rect 13373 -328 13419 -316
rect 13491 60 13537 72
rect 13491 -316 13497 60
rect 13531 -316 13537 60
rect 13491 -328 13537 -316
rect 13609 60 13655 72
rect 13609 -316 13615 60
rect 13649 -316 13655 60
rect 13609 -328 13655 -316
rect 13727 60 13773 72
rect 13727 -316 13733 60
rect 13767 -316 13773 60
rect 13727 -328 13773 -316
rect 13845 60 13891 72
rect 13845 -316 13851 60
rect 13885 -316 13891 60
rect 14251 60 14297 72
rect 14251 -116 14257 60
rect 14291 -116 14297 60
rect 14251 -128 14297 -116
rect 14369 60 14415 72
rect 14369 -116 14375 60
rect 14409 -116 14415 60
rect 14369 -128 14415 -116
rect 13845 -328 13891 -316
rect 13733 -422 13767 -328
rect 14257 -422 14290 -128
rect 13076 -454 14290 -422
rect 10296 -479 10447 -473
rect 9974 -515 10188 -491
rect 9934 -527 10188 -515
rect 8946 -531 9531 -529
rect 9940 -531 10188 -527
rect 8946 -559 9576 -531
rect 8946 -565 9813 -559
rect 8946 -599 9763 -565
rect 9797 -599 9813 -565
rect 8946 -615 9813 -599
rect 9865 -565 9931 -559
rect 9865 -599 9881 -565
rect 9915 -599 9931 -565
rect 10114 -575 10188 -531
rect 10435 -546 10447 -479
rect 11671 -539 11803 -454
rect 13569 -539 13701 -454
rect 10296 -552 10447 -546
rect 10188 -585 10296 -575
rect 8946 -631 9576 -615
rect 8946 -635 9531 -631
rect 8946 -636 9047 -635
rect 9476 -684 9576 -673
rect 9440 -790 9450 -684
rect 9562 -695 9576 -684
rect 9865 -695 9931 -599
rect 11661 -647 11671 -539
rect 11803 -647 11813 -539
rect 13559 -647 13569 -539
rect 13701 -647 13711 -539
rect 14490 -567 14557 816
rect 14618 387 14774 393
rect 14618 289 14630 387
rect 14762 289 14774 387
rect 14618 283 14774 289
rect 9562 -743 9931 -695
rect 9562 -773 9576 -743
rect 9562 -790 9572 -773
rect 9864 -846 9930 -743
rect 11694 -785 11700 -647
rect 11767 -785 11773 -647
rect 11694 -797 11773 -785
rect 14490 -846 14556 -567
rect 9862 -926 14556 -846
rect 12402 -1850 12481 -1838
rect 9921 -1903 10000 -1891
rect 9921 -2000 9927 -1903
rect 9849 -2020 9927 -2000
rect 9994 -2000 10000 -1903
rect 12402 -1966 12408 -1850
rect 12475 -1966 12481 -1850
rect 13550 -1850 13629 -1838
rect 13550 -1966 13556 -1850
rect 13623 -1966 13629 -1850
rect 9994 -2020 10069 -2000
rect 9849 -2128 9893 -2020
rect 10025 -2128 10069 -2020
rect 11646 -2062 11702 -2054
rect 9849 -2170 10069 -2128
rect 10720 -2070 11702 -2062
rect 10720 -2104 11662 -2070
rect 11696 -2104 11702 -2070
rect 12365 -2074 12375 -1966
rect 12507 -2029 12517 -1966
rect 12507 -2040 12519 -2029
rect 12507 -2074 12520 -2040
rect 12776 -2050 12832 -2048
rect 10720 -2120 11702 -2104
rect 12375 -2112 12520 -2074
rect 10720 -2121 11699 -2120
rect 9453 -2200 10430 -2170
rect 9453 -2306 9485 -2200
rect 9689 -2306 9721 -2200
rect 9925 -2306 9957 -2200
rect 10161 -2306 10193 -2200
rect 10396 -2306 10430 -2200
rect 9446 -2318 9492 -2306
rect 9446 -2494 9452 -2318
rect 9486 -2494 9492 -2318
rect 9446 -2506 9492 -2494
rect 9564 -2318 9610 -2306
rect 9564 -2494 9570 -2318
rect 9604 -2494 9610 -2318
rect 9564 -2506 9610 -2494
rect 9682 -2318 9728 -2306
rect 9682 -2494 9688 -2318
rect 9722 -2494 9728 -2318
rect 9682 -2506 9728 -2494
rect 9800 -2318 9846 -2306
rect 9800 -2494 9806 -2318
rect 9840 -2494 9846 -2318
rect 9800 -2506 9846 -2494
rect 9918 -2318 9964 -2306
rect 9918 -2494 9924 -2318
rect 9958 -2494 9964 -2318
rect 9918 -2506 9964 -2494
rect 10036 -2318 10082 -2306
rect 10036 -2494 10042 -2318
rect 10076 -2494 10082 -2318
rect 10036 -2506 10082 -2494
rect 10154 -2318 10200 -2306
rect 10154 -2494 10160 -2318
rect 10194 -2494 10200 -2318
rect 10154 -2506 10200 -2494
rect 10272 -2318 10318 -2306
rect 10272 -2494 10278 -2318
rect 10312 -2494 10318 -2318
rect 10272 -2506 10318 -2494
rect 10390 -2318 10436 -2306
rect 10390 -2494 10396 -2318
rect 10430 -2494 10436 -2318
rect 10390 -2506 10436 -2494
rect 10508 -2318 10554 -2306
rect 10508 -2494 10514 -2318
rect 10548 -2494 10554 -2318
rect 10508 -2506 10554 -2494
rect 9569 -2600 9605 -2506
rect 9805 -2600 9841 -2506
rect 10041 -2599 10077 -2506
rect 10203 -2554 10269 -2547
rect 10203 -2588 10219 -2554
rect 10253 -2588 10269 -2554
rect 10203 -2599 10269 -2588
rect 10041 -2600 10269 -2599
rect 9569 -2629 10269 -2600
rect 9569 -2630 10151 -2629
rect 9689 -2743 9723 -2630
rect 10085 -2671 10151 -2630
rect 10085 -2705 10101 -2671
rect 10135 -2705 10151 -2671
rect 10085 -2712 10151 -2705
rect 10513 -2711 10548 -2506
rect 10720 -2711 10787 -2121
rect 12479 -2144 12520 -2112
rect 12766 -2116 12776 -2050
rect 12832 -2116 12842 -2050
rect 13512 -2074 13522 -1966
rect 13654 -2029 13664 -1966
rect 13654 -2040 13666 -2029
rect 13654 -2074 13667 -2040
rect 13522 -2112 13667 -2074
rect 13626 -2140 13667 -2112
rect 11895 -2172 12165 -2144
rect 11636 -2238 11646 -2172
rect 11712 -2238 11722 -2172
rect 11895 -2234 11929 -2172
rect 12131 -2234 12165 -2172
rect 12249 -2172 12520 -2144
rect 13037 -2168 13307 -2140
rect 12249 -2234 12283 -2172
rect 12485 -2234 12520 -2172
rect 12661 -2184 12832 -2168
rect 12661 -2218 12792 -2184
rect 12826 -2218 12832 -2184
rect 12661 -2234 12832 -2218
rect 13037 -2230 13071 -2168
rect 13273 -2230 13307 -2168
rect 13391 -2168 13667 -2140
rect 13391 -2230 13425 -2168
rect 13627 -2230 13667 -2168
rect 11771 -2246 11817 -2234
rect 11771 -2622 11777 -2246
rect 11811 -2622 11817 -2246
rect 11771 -2634 11817 -2622
rect 11889 -2246 11935 -2234
rect 11889 -2622 11895 -2246
rect 11929 -2622 11935 -2246
rect 11889 -2634 11935 -2622
rect 12007 -2246 12053 -2234
rect 12007 -2622 12013 -2246
rect 12047 -2622 12053 -2246
rect 12007 -2634 12053 -2622
rect 12125 -2246 12171 -2234
rect 12125 -2622 12131 -2246
rect 12165 -2622 12171 -2246
rect 12125 -2634 12171 -2622
rect 12243 -2246 12289 -2234
rect 12243 -2622 12249 -2246
rect 12283 -2622 12289 -2246
rect 12243 -2634 12289 -2622
rect 12361 -2246 12407 -2234
rect 12361 -2622 12367 -2246
rect 12401 -2622 12407 -2246
rect 12361 -2634 12407 -2622
rect 12479 -2246 12525 -2234
rect 12479 -2622 12485 -2246
rect 12519 -2622 12525 -2246
rect 12479 -2634 12525 -2622
rect 10513 -2739 10787 -2711
rect 10159 -2743 10787 -2739
rect 8067 -2797 8422 -2796
rect 7076 -2865 7185 -2811
rect 6396 -2904 6623 -2868
rect 6396 -3011 6431 -2904
rect 6557 -2938 6623 -2904
rect 6557 -2972 6573 -2938
rect 6607 -2972 6623 -2938
rect 6904 -2880 7001 -2865
rect 6904 -2947 6961 -2880
rect 6557 -2978 6623 -2972
rect 6798 -2983 7067 -2947
rect 6798 -3011 6831 -2983
rect 7034 -3011 7067 -2983
rect 7151 -3011 7185 -2865
rect 8002 -2872 8012 -2797
rect 8080 -2872 8422 -2797
rect 8029 -2873 8422 -2872
rect 8067 -2874 8422 -2873
rect 9683 -2755 9729 -2743
rect 6272 -3023 6318 -3011
rect 6272 -3199 6278 -3023
rect 6312 -3199 6318 -3023
rect 6272 -3211 6318 -3199
rect 6390 -3023 6436 -3011
rect 6390 -3199 6396 -3023
rect 6430 -3199 6436 -3023
rect 6390 -3211 6436 -3199
rect 6508 -3023 6554 -3011
rect 6508 -3199 6514 -3023
rect 6548 -3199 6554 -3023
rect 6508 -3211 6554 -3199
rect 6626 -3023 6672 -3011
rect 6626 -3199 6632 -3023
rect 6666 -3078 6672 -3023
rect 6791 -3023 6837 -3011
rect 6791 -3078 6797 -3023
rect 6666 -3166 6797 -3078
rect 6666 -3199 6672 -3166
rect 6626 -3211 6672 -3199
rect 6791 -3199 6797 -3166
rect 6831 -3199 6837 -3023
rect 6791 -3211 6837 -3199
rect 6909 -3023 6955 -3011
rect 6909 -3199 6915 -3023
rect 6949 -3199 6955 -3023
rect 6909 -3211 6955 -3199
rect 7027 -3023 7073 -3011
rect 7027 -3199 7033 -3023
rect 7067 -3199 7073 -3023
rect 7027 -3211 7073 -3199
rect 7145 -3023 7191 -3011
rect 7145 -3199 7151 -3023
rect 7185 -3199 7191 -3023
rect 9683 -3131 9689 -2755
rect 9723 -3131 9729 -2755
rect 9683 -3143 9729 -3131
rect 9801 -2755 9847 -2743
rect 9801 -3131 9807 -2755
rect 9841 -3131 9847 -2755
rect 9801 -3143 9847 -3131
rect 9919 -2755 9965 -2743
rect 9919 -3131 9925 -2755
rect 9959 -3107 9965 -2755
rect 10036 -2755 10082 -2743
rect 10036 -2931 10042 -2755
rect 10076 -2931 10082 -2755
rect 10036 -2943 10082 -2931
rect 10154 -2755 10787 -2743
rect 10154 -2931 10160 -2755
rect 10194 -2768 10787 -2755
rect 11777 -2676 11811 -2634
rect 12013 -2676 12047 -2634
rect 11777 -2704 12047 -2676
rect 12131 -2675 12165 -2634
rect 12367 -2675 12401 -2634
rect 12131 -2704 12401 -2675
rect 11777 -2752 11811 -2704
rect 10194 -2931 10200 -2768
rect 11777 -2782 11840 -2752
rect 10154 -2943 10200 -2931
rect 11805 -2874 11840 -2782
rect 11805 -2910 12032 -2874
rect 12302 -2885 12312 -2788
rect 12411 -2885 12421 -2788
rect 12485 -2817 12519 -2634
rect 12485 -2871 12594 -2817
rect 10042 -3059 10077 -2943
rect 11805 -3017 11840 -2910
rect 11966 -2944 12032 -2910
rect 11966 -2978 11982 -2944
rect 12016 -2978 12032 -2944
rect 12313 -2886 12410 -2885
rect 12313 -2953 12370 -2886
rect 11966 -2984 12032 -2978
rect 12207 -2989 12476 -2953
rect 12207 -3017 12240 -2989
rect 12443 -3017 12476 -2989
rect 12560 -3017 12594 -2871
rect 11681 -3029 11727 -3017
rect 10173 -3059 10281 -3049
rect 10042 -3107 10173 -3059
rect 10281 -3103 10426 -3097
rect 9959 -3131 10173 -3107
rect 9919 -3143 10173 -3131
rect 9925 -3147 10173 -3143
rect 7145 -3211 7191 -3199
rect 8061 -3175 9561 -3148
rect 8061 -3181 9798 -3175
rect 6278 -3250 6312 -3211
rect 6514 -3250 6548 -3211
rect 6278 -3286 6548 -3250
rect 6915 -3249 6948 -3211
rect 7151 -3249 7184 -3211
rect 6915 -3285 7184 -3249
rect 8061 -3215 9748 -3181
rect 9782 -3215 9798 -3181
rect 8061 -3231 9798 -3215
rect 9850 -3181 9916 -3175
rect 9850 -3215 9866 -3181
rect 9900 -3215 9916 -3181
rect 10099 -3191 10173 -3147
rect 10414 -3170 10426 -3103
rect 10281 -3176 10426 -3170
rect 10173 -3201 10281 -3191
rect 8061 -3247 9561 -3231
rect 8061 -3248 9498 -3247
rect 8061 -3254 9033 -3248
rect 6278 -3287 6444 -3286
rect 6312 -3366 6444 -3287
rect 6302 -3474 6312 -3366
rect 6444 -3474 6454 -3366
rect 6339 -3612 6345 -3474
rect 6412 -3612 6418 -3474
rect 6339 -3624 6418 -3612
rect 2916 -3848 3893 -3818
rect 6110 -3820 6173 -3803
rect 6035 -3824 6173 -3820
rect 2916 -3954 2948 -3848
rect 3152 -3954 3184 -3848
rect 3388 -3954 3420 -3848
rect 3624 -3954 3656 -3848
rect 3859 -3954 3893 -3848
rect 4203 -3858 6173 -3824
rect 4201 -3887 6173 -3858
rect 4201 -3903 4247 -3887
rect 6035 -3889 6173 -3887
rect 2909 -3966 2955 -3954
rect 2909 -4142 2915 -3966
rect 2949 -4142 2955 -3966
rect 2909 -4154 2955 -4142
rect 3027 -3966 3073 -3954
rect 3027 -4142 3033 -3966
rect 3067 -4142 3073 -3966
rect 3027 -4154 3073 -4142
rect 3145 -3966 3191 -3954
rect 3145 -4142 3151 -3966
rect 3185 -4142 3191 -3966
rect 3145 -4154 3191 -4142
rect 3263 -3966 3309 -3954
rect 3263 -4142 3269 -3966
rect 3303 -4142 3309 -3966
rect 3263 -4154 3309 -4142
rect 3381 -3966 3427 -3954
rect 3381 -4142 3387 -3966
rect 3421 -4142 3427 -3966
rect 3381 -4154 3427 -4142
rect 3499 -3966 3545 -3954
rect 3499 -4142 3505 -3966
rect 3539 -4142 3545 -3966
rect 3499 -4154 3545 -4142
rect 3617 -3966 3663 -3954
rect 3617 -4142 3623 -3966
rect 3657 -4142 3663 -3966
rect 3617 -4154 3663 -4142
rect 3735 -3966 3781 -3954
rect 3735 -4142 3741 -3966
rect 3775 -4142 3781 -3966
rect 3735 -4154 3781 -4142
rect 3853 -3966 3899 -3954
rect 3853 -4142 3859 -3966
rect 3893 -4142 3899 -3966
rect 3853 -4154 3899 -4142
rect 3971 -3966 4017 -3954
rect 3971 -4142 3977 -3966
rect 4011 -4142 4017 -3966
rect 3971 -4154 4017 -4142
rect 3032 -4248 3068 -4154
rect 3268 -4248 3304 -4154
rect 3504 -4247 3540 -4154
rect 3666 -4202 3732 -4195
rect 3666 -4236 3682 -4202
rect 3716 -4236 3732 -4202
rect 3666 -4247 3732 -4236
rect 3504 -4248 3732 -4247
rect 3032 -4277 3732 -4248
rect 3032 -4278 3614 -4277
rect 3152 -4391 3186 -4278
rect 3548 -4319 3614 -4278
rect 3548 -4353 3564 -4319
rect 3598 -4353 3614 -4319
rect 3548 -4360 3614 -4353
rect 3976 -4372 4011 -4154
rect 4200 -4355 4247 -3903
rect 7093 -3895 7172 -3883
rect 7093 -4011 7099 -3895
rect 7166 -4011 7172 -3895
rect 5159 -4119 5169 -4011
rect 5301 -4119 5311 -4011
rect 7057 -4119 7067 -4011
rect 7199 -4119 7209 -4011
rect 5169 -4159 5301 -4119
rect 7067 -4159 7199 -4119
rect 5168 -4225 5301 -4159
rect 7066 -4225 7199 -4159
rect 4497 -4268 5970 -4225
rect 4200 -4371 4246 -4355
rect 4165 -4372 4246 -4371
rect 3976 -4387 4246 -4372
rect 3622 -4391 4246 -4387
rect 3146 -4403 3192 -4391
rect 2881 -4881 2891 -4763
rect 3009 -4795 3019 -4763
rect 3146 -4779 3152 -4403
rect 3186 -4779 3192 -4403
rect 3146 -4791 3192 -4779
rect 3264 -4403 3310 -4391
rect 3264 -4779 3270 -4403
rect 3304 -4779 3310 -4403
rect 3264 -4791 3310 -4779
rect 3382 -4403 3428 -4391
rect 3382 -4779 3388 -4403
rect 3422 -4755 3428 -4403
rect 3499 -4403 3545 -4391
rect 3499 -4579 3505 -4403
rect 3539 -4579 3545 -4403
rect 3499 -4591 3545 -4579
rect 3617 -4403 4246 -4391
rect 3617 -4579 3623 -4403
rect 3657 -4415 4246 -4403
rect 3657 -4416 3899 -4415
rect 3657 -4579 3663 -4416
rect 4165 -4417 4246 -4415
rect 4497 -4571 4531 -4268
rect 4863 -4371 4897 -4268
rect 5099 -4371 5133 -4268
rect 5335 -4371 5369 -4268
rect 5571 -4371 5605 -4268
rect 4857 -4383 4903 -4371
rect 3617 -4591 3663 -4579
rect 4373 -4583 4419 -4571
rect 3505 -4707 3540 -4591
rect 3636 -4707 3744 -4697
rect 3505 -4755 3636 -4707
rect 3744 -4747 3884 -4741
rect 3422 -4779 3636 -4755
rect 3382 -4791 3636 -4779
rect 3388 -4795 3636 -4791
rect 3009 -4823 3024 -4795
rect 3009 -4829 3261 -4823
rect 3009 -4863 3211 -4829
rect 3245 -4863 3261 -4829
rect 3009 -4879 3261 -4863
rect 3313 -4829 3379 -4823
rect 3313 -4863 3329 -4829
rect 3363 -4863 3379 -4829
rect 3562 -4839 3636 -4795
rect 3872 -4814 3884 -4747
rect 4373 -4759 4379 -4583
rect 4413 -4759 4419 -4583
rect 4373 -4771 4419 -4759
rect 4491 -4583 4537 -4571
rect 4491 -4759 4497 -4583
rect 4531 -4759 4537 -4583
rect 4491 -4771 4537 -4759
rect 4609 -4583 4655 -4571
rect 4609 -4759 4615 -4583
rect 4649 -4759 4655 -4583
rect 4609 -4771 4655 -4759
rect 4727 -4583 4773 -4571
rect 4857 -4583 4863 -4383
rect 4727 -4759 4733 -4583
rect 4767 -4759 4863 -4583
rect 4897 -4759 4903 -4383
rect 4727 -4771 4773 -4759
rect 4857 -4771 4903 -4759
rect 4975 -4383 5021 -4371
rect 4975 -4759 4981 -4383
rect 5015 -4759 5021 -4383
rect 4975 -4771 5021 -4759
rect 5093 -4383 5139 -4371
rect 5093 -4759 5099 -4383
rect 5133 -4759 5139 -4383
rect 5093 -4771 5139 -4759
rect 5211 -4383 5257 -4371
rect 5211 -4759 5217 -4383
rect 5251 -4759 5257 -4383
rect 5211 -4771 5257 -4759
rect 5329 -4383 5375 -4371
rect 5329 -4759 5335 -4383
rect 5369 -4759 5375 -4383
rect 5329 -4771 5375 -4759
rect 5447 -4383 5493 -4371
rect 5447 -4759 5453 -4383
rect 5487 -4759 5493 -4383
rect 5447 -4771 5493 -4759
rect 5565 -4383 5611 -4371
rect 5565 -4759 5571 -4383
rect 5605 -4583 5611 -4383
rect 5936 -4571 5970 -4268
rect 6395 -4268 7868 -4225
rect 6395 -4571 6429 -4268
rect 6761 -4371 6795 -4268
rect 6997 -4371 7031 -4268
rect 7233 -4371 7267 -4268
rect 7469 -4371 7503 -4268
rect 6755 -4383 6801 -4371
rect 5694 -4583 5740 -4571
rect 5605 -4759 5700 -4583
rect 5734 -4759 5740 -4583
rect 5565 -4771 5611 -4759
rect 5694 -4771 5740 -4759
rect 5812 -4583 5858 -4571
rect 5812 -4759 5818 -4583
rect 5852 -4759 5858 -4583
rect 5812 -4771 5858 -4759
rect 5930 -4583 5976 -4571
rect 5930 -4759 5936 -4583
rect 5970 -4759 5976 -4583
rect 5930 -4771 5976 -4759
rect 6048 -4583 6094 -4571
rect 6048 -4759 6054 -4583
rect 6088 -4759 6094 -4583
rect 6048 -4771 6094 -4759
rect 6271 -4583 6317 -4571
rect 6271 -4759 6277 -4583
rect 6311 -4759 6317 -4583
rect 6271 -4771 6317 -4759
rect 6389 -4583 6435 -4571
rect 6389 -4759 6395 -4583
rect 6429 -4759 6435 -4583
rect 6389 -4771 6435 -4759
rect 6507 -4583 6553 -4571
rect 6507 -4759 6513 -4583
rect 6547 -4759 6553 -4583
rect 6507 -4771 6553 -4759
rect 6625 -4583 6671 -4571
rect 6755 -4583 6761 -4383
rect 6625 -4759 6631 -4583
rect 6665 -4759 6761 -4583
rect 6795 -4759 6801 -4383
rect 6625 -4771 6671 -4759
rect 6755 -4771 6801 -4759
rect 6873 -4383 6919 -4371
rect 6873 -4759 6879 -4383
rect 6913 -4759 6919 -4383
rect 6873 -4771 6919 -4759
rect 6991 -4383 7037 -4371
rect 6991 -4759 6997 -4383
rect 7031 -4759 7037 -4383
rect 6991 -4771 7037 -4759
rect 7109 -4383 7155 -4371
rect 7109 -4759 7115 -4383
rect 7149 -4759 7155 -4383
rect 7109 -4771 7155 -4759
rect 7227 -4383 7273 -4371
rect 7227 -4759 7233 -4383
rect 7267 -4759 7273 -4383
rect 7227 -4771 7273 -4759
rect 7345 -4383 7391 -4371
rect 7345 -4759 7351 -4383
rect 7385 -4759 7391 -4383
rect 7345 -4771 7391 -4759
rect 7463 -4383 7509 -4371
rect 7463 -4759 7469 -4383
rect 7503 -4583 7509 -4383
rect 7834 -4571 7868 -4268
rect 7592 -4583 7638 -4571
rect 7503 -4759 7598 -4583
rect 7632 -4759 7638 -4583
rect 7463 -4771 7509 -4759
rect 7592 -4771 7638 -4759
rect 7710 -4583 7756 -4571
rect 7710 -4759 7716 -4583
rect 7750 -4759 7756 -4583
rect 7710 -4771 7756 -4759
rect 7828 -4583 7874 -4571
rect 7828 -4759 7834 -4583
rect 7868 -4759 7874 -4583
rect 7828 -4771 7874 -4759
rect 7946 -4583 7992 -4571
rect 7946 -4759 7952 -4583
rect 7986 -4759 7992 -4583
rect 7946 -4771 7992 -4759
rect 3744 -4820 3884 -4814
rect 4379 -4805 4413 -4771
rect 4981 -4805 5015 -4771
rect 5217 -4805 5251 -4771
rect 3636 -4849 3744 -4839
rect 4379 -4840 4538 -4805
rect 4981 -4840 5251 -4805
rect 5818 -4805 5852 -4771
rect 6054 -4805 6088 -4771
rect 5818 -4840 6088 -4805
rect 6277 -4805 6311 -4771
rect 6879 -4805 6913 -4771
rect 7115 -4805 7149 -4771
rect 6277 -4840 6436 -4805
rect 6879 -4840 7149 -4805
rect 7716 -4805 7750 -4771
rect 7952 -4805 7986 -4771
rect 7716 -4840 7986 -4805
rect 3009 -4881 3024 -4879
rect 2924 -4895 3024 -4881
rect 2924 -4938 3024 -4937
rect 2545 -4959 3024 -4938
rect 3313 -4959 3379 -4863
rect 2545 -5007 3379 -4959
rect 2545 -5036 3024 -5007
rect 2545 -5038 2650 -5036
rect 2924 -5037 3024 -5036
rect 2378 -5223 2388 -5144
rect 2481 -5223 2491 -5144
rect 3376 -5153 3455 -5141
rect 715 -5317 1421 -5313
rect 239 -5329 285 -5317
rect -1124 -5474 199 -5457
rect -1124 -5537 -760 -5474
rect -679 -5537 199 -5474
rect -1124 -5555 199 -5537
rect 123 -5557 199 -5555
rect -1121 -5585 23 -5584
rect -1121 -5593 87 -5585
rect -1121 -5674 -630 -5593
rect -528 -5674 87 -5593
rect -1121 -5685 87 -5674
rect -357 -8565 -239 -5685
rect 9 -5834 63 -5685
rect 123 -5749 177 -5557
rect 239 -5705 245 -5329
rect 279 -5705 285 -5329
rect 239 -5717 285 -5705
rect 357 -5329 403 -5317
rect 357 -5705 363 -5329
rect 397 -5705 403 -5329
rect 357 -5717 403 -5705
rect 475 -5329 521 -5317
rect 475 -5705 481 -5329
rect 515 -5678 521 -5329
rect 592 -5329 638 -5317
rect 592 -5505 598 -5329
rect 632 -5505 638 -5329
rect 592 -5512 638 -5505
rect 710 -5329 1421 -5317
rect 710 -5505 716 -5329
rect 750 -5342 1421 -5329
rect 750 -5505 756 -5342
rect 1000 -5421 1421 -5342
rect 1000 -5422 1104 -5421
rect 592 -5517 641 -5512
rect 710 -5517 756 -5505
rect 598 -5678 641 -5517
rect 515 -5705 641 -5678
rect 475 -5717 641 -5705
rect 481 -5721 641 -5717
rect 123 -5755 354 -5749
rect 123 -5789 304 -5755
rect 338 -5789 354 -5755
rect 123 -5805 354 -5789
rect 406 -5755 472 -5749
rect 406 -5789 422 -5755
rect 456 -5789 472 -5755
rect 406 -5834 472 -5789
rect 9 -5842 472 -5834
rect 9 -5874 473 -5842
rect 565 -5858 641 -5721
rect 561 -5918 571 -5858
rect 633 -5918 643 -5858
rect 2389 -6397 2482 -5223
rect 3376 -5252 3382 -5153
rect 3307 -5272 3382 -5252
rect 3449 -5252 3455 -5153
rect 3449 -5272 3527 -5252
rect 3307 -5380 3351 -5272
rect 3483 -5380 3527 -5272
rect 3307 -5422 3527 -5380
rect 2911 -5452 3888 -5422
rect 2911 -5558 2943 -5452
rect 3147 -5558 3179 -5452
rect 3383 -5558 3415 -5452
rect 3619 -5558 3651 -5452
rect 3854 -5558 3888 -5452
rect 2904 -5570 2950 -5558
rect 2904 -5746 2910 -5570
rect 2944 -5746 2950 -5570
rect 2904 -5758 2950 -5746
rect 3022 -5570 3068 -5558
rect 3022 -5746 3028 -5570
rect 3062 -5746 3068 -5570
rect 3022 -5758 3068 -5746
rect 3140 -5570 3186 -5558
rect 3140 -5746 3146 -5570
rect 3180 -5746 3186 -5570
rect 3140 -5758 3186 -5746
rect 3258 -5570 3304 -5558
rect 3258 -5746 3264 -5570
rect 3298 -5746 3304 -5570
rect 3258 -5758 3304 -5746
rect 3376 -5570 3422 -5558
rect 3376 -5746 3382 -5570
rect 3416 -5746 3422 -5570
rect 3376 -5758 3422 -5746
rect 3494 -5570 3540 -5558
rect 3494 -5746 3500 -5570
rect 3534 -5746 3540 -5570
rect 3494 -5758 3540 -5746
rect 3612 -5570 3658 -5558
rect 3612 -5746 3618 -5570
rect 3652 -5746 3658 -5570
rect 3612 -5758 3658 -5746
rect 3730 -5570 3776 -5558
rect 3730 -5746 3736 -5570
rect 3770 -5746 3776 -5570
rect 3730 -5758 3776 -5746
rect 3848 -5570 3894 -5558
rect 3848 -5746 3854 -5570
rect 3888 -5746 3894 -5570
rect 3848 -5758 3894 -5746
rect 3966 -5570 4012 -5558
rect 3966 -5746 3972 -5570
rect 4006 -5746 4012 -5570
rect 3966 -5758 4012 -5746
rect 4504 -5624 4538 -4840
rect 5217 -4902 5251 -4840
rect 4806 -4940 5548 -4902
rect 4806 -5064 4840 -4940
rect 5042 -5064 5076 -4940
rect 5278 -5064 5312 -4940
rect 5514 -5064 5548 -4940
rect 5804 -5047 5814 -4981
rect 5877 -5047 5887 -4981
rect 4800 -5076 4846 -5064
rect 4800 -5452 4806 -5076
rect 4840 -5452 4846 -5076
rect 4800 -5464 4846 -5452
rect 4918 -5076 4964 -5064
rect 4918 -5452 4924 -5076
rect 4958 -5452 4964 -5076
rect 4918 -5464 4964 -5452
rect 5036 -5076 5082 -5064
rect 5036 -5452 5042 -5076
rect 5076 -5452 5082 -5076
rect 5036 -5464 5082 -5452
rect 5154 -5076 5200 -5064
rect 5154 -5452 5160 -5076
rect 5194 -5452 5200 -5076
rect 5154 -5464 5200 -5452
rect 5272 -5076 5318 -5064
rect 5272 -5452 5278 -5076
rect 5312 -5452 5318 -5076
rect 5272 -5464 5318 -5452
rect 5390 -5076 5436 -5064
rect 5390 -5452 5396 -5076
rect 5430 -5452 5436 -5076
rect 5390 -5464 5436 -5452
rect 5508 -5076 5554 -5064
rect 5508 -5452 5514 -5076
rect 5548 -5452 5554 -5076
rect 5508 -5464 5554 -5452
rect 5920 -5623 5954 -4840
rect 5647 -5624 5954 -5623
rect 4504 -5629 4820 -5624
rect 5534 -5629 5954 -5624
rect 4504 -5640 4887 -5629
rect 4504 -5667 4836 -5640
rect 3027 -5852 3063 -5758
rect 3263 -5852 3299 -5758
rect 3499 -5851 3535 -5758
rect 3661 -5806 3727 -5799
rect 3661 -5840 3677 -5806
rect 3711 -5840 3727 -5806
rect 3661 -5851 3727 -5840
rect 3499 -5852 3727 -5851
rect 3027 -5881 3727 -5852
rect 3027 -5882 3609 -5881
rect 3147 -5995 3181 -5882
rect 3543 -5923 3609 -5882
rect 3543 -5957 3559 -5923
rect 3593 -5957 3609 -5923
rect 3543 -5964 3609 -5957
rect 3971 -5991 4006 -5758
rect 4504 -5796 4538 -5667
rect 4820 -5674 4836 -5667
rect 4870 -5674 4887 -5640
rect 4820 -5680 4887 -5674
rect 5467 -5640 5954 -5629
rect 5467 -5674 5484 -5640
rect 5518 -5667 5954 -5640
rect 5518 -5674 5534 -5667
rect 5647 -5668 5954 -5667
rect 5467 -5680 5534 -5674
rect 4645 -5707 4701 -5695
rect 4645 -5741 4651 -5707
rect 4685 -5708 4701 -5707
rect 5758 -5708 5814 -5696
rect 4685 -5724 5152 -5708
rect 4685 -5741 5102 -5724
rect 4645 -5757 5102 -5741
rect 5086 -5758 5102 -5757
rect 5136 -5758 5152 -5724
rect 5086 -5765 5152 -5758
rect 5204 -5723 5774 -5708
rect 5204 -5757 5220 -5723
rect 5254 -5742 5774 -5723
rect 5808 -5742 5814 -5708
rect 5254 -5757 5814 -5742
rect 5204 -5767 5271 -5757
rect 5758 -5758 5814 -5757
rect 5920 -5796 5954 -5668
rect 6402 -5624 6436 -4840
rect 7115 -4902 7149 -4840
rect 6704 -4940 7446 -4902
rect 6704 -5064 6738 -4940
rect 6940 -5064 6974 -4940
rect 7176 -5064 7210 -4940
rect 7412 -5064 7446 -4940
rect 6698 -5076 6744 -5064
rect 6698 -5452 6704 -5076
rect 6738 -5452 6744 -5076
rect 6698 -5464 6744 -5452
rect 6816 -5076 6862 -5064
rect 6816 -5452 6822 -5076
rect 6856 -5452 6862 -5076
rect 6816 -5464 6862 -5452
rect 6934 -5076 6980 -5064
rect 6934 -5452 6940 -5076
rect 6974 -5452 6980 -5076
rect 6934 -5464 6980 -5452
rect 7052 -5076 7098 -5064
rect 7052 -5452 7058 -5076
rect 7092 -5452 7098 -5076
rect 7052 -5464 7098 -5452
rect 7170 -5076 7216 -5064
rect 7170 -5452 7176 -5076
rect 7210 -5452 7216 -5076
rect 7170 -5464 7216 -5452
rect 7288 -5076 7334 -5064
rect 7288 -5452 7294 -5076
rect 7328 -5452 7334 -5076
rect 7288 -5464 7334 -5452
rect 7406 -5076 7452 -5064
rect 7406 -5452 7412 -5076
rect 7446 -5452 7452 -5076
rect 7406 -5464 7452 -5452
rect 7818 -5623 7852 -4840
rect 7430 -5624 7499 -5623
rect 7545 -5624 7852 -5623
rect 6402 -5629 6718 -5624
rect 7430 -5628 7852 -5624
rect 6402 -5640 6785 -5629
rect 6402 -5667 6734 -5640
rect 6402 -5796 6436 -5667
rect 6718 -5674 6734 -5667
rect 6768 -5674 6785 -5640
rect 6718 -5680 6785 -5674
rect 7363 -5639 7852 -5628
rect 7363 -5673 7380 -5639
rect 7414 -5667 7852 -5639
rect 7414 -5673 7430 -5667
rect 7545 -5668 7852 -5667
rect 7363 -5679 7430 -5673
rect 6543 -5707 6599 -5695
rect 6543 -5741 6549 -5707
rect 6583 -5708 6599 -5707
rect 7656 -5708 7712 -5696
rect 6583 -5724 7050 -5708
rect 6583 -5741 7000 -5724
rect 6543 -5757 7000 -5741
rect 6984 -5758 7000 -5757
rect 7034 -5758 7050 -5724
rect 6984 -5765 7050 -5758
rect 7102 -5723 7672 -5708
rect 7102 -5757 7118 -5723
rect 7152 -5742 7672 -5723
rect 7706 -5742 7712 -5708
rect 7152 -5757 7712 -5742
rect 7102 -5767 7169 -5757
rect 7656 -5758 7712 -5757
rect 7818 -5796 7852 -5668
rect 7933 -5018 8000 -4994
rect 7933 -5052 7950 -5018
rect 7984 -5052 8000 -5018
rect 3617 -5995 4006 -5991
rect 3141 -6007 3187 -5995
rect 3141 -6383 3147 -6007
rect 3181 -6383 3187 -6007
rect 3141 -6395 3187 -6383
rect 3259 -6007 3305 -5995
rect 3259 -6383 3265 -6007
rect 3299 -6383 3305 -6007
rect 3259 -6395 3305 -6383
rect 3377 -6007 3423 -5995
rect 3377 -6383 3383 -6007
rect 3417 -6359 3423 -6007
rect 3494 -6007 3540 -5995
rect 3494 -6183 3500 -6007
rect 3534 -6183 3540 -6007
rect 3494 -6195 3540 -6183
rect 3612 -6007 4006 -5995
rect 4498 -5808 4544 -5796
rect 4498 -5984 4504 -5808
rect 4538 -5984 4544 -5808
rect 4498 -5996 4544 -5984
rect 4616 -5808 4662 -5796
rect 4616 -5984 4622 -5808
rect 4656 -5984 4662 -5808
rect 4616 -5996 4662 -5984
rect 4918 -5808 4964 -5796
rect 3612 -6183 3618 -6007
rect 3652 -6020 4006 -6007
rect 3652 -6183 3658 -6020
rect 3928 -6023 4006 -6020
rect 3928 -6075 3938 -6023
rect 4001 -6075 4011 -6023
rect 3933 -6081 4006 -6075
rect 3612 -6195 3658 -6183
rect 3500 -6311 3535 -6195
rect 4621 -6290 4655 -5996
rect 4918 -6184 4924 -5808
rect 4958 -6184 4964 -5808
rect 4918 -6196 4964 -6184
rect 5036 -5808 5082 -5796
rect 5036 -6184 5042 -5808
rect 5076 -6184 5082 -5808
rect 5036 -6196 5082 -6184
rect 5154 -5808 5200 -5796
rect 5154 -6184 5160 -5808
rect 5194 -6184 5200 -5808
rect 5154 -6196 5200 -6184
rect 5272 -5808 5318 -5796
rect 5272 -6184 5278 -5808
rect 5312 -6184 5318 -5808
rect 5272 -6196 5318 -6184
rect 5390 -5808 5436 -5796
rect 5390 -6184 5396 -5808
rect 5430 -6184 5436 -5808
rect 5796 -5808 5842 -5796
rect 5796 -5984 5802 -5808
rect 5836 -5984 5842 -5808
rect 5796 -5996 5842 -5984
rect 5914 -5808 5960 -5796
rect 5914 -5984 5920 -5808
rect 5954 -5984 5960 -5808
rect 5914 -5996 5960 -5984
rect 6396 -5808 6442 -5796
rect 6396 -5984 6402 -5808
rect 6436 -5984 6442 -5808
rect 6396 -5996 6442 -5984
rect 6514 -5808 6560 -5796
rect 6514 -5984 6520 -5808
rect 6554 -5984 6560 -5808
rect 6514 -5996 6560 -5984
rect 6816 -5808 6862 -5796
rect 5390 -6196 5436 -6184
rect 5278 -6290 5312 -6196
rect 5802 -6290 5835 -5996
rect 3631 -6311 3739 -6301
rect 3500 -6359 3631 -6311
rect 4621 -6322 5835 -6290
rect 6519 -6290 6553 -5996
rect 6816 -6184 6822 -5808
rect 6856 -6184 6862 -5808
rect 6816 -6196 6862 -6184
rect 6934 -5808 6980 -5796
rect 6934 -6184 6940 -5808
rect 6974 -6184 6980 -5808
rect 6934 -6196 6980 -6184
rect 7052 -5808 7098 -5796
rect 7052 -6184 7058 -5808
rect 7092 -6184 7098 -5808
rect 7052 -6196 7098 -6184
rect 7170 -5808 7216 -5796
rect 7170 -6184 7176 -5808
rect 7210 -6184 7216 -5808
rect 7170 -6196 7216 -6184
rect 7288 -5808 7334 -5796
rect 7288 -6184 7294 -5808
rect 7328 -6184 7334 -5808
rect 7694 -5808 7740 -5796
rect 7694 -5984 7700 -5808
rect 7734 -5984 7740 -5808
rect 7694 -5996 7740 -5984
rect 7812 -5808 7858 -5796
rect 7812 -5984 7818 -5808
rect 7852 -5984 7858 -5808
rect 7812 -5996 7858 -5984
rect 7288 -6196 7334 -6184
rect 7176 -6290 7210 -6196
rect 7700 -6290 7733 -5996
rect 6519 -6322 7733 -6290
rect 3739 -6339 3884 -6333
rect 3417 -6383 3631 -6359
rect 3377 -6395 3631 -6383
rect 2389 -6399 2974 -6397
rect 3383 -6399 3631 -6395
rect 2389 -6427 3019 -6399
rect 2389 -6433 3256 -6427
rect 2389 -6467 3206 -6433
rect 3240 -6467 3256 -6433
rect 2389 -6483 3256 -6467
rect 3308 -6433 3374 -6427
rect 3308 -6467 3324 -6433
rect 3358 -6467 3374 -6433
rect 3557 -6443 3631 -6399
rect 3872 -6406 3884 -6339
rect 3739 -6412 3884 -6406
rect 5114 -6407 5246 -6322
rect 7012 -6407 7144 -6322
rect 3631 -6453 3739 -6443
rect 2389 -6499 3019 -6483
rect 2389 -6503 2974 -6499
rect 2389 -6504 2490 -6503
rect 2919 -6552 3019 -6541
rect 2883 -6658 2893 -6552
rect 3005 -6563 3019 -6552
rect 3308 -6563 3374 -6467
rect 5104 -6515 5114 -6407
rect 5246 -6515 5256 -6407
rect 7002 -6515 7012 -6407
rect 7144 -6515 7154 -6407
rect 7933 -6435 8000 -5052
rect 8061 -5481 8219 -3254
rect 8061 -5579 8073 -5481
rect 8205 -5556 8219 -5481
rect 8303 -3663 8817 -3639
rect 8303 -3769 8665 -3663
rect 8777 -3676 8817 -3663
rect 8777 -3769 8819 -3676
rect 8303 -3780 8819 -3769
rect 8303 -3781 8817 -3780
rect 8205 -5579 8217 -5556
rect 8061 -5585 8217 -5579
rect 3005 -6611 3374 -6563
rect 3005 -6641 3019 -6611
rect 3005 -6658 3015 -6641
rect 3307 -6714 3373 -6611
rect 5138 -6656 5144 -6515
rect 5211 -6656 5217 -6515
rect 5138 -6668 5217 -6656
rect 7933 -6714 7999 -6435
rect 3305 -6794 7999 -6714
rect 6719 -7299 7183 -7267
rect 7271 -7283 7281 -7223
rect 7343 -7283 7353 -7223
rect 6719 -7307 7182 -7299
rect 6719 -7456 6773 -7307
rect 6334 -7462 6773 -7456
rect 6332 -7548 6342 -7462
rect 6418 -7548 6773 -7462
rect 6334 -7556 6773 -7548
rect 6833 -7352 7064 -7336
rect 6833 -7386 7014 -7352
rect 7048 -7386 7064 -7352
rect 6833 -7392 7064 -7386
rect 7116 -7352 7182 -7307
rect 7116 -7386 7132 -7352
rect 7166 -7386 7182 -7352
rect 7116 -7392 7182 -7386
rect 6833 -7584 6887 -7392
rect 7275 -7420 7351 -7283
rect 7191 -7424 7351 -7420
rect 6569 -7589 6887 -7584
rect 6563 -7680 6573 -7589
rect 6702 -7680 6887 -7589
rect 6569 -7684 6887 -7680
rect 6949 -7436 6995 -7424
rect 6949 -7812 6955 -7436
rect 6989 -7812 6995 -7436
rect 6949 -7824 6995 -7812
rect 7067 -7436 7113 -7424
rect 7067 -7812 7073 -7436
rect 7107 -7812 7113 -7436
rect 7067 -7824 7113 -7812
rect 7185 -7436 7351 -7424
rect 7185 -7812 7191 -7436
rect 7225 -7463 7351 -7436
rect 7225 -7812 7231 -7463
rect 7308 -7624 7351 -7463
rect 7185 -7824 7231 -7812
rect 7302 -7629 7351 -7624
rect 7302 -7636 7348 -7629
rect 7302 -7812 7308 -7636
rect 7342 -7812 7348 -7636
rect 7302 -7824 7348 -7812
rect 7420 -7636 7466 -7624
rect 7420 -7812 7426 -7636
rect 7460 -7799 7466 -7636
rect 8303 -7719 8439 -3781
rect 8940 -5146 9033 -3254
rect 9096 -3311 9562 -3289
rect 9850 -3311 9916 -3215
rect 11681 -3205 11687 -3029
rect 11721 -3205 11727 -3029
rect 11681 -3217 11727 -3205
rect 11799 -3029 11845 -3017
rect 11799 -3205 11805 -3029
rect 11839 -3205 11845 -3029
rect 11799 -3217 11845 -3205
rect 11917 -3029 11963 -3017
rect 11917 -3205 11923 -3029
rect 11957 -3205 11963 -3029
rect 11917 -3217 11963 -3205
rect 12035 -3029 12081 -3017
rect 12035 -3205 12041 -3029
rect 12075 -3084 12081 -3029
rect 12200 -3029 12246 -3017
rect 12200 -3084 12206 -3029
rect 12075 -3172 12206 -3084
rect 12075 -3205 12081 -3172
rect 12035 -3217 12081 -3205
rect 12200 -3205 12206 -3172
rect 12240 -3205 12246 -3029
rect 12200 -3217 12246 -3205
rect 12318 -3029 12364 -3017
rect 12318 -3205 12324 -3029
rect 12358 -3205 12364 -3029
rect 12318 -3217 12364 -3205
rect 12436 -3029 12482 -3017
rect 12436 -3205 12442 -3029
rect 12476 -3205 12482 -3029
rect 12436 -3217 12482 -3205
rect 12554 -3029 12600 -3017
rect 12554 -3205 12560 -3029
rect 12594 -3205 12600 -3029
rect 12554 -3217 12600 -3205
rect 11687 -3256 11721 -3217
rect 11923 -3256 11957 -3217
rect 11687 -3291 11957 -3256
rect 12324 -3255 12357 -3217
rect 12560 -3255 12593 -3217
rect 12324 -3291 12593 -3255
rect 9096 -3359 9916 -3311
rect 11721 -3292 11957 -3291
rect 9096 -3390 9562 -3359
rect 11721 -3366 11853 -3292
rect 9096 -3646 9201 -3390
rect 11711 -3474 11721 -3366
rect 11853 -3474 11863 -3366
rect 9932 -3547 10011 -3535
rect 9096 -3752 9159 -3646
rect 9271 -3752 9281 -3646
rect 9932 -3650 9938 -3547
rect 9863 -3670 9938 -3650
rect 10005 -3650 10011 -3547
rect 11744 -3610 11750 -3474
rect 11817 -3610 11823 -3474
rect 11744 -3622 11823 -3610
rect 10005 -3670 10083 -3650
rect 9096 -3763 9245 -3752
rect 9096 -4940 9201 -3763
rect 9863 -3778 9907 -3670
rect 10039 -3778 10083 -3670
rect 9863 -3820 10083 -3778
rect 12661 -3805 12723 -2234
rect 12913 -2242 12959 -2230
rect 12913 -2618 12919 -2242
rect 12953 -2618 12959 -2242
rect 12913 -2630 12959 -2618
rect 13031 -2242 13077 -2230
rect 13031 -2618 13037 -2242
rect 13071 -2618 13077 -2242
rect 13031 -2630 13077 -2618
rect 13149 -2242 13195 -2230
rect 13149 -2618 13155 -2242
rect 13189 -2618 13195 -2242
rect 13149 -2630 13195 -2618
rect 13267 -2242 13313 -2230
rect 13267 -2618 13273 -2242
rect 13307 -2618 13313 -2242
rect 13267 -2630 13313 -2618
rect 13385 -2242 13431 -2230
rect 13385 -2618 13391 -2242
rect 13425 -2618 13431 -2242
rect 13385 -2630 13431 -2618
rect 13503 -2242 13549 -2230
rect 13503 -2618 13509 -2242
rect 13543 -2618 13549 -2242
rect 13503 -2630 13549 -2618
rect 13621 -2242 13667 -2230
rect 13621 -2618 13627 -2242
rect 13661 -2618 13667 -2242
rect 13621 -2630 13667 -2618
rect 12919 -2672 12953 -2630
rect 13155 -2672 13189 -2630
rect 12919 -2700 13189 -2672
rect 13273 -2671 13307 -2630
rect 13509 -2671 13543 -2630
rect 13273 -2700 13543 -2671
rect 12919 -2748 12953 -2700
rect 12919 -2778 12982 -2748
rect 12947 -2870 12982 -2778
rect 13454 -2808 13554 -2787
rect 13454 -2862 13468 -2808
rect 13533 -2862 13554 -2808
rect 13454 -2867 13554 -2862
rect 13627 -2813 13661 -2630
rect 13627 -2867 13736 -2813
rect 12947 -2906 13174 -2870
rect 12947 -3013 12982 -2906
rect 13108 -2940 13174 -2906
rect 13108 -2974 13124 -2940
rect 13158 -2974 13174 -2940
rect 13455 -2882 13552 -2867
rect 13455 -2949 13512 -2882
rect 13108 -2980 13174 -2974
rect 13349 -2985 13618 -2949
rect 13349 -3013 13382 -2985
rect 13585 -3013 13618 -2985
rect 13702 -3013 13736 -2867
rect 12823 -3025 12869 -3013
rect 12823 -3201 12829 -3025
rect 12863 -3201 12869 -3025
rect 12823 -3213 12869 -3201
rect 12941 -3025 12987 -3013
rect 12941 -3201 12947 -3025
rect 12981 -3201 12987 -3025
rect 12941 -3213 12987 -3201
rect 13059 -3025 13105 -3013
rect 13059 -3201 13065 -3025
rect 13099 -3201 13105 -3025
rect 13059 -3213 13105 -3201
rect 13177 -3025 13223 -3013
rect 13177 -3201 13183 -3025
rect 13217 -3080 13223 -3025
rect 13342 -3025 13388 -3013
rect 13342 -3080 13348 -3025
rect 13217 -3168 13348 -3080
rect 13217 -3201 13223 -3168
rect 13177 -3213 13223 -3201
rect 13342 -3201 13348 -3168
rect 13382 -3201 13388 -3025
rect 13342 -3213 13388 -3201
rect 13460 -3025 13506 -3013
rect 13460 -3201 13466 -3025
rect 13500 -3201 13506 -3025
rect 13460 -3213 13506 -3201
rect 13578 -3025 13624 -3013
rect 13578 -3201 13584 -3025
rect 13618 -3201 13624 -3025
rect 13578 -3213 13624 -3201
rect 13696 -3025 13742 -3013
rect 13696 -3201 13702 -3025
rect 13736 -3201 13742 -3025
rect 13696 -3213 13742 -3201
rect 14891 -3146 15031 2995
rect 15460 2703 15642 4191
rect 19061 3953 19140 3965
rect 16580 3897 16659 3909
rect 16580 3802 16586 3897
rect 16509 3782 16586 3802
rect 16653 3802 16659 3897
rect 19061 3836 19067 3953
rect 19134 3836 19140 3953
rect 20208 3952 20287 3964
rect 20208 3836 20214 3952
rect 20281 3836 20287 3952
rect 16653 3782 16729 3802
rect 16509 3674 16553 3782
rect 16685 3674 16729 3782
rect 18306 3740 18362 3748
rect 16509 3632 16729 3674
rect 17380 3732 18362 3740
rect 17380 3698 18322 3732
rect 18356 3698 18362 3732
rect 19025 3728 19035 3836
rect 19167 3773 19177 3836
rect 19167 3762 19179 3773
rect 19167 3728 19180 3762
rect 19436 3752 19492 3754
rect 17380 3682 18362 3698
rect 19035 3690 19180 3728
rect 17380 3681 18359 3682
rect 16113 3602 17090 3632
rect 16113 3496 16145 3602
rect 16349 3496 16381 3602
rect 16585 3496 16617 3602
rect 16821 3496 16853 3602
rect 17056 3496 17090 3602
rect 16106 3484 16152 3496
rect 16106 3308 16112 3484
rect 16146 3308 16152 3484
rect 16106 3296 16152 3308
rect 16224 3484 16270 3496
rect 16224 3308 16230 3484
rect 16264 3308 16270 3484
rect 16224 3296 16270 3308
rect 16342 3484 16388 3496
rect 16342 3308 16348 3484
rect 16382 3308 16388 3484
rect 16342 3296 16388 3308
rect 16460 3484 16506 3496
rect 16460 3308 16466 3484
rect 16500 3308 16506 3484
rect 16460 3296 16506 3308
rect 16578 3484 16624 3496
rect 16578 3308 16584 3484
rect 16618 3308 16624 3484
rect 16578 3296 16624 3308
rect 16696 3484 16742 3496
rect 16696 3308 16702 3484
rect 16736 3308 16742 3484
rect 16696 3296 16742 3308
rect 16814 3484 16860 3496
rect 16814 3308 16820 3484
rect 16854 3308 16860 3484
rect 16814 3296 16860 3308
rect 16932 3484 16978 3496
rect 16932 3308 16938 3484
rect 16972 3308 16978 3484
rect 16932 3296 16978 3308
rect 17050 3484 17096 3496
rect 17050 3308 17056 3484
rect 17090 3308 17096 3484
rect 17050 3296 17096 3308
rect 17168 3484 17214 3496
rect 17168 3308 17174 3484
rect 17208 3308 17214 3484
rect 17168 3296 17214 3308
rect 16229 3202 16265 3296
rect 16465 3202 16501 3296
rect 16701 3203 16737 3296
rect 16863 3248 16929 3255
rect 16863 3214 16879 3248
rect 16913 3214 16929 3248
rect 16863 3203 16929 3214
rect 16701 3202 16929 3203
rect 16229 3173 16929 3202
rect 16229 3172 16811 3173
rect 16349 3059 16383 3172
rect 16745 3131 16811 3172
rect 16745 3097 16761 3131
rect 16795 3097 16811 3131
rect 16745 3090 16811 3097
rect 17173 3091 17208 3296
rect 17380 3091 17447 3681
rect 19139 3658 19180 3690
rect 19426 3686 19436 3752
rect 19492 3686 19502 3752
rect 20172 3728 20182 3836
rect 20314 3773 20324 3836
rect 20314 3762 20326 3773
rect 20314 3728 20327 3762
rect 20182 3690 20327 3728
rect 20286 3662 20327 3690
rect 18555 3630 18825 3658
rect 18296 3564 18306 3630
rect 18372 3564 18382 3630
rect 18555 3568 18589 3630
rect 18791 3568 18825 3630
rect 18909 3630 19180 3658
rect 19697 3634 19967 3662
rect 18909 3568 18943 3630
rect 19145 3568 19180 3630
rect 19321 3618 19492 3634
rect 19321 3584 19452 3618
rect 19486 3584 19492 3618
rect 19321 3568 19492 3584
rect 19697 3572 19731 3634
rect 19933 3572 19967 3634
rect 20051 3634 20327 3662
rect 20051 3572 20085 3634
rect 20287 3572 20327 3634
rect 18431 3556 18477 3568
rect 18431 3180 18437 3556
rect 18471 3180 18477 3556
rect 18431 3168 18477 3180
rect 18549 3556 18595 3568
rect 18549 3180 18555 3556
rect 18589 3180 18595 3556
rect 18549 3168 18595 3180
rect 18667 3556 18713 3568
rect 18667 3180 18673 3556
rect 18707 3180 18713 3556
rect 18667 3168 18713 3180
rect 18785 3556 18831 3568
rect 18785 3180 18791 3556
rect 18825 3180 18831 3556
rect 18785 3168 18831 3180
rect 18903 3556 18949 3568
rect 18903 3180 18909 3556
rect 18943 3180 18949 3556
rect 18903 3168 18949 3180
rect 19021 3556 19067 3568
rect 19021 3180 19027 3556
rect 19061 3180 19067 3556
rect 19021 3168 19067 3180
rect 19139 3556 19185 3568
rect 19139 3180 19145 3556
rect 19179 3180 19185 3556
rect 19139 3168 19185 3180
rect 17173 3063 17447 3091
rect 16819 3059 17447 3063
rect 15459 2654 15642 2703
rect 16343 3047 16389 3059
rect 16343 2671 16349 3047
rect 16383 2671 16389 3047
rect 16343 2659 16389 2671
rect 16461 3047 16507 3059
rect 16461 2671 16467 3047
rect 16501 2671 16507 3047
rect 16461 2659 16507 2671
rect 16579 3047 16625 3059
rect 16579 2671 16585 3047
rect 16619 2695 16625 3047
rect 16696 3047 16742 3059
rect 16696 2871 16702 3047
rect 16736 2871 16742 3047
rect 16696 2859 16742 2871
rect 16814 3047 17447 3059
rect 16814 2871 16820 3047
rect 16854 3034 17447 3047
rect 18437 3126 18471 3168
rect 18673 3126 18707 3168
rect 18437 3098 18707 3126
rect 18791 3127 18825 3168
rect 19027 3127 19061 3168
rect 18791 3098 19061 3127
rect 18437 3050 18471 3098
rect 16854 2871 16860 3034
rect 18437 3020 18500 3050
rect 16814 2859 16860 2871
rect 18465 2928 18500 3020
rect 18465 2892 18692 2928
rect 18962 2917 18972 3014
rect 19071 2917 19081 3014
rect 19145 2985 19179 3168
rect 19145 2931 19254 2985
rect 16702 2743 16737 2859
rect 18465 2785 18500 2892
rect 18626 2858 18692 2892
rect 18626 2824 18642 2858
rect 18676 2824 18692 2858
rect 18973 2916 19070 2917
rect 18973 2849 19030 2916
rect 18626 2818 18692 2824
rect 18867 2813 19136 2849
rect 18867 2785 18900 2813
rect 19103 2785 19136 2813
rect 19220 2785 19254 2931
rect 18341 2773 18387 2785
rect 16833 2743 16941 2753
rect 16702 2695 16833 2743
rect 16941 2706 17082 2712
rect 16619 2671 16833 2695
rect 16579 2659 16833 2671
rect 16585 2655 16833 2659
rect 15459 2627 16221 2654
rect 15459 2621 16458 2627
rect 15459 2587 16408 2621
rect 16442 2587 16458 2621
rect 15459 2571 16458 2587
rect 16510 2621 16576 2627
rect 16510 2587 16526 2621
rect 16560 2587 16576 2621
rect 16759 2611 16833 2655
rect 17070 2639 17082 2706
rect 16941 2633 17082 2639
rect 16833 2601 16941 2611
rect 15459 2555 16221 2571
rect 15459 2554 16158 2555
rect 15459 2550 15693 2554
rect 15311 1037 15476 1057
rect 15311 920 15323 1037
rect 15462 1014 15476 1037
rect 15462 920 15477 1014
rect 15311 919 15330 920
rect 15442 919 15477 920
rect 15311 910 15477 919
rect 15311 909 15476 910
rect 15311 908 15444 909
rect 15600 656 15693 2550
rect 15756 2491 16222 2513
rect 16510 2491 16576 2587
rect 18341 2597 18347 2773
rect 18381 2597 18387 2773
rect 18341 2585 18387 2597
rect 18459 2773 18505 2785
rect 18459 2597 18465 2773
rect 18499 2597 18505 2773
rect 18459 2585 18505 2597
rect 18577 2773 18623 2785
rect 18577 2597 18583 2773
rect 18617 2597 18623 2773
rect 18577 2585 18623 2597
rect 18695 2773 18741 2785
rect 18695 2597 18701 2773
rect 18735 2718 18741 2773
rect 18860 2773 18906 2785
rect 18860 2718 18866 2773
rect 18735 2630 18866 2718
rect 18735 2597 18741 2630
rect 18695 2585 18741 2597
rect 18860 2597 18866 2630
rect 18900 2597 18906 2773
rect 18860 2585 18906 2597
rect 18978 2773 19024 2785
rect 18978 2597 18984 2773
rect 19018 2597 19024 2773
rect 18978 2585 19024 2597
rect 19096 2773 19142 2785
rect 19096 2597 19102 2773
rect 19136 2597 19142 2773
rect 19096 2585 19142 2597
rect 19214 2773 19260 2785
rect 19214 2597 19220 2773
rect 19254 2597 19260 2773
rect 19214 2585 19260 2597
rect 18347 2546 18381 2585
rect 18583 2546 18617 2585
rect 18347 2511 18617 2546
rect 18984 2547 19017 2585
rect 19220 2547 19253 2585
rect 18984 2511 19253 2547
rect 15756 2443 16576 2491
rect 18381 2510 18617 2511
rect 15756 2412 16222 2443
rect 18381 2436 18513 2510
rect 15756 2156 15861 2412
rect 18371 2328 18381 2436
rect 18513 2328 18523 2436
rect 16595 2249 16674 2261
rect 15756 2050 15819 2156
rect 15931 2050 15941 2156
rect 16595 2152 16601 2249
rect 16523 2132 16601 2152
rect 16668 2152 16674 2249
rect 18403 2194 18409 2328
rect 18476 2194 18482 2328
rect 18403 2182 18482 2194
rect 16668 2132 16743 2152
rect 15756 2039 15905 2050
rect 15756 862 15861 2039
rect 16523 2024 16567 2132
rect 16699 2024 16743 2132
rect 16523 1982 16743 2024
rect 19321 1997 19383 3568
rect 19573 3560 19619 3572
rect 19573 3184 19579 3560
rect 19613 3184 19619 3560
rect 19573 3172 19619 3184
rect 19691 3560 19737 3572
rect 19691 3184 19697 3560
rect 19731 3184 19737 3560
rect 19691 3172 19737 3184
rect 19809 3560 19855 3572
rect 19809 3184 19815 3560
rect 19849 3184 19855 3560
rect 19809 3172 19855 3184
rect 19927 3560 19973 3572
rect 19927 3184 19933 3560
rect 19967 3184 19973 3560
rect 19927 3172 19973 3184
rect 20045 3560 20091 3572
rect 20045 3184 20051 3560
rect 20085 3184 20091 3560
rect 20045 3172 20091 3184
rect 20163 3560 20209 3572
rect 20163 3184 20169 3560
rect 20203 3184 20209 3560
rect 20163 3172 20209 3184
rect 20281 3560 20327 3572
rect 20281 3184 20287 3560
rect 20321 3184 20327 3560
rect 20281 3172 20327 3184
rect 19579 3130 19613 3172
rect 19815 3130 19849 3172
rect 19579 3102 19849 3130
rect 19933 3131 19967 3172
rect 20169 3131 20203 3172
rect 19933 3102 20203 3131
rect 19579 3054 19613 3102
rect 19579 3024 19642 3054
rect 19607 2932 19642 3024
rect 20114 2994 20214 3015
rect 20114 2940 20128 2994
rect 20193 2940 20214 2994
rect 20114 2935 20214 2940
rect 20287 2989 20321 3172
rect 20287 2935 20396 2989
rect 19607 2896 19834 2932
rect 19607 2789 19642 2896
rect 19768 2862 19834 2896
rect 19768 2828 19784 2862
rect 19818 2828 19834 2862
rect 20115 2920 20212 2935
rect 20115 2853 20172 2920
rect 19768 2822 19834 2828
rect 20009 2817 20278 2853
rect 20009 2789 20042 2817
rect 20245 2789 20278 2817
rect 20362 2789 20396 2935
rect 19483 2777 19529 2789
rect 19483 2601 19489 2777
rect 19523 2601 19529 2777
rect 19483 2589 19529 2601
rect 19601 2777 19647 2789
rect 19601 2601 19607 2777
rect 19641 2601 19647 2777
rect 19601 2589 19647 2601
rect 19719 2777 19765 2789
rect 19719 2601 19725 2777
rect 19759 2601 19765 2777
rect 19719 2589 19765 2601
rect 19837 2777 19883 2789
rect 19837 2601 19843 2777
rect 19877 2722 19883 2777
rect 20002 2777 20048 2789
rect 20002 2722 20008 2777
rect 19877 2634 20008 2722
rect 19877 2601 19883 2634
rect 19837 2589 19883 2601
rect 20002 2601 20008 2634
rect 20042 2601 20048 2777
rect 20002 2589 20048 2601
rect 20120 2777 20166 2789
rect 20120 2601 20126 2777
rect 20160 2601 20166 2777
rect 20120 2589 20166 2601
rect 20238 2777 20284 2789
rect 20238 2601 20244 2777
rect 20278 2601 20284 2777
rect 20238 2589 20284 2601
rect 20356 2777 20402 2789
rect 20356 2601 20362 2777
rect 20396 2601 20402 2777
rect 22086 2722 22268 4259
rect 25684 4018 25763 4030
rect 23200 3966 23279 3978
rect 23200 3870 23206 3966
rect 23134 3850 23206 3870
rect 23273 3870 23279 3966
rect 25684 3904 25690 4018
rect 25757 3904 25763 4018
rect 26833 4024 26912 4036
rect 26833 3904 26839 4024
rect 26906 3904 26912 4024
rect 23273 3850 23354 3870
rect 23134 3742 23178 3850
rect 23310 3742 23354 3850
rect 24931 3808 24987 3816
rect 23134 3700 23354 3742
rect 24005 3800 24987 3808
rect 24005 3766 24947 3800
rect 24981 3766 24987 3800
rect 25650 3796 25660 3904
rect 25792 3841 25802 3904
rect 25792 3830 25804 3841
rect 25792 3796 25805 3830
rect 26061 3820 26117 3822
rect 24005 3750 24987 3766
rect 25660 3758 25805 3796
rect 24005 3749 24984 3750
rect 22738 3670 23715 3700
rect 22738 3564 22770 3670
rect 22974 3564 23006 3670
rect 23210 3564 23242 3670
rect 23446 3564 23478 3670
rect 23681 3564 23715 3670
rect 22731 3552 22777 3564
rect 22731 3376 22737 3552
rect 22771 3376 22777 3552
rect 22731 3364 22777 3376
rect 22849 3552 22895 3564
rect 22849 3376 22855 3552
rect 22889 3376 22895 3552
rect 22849 3364 22895 3376
rect 22967 3552 23013 3564
rect 22967 3376 22973 3552
rect 23007 3376 23013 3552
rect 22967 3364 23013 3376
rect 23085 3552 23131 3564
rect 23085 3376 23091 3552
rect 23125 3376 23131 3552
rect 23085 3364 23131 3376
rect 23203 3552 23249 3564
rect 23203 3376 23209 3552
rect 23243 3376 23249 3552
rect 23203 3364 23249 3376
rect 23321 3552 23367 3564
rect 23321 3376 23327 3552
rect 23361 3376 23367 3552
rect 23321 3364 23367 3376
rect 23439 3552 23485 3564
rect 23439 3376 23445 3552
rect 23479 3376 23485 3552
rect 23439 3364 23485 3376
rect 23557 3552 23603 3564
rect 23557 3376 23563 3552
rect 23597 3376 23603 3552
rect 23557 3364 23603 3376
rect 23675 3552 23721 3564
rect 23675 3376 23681 3552
rect 23715 3376 23721 3552
rect 23675 3364 23721 3376
rect 23793 3552 23839 3564
rect 23793 3376 23799 3552
rect 23833 3376 23839 3552
rect 23793 3364 23839 3376
rect 22854 3270 22890 3364
rect 23090 3270 23126 3364
rect 23326 3271 23362 3364
rect 23488 3316 23554 3323
rect 23488 3282 23504 3316
rect 23538 3282 23554 3316
rect 23488 3271 23554 3282
rect 23326 3270 23554 3271
rect 22854 3241 23554 3270
rect 22854 3240 23436 3241
rect 22974 3127 23008 3240
rect 23370 3199 23436 3240
rect 23370 3165 23386 3199
rect 23420 3165 23436 3199
rect 23370 3158 23436 3165
rect 23798 3159 23833 3364
rect 24005 3159 24072 3749
rect 25764 3726 25805 3758
rect 26051 3754 26061 3820
rect 26117 3754 26127 3820
rect 26797 3796 26807 3904
rect 26939 3841 26949 3904
rect 26939 3830 26951 3841
rect 26939 3796 26952 3830
rect 26807 3758 26952 3796
rect 26911 3730 26952 3758
rect 25180 3698 25450 3726
rect 24921 3632 24931 3698
rect 24997 3632 25007 3698
rect 25180 3636 25214 3698
rect 25416 3636 25450 3698
rect 25534 3698 25805 3726
rect 26322 3702 26592 3730
rect 25534 3636 25568 3698
rect 25770 3636 25805 3698
rect 25946 3686 26117 3702
rect 25946 3652 26077 3686
rect 26111 3652 26117 3686
rect 25946 3636 26117 3652
rect 26322 3640 26356 3702
rect 26558 3640 26592 3702
rect 26676 3702 26952 3730
rect 26676 3640 26710 3702
rect 26912 3640 26952 3702
rect 25056 3624 25102 3636
rect 25056 3248 25062 3624
rect 25096 3248 25102 3624
rect 25056 3236 25102 3248
rect 25174 3624 25220 3636
rect 25174 3248 25180 3624
rect 25214 3248 25220 3624
rect 25174 3236 25220 3248
rect 25292 3624 25338 3636
rect 25292 3248 25298 3624
rect 25332 3248 25338 3624
rect 25292 3236 25338 3248
rect 25410 3624 25456 3636
rect 25410 3248 25416 3624
rect 25450 3248 25456 3624
rect 25410 3236 25456 3248
rect 25528 3624 25574 3636
rect 25528 3248 25534 3624
rect 25568 3248 25574 3624
rect 25528 3236 25574 3248
rect 25646 3624 25692 3636
rect 25646 3248 25652 3624
rect 25686 3248 25692 3624
rect 25646 3236 25692 3248
rect 25764 3624 25810 3636
rect 25764 3248 25770 3624
rect 25804 3248 25810 3624
rect 25764 3236 25810 3248
rect 23798 3131 24072 3159
rect 23444 3127 24072 3131
rect 22968 3115 23014 3127
rect 22968 2739 22974 3115
rect 23008 2739 23014 3115
rect 22968 2727 23014 2739
rect 23086 3115 23132 3127
rect 23086 2739 23092 3115
rect 23126 2739 23132 3115
rect 23086 2727 23132 2739
rect 23204 3115 23250 3127
rect 23204 2739 23210 3115
rect 23244 2763 23250 3115
rect 23321 3115 23367 3127
rect 23321 2939 23327 3115
rect 23361 2939 23367 3115
rect 23321 2927 23367 2939
rect 23439 3115 24072 3127
rect 23439 2939 23445 3115
rect 23479 3102 24072 3115
rect 25062 3194 25096 3236
rect 25298 3194 25332 3236
rect 25062 3166 25332 3194
rect 25416 3195 25450 3236
rect 25652 3195 25686 3236
rect 25416 3166 25686 3195
rect 25062 3118 25096 3166
rect 23479 2939 23485 3102
rect 25062 3088 25125 3118
rect 23439 2927 23485 2939
rect 25090 2996 25125 3088
rect 25090 2960 25317 2996
rect 25587 2985 25597 3082
rect 25696 2985 25706 3082
rect 25770 3053 25804 3236
rect 25770 2999 25879 3053
rect 23327 2811 23362 2927
rect 25090 2853 25125 2960
rect 25251 2926 25317 2960
rect 25251 2892 25267 2926
rect 25301 2892 25317 2926
rect 25598 2984 25695 2985
rect 25598 2917 25655 2984
rect 25251 2886 25317 2892
rect 25492 2881 25761 2917
rect 25492 2853 25525 2881
rect 25728 2853 25761 2881
rect 25845 2853 25879 2999
rect 24966 2841 25012 2853
rect 23458 2811 23566 2821
rect 23327 2763 23458 2811
rect 23566 2782 23714 2788
rect 23244 2739 23458 2763
rect 23204 2727 23458 2739
rect 23210 2723 23458 2727
rect 22086 2695 22846 2722
rect 22086 2689 23083 2695
rect 22086 2655 23033 2689
rect 23067 2655 23083 2689
rect 22086 2639 23083 2655
rect 23135 2689 23201 2695
rect 23135 2655 23151 2689
rect 23185 2655 23201 2689
rect 23384 2679 23458 2723
rect 23702 2715 23714 2782
rect 23566 2709 23714 2715
rect 23458 2669 23566 2679
rect 22086 2623 22846 2639
rect 22086 2622 22783 2623
rect 22086 2618 22318 2622
rect 20356 2589 20402 2601
rect 19489 2550 19523 2589
rect 19725 2550 19759 2589
rect 19489 2514 19759 2550
rect 20126 2551 20159 2589
rect 20362 2551 20395 2589
rect 20126 2515 20395 2551
rect 19489 2513 19655 2514
rect 19523 2434 19655 2513
rect 19513 2326 19523 2434
rect 19655 2326 19665 2434
rect 19549 2197 19555 2326
rect 19622 2197 19628 2326
rect 19549 2185 19628 2197
rect 21498 2207 22102 2235
rect 21498 2101 21950 2207
rect 22062 2194 22102 2207
rect 22062 2101 22104 2194
rect 21498 2090 22104 2101
rect 16127 1952 17104 1982
rect 19321 1980 19384 1997
rect 19246 1976 19384 1980
rect 16127 1846 16159 1952
rect 16363 1846 16395 1952
rect 16599 1846 16631 1952
rect 16835 1846 16867 1952
rect 17070 1846 17104 1952
rect 17414 1942 19384 1976
rect 17412 1913 19384 1942
rect 17412 1897 17458 1913
rect 19246 1911 19384 1913
rect 16120 1834 16166 1846
rect 16120 1658 16126 1834
rect 16160 1658 16166 1834
rect 16120 1646 16166 1658
rect 16238 1834 16284 1846
rect 16238 1658 16244 1834
rect 16278 1658 16284 1834
rect 16238 1646 16284 1658
rect 16356 1834 16402 1846
rect 16356 1658 16362 1834
rect 16396 1658 16402 1834
rect 16356 1646 16402 1658
rect 16474 1834 16520 1846
rect 16474 1658 16480 1834
rect 16514 1658 16520 1834
rect 16474 1646 16520 1658
rect 16592 1834 16638 1846
rect 16592 1658 16598 1834
rect 16632 1658 16638 1834
rect 16592 1646 16638 1658
rect 16710 1834 16756 1846
rect 16710 1658 16716 1834
rect 16750 1658 16756 1834
rect 16710 1646 16756 1658
rect 16828 1834 16874 1846
rect 16828 1658 16834 1834
rect 16868 1658 16874 1834
rect 16828 1646 16874 1658
rect 16946 1834 16992 1846
rect 16946 1658 16952 1834
rect 16986 1658 16992 1834
rect 16946 1646 16992 1658
rect 17064 1834 17110 1846
rect 17064 1658 17070 1834
rect 17104 1658 17110 1834
rect 17064 1646 17110 1658
rect 17182 1834 17228 1846
rect 17182 1658 17188 1834
rect 17222 1658 17228 1834
rect 17182 1646 17228 1658
rect 16243 1552 16279 1646
rect 16479 1552 16515 1646
rect 16715 1553 16751 1646
rect 16877 1598 16943 1605
rect 16877 1564 16893 1598
rect 16927 1564 16943 1598
rect 16877 1553 16943 1564
rect 16715 1552 16943 1553
rect 16243 1523 16943 1552
rect 16243 1522 16825 1523
rect 16363 1409 16397 1522
rect 16759 1481 16825 1522
rect 16759 1447 16775 1481
rect 16809 1447 16825 1481
rect 16759 1440 16825 1447
rect 17187 1428 17222 1646
rect 17411 1445 17458 1897
rect 20302 1901 20381 1913
rect 20302 1789 20308 1901
rect 20375 1789 20381 1901
rect 18370 1681 18380 1789
rect 18512 1681 18522 1789
rect 20268 1681 20278 1789
rect 20410 1681 20420 1789
rect 18380 1641 18512 1681
rect 20278 1641 20410 1681
rect 18379 1575 18512 1641
rect 20277 1575 20410 1641
rect 21498 1590 21648 2090
rect 21709 2089 22102 2090
rect 17708 1532 19181 1575
rect 17411 1429 17457 1445
rect 17376 1428 17457 1429
rect 17187 1413 17457 1428
rect 16833 1409 17457 1413
rect 16357 1397 16403 1409
rect 16092 919 16102 1037
rect 16220 1005 16230 1037
rect 16357 1021 16363 1397
rect 16397 1021 16403 1397
rect 16357 1009 16403 1021
rect 16475 1397 16521 1409
rect 16475 1021 16481 1397
rect 16515 1021 16521 1397
rect 16475 1009 16521 1021
rect 16593 1397 16639 1409
rect 16593 1021 16599 1397
rect 16633 1045 16639 1397
rect 16710 1397 16756 1409
rect 16710 1221 16716 1397
rect 16750 1221 16756 1397
rect 16710 1209 16756 1221
rect 16828 1397 17457 1409
rect 16828 1221 16834 1397
rect 16868 1385 17457 1397
rect 16868 1384 17110 1385
rect 16868 1221 16874 1384
rect 17376 1383 17457 1385
rect 17708 1229 17742 1532
rect 18074 1429 18108 1532
rect 18310 1429 18344 1532
rect 18546 1429 18580 1532
rect 18782 1429 18816 1532
rect 18068 1417 18114 1429
rect 16828 1209 16874 1221
rect 17584 1217 17630 1229
rect 16716 1093 16751 1209
rect 16847 1093 16955 1103
rect 16716 1045 16847 1093
rect 16955 1055 17099 1061
rect 16633 1021 16847 1045
rect 16593 1009 16847 1021
rect 16599 1005 16847 1009
rect 16220 977 16235 1005
rect 16220 971 16472 977
rect 16220 937 16422 971
rect 16456 937 16472 971
rect 16220 921 16472 937
rect 16524 971 16590 977
rect 16524 937 16540 971
rect 16574 937 16590 971
rect 16773 961 16847 1005
rect 17087 988 17099 1055
rect 17584 1041 17590 1217
rect 17624 1041 17630 1217
rect 17584 1029 17630 1041
rect 17702 1217 17748 1229
rect 17702 1041 17708 1217
rect 17742 1041 17748 1217
rect 17702 1029 17748 1041
rect 17820 1217 17866 1229
rect 17820 1041 17826 1217
rect 17860 1041 17866 1217
rect 17820 1029 17866 1041
rect 17938 1217 17984 1229
rect 18068 1217 18074 1417
rect 17938 1041 17944 1217
rect 17978 1041 18074 1217
rect 18108 1041 18114 1417
rect 17938 1029 17984 1041
rect 18068 1029 18114 1041
rect 18186 1417 18232 1429
rect 18186 1041 18192 1417
rect 18226 1041 18232 1417
rect 18186 1029 18232 1041
rect 18304 1417 18350 1429
rect 18304 1041 18310 1417
rect 18344 1041 18350 1417
rect 18304 1029 18350 1041
rect 18422 1417 18468 1429
rect 18422 1041 18428 1417
rect 18462 1041 18468 1417
rect 18422 1029 18468 1041
rect 18540 1417 18586 1429
rect 18540 1041 18546 1417
rect 18580 1041 18586 1417
rect 18540 1029 18586 1041
rect 18658 1417 18704 1429
rect 18658 1041 18664 1417
rect 18698 1041 18704 1417
rect 18658 1029 18704 1041
rect 18776 1417 18822 1429
rect 18776 1041 18782 1417
rect 18816 1217 18822 1417
rect 19147 1229 19181 1532
rect 19606 1532 21079 1575
rect 19606 1229 19640 1532
rect 19972 1429 20006 1532
rect 20208 1429 20242 1532
rect 20444 1429 20478 1532
rect 20680 1429 20714 1532
rect 19966 1417 20012 1429
rect 18905 1217 18951 1229
rect 18816 1041 18911 1217
rect 18945 1041 18951 1217
rect 18776 1029 18822 1041
rect 18905 1029 18951 1041
rect 19023 1217 19069 1229
rect 19023 1041 19029 1217
rect 19063 1041 19069 1217
rect 19023 1029 19069 1041
rect 19141 1217 19187 1229
rect 19141 1041 19147 1217
rect 19181 1041 19187 1217
rect 19141 1029 19187 1041
rect 19259 1217 19305 1229
rect 19259 1041 19265 1217
rect 19299 1041 19305 1217
rect 19259 1029 19305 1041
rect 19482 1217 19528 1229
rect 19482 1041 19488 1217
rect 19522 1041 19528 1217
rect 19482 1029 19528 1041
rect 19600 1217 19646 1229
rect 19600 1041 19606 1217
rect 19640 1041 19646 1217
rect 19600 1029 19646 1041
rect 19718 1217 19764 1229
rect 19718 1041 19724 1217
rect 19758 1041 19764 1217
rect 19718 1029 19764 1041
rect 19836 1217 19882 1229
rect 19966 1217 19972 1417
rect 19836 1041 19842 1217
rect 19876 1041 19972 1217
rect 20006 1041 20012 1417
rect 19836 1029 19882 1041
rect 19966 1029 20012 1041
rect 20084 1417 20130 1429
rect 20084 1041 20090 1417
rect 20124 1041 20130 1417
rect 20084 1029 20130 1041
rect 20202 1417 20248 1429
rect 20202 1041 20208 1417
rect 20242 1041 20248 1417
rect 20202 1029 20248 1041
rect 20320 1417 20366 1429
rect 20320 1041 20326 1417
rect 20360 1041 20366 1417
rect 20320 1029 20366 1041
rect 20438 1417 20484 1429
rect 20438 1041 20444 1417
rect 20478 1041 20484 1417
rect 20438 1029 20484 1041
rect 20556 1417 20602 1429
rect 20556 1041 20562 1417
rect 20596 1041 20602 1417
rect 20556 1029 20602 1041
rect 20674 1417 20720 1429
rect 20674 1041 20680 1417
rect 20714 1217 20720 1417
rect 21045 1229 21079 1532
rect 21497 1524 21648 1590
rect 20803 1217 20849 1229
rect 20714 1041 20809 1217
rect 20843 1041 20849 1217
rect 20674 1029 20720 1041
rect 20803 1029 20849 1041
rect 20921 1217 20967 1229
rect 20921 1041 20927 1217
rect 20961 1041 20967 1217
rect 20921 1029 20967 1041
rect 21039 1217 21085 1229
rect 21039 1041 21045 1217
rect 21079 1041 21085 1217
rect 21039 1029 21085 1041
rect 21157 1217 21203 1229
rect 21157 1041 21163 1217
rect 21197 1041 21203 1217
rect 21157 1029 21203 1041
rect 16955 982 17099 988
rect 17590 995 17624 1029
rect 18192 995 18226 1029
rect 18428 995 18462 1029
rect 16847 951 16955 961
rect 17590 960 17749 995
rect 18192 960 18462 995
rect 19029 995 19063 1029
rect 19265 995 19299 1029
rect 19029 960 19299 995
rect 19488 995 19522 1029
rect 20090 995 20124 1029
rect 20326 995 20360 1029
rect 19488 960 19647 995
rect 20090 960 20360 995
rect 20927 995 20961 1029
rect 21163 995 21197 1029
rect 20927 960 21197 995
rect 16220 919 16235 921
rect 16135 905 16235 919
rect 16135 862 16235 863
rect 15756 841 16235 862
rect 16524 841 16590 937
rect 15756 793 16590 841
rect 15756 764 16235 793
rect 15756 762 15861 764
rect 16135 763 16235 764
rect 15589 577 15599 656
rect 15692 577 15702 656
rect 16590 646 16669 658
rect 15600 -597 15693 577
rect 16590 548 16596 646
rect 16518 528 16596 548
rect 16663 548 16669 646
rect 16663 528 16738 548
rect 16518 420 16562 528
rect 16694 420 16738 528
rect 16518 378 16738 420
rect 16122 348 17099 378
rect 16122 242 16154 348
rect 16358 242 16390 348
rect 16594 242 16626 348
rect 16830 242 16862 348
rect 17065 242 17099 348
rect 16115 230 16161 242
rect 16115 54 16121 230
rect 16155 54 16161 230
rect 16115 42 16161 54
rect 16233 230 16279 242
rect 16233 54 16239 230
rect 16273 54 16279 230
rect 16233 42 16279 54
rect 16351 230 16397 242
rect 16351 54 16357 230
rect 16391 54 16397 230
rect 16351 42 16397 54
rect 16469 230 16515 242
rect 16469 54 16475 230
rect 16509 54 16515 230
rect 16469 42 16515 54
rect 16587 230 16633 242
rect 16587 54 16593 230
rect 16627 54 16633 230
rect 16587 42 16633 54
rect 16705 230 16751 242
rect 16705 54 16711 230
rect 16745 54 16751 230
rect 16705 42 16751 54
rect 16823 230 16869 242
rect 16823 54 16829 230
rect 16863 54 16869 230
rect 16823 42 16869 54
rect 16941 230 16987 242
rect 16941 54 16947 230
rect 16981 54 16987 230
rect 16941 42 16987 54
rect 17059 230 17105 242
rect 17059 54 17065 230
rect 17099 54 17105 230
rect 17059 42 17105 54
rect 17177 230 17223 242
rect 17177 54 17183 230
rect 17217 54 17223 230
rect 17177 42 17223 54
rect 17715 176 17749 960
rect 18428 898 18462 960
rect 18017 860 18759 898
rect 18017 736 18051 860
rect 18253 736 18287 860
rect 18489 736 18523 860
rect 18725 736 18759 860
rect 19015 753 19025 819
rect 19088 753 19098 819
rect 18011 724 18057 736
rect 18011 348 18017 724
rect 18051 348 18057 724
rect 18011 336 18057 348
rect 18129 724 18175 736
rect 18129 348 18135 724
rect 18169 348 18175 724
rect 18129 336 18175 348
rect 18247 724 18293 736
rect 18247 348 18253 724
rect 18287 348 18293 724
rect 18247 336 18293 348
rect 18365 724 18411 736
rect 18365 348 18371 724
rect 18405 348 18411 724
rect 18365 336 18411 348
rect 18483 724 18529 736
rect 18483 348 18489 724
rect 18523 348 18529 724
rect 18483 336 18529 348
rect 18601 724 18647 736
rect 18601 348 18607 724
rect 18641 348 18647 724
rect 18601 336 18647 348
rect 18719 724 18765 736
rect 18719 348 18725 724
rect 18759 348 18765 724
rect 18719 336 18765 348
rect 19131 177 19165 960
rect 18858 176 19165 177
rect 17715 171 18031 176
rect 18745 171 19165 176
rect 17715 160 18098 171
rect 17715 133 18047 160
rect 16238 -52 16274 42
rect 16474 -52 16510 42
rect 16710 -51 16746 42
rect 16872 -6 16938 1
rect 16872 -40 16888 -6
rect 16922 -40 16938 -6
rect 16872 -51 16938 -40
rect 16710 -52 16938 -51
rect 16238 -81 16938 -52
rect 16238 -82 16820 -81
rect 16358 -195 16392 -82
rect 16754 -123 16820 -82
rect 16754 -157 16770 -123
rect 16804 -157 16820 -123
rect 16754 -164 16820 -157
rect 17182 -191 17217 42
rect 17715 4 17749 133
rect 18031 126 18047 133
rect 18081 126 18098 160
rect 18031 120 18098 126
rect 18678 160 19165 171
rect 18678 126 18695 160
rect 18729 133 19165 160
rect 18729 126 18745 133
rect 18858 132 19165 133
rect 18678 120 18745 126
rect 17856 93 17912 105
rect 17856 59 17862 93
rect 17896 92 17912 93
rect 18969 92 19025 104
rect 17896 76 18363 92
rect 17896 59 18313 76
rect 17856 43 18313 59
rect 18297 42 18313 43
rect 18347 42 18363 76
rect 18297 35 18363 42
rect 18415 77 18985 92
rect 18415 43 18431 77
rect 18465 58 18985 77
rect 19019 58 19025 92
rect 18465 43 19025 58
rect 18415 33 18482 43
rect 18969 42 19025 43
rect 19131 4 19165 132
rect 19613 176 19647 960
rect 20326 898 20360 960
rect 19915 860 20657 898
rect 19915 736 19949 860
rect 20151 736 20185 860
rect 20387 736 20421 860
rect 20623 736 20657 860
rect 19909 724 19955 736
rect 19909 348 19915 724
rect 19949 348 19955 724
rect 19909 336 19955 348
rect 20027 724 20073 736
rect 20027 348 20033 724
rect 20067 348 20073 724
rect 20027 336 20073 348
rect 20145 724 20191 736
rect 20145 348 20151 724
rect 20185 348 20191 724
rect 20145 336 20191 348
rect 20263 724 20309 736
rect 20263 348 20269 724
rect 20303 348 20309 724
rect 20263 336 20309 348
rect 20381 724 20427 736
rect 20381 348 20387 724
rect 20421 348 20427 724
rect 20381 336 20427 348
rect 20499 724 20545 736
rect 20499 348 20505 724
rect 20539 348 20545 724
rect 20499 336 20545 348
rect 20617 724 20663 736
rect 20617 348 20623 724
rect 20657 348 20663 724
rect 20617 336 20663 348
rect 21029 177 21063 960
rect 20641 176 20710 177
rect 20756 176 21063 177
rect 19613 171 19929 176
rect 20641 172 21063 176
rect 19613 160 19996 171
rect 19613 133 19945 160
rect 19613 4 19647 133
rect 19929 126 19945 133
rect 19979 126 19996 160
rect 19929 120 19996 126
rect 20574 161 21063 172
rect 20574 127 20591 161
rect 20625 133 21063 161
rect 20625 127 20641 133
rect 20756 132 21063 133
rect 20574 121 20641 127
rect 19754 93 19810 105
rect 19754 59 19760 93
rect 19794 92 19810 93
rect 20867 92 20923 104
rect 19794 76 20261 92
rect 19794 59 20211 76
rect 19754 43 20211 59
rect 20195 42 20211 43
rect 20245 42 20261 76
rect 20195 35 20261 42
rect 20313 77 20883 92
rect 20313 43 20329 77
rect 20363 58 20883 77
rect 20917 58 20923 92
rect 20363 43 20923 58
rect 20313 33 20380 43
rect 20867 42 20923 43
rect 21029 4 21063 132
rect 21144 782 21211 806
rect 21144 748 21161 782
rect 21195 748 21211 782
rect 16828 -195 17217 -191
rect 16352 -207 16398 -195
rect 16352 -583 16358 -207
rect 16392 -583 16398 -207
rect 16352 -595 16398 -583
rect 16470 -207 16516 -195
rect 16470 -583 16476 -207
rect 16510 -583 16516 -207
rect 16470 -595 16516 -583
rect 16588 -207 16634 -195
rect 16588 -583 16594 -207
rect 16628 -559 16634 -207
rect 16705 -207 16751 -195
rect 16705 -383 16711 -207
rect 16745 -383 16751 -207
rect 16705 -395 16751 -383
rect 16823 -207 17217 -195
rect 17709 -8 17755 4
rect 17709 -184 17715 -8
rect 17749 -184 17755 -8
rect 17709 -196 17755 -184
rect 17827 -8 17873 4
rect 17827 -184 17833 -8
rect 17867 -184 17873 -8
rect 17827 -196 17873 -184
rect 18129 -8 18175 4
rect 16823 -383 16829 -207
rect 16863 -220 17217 -207
rect 16863 -383 16869 -220
rect 17139 -223 17217 -220
rect 17139 -275 17149 -223
rect 17212 -275 17222 -223
rect 17144 -281 17217 -275
rect 16823 -395 16869 -383
rect 16711 -511 16746 -395
rect 17832 -490 17866 -196
rect 18129 -384 18135 -8
rect 18169 -384 18175 -8
rect 18129 -396 18175 -384
rect 18247 -8 18293 4
rect 18247 -384 18253 -8
rect 18287 -384 18293 -8
rect 18247 -396 18293 -384
rect 18365 -8 18411 4
rect 18365 -384 18371 -8
rect 18405 -384 18411 -8
rect 18365 -396 18411 -384
rect 18483 -8 18529 4
rect 18483 -384 18489 -8
rect 18523 -384 18529 -8
rect 18483 -396 18529 -384
rect 18601 -8 18647 4
rect 18601 -384 18607 -8
rect 18641 -384 18647 -8
rect 19007 -8 19053 4
rect 19007 -184 19013 -8
rect 19047 -184 19053 -8
rect 19007 -196 19053 -184
rect 19125 -8 19171 4
rect 19125 -184 19131 -8
rect 19165 -184 19171 -8
rect 19125 -196 19171 -184
rect 19607 -8 19653 4
rect 19607 -184 19613 -8
rect 19647 -184 19653 -8
rect 19607 -196 19653 -184
rect 19725 -8 19771 4
rect 19725 -184 19731 -8
rect 19765 -184 19771 -8
rect 19725 -196 19771 -184
rect 20027 -8 20073 4
rect 18601 -396 18647 -384
rect 18489 -490 18523 -396
rect 19013 -490 19046 -196
rect 16842 -511 16950 -501
rect 16711 -559 16842 -511
rect 17832 -522 19046 -490
rect 19730 -490 19764 -196
rect 20027 -384 20033 -8
rect 20067 -384 20073 -8
rect 20027 -396 20073 -384
rect 20145 -8 20191 4
rect 20145 -384 20151 -8
rect 20185 -384 20191 -8
rect 20145 -396 20191 -384
rect 20263 -8 20309 4
rect 20263 -384 20269 -8
rect 20303 -384 20309 -8
rect 20263 -396 20309 -384
rect 20381 -8 20427 4
rect 20381 -384 20387 -8
rect 20421 -384 20427 -8
rect 20381 -396 20427 -384
rect 20499 -8 20545 4
rect 20499 -384 20505 -8
rect 20539 -384 20545 -8
rect 20905 -8 20951 4
rect 20905 -184 20911 -8
rect 20945 -184 20951 -8
rect 20905 -196 20951 -184
rect 21023 -8 21069 4
rect 21023 -184 21029 -8
rect 21063 -184 21069 -8
rect 21023 -196 21069 -184
rect 20499 -396 20545 -384
rect 20387 -490 20421 -396
rect 20911 -490 20944 -196
rect 19730 -522 20944 -490
rect 16950 -550 17101 -544
rect 16628 -583 16842 -559
rect 16588 -595 16842 -583
rect 15600 -599 16185 -597
rect 16594 -599 16842 -595
rect 15600 -627 16230 -599
rect 15600 -633 16467 -627
rect 15600 -667 16417 -633
rect 16451 -667 16467 -633
rect 15600 -683 16467 -667
rect 16519 -633 16585 -627
rect 16519 -667 16535 -633
rect 16569 -667 16585 -633
rect 16768 -643 16842 -599
rect 17089 -617 17101 -550
rect 18325 -607 18457 -522
rect 20223 -607 20355 -522
rect 16950 -623 17101 -617
rect 16842 -653 16950 -643
rect 15600 -699 16230 -683
rect 15600 -703 16185 -699
rect 15600 -704 15701 -703
rect 16130 -752 16230 -741
rect 16094 -858 16104 -752
rect 16216 -763 16230 -752
rect 16519 -763 16585 -667
rect 18315 -715 18325 -607
rect 18457 -715 18467 -607
rect 20213 -715 20223 -607
rect 20355 -715 20365 -607
rect 21144 -635 21211 748
rect 16216 -811 16585 -763
rect 16216 -841 16230 -811
rect 16216 -858 16226 -841
rect 16518 -914 16584 -811
rect 18343 -851 18349 -715
rect 18416 -851 18422 -715
rect 18343 -863 18422 -851
rect 21144 -914 21210 -635
rect 16516 -994 21210 -914
rect 15258 -1028 15421 -1014
rect 15258 -1096 15302 -1028
rect 15372 -1096 15421 -1028
rect 15258 -1815 15421 -1096
rect 21266 -1108 21276 -994
rect 21399 -1108 21409 -994
rect 15258 -1845 15422 -1815
rect 15258 -1913 15301 -1845
rect 15371 -1913 15422 -1845
rect 19057 -1846 19136 -1834
rect 15258 -1927 15422 -1913
rect 16572 -1906 16651 -1894
rect 16572 -1999 16578 -1906
rect 16504 -2019 16578 -1999
rect 16645 -1999 16651 -1906
rect 19057 -1965 19063 -1846
rect 19130 -1965 19136 -1846
rect 20206 -1849 20285 -1837
rect 20206 -1965 20212 -1849
rect 20279 -1965 20285 -1849
rect 16645 -2019 16724 -1999
rect 16504 -2127 16548 -2019
rect 16680 -2127 16724 -2019
rect 18301 -2061 18357 -2053
rect 16504 -2169 16724 -2127
rect 17375 -2069 18357 -2061
rect 17375 -2103 18317 -2069
rect 18351 -2103 18357 -2069
rect 19020 -2073 19030 -1965
rect 19162 -2028 19172 -1965
rect 19162 -2039 19174 -2028
rect 19162 -2073 19175 -2039
rect 19431 -2049 19487 -2047
rect 17375 -2119 18357 -2103
rect 19030 -2111 19175 -2073
rect 17375 -2120 18354 -2119
rect 16108 -2199 17085 -2169
rect 16108 -2305 16140 -2199
rect 16344 -2305 16376 -2199
rect 16580 -2305 16612 -2199
rect 16816 -2305 16848 -2199
rect 17051 -2305 17085 -2199
rect 16101 -2317 16147 -2305
rect 16101 -2493 16107 -2317
rect 16141 -2493 16147 -2317
rect 16101 -2505 16147 -2493
rect 16219 -2317 16265 -2305
rect 16219 -2493 16225 -2317
rect 16259 -2493 16265 -2317
rect 16219 -2505 16265 -2493
rect 16337 -2317 16383 -2305
rect 16337 -2493 16343 -2317
rect 16377 -2493 16383 -2317
rect 16337 -2505 16383 -2493
rect 16455 -2317 16501 -2305
rect 16455 -2493 16461 -2317
rect 16495 -2493 16501 -2317
rect 16455 -2505 16501 -2493
rect 16573 -2317 16619 -2305
rect 16573 -2493 16579 -2317
rect 16613 -2493 16619 -2317
rect 16573 -2505 16619 -2493
rect 16691 -2317 16737 -2305
rect 16691 -2493 16697 -2317
rect 16731 -2493 16737 -2317
rect 16691 -2505 16737 -2493
rect 16809 -2317 16855 -2305
rect 16809 -2493 16815 -2317
rect 16849 -2493 16855 -2317
rect 16809 -2505 16855 -2493
rect 16927 -2317 16973 -2305
rect 16927 -2493 16933 -2317
rect 16967 -2493 16973 -2317
rect 16927 -2505 16973 -2493
rect 17045 -2317 17091 -2305
rect 17045 -2493 17051 -2317
rect 17085 -2493 17091 -2317
rect 17045 -2505 17091 -2493
rect 17163 -2317 17209 -2305
rect 17163 -2493 17169 -2317
rect 17203 -2493 17209 -2317
rect 17163 -2505 17209 -2493
rect 16224 -2599 16260 -2505
rect 16460 -2599 16496 -2505
rect 16696 -2598 16732 -2505
rect 16858 -2553 16924 -2546
rect 16858 -2587 16874 -2553
rect 16908 -2587 16924 -2553
rect 16858 -2598 16924 -2587
rect 16696 -2599 16924 -2598
rect 16224 -2628 16924 -2599
rect 16224 -2629 16806 -2628
rect 16344 -2742 16378 -2629
rect 16740 -2670 16806 -2629
rect 16740 -2704 16756 -2670
rect 16790 -2704 16806 -2670
rect 16740 -2711 16806 -2704
rect 17168 -2710 17203 -2505
rect 17375 -2710 17442 -2120
rect 19134 -2143 19175 -2111
rect 19421 -2115 19431 -2049
rect 19487 -2115 19497 -2049
rect 20167 -2073 20177 -1965
rect 20309 -2028 20319 -1965
rect 20309 -2039 20321 -2028
rect 20309 -2073 20322 -2039
rect 20177 -2111 20322 -2073
rect 20281 -2139 20322 -2111
rect 18550 -2171 18820 -2143
rect 18291 -2237 18301 -2171
rect 18367 -2237 18377 -2171
rect 18550 -2233 18584 -2171
rect 18786 -2233 18820 -2171
rect 18904 -2171 19175 -2143
rect 19692 -2167 19962 -2139
rect 18904 -2233 18938 -2171
rect 19140 -2233 19175 -2171
rect 19316 -2183 19487 -2167
rect 19316 -2217 19447 -2183
rect 19481 -2217 19487 -2183
rect 19316 -2233 19487 -2217
rect 19692 -2229 19726 -2167
rect 19928 -2229 19962 -2167
rect 20046 -2167 20322 -2139
rect 20046 -2229 20080 -2167
rect 20282 -2229 20322 -2167
rect 18426 -2245 18472 -2233
rect 18426 -2621 18432 -2245
rect 18466 -2621 18472 -2245
rect 18426 -2633 18472 -2621
rect 18544 -2245 18590 -2233
rect 18544 -2621 18550 -2245
rect 18584 -2621 18590 -2245
rect 18544 -2633 18590 -2621
rect 18662 -2245 18708 -2233
rect 18662 -2621 18668 -2245
rect 18702 -2621 18708 -2245
rect 18662 -2633 18708 -2621
rect 18780 -2245 18826 -2233
rect 18780 -2621 18786 -2245
rect 18820 -2621 18826 -2245
rect 18780 -2633 18826 -2621
rect 18898 -2245 18944 -2233
rect 18898 -2621 18904 -2245
rect 18938 -2621 18944 -2245
rect 18898 -2633 18944 -2621
rect 19016 -2245 19062 -2233
rect 19016 -2621 19022 -2245
rect 19056 -2621 19062 -2245
rect 19016 -2633 19062 -2621
rect 19134 -2245 19180 -2233
rect 19134 -2621 19140 -2245
rect 19174 -2621 19180 -2245
rect 19134 -2633 19180 -2621
rect 17168 -2738 17442 -2710
rect 16814 -2742 17442 -2738
rect 16338 -2754 16384 -2742
rect 16338 -3130 16344 -2754
rect 16378 -3130 16384 -2754
rect 16338 -3142 16384 -3130
rect 16456 -2754 16502 -2742
rect 16456 -3130 16462 -2754
rect 16496 -3130 16502 -2754
rect 16456 -3142 16502 -3130
rect 16574 -2754 16620 -2742
rect 16574 -3130 16580 -2754
rect 16614 -3106 16620 -2754
rect 16691 -2754 16737 -2742
rect 16691 -2930 16697 -2754
rect 16731 -2930 16737 -2754
rect 16691 -2942 16737 -2930
rect 16809 -2754 17442 -2742
rect 16809 -2930 16815 -2754
rect 16849 -2767 17442 -2754
rect 18432 -2675 18466 -2633
rect 18668 -2675 18702 -2633
rect 18432 -2703 18702 -2675
rect 18786 -2674 18820 -2633
rect 19022 -2674 19056 -2633
rect 18786 -2703 19056 -2674
rect 18432 -2751 18466 -2703
rect 16849 -2930 16855 -2767
rect 18432 -2781 18495 -2751
rect 16809 -2942 16855 -2930
rect 18460 -2873 18495 -2781
rect 18460 -2909 18687 -2873
rect 18957 -2884 18967 -2787
rect 19066 -2884 19076 -2787
rect 19140 -2816 19174 -2633
rect 19140 -2870 19249 -2816
rect 16697 -3058 16732 -2942
rect 18460 -3016 18495 -2909
rect 18621 -2943 18687 -2909
rect 18621 -2977 18637 -2943
rect 18671 -2977 18687 -2943
rect 18968 -2885 19065 -2884
rect 18968 -2952 19025 -2885
rect 18621 -2983 18687 -2977
rect 18862 -2988 19131 -2952
rect 18862 -3016 18895 -2988
rect 19098 -3016 19131 -2988
rect 19215 -3016 19249 -2870
rect 18336 -3028 18382 -3016
rect 16828 -3058 16936 -3048
rect 16697 -3106 16828 -3058
rect 16936 -3094 17087 -3088
rect 16614 -3130 16828 -3106
rect 16574 -3142 16828 -3130
rect 16580 -3146 16828 -3142
rect 14891 -3147 15514 -3146
rect 14891 -3174 16216 -3147
rect 14891 -3180 16453 -3174
rect 12829 -3252 12863 -3213
rect 13065 -3252 13099 -3213
rect 12829 -3288 13099 -3252
rect 13466 -3251 13499 -3213
rect 13702 -3251 13735 -3213
rect 13466 -3287 13735 -3251
rect 14891 -3214 16403 -3180
rect 16437 -3214 16453 -3180
rect 14891 -3230 16453 -3214
rect 16505 -3180 16571 -3174
rect 16505 -3214 16521 -3180
rect 16555 -3214 16571 -3180
rect 16754 -3190 16828 -3146
rect 17075 -3161 17087 -3094
rect 16936 -3167 17087 -3161
rect 16828 -3200 16936 -3190
rect 14891 -3246 16216 -3230
rect 14891 -3247 16153 -3246
rect 14891 -3251 15688 -3247
rect 14891 -3252 15514 -3251
rect 12829 -3289 12995 -3288
rect 12863 -3368 12995 -3289
rect 12853 -3476 12863 -3368
rect 12995 -3476 13005 -3368
rect 12885 -3621 12891 -3476
rect 12958 -3621 12964 -3476
rect 12885 -3633 12964 -3621
rect 14892 -3639 15473 -3631
rect 14891 -3657 15473 -3639
rect 14891 -3770 15253 -3657
rect 15457 -3675 15473 -3657
rect 14891 -3771 15405 -3770
rect 15457 -3771 15474 -3675
rect 14891 -3781 15474 -3771
rect 9467 -3850 10444 -3820
rect 12661 -3822 12724 -3805
rect 12586 -3826 12724 -3822
rect 9467 -3956 9499 -3850
rect 9703 -3956 9735 -3850
rect 9939 -3956 9971 -3850
rect 10175 -3956 10207 -3850
rect 10410 -3956 10444 -3850
rect 10754 -3860 12724 -3826
rect 10752 -3889 12724 -3860
rect 10752 -3905 10798 -3889
rect 12586 -3891 12724 -3889
rect 9460 -3968 9506 -3956
rect 9460 -4144 9466 -3968
rect 9500 -4144 9506 -3968
rect 9460 -4156 9506 -4144
rect 9578 -3968 9624 -3956
rect 9578 -4144 9584 -3968
rect 9618 -4144 9624 -3968
rect 9578 -4156 9624 -4144
rect 9696 -3968 9742 -3956
rect 9696 -4144 9702 -3968
rect 9736 -4144 9742 -3968
rect 9696 -4156 9742 -4144
rect 9814 -3968 9860 -3956
rect 9814 -4144 9820 -3968
rect 9854 -4144 9860 -3968
rect 9814 -4156 9860 -4144
rect 9932 -3968 9978 -3956
rect 9932 -4144 9938 -3968
rect 9972 -4144 9978 -3968
rect 9932 -4156 9978 -4144
rect 10050 -3968 10096 -3956
rect 10050 -4144 10056 -3968
rect 10090 -4144 10096 -3968
rect 10050 -4156 10096 -4144
rect 10168 -3968 10214 -3956
rect 10168 -4144 10174 -3968
rect 10208 -4144 10214 -3968
rect 10168 -4156 10214 -4144
rect 10286 -3968 10332 -3956
rect 10286 -4144 10292 -3968
rect 10326 -4144 10332 -3968
rect 10286 -4156 10332 -4144
rect 10404 -3968 10450 -3956
rect 10404 -4144 10410 -3968
rect 10444 -4144 10450 -3968
rect 10404 -4156 10450 -4144
rect 10522 -3968 10568 -3956
rect 10522 -4144 10528 -3968
rect 10562 -4144 10568 -3968
rect 10522 -4156 10568 -4144
rect 9583 -4250 9619 -4156
rect 9819 -4250 9855 -4156
rect 10055 -4249 10091 -4156
rect 10217 -4204 10283 -4197
rect 10217 -4238 10233 -4204
rect 10267 -4238 10283 -4204
rect 10217 -4249 10283 -4238
rect 10055 -4250 10283 -4249
rect 9583 -4279 10283 -4250
rect 9583 -4280 10165 -4279
rect 9703 -4393 9737 -4280
rect 10099 -4321 10165 -4280
rect 10099 -4355 10115 -4321
rect 10149 -4355 10165 -4321
rect 10099 -4362 10165 -4355
rect 10527 -4374 10562 -4156
rect 10751 -4357 10798 -3905
rect 13649 -3896 13728 -3884
rect 13649 -4013 13655 -3896
rect 13722 -4013 13728 -3896
rect 11710 -4121 11720 -4013
rect 11852 -4121 11862 -4013
rect 13608 -4121 13618 -4013
rect 13750 -4121 13760 -4013
rect 11720 -4161 11852 -4121
rect 13618 -4161 13750 -4121
rect 11719 -4227 11852 -4161
rect 13617 -4227 13750 -4161
rect 11048 -4270 12521 -4227
rect 10751 -4373 10797 -4357
rect 10716 -4374 10797 -4373
rect 10527 -4389 10797 -4374
rect 10173 -4393 10797 -4389
rect 9697 -4405 9743 -4393
rect 9432 -4883 9442 -4765
rect 9560 -4797 9570 -4765
rect 9697 -4781 9703 -4405
rect 9737 -4781 9743 -4405
rect 9697 -4793 9743 -4781
rect 9815 -4405 9861 -4393
rect 9815 -4781 9821 -4405
rect 9855 -4781 9861 -4405
rect 9815 -4793 9861 -4781
rect 9933 -4405 9979 -4393
rect 9933 -4781 9939 -4405
rect 9973 -4757 9979 -4405
rect 10050 -4405 10096 -4393
rect 10050 -4581 10056 -4405
rect 10090 -4581 10096 -4405
rect 10050 -4593 10096 -4581
rect 10168 -4405 10797 -4393
rect 10168 -4581 10174 -4405
rect 10208 -4417 10797 -4405
rect 10208 -4418 10450 -4417
rect 10208 -4581 10214 -4418
rect 10716 -4419 10797 -4417
rect 11048 -4573 11082 -4270
rect 11414 -4373 11448 -4270
rect 11650 -4373 11684 -4270
rect 11886 -4373 11920 -4270
rect 12122 -4373 12156 -4270
rect 11408 -4385 11454 -4373
rect 10168 -4593 10214 -4581
rect 10924 -4585 10970 -4573
rect 10056 -4709 10091 -4593
rect 10187 -4709 10295 -4699
rect 10056 -4757 10187 -4709
rect 10295 -4748 10442 -4742
rect 9973 -4781 10187 -4757
rect 9933 -4793 10187 -4781
rect 9939 -4797 10187 -4793
rect 9560 -4825 9575 -4797
rect 9560 -4831 9812 -4825
rect 9560 -4865 9762 -4831
rect 9796 -4865 9812 -4831
rect 9560 -4881 9812 -4865
rect 9864 -4831 9930 -4825
rect 9864 -4865 9880 -4831
rect 9914 -4865 9930 -4831
rect 10113 -4841 10187 -4797
rect 10430 -4815 10442 -4748
rect 10924 -4761 10930 -4585
rect 10964 -4761 10970 -4585
rect 10924 -4773 10970 -4761
rect 11042 -4585 11088 -4573
rect 11042 -4761 11048 -4585
rect 11082 -4761 11088 -4585
rect 11042 -4773 11088 -4761
rect 11160 -4585 11206 -4573
rect 11160 -4761 11166 -4585
rect 11200 -4761 11206 -4585
rect 11160 -4773 11206 -4761
rect 11278 -4585 11324 -4573
rect 11408 -4585 11414 -4385
rect 11278 -4761 11284 -4585
rect 11318 -4761 11414 -4585
rect 11448 -4761 11454 -4385
rect 11278 -4773 11324 -4761
rect 11408 -4773 11454 -4761
rect 11526 -4385 11572 -4373
rect 11526 -4761 11532 -4385
rect 11566 -4761 11572 -4385
rect 11526 -4773 11572 -4761
rect 11644 -4385 11690 -4373
rect 11644 -4761 11650 -4385
rect 11684 -4761 11690 -4385
rect 11644 -4773 11690 -4761
rect 11762 -4385 11808 -4373
rect 11762 -4761 11768 -4385
rect 11802 -4761 11808 -4385
rect 11762 -4773 11808 -4761
rect 11880 -4385 11926 -4373
rect 11880 -4761 11886 -4385
rect 11920 -4761 11926 -4385
rect 11880 -4773 11926 -4761
rect 11998 -4385 12044 -4373
rect 11998 -4761 12004 -4385
rect 12038 -4761 12044 -4385
rect 11998 -4773 12044 -4761
rect 12116 -4385 12162 -4373
rect 12116 -4761 12122 -4385
rect 12156 -4585 12162 -4385
rect 12487 -4573 12521 -4270
rect 12946 -4270 14419 -4227
rect 12946 -4573 12980 -4270
rect 13312 -4373 13346 -4270
rect 13548 -4373 13582 -4270
rect 13784 -4373 13818 -4270
rect 14020 -4373 14054 -4270
rect 13306 -4385 13352 -4373
rect 12245 -4585 12291 -4573
rect 12156 -4761 12251 -4585
rect 12285 -4761 12291 -4585
rect 12116 -4773 12162 -4761
rect 12245 -4773 12291 -4761
rect 12363 -4585 12409 -4573
rect 12363 -4761 12369 -4585
rect 12403 -4761 12409 -4585
rect 12363 -4773 12409 -4761
rect 12481 -4585 12527 -4573
rect 12481 -4761 12487 -4585
rect 12521 -4761 12527 -4585
rect 12481 -4773 12527 -4761
rect 12599 -4585 12645 -4573
rect 12599 -4761 12605 -4585
rect 12639 -4761 12645 -4585
rect 12599 -4773 12645 -4761
rect 12822 -4585 12868 -4573
rect 12822 -4761 12828 -4585
rect 12862 -4761 12868 -4585
rect 12822 -4773 12868 -4761
rect 12940 -4585 12986 -4573
rect 12940 -4761 12946 -4585
rect 12980 -4761 12986 -4585
rect 12940 -4773 12986 -4761
rect 13058 -4585 13104 -4573
rect 13058 -4761 13064 -4585
rect 13098 -4761 13104 -4585
rect 13058 -4773 13104 -4761
rect 13176 -4585 13222 -4573
rect 13306 -4585 13312 -4385
rect 13176 -4761 13182 -4585
rect 13216 -4761 13312 -4585
rect 13346 -4761 13352 -4385
rect 13176 -4773 13222 -4761
rect 13306 -4773 13352 -4761
rect 13424 -4385 13470 -4373
rect 13424 -4761 13430 -4385
rect 13464 -4761 13470 -4385
rect 13424 -4773 13470 -4761
rect 13542 -4385 13588 -4373
rect 13542 -4761 13548 -4385
rect 13582 -4761 13588 -4385
rect 13542 -4773 13588 -4761
rect 13660 -4385 13706 -4373
rect 13660 -4761 13666 -4385
rect 13700 -4761 13706 -4385
rect 13660 -4773 13706 -4761
rect 13778 -4385 13824 -4373
rect 13778 -4761 13784 -4385
rect 13818 -4761 13824 -4385
rect 13778 -4773 13824 -4761
rect 13896 -4385 13942 -4373
rect 13896 -4761 13902 -4385
rect 13936 -4761 13942 -4385
rect 13896 -4773 13942 -4761
rect 14014 -4385 14060 -4373
rect 14014 -4761 14020 -4385
rect 14054 -4585 14060 -4385
rect 14385 -4573 14419 -4270
rect 14143 -4585 14189 -4573
rect 14054 -4761 14149 -4585
rect 14183 -4761 14189 -4585
rect 14014 -4773 14060 -4761
rect 14143 -4773 14189 -4761
rect 14261 -4585 14307 -4573
rect 14261 -4761 14267 -4585
rect 14301 -4761 14307 -4585
rect 14261 -4773 14307 -4761
rect 14379 -4585 14425 -4573
rect 14379 -4761 14385 -4585
rect 14419 -4761 14425 -4585
rect 14379 -4773 14425 -4761
rect 14497 -4585 14543 -4573
rect 14497 -4761 14503 -4585
rect 14537 -4761 14543 -4585
rect 14497 -4773 14543 -4761
rect 10295 -4821 10442 -4815
rect 10930 -4807 10964 -4773
rect 11532 -4807 11566 -4773
rect 11768 -4807 11802 -4773
rect 10187 -4851 10295 -4841
rect 10930 -4842 11089 -4807
rect 11532 -4842 11802 -4807
rect 12369 -4807 12403 -4773
rect 12605 -4807 12639 -4773
rect 12369 -4842 12639 -4807
rect 12828 -4807 12862 -4773
rect 13430 -4807 13464 -4773
rect 13666 -4807 13700 -4773
rect 12828 -4842 12987 -4807
rect 13430 -4842 13700 -4807
rect 14267 -4807 14301 -4773
rect 14503 -4807 14537 -4773
rect 14267 -4842 14537 -4807
rect 9560 -4883 9575 -4881
rect 9475 -4897 9575 -4883
rect 9475 -4940 9575 -4939
rect 9096 -4961 9575 -4940
rect 9864 -4961 9930 -4865
rect 9096 -5009 9930 -4961
rect 9096 -5038 9575 -5009
rect 9096 -5040 9201 -5038
rect 9475 -5039 9575 -5038
rect 8929 -5225 8939 -5146
rect 9032 -5225 9042 -5146
rect 9932 -5158 10011 -5146
rect 8940 -6399 9033 -5225
rect 9932 -5254 9938 -5158
rect 9858 -5274 9938 -5254
rect 10005 -5254 10011 -5158
rect 10005 -5274 10078 -5254
rect 9858 -5382 9902 -5274
rect 10034 -5382 10078 -5274
rect 9858 -5424 10078 -5382
rect 9462 -5454 10439 -5424
rect 9462 -5560 9494 -5454
rect 9698 -5560 9730 -5454
rect 9934 -5560 9966 -5454
rect 10170 -5560 10202 -5454
rect 10405 -5560 10439 -5454
rect 9455 -5572 9501 -5560
rect 9455 -5748 9461 -5572
rect 9495 -5748 9501 -5572
rect 9455 -5760 9501 -5748
rect 9573 -5572 9619 -5560
rect 9573 -5748 9579 -5572
rect 9613 -5748 9619 -5572
rect 9573 -5760 9619 -5748
rect 9691 -5572 9737 -5560
rect 9691 -5748 9697 -5572
rect 9731 -5748 9737 -5572
rect 9691 -5760 9737 -5748
rect 9809 -5572 9855 -5560
rect 9809 -5748 9815 -5572
rect 9849 -5748 9855 -5572
rect 9809 -5760 9855 -5748
rect 9927 -5572 9973 -5560
rect 9927 -5748 9933 -5572
rect 9967 -5748 9973 -5572
rect 9927 -5760 9973 -5748
rect 10045 -5572 10091 -5560
rect 10045 -5748 10051 -5572
rect 10085 -5748 10091 -5572
rect 10045 -5760 10091 -5748
rect 10163 -5572 10209 -5560
rect 10163 -5748 10169 -5572
rect 10203 -5748 10209 -5572
rect 10163 -5760 10209 -5748
rect 10281 -5572 10327 -5560
rect 10281 -5748 10287 -5572
rect 10321 -5748 10327 -5572
rect 10281 -5760 10327 -5748
rect 10399 -5572 10445 -5560
rect 10399 -5748 10405 -5572
rect 10439 -5748 10445 -5572
rect 10399 -5760 10445 -5748
rect 10517 -5572 10563 -5560
rect 10517 -5748 10523 -5572
rect 10557 -5748 10563 -5572
rect 10517 -5760 10563 -5748
rect 11055 -5626 11089 -4842
rect 11768 -4904 11802 -4842
rect 11357 -4942 12099 -4904
rect 11357 -5066 11391 -4942
rect 11593 -5066 11627 -4942
rect 11829 -5066 11863 -4942
rect 12065 -5066 12099 -4942
rect 12355 -5049 12365 -4983
rect 12428 -5049 12438 -4983
rect 11351 -5078 11397 -5066
rect 11351 -5454 11357 -5078
rect 11391 -5454 11397 -5078
rect 11351 -5466 11397 -5454
rect 11469 -5078 11515 -5066
rect 11469 -5454 11475 -5078
rect 11509 -5454 11515 -5078
rect 11469 -5466 11515 -5454
rect 11587 -5078 11633 -5066
rect 11587 -5454 11593 -5078
rect 11627 -5454 11633 -5078
rect 11587 -5466 11633 -5454
rect 11705 -5078 11751 -5066
rect 11705 -5454 11711 -5078
rect 11745 -5454 11751 -5078
rect 11705 -5466 11751 -5454
rect 11823 -5078 11869 -5066
rect 11823 -5454 11829 -5078
rect 11863 -5454 11869 -5078
rect 11823 -5466 11869 -5454
rect 11941 -5078 11987 -5066
rect 11941 -5454 11947 -5078
rect 11981 -5454 11987 -5078
rect 11941 -5466 11987 -5454
rect 12059 -5078 12105 -5066
rect 12059 -5454 12065 -5078
rect 12099 -5454 12105 -5078
rect 12059 -5466 12105 -5454
rect 12471 -5625 12505 -4842
rect 12198 -5626 12505 -5625
rect 11055 -5631 11371 -5626
rect 12085 -5631 12505 -5626
rect 11055 -5642 11438 -5631
rect 11055 -5669 11387 -5642
rect 9578 -5854 9614 -5760
rect 9814 -5854 9850 -5760
rect 10050 -5853 10086 -5760
rect 10212 -5808 10278 -5801
rect 10212 -5842 10228 -5808
rect 10262 -5842 10278 -5808
rect 10212 -5853 10278 -5842
rect 10050 -5854 10278 -5853
rect 9578 -5883 10278 -5854
rect 9578 -5884 10160 -5883
rect 9698 -5997 9732 -5884
rect 10094 -5925 10160 -5884
rect 10094 -5959 10110 -5925
rect 10144 -5959 10160 -5925
rect 10094 -5966 10160 -5959
rect 10522 -5993 10557 -5760
rect 11055 -5798 11089 -5669
rect 11371 -5676 11387 -5669
rect 11421 -5676 11438 -5642
rect 11371 -5682 11438 -5676
rect 12018 -5642 12505 -5631
rect 12018 -5676 12035 -5642
rect 12069 -5669 12505 -5642
rect 12069 -5676 12085 -5669
rect 12198 -5670 12505 -5669
rect 12018 -5682 12085 -5676
rect 11196 -5709 11252 -5697
rect 11196 -5743 11202 -5709
rect 11236 -5710 11252 -5709
rect 12309 -5710 12365 -5698
rect 11236 -5726 11703 -5710
rect 11236 -5743 11653 -5726
rect 11196 -5759 11653 -5743
rect 11637 -5760 11653 -5759
rect 11687 -5760 11703 -5726
rect 11637 -5767 11703 -5760
rect 11755 -5725 12325 -5710
rect 11755 -5759 11771 -5725
rect 11805 -5744 12325 -5725
rect 12359 -5744 12365 -5710
rect 11805 -5759 12365 -5744
rect 11755 -5769 11822 -5759
rect 12309 -5760 12365 -5759
rect 12471 -5798 12505 -5670
rect 12953 -5626 12987 -4842
rect 13666 -4904 13700 -4842
rect 13255 -4942 13997 -4904
rect 13255 -5066 13289 -4942
rect 13491 -5066 13525 -4942
rect 13727 -5066 13761 -4942
rect 13963 -5066 13997 -4942
rect 13249 -5078 13295 -5066
rect 13249 -5454 13255 -5078
rect 13289 -5454 13295 -5078
rect 13249 -5466 13295 -5454
rect 13367 -5078 13413 -5066
rect 13367 -5454 13373 -5078
rect 13407 -5454 13413 -5078
rect 13367 -5466 13413 -5454
rect 13485 -5078 13531 -5066
rect 13485 -5454 13491 -5078
rect 13525 -5454 13531 -5078
rect 13485 -5466 13531 -5454
rect 13603 -5078 13649 -5066
rect 13603 -5454 13609 -5078
rect 13643 -5454 13649 -5078
rect 13603 -5466 13649 -5454
rect 13721 -5078 13767 -5066
rect 13721 -5454 13727 -5078
rect 13761 -5454 13767 -5078
rect 13721 -5466 13767 -5454
rect 13839 -5078 13885 -5066
rect 13839 -5454 13845 -5078
rect 13879 -5454 13885 -5078
rect 13839 -5466 13885 -5454
rect 13957 -5078 14003 -5066
rect 13957 -5454 13963 -5078
rect 13997 -5454 14003 -5078
rect 13957 -5466 14003 -5454
rect 14369 -5625 14403 -4842
rect 13981 -5626 14050 -5625
rect 14096 -5626 14403 -5625
rect 12953 -5631 13269 -5626
rect 13981 -5630 14403 -5626
rect 12953 -5642 13336 -5631
rect 12953 -5669 13285 -5642
rect 12953 -5798 12987 -5669
rect 13269 -5676 13285 -5669
rect 13319 -5676 13336 -5642
rect 13269 -5682 13336 -5676
rect 13914 -5641 14403 -5630
rect 13914 -5675 13931 -5641
rect 13965 -5669 14403 -5641
rect 13965 -5675 13981 -5669
rect 14096 -5670 14403 -5669
rect 13914 -5681 13981 -5675
rect 13094 -5709 13150 -5697
rect 13094 -5743 13100 -5709
rect 13134 -5710 13150 -5709
rect 14207 -5710 14263 -5698
rect 13134 -5726 13601 -5710
rect 13134 -5743 13551 -5726
rect 13094 -5759 13551 -5743
rect 13535 -5760 13551 -5759
rect 13585 -5760 13601 -5726
rect 13535 -5767 13601 -5760
rect 13653 -5725 14223 -5710
rect 13653 -5759 13669 -5725
rect 13703 -5744 14223 -5725
rect 14257 -5744 14263 -5710
rect 13703 -5759 14263 -5744
rect 13653 -5769 13720 -5759
rect 14207 -5760 14263 -5759
rect 14369 -5798 14403 -5670
rect 14484 -5020 14551 -4996
rect 14484 -5054 14501 -5020
rect 14535 -5054 14551 -5020
rect 10168 -5997 10557 -5993
rect 9692 -6009 9738 -5997
rect 9692 -6385 9698 -6009
rect 9732 -6385 9738 -6009
rect 9692 -6397 9738 -6385
rect 9810 -6009 9856 -5997
rect 9810 -6385 9816 -6009
rect 9850 -6385 9856 -6009
rect 9810 -6397 9856 -6385
rect 9928 -6009 9974 -5997
rect 9928 -6385 9934 -6009
rect 9968 -6361 9974 -6009
rect 10045 -6009 10091 -5997
rect 10045 -6185 10051 -6009
rect 10085 -6185 10091 -6009
rect 10045 -6197 10091 -6185
rect 10163 -6009 10557 -5997
rect 11049 -5810 11095 -5798
rect 11049 -5986 11055 -5810
rect 11089 -5986 11095 -5810
rect 11049 -5998 11095 -5986
rect 11167 -5810 11213 -5798
rect 11167 -5986 11173 -5810
rect 11207 -5986 11213 -5810
rect 11167 -5998 11213 -5986
rect 11469 -5810 11515 -5798
rect 10163 -6185 10169 -6009
rect 10203 -6022 10557 -6009
rect 10203 -6185 10209 -6022
rect 10479 -6025 10557 -6022
rect 10479 -6077 10489 -6025
rect 10552 -6077 10562 -6025
rect 10484 -6083 10557 -6077
rect 10163 -6197 10209 -6185
rect 10051 -6313 10086 -6197
rect 11172 -6292 11206 -5998
rect 11469 -6186 11475 -5810
rect 11509 -6186 11515 -5810
rect 11469 -6198 11515 -6186
rect 11587 -5810 11633 -5798
rect 11587 -6186 11593 -5810
rect 11627 -6186 11633 -5810
rect 11587 -6198 11633 -6186
rect 11705 -5810 11751 -5798
rect 11705 -6186 11711 -5810
rect 11745 -6186 11751 -5810
rect 11705 -6198 11751 -6186
rect 11823 -5810 11869 -5798
rect 11823 -6186 11829 -5810
rect 11863 -6186 11869 -5810
rect 11823 -6198 11869 -6186
rect 11941 -5810 11987 -5798
rect 11941 -6186 11947 -5810
rect 11981 -6186 11987 -5810
rect 12347 -5810 12393 -5798
rect 12347 -5986 12353 -5810
rect 12387 -5986 12393 -5810
rect 12347 -5998 12393 -5986
rect 12465 -5810 12511 -5798
rect 12465 -5986 12471 -5810
rect 12505 -5986 12511 -5810
rect 12465 -5998 12511 -5986
rect 12947 -5810 12993 -5798
rect 12947 -5986 12953 -5810
rect 12987 -5986 12993 -5810
rect 12947 -5998 12993 -5986
rect 13065 -5810 13111 -5798
rect 13065 -5986 13071 -5810
rect 13105 -5986 13111 -5810
rect 13065 -5998 13111 -5986
rect 13367 -5810 13413 -5798
rect 11941 -6198 11987 -6186
rect 11829 -6292 11863 -6198
rect 12353 -6292 12386 -5998
rect 10182 -6313 10290 -6303
rect 10051 -6361 10182 -6313
rect 11172 -6324 12386 -6292
rect 13070 -6292 13104 -5998
rect 13367 -6186 13373 -5810
rect 13407 -6186 13413 -5810
rect 13367 -6198 13413 -6186
rect 13485 -5810 13531 -5798
rect 13485 -6186 13491 -5810
rect 13525 -6186 13531 -5810
rect 13485 -6198 13531 -6186
rect 13603 -5810 13649 -5798
rect 13603 -6186 13609 -5810
rect 13643 -6186 13649 -5810
rect 13603 -6198 13649 -6186
rect 13721 -5810 13767 -5798
rect 13721 -6186 13727 -5810
rect 13761 -6186 13767 -5810
rect 13721 -6198 13767 -6186
rect 13839 -5810 13885 -5798
rect 13839 -6186 13845 -5810
rect 13879 -6186 13885 -5810
rect 14245 -5810 14291 -5798
rect 14245 -5986 14251 -5810
rect 14285 -5986 14291 -5810
rect 14245 -5998 14291 -5986
rect 14363 -5810 14409 -5798
rect 14363 -5986 14369 -5810
rect 14403 -5986 14409 -5810
rect 14363 -5998 14409 -5986
rect 13839 -6198 13885 -6186
rect 13727 -6292 13761 -6198
rect 14251 -6292 14284 -5998
rect 13070 -6324 14284 -6292
rect 10290 -6348 10431 -6342
rect 9968 -6385 10182 -6361
rect 9928 -6397 10182 -6385
rect 8940 -6401 9525 -6399
rect 9934 -6401 10182 -6397
rect 8940 -6429 9570 -6401
rect 8940 -6435 9807 -6429
rect 8940 -6469 9757 -6435
rect 9791 -6469 9807 -6435
rect 8940 -6485 9807 -6469
rect 9859 -6435 9925 -6429
rect 9859 -6469 9875 -6435
rect 9909 -6469 9925 -6435
rect 10108 -6445 10182 -6401
rect 10419 -6415 10431 -6348
rect 11665 -6409 11797 -6324
rect 13563 -6409 13695 -6324
rect 10290 -6421 10431 -6415
rect 10182 -6455 10290 -6445
rect 8940 -6501 9570 -6485
rect 8940 -6505 9525 -6501
rect 8940 -6506 9041 -6505
rect 9470 -6554 9570 -6543
rect 9434 -6660 9444 -6554
rect 9556 -6565 9570 -6554
rect 9859 -6565 9925 -6469
rect 11655 -6517 11665 -6409
rect 11797 -6517 11807 -6409
rect 13553 -6517 13563 -6409
rect 13695 -6517 13705 -6409
rect 14484 -6437 14551 -5054
rect 9556 -6613 9925 -6565
rect 9556 -6643 9570 -6613
rect 9556 -6660 9566 -6643
rect 9858 -6716 9924 -6613
rect 11686 -6657 11692 -6517
rect 11759 -6657 11765 -6517
rect 11686 -6669 11765 -6657
rect 14484 -6716 14550 -6437
rect 9856 -6796 14550 -6716
rect 13273 -7294 13737 -7262
rect 13825 -7278 13835 -7218
rect 13897 -7278 13907 -7218
rect 13273 -7302 13736 -7294
rect 13273 -7451 13327 -7302
rect 7710 -7799 8439 -7719
rect 7460 -7812 8439 -7799
rect 7420 -7824 8439 -7812
rect 6955 -7937 6989 -7824
rect 7425 -7828 8439 -7824
rect 12953 -7551 13327 -7451
rect 13387 -7347 13618 -7331
rect 13387 -7381 13568 -7347
rect 13602 -7381 13618 -7347
rect 13387 -7387 13618 -7381
rect 13670 -7347 13736 -7302
rect 13670 -7381 13686 -7347
rect 13720 -7381 13736 -7347
rect 13670 -7387 13736 -7381
rect 7351 -7862 7417 -7855
rect 7351 -7896 7367 -7862
rect 7401 -7896 7417 -7862
rect 7351 -7937 7417 -7896
rect 6835 -7938 7417 -7937
rect 6835 -7967 7535 -7938
rect 6835 -8061 6871 -7967
rect 7071 -8061 7107 -7967
rect 7307 -7968 7535 -7967
rect 7307 -8061 7343 -7968
rect 7469 -7979 7535 -7968
rect 7469 -8013 7485 -7979
rect 7519 -8013 7535 -7979
rect 7469 -8020 7535 -8013
rect 7779 -8061 7814 -7828
rect 6712 -8073 6758 -8061
rect 6712 -8249 6718 -8073
rect 6752 -8249 6758 -8073
rect 6712 -8261 6758 -8249
rect 6830 -8073 6876 -8061
rect 6830 -8249 6836 -8073
rect 6870 -8249 6876 -8073
rect 6830 -8261 6876 -8249
rect 6948 -8073 6994 -8061
rect 6948 -8249 6954 -8073
rect 6988 -8249 6994 -8073
rect 6948 -8261 6994 -8249
rect 7066 -8073 7112 -8061
rect 7066 -8249 7072 -8073
rect 7106 -8249 7112 -8073
rect 7066 -8261 7112 -8249
rect 7184 -8073 7230 -8061
rect 7184 -8249 7190 -8073
rect 7224 -8249 7230 -8073
rect 7184 -8261 7230 -8249
rect 7302 -8073 7348 -8061
rect 7302 -8249 7308 -8073
rect 7342 -8249 7348 -8073
rect 7302 -8261 7348 -8249
rect 7420 -8073 7466 -8061
rect 7420 -8249 7426 -8073
rect 7460 -8249 7466 -8073
rect 7420 -8261 7466 -8249
rect 7538 -8073 7584 -8061
rect 7538 -8249 7544 -8073
rect 7578 -8249 7584 -8073
rect 7538 -8261 7584 -8249
rect 7656 -8073 7702 -8061
rect 7656 -8249 7662 -8073
rect 7696 -8249 7702 -8073
rect 7656 -8261 7702 -8249
rect 7774 -8073 7820 -8061
rect 7774 -8249 7780 -8073
rect 7814 -8249 7820 -8073
rect 7774 -8261 7820 -8249
rect 6719 -8367 6751 -8261
rect 6955 -8367 6987 -8261
rect 7191 -8367 7223 -8261
rect 7427 -8367 7459 -8261
rect 7662 -8367 7696 -8261
rect 6719 -8397 7696 -8367
rect 7023 -8425 7159 -8397
rect 7023 -8487 7059 -8425
rect 7119 -8487 7159 -8425
rect 7023 -8507 7159 -8487
rect -357 -8566 416 -8565
rect 12953 -8566 13076 -7551
rect 13387 -7580 13441 -7387
rect 13829 -7415 13905 -7278
rect 13745 -7419 13905 -7415
rect -357 -8665 13076 -8566
rect 13114 -7679 13441 -7580
rect 13503 -7431 13549 -7419
rect -258 -8666 12677 -8665
rect -1124 -8695 -999 -8684
rect 13114 -8695 13219 -7679
rect 13503 -7807 13509 -7431
rect 13543 -7807 13549 -7431
rect 13503 -7819 13549 -7807
rect 13621 -7431 13667 -7419
rect 13621 -7807 13627 -7431
rect 13661 -7807 13667 -7431
rect 13621 -7819 13667 -7807
rect 13739 -7431 13905 -7419
rect 13739 -7807 13745 -7431
rect 13779 -7458 13905 -7431
rect 13779 -7807 13785 -7458
rect 13862 -7619 13905 -7458
rect 13739 -7819 13785 -7807
rect 13856 -7624 13905 -7619
rect 13856 -7631 13902 -7624
rect 13856 -7807 13862 -7631
rect 13896 -7807 13902 -7631
rect 13856 -7819 13902 -7807
rect 13974 -7631 14020 -7619
rect 13974 -7807 13980 -7631
rect 14014 -7794 14020 -7631
rect 14891 -7714 15027 -3781
rect 15595 -5145 15688 -3251
rect 15751 -3310 16217 -3288
rect 16505 -3310 16571 -3214
rect 18336 -3204 18342 -3028
rect 18376 -3204 18382 -3028
rect 18336 -3216 18382 -3204
rect 18454 -3028 18500 -3016
rect 18454 -3204 18460 -3028
rect 18494 -3204 18500 -3028
rect 18454 -3216 18500 -3204
rect 18572 -3028 18618 -3016
rect 18572 -3204 18578 -3028
rect 18612 -3204 18618 -3028
rect 18572 -3216 18618 -3204
rect 18690 -3028 18736 -3016
rect 18690 -3204 18696 -3028
rect 18730 -3083 18736 -3028
rect 18855 -3028 18901 -3016
rect 18855 -3083 18861 -3028
rect 18730 -3171 18861 -3083
rect 18730 -3204 18736 -3171
rect 18690 -3216 18736 -3204
rect 18855 -3204 18861 -3171
rect 18895 -3204 18901 -3028
rect 18855 -3216 18901 -3204
rect 18973 -3028 19019 -3016
rect 18973 -3204 18979 -3028
rect 19013 -3204 19019 -3028
rect 18973 -3216 19019 -3204
rect 19091 -3028 19137 -3016
rect 19091 -3204 19097 -3028
rect 19131 -3204 19137 -3028
rect 19091 -3216 19137 -3204
rect 19209 -3028 19255 -3016
rect 19209 -3204 19215 -3028
rect 19249 -3204 19255 -3028
rect 19209 -3216 19255 -3204
rect 18342 -3255 18376 -3216
rect 18578 -3255 18612 -3216
rect 18342 -3290 18612 -3255
rect 18979 -3254 19012 -3216
rect 19215 -3254 19248 -3216
rect 18979 -3290 19248 -3254
rect 15751 -3358 16571 -3310
rect 18376 -3291 18612 -3290
rect 15751 -3389 16217 -3358
rect 18376 -3365 18508 -3291
rect 15751 -3645 15856 -3389
rect 18366 -3473 18376 -3365
rect 18508 -3473 18518 -3365
rect 16592 -3552 16671 -3540
rect 15751 -3751 15814 -3645
rect 15926 -3751 15936 -3645
rect 16592 -3649 16598 -3552
rect 16518 -3669 16598 -3649
rect 16665 -3649 16671 -3552
rect 18396 -3606 18402 -3473
rect 18469 -3606 18475 -3473
rect 18396 -3618 18475 -3606
rect 16665 -3669 16738 -3649
rect 15751 -3762 15900 -3751
rect 15751 -4939 15856 -3762
rect 16518 -3777 16562 -3669
rect 16694 -3777 16738 -3669
rect 16518 -3819 16738 -3777
rect 19316 -3804 19378 -2233
rect 19568 -2241 19614 -2229
rect 19568 -2617 19574 -2241
rect 19608 -2617 19614 -2241
rect 19568 -2629 19614 -2617
rect 19686 -2241 19732 -2229
rect 19686 -2617 19692 -2241
rect 19726 -2617 19732 -2241
rect 19686 -2629 19732 -2617
rect 19804 -2241 19850 -2229
rect 19804 -2617 19810 -2241
rect 19844 -2617 19850 -2241
rect 19804 -2629 19850 -2617
rect 19922 -2241 19968 -2229
rect 19922 -2617 19928 -2241
rect 19962 -2617 19968 -2241
rect 19922 -2629 19968 -2617
rect 20040 -2241 20086 -2229
rect 20040 -2617 20046 -2241
rect 20080 -2617 20086 -2241
rect 20040 -2629 20086 -2617
rect 20158 -2241 20204 -2229
rect 20158 -2617 20164 -2241
rect 20198 -2617 20204 -2241
rect 20158 -2629 20204 -2617
rect 20276 -2241 20322 -2229
rect 20276 -2617 20282 -2241
rect 20316 -2617 20322 -2241
rect 20276 -2629 20322 -2617
rect 19574 -2671 19608 -2629
rect 19810 -2671 19844 -2629
rect 19574 -2699 19844 -2671
rect 19928 -2670 19962 -2629
rect 20164 -2670 20198 -2629
rect 19928 -2699 20198 -2670
rect 19574 -2747 19608 -2699
rect 19574 -2777 19637 -2747
rect 19602 -2869 19637 -2777
rect 20109 -2807 20209 -2786
rect 20109 -2861 20123 -2807
rect 20188 -2861 20209 -2807
rect 20109 -2866 20209 -2861
rect 20282 -2812 20316 -2629
rect 21497 -2660 21649 1524
rect 22225 724 22318 2618
rect 22381 2559 22847 2581
rect 23135 2559 23201 2655
rect 24966 2665 24972 2841
rect 25006 2665 25012 2841
rect 24966 2653 25012 2665
rect 25084 2841 25130 2853
rect 25084 2665 25090 2841
rect 25124 2665 25130 2841
rect 25084 2653 25130 2665
rect 25202 2841 25248 2853
rect 25202 2665 25208 2841
rect 25242 2665 25248 2841
rect 25202 2653 25248 2665
rect 25320 2841 25366 2853
rect 25320 2665 25326 2841
rect 25360 2786 25366 2841
rect 25485 2841 25531 2853
rect 25485 2786 25491 2841
rect 25360 2698 25491 2786
rect 25360 2665 25366 2698
rect 25320 2653 25366 2665
rect 25485 2665 25491 2698
rect 25525 2665 25531 2841
rect 25485 2653 25531 2665
rect 25603 2841 25649 2853
rect 25603 2665 25609 2841
rect 25643 2665 25649 2841
rect 25603 2653 25649 2665
rect 25721 2841 25767 2853
rect 25721 2665 25727 2841
rect 25761 2665 25767 2841
rect 25721 2653 25767 2665
rect 25839 2841 25885 2853
rect 25839 2665 25845 2841
rect 25879 2665 25885 2841
rect 25839 2653 25885 2665
rect 24972 2614 25006 2653
rect 25208 2614 25242 2653
rect 24972 2579 25242 2614
rect 25609 2615 25642 2653
rect 25845 2615 25878 2653
rect 25609 2579 25878 2615
rect 22381 2511 23201 2559
rect 25006 2578 25242 2579
rect 22381 2480 22847 2511
rect 25006 2504 25138 2578
rect 22381 2224 22486 2480
rect 24996 2396 25006 2504
rect 25138 2396 25148 2504
rect 23223 2315 23302 2327
rect 22381 2118 22444 2224
rect 22556 2118 22566 2224
rect 23223 2220 23229 2315
rect 23148 2200 23229 2220
rect 23296 2220 23302 2315
rect 25024 2253 25030 2396
rect 25097 2253 25103 2396
rect 25024 2241 25103 2253
rect 23296 2200 23368 2220
rect 22381 2107 22530 2118
rect 22381 930 22486 2107
rect 23148 2092 23192 2200
rect 23324 2092 23368 2200
rect 23148 2050 23368 2092
rect 25946 2065 26008 3636
rect 26198 3628 26244 3640
rect 26198 3252 26204 3628
rect 26238 3252 26244 3628
rect 26198 3240 26244 3252
rect 26316 3628 26362 3640
rect 26316 3252 26322 3628
rect 26356 3252 26362 3628
rect 26316 3240 26362 3252
rect 26434 3628 26480 3640
rect 26434 3252 26440 3628
rect 26474 3252 26480 3628
rect 26434 3240 26480 3252
rect 26552 3628 26598 3640
rect 26552 3252 26558 3628
rect 26592 3252 26598 3628
rect 26552 3240 26598 3252
rect 26670 3628 26716 3640
rect 26670 3252 26676 3628
rect 26710 3252 26716 3628
rect 26670 3240 26716 3252
rect 26788 3628 26834 3640
rect 26788 3252 26794 3628
rect 26828 3252 26834 3628
rect 26788 3240 26834 3252
rect 26906 3628 26952 3640
rect 26906 3252 26912 3628
rect 26946 3252 26952 3628
rect 26906 3240 26952 3252
rect 26204 3198 26238 3240
rect 26440 3198 26474 3240
rect 26204 3170 26474 3198
rect 26558 3199 26592 3240
rect 26794 3199 26828 3240
rect 26558 3170 26828 3199
rect 26204 3122 26238 3170
rect 26204 3092 26267 3122
rect 26232 3000 26267 3092
rect 26739 3062 26839 3083
rect 26739 3008 26753 3062
rect 26818 3008 26839 3062
rect 26739 3003 26839 3008
rect 26912 3057 26946 3240
rect 26912 3003 27021 3057
rect 26232 2964 26459 3000
rect 26232 2857 26267 2964
rect 26393 2930 26459 2964
rect 26393 2896 26409 2930
rect 26443 2896 26459 2930
rect 26740 2988 26837 3003
rect 26740 2921 26797 2988
rect 26393 2890 26459 2896
rect 26634 2885 26903 2921
rect 26634 2857 26667 2885
rect 26870 2857 26903 2885
rect 26987 2857 27021 3003
rect 27721 2996 27731 3071
rect 27799 2996 27911 5939
rect 27748 2995 27911 2996
rect 27800 2985 27911 2995
rect 26108 2845 26154 2857
rect 26108 2669 26114 2845
rect 26148 2669 26154 2845
rect 26108 2657 26154 2669
rect 26226 2845 26272 2857
rect 26226 2669 26232 2845
rect 26266 2669 26272 2845
rect 26226 2657 26272 2669
rect 26344 2845 26390 2857
rect 26344 2669 26350 2845
rect 26384 2669 26390 2845
rect 26344 2657 26390 2669
rect 26462 2845 26508 2857
rect 26462 2669 26468 2845
rect 26502 2790 26508 2845
rect 26627 2845 26673 2857
rect 26627 2790 26633 2845
rect 26502 2702 26633 2790
rect 26502 2669 26508 2702
rect 26462 2657 26508 2669
rect 26627 2669 26633 2702
rect 26667 2669 26673 2845
rect 26627 2657 26673 2669
rect 26745 2845 26791 2857
rect 26745 2669 26751 2845
rect 26785 2669 26791 2845
rect 26745 2657 26791 2669
rect 26863 2845 26909 2857
rect 26863 2669 26869 2845
rect 26903 2669 26909 2845
rect 26863 2657 26909 2669
rect 26981 2845 27027 2857
rect 26981 2669 26987 2845
rect 27021 2669 27027 2845
rect 26981 2657 27027 2669
rect 26114 2618 26148 2657
rect 26350 2618 26384 2657
rect 26114 2582 26384 2618
rect 26751 2619 26784 2657
rect 26987 2619 27020 2657
rect 26751 2583 27020 2619
rect 26114 2581 26280 2582
rect 26148 2502 26280 2581
rect 26138 2394 26148 2502
rect 26280 2394 26290 2502
rect 26167 2255 26173 2394
rect 26240 2255 26246 2394
rect 26167 2243 26246 2255
rect 22752 2020 23729 2050
rect 25946 2048 26009 2065
rect 25871 2044 26009 2048
rect 22752 1914 22784 2020
rect 22988 1914 23020 2020
rect 23224 1914 23256 2020
rect 23460 1914 23492 2020
rect 23695 1914 23729 2020
rect 24039 2010 26009 2044
rect 24037 1981 26009 2010
rect 24037 1965 24083 1981
rect 25871 1979 26009 1981
rect 22745 1902 22791 1914
rect 22745 1726 22751 1902
rect 22785 1726 22791 1902
rect 22745 1714 22791 1726
rect 22863 1902 22909 1914
rect 22863 1726 22869 1902
rect 22903 1726 22909 1902
rect 22863 1714 22909 1726
rect 22981 1902 23027 1914
rect 22981 1726 22987 1902
rect 23021 1726 23027 1902
rect 22981 1714 23027 1726
rect 23099 1902 23145 1914
rect 23099 1726 23105 1902
rect 23139 1726 23145 1902
rect 23099 1714 23145 1726
rect 23217 1902 23263 1914
rect 23217 1726 23223 1902
rect 23257 1726 23263 1902
rect 23217 1714 23263 1726
rect 23335 1902 23381 1914
rect 23335 1726 23341 1902
rect 23375 1726 23381 1902
rect 23335 1714 23381 1726
rect 23453 1902 23499 1914
rect 23453 1726 23459 1902
rect 23493 1726 23499 1902
rect 23453 1714 23499 1726
rect 23571 1902 23617 1914
rect 23571 1726 23577 1902
rect 23611 1726 23617 1902
rect 23571 1714 23617 1726
rect 23689 1902 23735 1914
rect 23689 1726 23695 1902
rect 23729 1726 23735 1902
rect 23689 1714 23735 1726
rect 23807 1902 23853 1914
rect 23807 1726 23813 1902
rect 23847 1726 23853 1902
rect 23807 1714 23853 1726
rect 22868 1620 22904 1714
rect 23104 1620 23140 1714
rect 23340 1621 23376 1714
rect 23502 1666 23568 1673
rect 23502 1632 23518 1666
rect 23552 1632 23568 1666
rect 23502 1621 23568 1632
rect 23340 1620 23568 1621
rect 22868 1591 23568 1620
rect 22868 1590 23450 1591
rect 22988 1477 23022 1590
rect 23384 1549 23450 1590
rect 23384 1515 23400 1549
rect 23434 1515 23450 1549
rect 23384 1508 23450 1515
rect 23812 1496 23847 1714
rect 24036 1513 24083 1965
rect 26930 1970 27009 1982
rect 26930 1857 26936 1970
rect 27003 1857 27009 1970
rect 24995 1749 25005 1857
rect 25137 1749 25147 1857
rect 26893 1749 26903 1857
rect 27035 1749 27045 1857
rect 25005 1709 25137 1749
rect 26903 1709 27035 1749
rect 25004 1643 25137 1709
rect 26902 1643 27035 1709
rect 24333 1600 25806 1643
rect 24036 1497 24082 1513
rect 24001 1496 24082 1497
rect 23812 1481 24082 1496
rect 23458 1477 24082 1481
rect 22982 1465 23028 1477
rect 22717 987 22727 1105
rect 22845 1073 22855 1105
rect 22982 1089 22988 1465
rect 23022 1089 23028 1465
rect 22982 1077 23028 1089
rect 23100 1465 23146 1477
rect 23100 1089 23106 1465
rect 23140 1089 23146 1465
rect 23100 1077 23146 1089
rect 23218 1465 23264 1477
rect 23218 1089 23224 1465
rect 23258 1113 23264 1465
rect 23335 1465 23381 1477
rect 23335 1289 23341 1465
rect 23375 1289 23381 1465
rect 23335 1277 23381 1289
rect 23453 1465 24082 1477
rect 23453 1289 23459 1465
rect 23493 1453 24082 1465
rect 23493 1452 23735 1453
rect 23493 1289 23499 1452
rect 24001 1451 24082 1453
rect 24333 1297 24367 1600
rect 24699 1497 24733 1600
rect 24935 1497 24969 1600
rect 25171 1497 25205 1600
rect 25407 1497 25441 1600
rect 24693 1485 24739 1497
rect 23453 1277 23499 1289
rect 24209 1285 24255 1297
rect 23341 1161 23376 1277
rect 23472 1161 23580 1171
rect 23341 1113 23472 1161
rect 23580 1121 23719 1127
rect 23258 1089 23472 1113
rect 23218 1077 23472 1089
rect 23224 1073 23472 1077
rect 22845 1045 22860 1073
rect 22845 1039 23097 1045
rect 22845 1005 23047 1039
rect 23081 1005 23097 1039
rect 22845 989 23097 1005
rect 23149 1039 23215 1045
rect 23149 1005 23165 1039
rect 23199 1005 23215 1039
rect 23398 1029 23472 1073
rect 23707 1054 23719 1121
rect 24209 1109 24215 1285
rect 24249 1109 24255 1285
rect 24209 1097 24255 1109
rect 24327 1285 24373 1297
rect 24327 1109 24333 1285
rect 24367 1109 24373 1285
rect 24327 1097 24373 1109
rect 24445 1285 24491 1297
rect 24445 1109 24451 1285
rect 24485 1109 24491 1285
rect 24445 1097 24491 1109
rect 24563 1285 24609 1297
rect 24693 1285 24699 1485
rect 24563 1109 24569 1285
rect 24603 1109 24699 1285
rect 24733 1109 24739 1485
rect 24563 1097 24609 1109
rect 24693 1097 24739 1109
rect 24811 1485 24857 1497
rect 24811 1109 24817 1485
rect 24851 1109 24857 1485
rect 24811 1097 24857 1109
rect 24929 1485 24975 1497
rect 24929 1109 24935 1485
rect 24969 1109 24975 1485
rect 24929 1097 24975 1109
rect 25047 1485 25093 1497
rect 25047 1109 25053 1485
rect 25087 1109 25093 1485
rect 25047 1097 25093 1109
rect 25165 1485 25211 1497
rect 25165 1109 25171 1485
rect 25205 1109 25211 1485
rect 25165 1097 25211 1109
rect 25283 1485 25329 1497
rect 25283 1109 25289 1485
rect 25323 1109 25329 1485
rect 25283 1097 25329 1109
rect 25401 1485 25447 1497
rect 25401 1109 25407 1485
rect 25441 1285 25447 1485
rect 25772 1297 25806 1600
rect 26231 1600 27704 1643
rect 26231 1297 26265 1600
rect 26597 1497 26631 1600
rect 26833 1497 26867 1600
rect 27069 1497 27103 1600
rect 27305 1497 27339 1600
rect 26591 1485 26637 1497
rect 25530 1285 25576 1297
rect 25441 1109 25536 1285
rect 25570 1109 25576 1285
rect 25401 1097 25447 1109
rect 25530 1097 25576 1109
rect 25648 1285 25694 1297
rect 25648 1109 25654 1285
rect 25688 1109 25694 1285
rect 25648 1097 25694 1109
rect 25766 1285 25812 1297
rect 25766 1109 25772 1285
rect 25806 1109 25812 1285
rect 25766 1097 25812 1109
rect 25884 1285 25930 1297
rect 25884 1109 25890 1285
rect 25924 1109 25930 1285
rect 25884 1097 25930 1109
rect 26107 1285 26153 1297
rect 26107 1109 26113 1285
rect 26147 1109 26153 1285
rect 26107 1097 26153 1109
rect 26225 1285 26271 1297
rect 26225 1109 26231 1285
rect 26265 1109 26271 1285
rect 26225 1097 26271 1109
rect 26343 1285 26389 1297
rect 26343 1109 26349 1285
rect 26383 1109 26389 1285
rect 26343 1097 26389 1109
rect 26461 1285 26507 1297
rect 26591 1285 26597 1485
rect 26461 1109 26467 1285
rect 26501 1109 26597 1285
rect 26631 1109 26637 1485
rect 26461 1097 26507 1109
rect 26591 1097 26637 1109
rect 26709 1485 26755 1497
rect 26709 1109 26715 1485
rect 26749 1109 26755 1485
rect 26709 1097 26755 1109
rect 26827 1485 26873 1497
rect 26827 1109 26833 1485
rect 26867 1109 26873 1485
rect 26827 1097 26873 1109
rect 26945 1485 26991 1497
rect 26945 1109 26951 1485
rect 26985 1109 26991 1485
rect 26945 1097 26991 1109
rect 27063 1485 27109 1497
rect 27063 1109 27069 1485
rect 27103 1109 27109 1485
rect 27063 1097 27109 1109
rect 27181 1485 27227 1497
rect 27181 1109 27187 1485
rect 27221 1109 27227 1485
rect 27181 1097 27227 1109
rect 27299 1485 27345 1497
rect 27299 1109 27305 1485
rect 27339 1285 27345 1485
rect 27670 1297 27704 1600
rect 27428 1285 27474 1297
rect 27339 1109 27434 1285
rect 27468 1109 27474 1285
rect 27299 1097 27345 1109
rect 27428 1097 27474 1109
rect 27546 1285 27592 1297
rect 27546 1109 27552 1285
rect 27586 1109 27592 1285
rect 27546 1097 27592 1109
rect 27664 1285 27710 1297
rect 27664 1109 27670 1285
rect 27704 1109 27710 1285
rect 27664 1097 27710 1109
rect 27782 1285 27828 1297
rect 27782 1109 27788 1285
rect 27822 1109 27828 1285
rect 27782 1097 27828 1109
rect 23580 1048 23719 1054
rect 24215 1063 24249 1097
rect 24817 1063 24851 1097
rect 25053 1063 25087 1097
rect 23472 1019 23580 1029
rect 24215 1028 24374 1063
rect 24817 1028 25087 1063
rect 25654 1063 25688 1097
rect 25890 1063 25924 1097
rect 25654 1028 25924 1063
rect 26113 1063 26147 1097
rect 26715 1063 26749 1097
rect 26951 1063 26985 1097
rect 26113 1028 26272 1063
rect 26715 1028 26985 1063
rect 27552 1063 27586 1097
rect 27788 1063 27822 1097
rect 27552 1028 27822 1063
rect 22845 987 22860 989
rect 22760 973 22860 987
rect 22760 930 22860 931
rect 22381 909 22860 930
rect 23149 909 23215 1005
rect 22381 861 23215 909
rect 22381 832 22860 861
rect 22381 830 22486 832
rect 22760 831 22860 832
rect 22214 645 22224 724
rect 22317 645 22327 724
rect 23215 707 23294 719
rect 21739 318 21847 330
rect 21735 218 21745 318
rect 21841 218 21851 318
rect 21739 206 21847 218
rect 22225 -529 22318 645
rect 23215 616 23221 707
rect 23143 596 23221 616
rect 23288 616 23294 707
rect 23288 596 23363 616
rect 23143 488 23187 596
rect 23319 488 23363 596
rect 23143 446 23363 488
rect 22747 416 23724 446
rect 22747 310 22779 416
rect 22983 310 23015 416
rect 23219 310 23251 416
rect 23455 310 23487 416
rect 23690 310 23724 416
rect 22740 298 22786 310
rect 22740 122 22746 298
rect 22780 122 22786 298
rect 22740 110 22786 122
rect 22858 298 22904 310
rect 22858 122 22864 298
rect 22898 122 22904 298
rect 22858 110 22904 122
rect 22976 298 23022 310
rect 22976 122 22982 298
rect 23016 122 23022 298
rect 22976 110 23022 122
rect 23094 298 23140 310
rect 23094 122 23100 298
rect 23134 122 23140 298
rect 23094 110 23140 122
rect 23212 298 23258 310
rect 23212 122 23218 298
rect 23252 122 23258 298
rect 23212 110 23258 122
rect 23330 298 23376 310
rect 23330 122 23336 298
rect 23370 122 23376 298
rect 23330 110 23376 122
rect 23448 298 23494 310
rect 23448 122 23454 298
rect 23488 122 23494 298
rect 23448 110 23494 122
rect 23566 298 23612 310
rect 23566 122 23572 298
rect 23606 122 23612 298
rect 23566 110 23612 122
rect 23684 298 23730 310
rect 23684 122 23690 298
rect 23724 122 23730 298
rect 23684 110 23730 122
rect 23802 298 23848 310
rect 23802 122 23808 298
rect 23842 122 23848 298
rect 23802 110 23848 122
rect 24340 244 24374 1028
rect 25053 966 25087 1028
rect 24642 928 25384 966
rect 24642 804 24676 928
rect 24878 804 24912 928
rect 25114 804 25148 928
rect 25350 804 25384 928
rect 25640 821 25650 887
rect 25713 821 25723 887
rect 24636 792 24682 804
rect 24636 416 24642 792
rect 24676 416 24682 792
rect 24636 404 24682 416
rect 24754 792 24800 804
rect 24754 416 24760 792
rect 24794 416 24800 792
rect 24754 404 24800 416
rect 24872 792 24918 804
rect 24872 416 24878 792
rect 24912 416 24918 792
rect 24872 404 24918 416
rect 24990 792 25036 804
rect 24990 416 24996 792
rect 25030 416 25036 792
rect 24990 404 25036 416
rect 25108 792 25154 804
rect 25108 416 25114 792
rect 25148 416 25154 792
rect 25108 404 25154 416
rect 25226 792 25272 804
rect 25226 416 25232 792
rect 25266 416 25272 792
rect 25226 404 25272 416
rect 25344 792 25390 804
rect 25344 416 25350 792
rect 25384 416 25390 792
rect 25344 404 25390 416
rect 25756 245 25790 1028
rect 25483 244 25790 245
rect 24340 239 24656 244
rect 25370 239 25790 244
rect 24340 228 24723 239
rect 24340 201 24672 228
rect 22863 16 22899 110
rect 23099 16 23135 110
rect 23335 17 23371 110
rect 23497 62 23563 69
rect 23497 28 23513 62
rect 23547 28 23563 62
rect 23497 17 23563 28
rect 23335 16 23563 17
rect 22863 -13 23563 16
rect 22863 -14 23445 -13
rect 22983 -127 23017 -14
rect 23379 -55 23445 -14
rect 23379 -89 23395 -55
rect 23429 -89 23445 -55
rect 23379 -96 23445 -89
rect 23807 -123 23842 110
rect 24340 72 24374 201
rect 24656 194 24672 201
rect 24706 194 24723 228
rect 24656 188 24723 194
rect 25303 228 25790 239
rect 25303 194 25320 228
rect 25354 201 25790 228
rect 25354 194 25370 201
rect 25483 200 25790 201
rect 25303 188 25370 194
rect 24481 161 24537 173
rect 24481 127 24487 161
rect 24521 160 24537 161
rect 25594 160 25650 172
rect 24521 144 24988 160
rect 24521 127 24938 144
rect 24481 111 24938 127
rect 24922 110 24938 111
rect 24972 110 24988 144
rect 24922 103 24988 110
rect 25040 145 25610 160
rect 25040 111 25056 145
rect 25090 126 25610 145
rect 25644 126 25650 160
rect 25090 111 25650 126
rect 25040 101 25107 111
rect 25594 110 25650 111
rect 25756 72 25790 200
rect 26238 244 26272 1028
rect 26951 966 26985 1028
rect 26540 928 27282 966
rect 26540 804 26574 928
rect 26776 804 26810 928
rect 27012 804 27046 928
rect 27248 804 27282 928
rect 26534 792 26580 804
rect 26534 416 26540 792
rect 26574 416 26580 792
rect 26534 404 26580 416
rect 26652 792 26698 804
rect 26652 416 26658 792
rect 26692 416 26698 792
rect 26652 404 26698 416
rect 26770 792 26816 804
rect 26770 416 26776 792
rect 26810 416 26816 792
rect 26770 404 26816 416
rect 26888 792 26934 804
rect 26888 416 26894 792
rect 26928 416 26934 792
rect 26888 404 26934 416
rect 27006 792 27052 804
rect 27006 416 27012 792
rect 27046 416 27052 792
rect 27006 404 27052 416
rect 27124 792 27170 804
rect 27124 416 27130 792
rect 27164 416 27170 792
rect 27124 404 27170 416
rect 27242 792 27288 804
rect 27242 416 27248 792
rect 27282 416 27288 792
rect 27242 404 27288 416
rect 27654 245 27688 1028
rect 27266 244 27335 245
rect 27381 244 27688 245
rect 26238 239 26554 244
rect 27266 240 27688 244
rect 26238 228 26621 239
rect 26238 201 26570 228
rect 26238 72 26272 201
rect 26554 194 26570 201
rect 26604 194 26621 228
rect 26554 188 26621 194
rect 27199 229 27688 240
rect 27199 195 27216 229
rect 27250 201 27688 229
rect 27250 195 27266 201
rect 27381 200 27688 201
rect 27199 189 27266 195
rect 26379 161 26435 173
rect 26379 127 26385 161
rect 26419 160 26435 161
rect 27492 160 27548 172
rect 26419 144 26886 160
rect 26419 127 26836 144
rect 26379 111 26836 127
rect 26820 110 26836 111
rect 26870 110 26886 144
rect 26820 103 26886 110
rect 26938 145 27508 160
rect 26938 111 26954 145
rect 26988 126 27508 145
rect 27542 126 27548 160
rect 26988 111 27548 126
rect 26938 101 27005 111
rect 27492 110 27548 111
rect 27654 72 27688 200
rect 27769 850 27836 874
rect 27769 816 27786 850
rect 27820 816 27836 850
rect 23453 -127 23842 -123
rect 22977 -139 23023 -127
rect 22977 -515 22983 -139
rect 23017 -515 23023 -139
rect 22977 -527 23023 -515
rect 23095 -139 23141 -127
rect 23095 -515 23101 -139
rect 23135 -515 23141 -139
rect 23095 -527 23141 -515
rect 23213 -139 23259 -127
rect 23213 -515 23219 -139
rect 23253 -491 23259 -139
rect 23330 -139 23376 -127
rect 23330 -315 23336 -139
rect 23370 -315 23376 -139
rect 23330 -327 23376 -315
rect 23448 -139 23842 -127
rect 24334 60 24380 72
rect 24334 -116 24340 60
rect 24374 -116 24380 60
rect 24334 -128 24380 -116
rect 24452 60 24498 72
rect 24452 -116 24458 60
rect 24492 -116 24498 60
rect 24452 -128 24498 -116
rect 24754 60 24800 72
rect 23448 -315 23454 -139
rect 23488 -152 23842 -139
rect 23488 -315 23494 -152
rect 23764 -155 23842 -152
rect 23764 -207 23774 -155
rect 23837 -207 23847 -155
rect 23769 -213 23842 -207
rect 23448 -327 23494 -315
rect 23336 -443 23371 -327
rect 24457 -422 24491 -128
rect 24754 -316 24760 60
rect 24794 -316 24800 60
rect 24754 -328 24800 -316
rect 24872 60 24918 72
rect 24872 -316 24878 60
rect 24912 -316 24918 60
rect 24872 -328 24918 -316
rect 24990 60 25036 72
rect 24990 -316 24996 60
rect 25030 -316 25036 60
rect 24990 -328 25036 -316
rect 25108 60 25154 72
rect 25108 -316 25114 60
rect 25148 -316 25154 60
rect 25108 -328 25154 -316
rect 25226 60 25272 72
rect 25226 -316 25232 60
rect 25266 -316 25272 60
rect 25632 60 25678 72
rect 25632 -116 25638 60
rect 25672 -116 25678 60
rect 25632 -128 25678 -116
rect 25750 60 25796 72
rect 25750 -116 25756 60
rect 25790 -116 25796 60
rect 25750 -128 25796 -116
rect 26232 60 26278 72
rect 26232 -116 26238 60
rect 26272 -116 26278 60
rect 26232 -128 26278 -116
rect 26350 60 26396 72
rect 26350 -116 26356 60
rect 26390 -116 26396 60
rect 26350 -128 26396 -116
rect 26652 60 26698 72
rect 25226 -328 25272 -316
rect 25114 -422 25148 -328
rect 25638 -422 25671 -128
rect 23467 -443 23575 -433
rect 23336 -491 23467 -443
rect 24457 -454 25671 -422
rect 26355 -422 26389 -128
rect 26652 -316 26658 60
rect 26692 -316 26698 60
rect 26652 -328 26698 -316
rect 26770 60 26816 72
rect 26770 -316 26776 60
rect 26810 -316 26816 60
rect 26770 -328 26816 -316
rect 26888 60 26934 72
rect 26888 -316 26894 60
rect 26928 -316 26934 60
rect 26888 -328 26934 -316
rect 27006 60 27052 72
rect 27006 -316 27012 60
rect 27046 -316 27052 60
rect 27006 -328 27052 -316
rect 27124 60 27170 72
rect 27124 -316 27130 60
rect 27164 -316 27170 60
rect 27530 60 27576 72
rect 27530 -116 27536 60
rect 27570 -116 27576 60
rect 27530 -128 27576 -116
rect 27648 60 27694 72
rect 27648 -116 27654 60
rect 27688 -116 27694 60
rect 27648 -128 27694 -116
rect 27124 -328 27170 -316
rect 27012 -422 27046 -328
rect 27536 -422 27569 -128
rect 26355 -454 27569 -422
rect 23575 -484 23725 -478
rect 23253 -515 23467 -491
rect 23213 -527 23467 -515
rect 22225 -531 22810 -529
rect 23219 -531 23467 -527
rect 22225 -559 22855 -531
rect 22225 -565 23092 -559
rect 22225 -599 23042 -565
rect 23076 -599 23092 -565
rect 22225 -615 23092 -599
rect 23144 -565 23210 -559
rect 23144 -599 23160 -565
rect 23194 -599 23210 -565
rect 23393 -575 23467 -531
rect 23713 -551 23725 -484
rect 24950 -539 25082 -454
rect 26848 -539 26980 -454
rect 23575 -557 23725 -551
rect 23467 -585 23575 -575
rect 22225 -631 22855 -615
rect 22225 -635 22810 -631
rect 22225 -636 22326 -635
rect 22755 -684 22855 -673
rect 22719 -790 22729 -684
rect 22841 -695 22855 -684
rect 23144 -695 23210 -599
rect 24940 -647 24950 -539
rect 25082 -647 25092 -539
rect 26838 -647 26848 -539
rect 26980 -647 26990 -539
rect 27769 -567 27836 816
rect 27982 393 28082 6232
rect 28844 5722 28980 5742
rect 28844 5660 28880 5722
rect 28940 5660 28980 5722
rect 28844 5632 28980 5660
rect 28540 5602 29517 5632
rect 28540 5496 28572 5602
rect 28776 5496 28808 5602
rect 29012 5496 29044 5602
rect 29248 5496 29280 5602
rect 29483 5496 29517 5602
rect 28533 5484 28579 5496
rect 28533 5308 28539 5484
rect 28573 5308 28579 5484
rect 28533 5296 28579 5308
rect 28651 5484 28697 5496
rect 28651 5308 28657 5484
rect 28691 5308 28697 5484
rect 28651 5296 28697 5308
rect 28769 5484 28815 5496
rect 28769 5308 28775 5484
rect 28809 5308 28815 5484
rect 28769 5296 28815 5308
rect 28887 5484 28933 5496
rect 28887 5308 28893 5484
rect 28927 5308 28933 5484
rect 28887 5296 28933 5308
rect 29005 5484 29051 5496
rect 29005 5308 29011 5484
rect 29045 5308 29051 5484
rect 29005 5296 29051 5308
rect 29123 5484 29169 5496
rect 29123 5308 29129 5484
rect 29163 5308 29169 5484
rect 29123 5296 29169 5308
rect 29241 5484 29287 5496
rect 29241 5308 29247 5484
rect 29281 5308 29287 5484
rect 29241 5296 29287 5308
rect 29359 5484 29405 5496
rect 29359 5308 29365 5484
rect 29399 5308 29405 5484
rect 29359 5296 29405 5308
rect 29477 5484 29523 5496
rect 29477 5308 29483 5484
rect 29517 5308 29523 5484
rect 29477 5296 29523 5308
rect 29595 5484 29641 5496
rect 29595 5308 29601 5484
rect 29635 5308 29641 5484
rect 29595 5296 29641 5308
rect 28656 5202 28692 5296
rect 28892 5202 28928 5296
rect 29128 5203 29164 5296
rect 29290 5248 29356 5255
rect 29290 5214 29306 5248
rect 29340 5214 29356 5248
rect 29290 5203 29356 5214
rect 29128 5202 29356 5203
rect 28656 5173 29356 5202
rect 28656 5172 29238 5173
rect 28776 5059 28810 5172
rect 29172 5131 29238 5172
rect 29172 5097 29188 5131
rect 29222 5097 29238 5131
rect 29172 5090 29238 5097
rect 29600 5064 29635 5296
rect 29716 5064 29811 6227
rect 30969 5817 31414 5823
rect 30969 5617 30981 5817
rect 31402 5617 31414 5817
rect 30969 5611 31137 5617
rect 31127 5543 31137 5611
rect 31269 5611 31414 5617
rect 31269 5543 31279 5611
rect 31137 5503 31269 5543
rect 31136 5437 31269 5503
rect 30465 5394 31938 5437
rect 30465 5091 30499 5394
rect 30831 5291 30865 5394
rect 31067 5291 31101 5394
rect 31303 5291 31337 5394
rect 31539 5291 31573 5394
rect 30825 5279 30871 5291
rect 29545 5063 29811 5064
rect 29246 5059 29811 5063
rect 28770 5047 28816 5059
rect 28770 4671 28776 5047
rect 28810 4671 28816 5047
rect 28770 4659 28816 4671
rect 28888 5047 28934 5059
rect 28888 4671 28894 5047
rect 28928 4671 28934 5047
rect 28888 4659 28934 4671
rect 29006 5047 29052 5059
rect 29006 4671 29012 5047
rect 29046 4698 29052 5047
rect 29123 5047 29169 5059
rect 29123 4871 29129 5047
rect 29163 4871 29169 5047
rect 29123 4864 29169 4871
rect 29241 5047 29811 5059
rect 29241 4871 29247 5047
rect 29281 5034 29811 5047
rect 29281 4871 29287 5034
rect 29531 4954 29811 5034
rect 29545 4953 29811 4954
rect 30341 5079 30387 5091
rect 30341 4903 30347 5079
rect 30381 4903 30387 5079
rect 30341 4891 30387 4903
rect 30459 5079 30505 5091
rect 30459 4903 30465 5079
rect 30499 4903 30505 5079
rect 30459 4891 30505 4903
rect 30577 5079 30623 5091
rect 30577 4903 30583 5079
rect 30617 4903 30623 5079
rect 30577 4891 30623 4903
rect 30695 5079 30741 5091
rect 30825 5079 30831 5279
rect 30695 4903 30701 5079
rect 30735 4903 30831 5079
rect 30865 4903 30871 5279
rect 30695 4891 30741 4903
rect 30825 4891 30871 4903
rect 30943 5279 30989 5291
rect 30943 4903 30949 5279
rect 30983 4903 30989 5279
rect 30943 4891 30989 4903
rect 31061 5279 31107 5291
rect 31061 4903 31067 5279
rect 31101 4903 31107 5279
rect 31061 4891 31107 4903
rect 31179 5279 31225 5291
rect 31179 4903 31185 5279
rect 31219 4903 31225 5279
rect 31179 4891 31225 4903
rect 31297 5279 31343 5291
rect 31297 4903 31303 5279
rect 31337 4903 31343 5279
rect 31297 4891 31343 4903
rect 31415 5279 31461 5291
rect 31415 4903 31421 5279
rect 31455 4903 31461 5279
rect 31415 4891 31461 4903
rect 31533 5279 31579 5291
rect 31533 4903 31539 5279
rect 31573 5079 31579 5279
rect 31904 5091 31938 5394
rect 32445 5314 32581 5334
rect 32445 5252 32481 5314
rect 32541 5252 32581 5314
rect 32445 5224 32581 5252
rect 32141 5194 33118 5224
rect 31662 5079 31708 5091
rect 31573 4903 31668 5079
rect 31702 4903 31708 5079
rect 31533 4891 31579 4903
rect 31662 4891 31708 4903
rect 31780 5079 31826 5091
rect 31780 4903 31786 5079
rect 31820 4903 31826 5079
rect 31780 4891 31826 4903
rect 31898 5079 31944 5091
rect 31898 4903 31904 5079
rect 31938 4903 31944 5079
rect 31898 4891 31944 4903
rect 32016 5079 32062 5091
rect 32141 5088 32173 5194
rect 32377 5088 32409 5194
rect 32613 5088 32645 5194
rect 32849 5088 32881 5194
rect 33084 5088 33118 5194
rect 32016 4903 32022 5079
rect 32056 4903 32062 5079
rect 32016 4891 32062 4903
rect 32134 5076 32180 5088
rect 32134 4900 32140 5076
rect 32174 4900 32180 5076
rect 29123 4859 29172 4864
rect 29241 4859 29287 4871
rect 29129 4698 29172 4859
rect 30347 4857 30381 4891
rect 30949 4857 30983 4891
rect 31185 4857 31219 4891
rect 30347 4822 30506 4857
rect 30949 4822 31219 4857
rect 31786 4857 31820 4891
rect 32022 4857 32056 4891
rect 32134 4888 32180 4900
rect 32252 5076 32298 5088
rect 32252 4900 32258 5076
rect 32292 4900 32298 5076
rect 32252 4888 32298 4900
rect 32370 5076 32416 5088
rect 32370 4900 32376 5076
rect 32410 4900 32416 5076
rect 32370 4888 32416 4900
rect 32488 5076 32534 5088
rect 32488 4900 32494 5076
rect 32528 4900 32534 5076
rect 32488 4888 32534 4900
rect 32606 5076 32652 5088
rect 32606 4900 32612 5076
rect 32646 4900 32652 5076
rect 32606 4888 32652 4900
rect 32724 5076 32770 5088
rect 32724 4900 32730 5076
rect 32764 4900 32770 5076
rect 32724 4888 32770 4900
rect 32842 5076 32888 5088
rect 32842 4900 32848 5076
rect 32882 4900 32888 5076
rect 32842 4888 32888 4900
rect 32960 5076 33006 5088
rect 32960 4900 32966 5076
rect 33000 4900 33006 5076
rect 32960 4888 33006 4900
rect 33078 5076 33124 5088
rect 33078 4900 33084 5076
rect 33118 4900 33124 5076
rect 33078 4888 33124 4900
rect 33196 5076 33242 5088
rect 33196 4900 33202 5076
rect 33236 4900 33242 5076
rect 33196 4888 33242 4900
rect 31786 4822 32056 4857
rect 30283 4740 30412 4741
rect 29046 4671 29172 4698
rect 29006 4659 29172 4671
rect 29012 4655 29172 4659
rect 28220 4653 28307 4654
rect 28220 4649 28603 4653
rect 28215 4575 28225 4649
rect 28304 4628 28603 4649
rect 28304 4627 28737 4628
rect 28304 4621 28885 4627
rect 28304 4587 28835 4621
rect 28869 4587 28885 4621
rect 28304 4575 28885 4587
rect 27897 387 28082 393
rect 27897 289 27909 387
rect 28041 289 28082 387
rect 27897 283 28082 289
rect 27982 282 28082 283
rect 28220 4571 28885 4575
rect 28937 4621 29003 4627
rect 28937 4587 28953 4621
rect 28987 4587 29003 4621
rect 22841 -743 23210 -695
rect 22841 -773 22855 -743
rect 22841 -790 22851 -773
rect 23143 -846 23209 -743
rect 24974 -785 24980 -647
rect 25047 -785 25053 -647
rect 24974 -797 25053 -785
rect 27769 -846 27835 -567
rect 23141 -926 27835 -846
rect 28220 -813 28310 4571
rect 28937 4542 29003 4587
rect 28370 4535 29003 4542
rect 28367 4439 28377 4535
rect 28458 4534 29003 4535
rect 28458 4502 29004 4534
rect 29096 4518 29172 4655
rect 29882 4737 30412 4740
rect 29882 4674 30334 4737
rect 30401 4674 30412 4737
rect 29882 4671 30412 4674
rect 28458 4439 28603 4502
rect 29092 4458 29102 4518
rect 29164 4458 29174 4518
rect 29882 4451 30024 4671
rect 30314 4615 30418 4621
rect 30314 4547 30326 4615
rect 30406 4547 30418 4615
rect 30314 4541 30418 4547
rect 28370 2348 28464 4439
rect 28839 3151 28975 3171
rect 28839 3089 28875 3151
rect 28935 3089 28975 3151
rect 28839 3061 28975 3089
rect 28535 3031 29512 3061
rect 28535 2925 28567 3031
rect 28771 2925 28803 3031
rect 29007 2925 29039 3031
rect 29243 2925 29275 3031
rect 29478 2925 29512 3031
rect 28528 2913 28574 2925
rect 28528 2737 28534 2913
rect 28568 2737 28574 2913
rect 28528 2725 28574 2737
rect 28646 2913 28692 2925
rect 28646 2737 28652 2913
rect 28686 2737 28692 2913
rect 28646 2725 28692 2737
rect 28764 2913 28810 2925
rect 28764 2737 28770 2913
rect 28804 2737 28810 2913
rect 28764 2725 28810 2737
rect 28882 2913 28928 2925
rect 28882 2737 28888 2913
rect 28922 2737 28928 2913
rect 28882 2725 28928 2737
rect 29000 2913 29046 2925
rect 29000 2737 29006 2913
rect 29040 2737 29046 2913
rect 29000 2725 29046 2737
rect 29118 2913 29164 2925
rect 29118 2737 29124 2913
rect 29158 2737 29164 2913
rect 29118 2725 29164 2737
rect 29236 2913 29282 2925
rect 29236 2737 29242 2913
rect 29276 2737 29282 2913
rect 29236 2725 29282 2737
rect 29354 2913 29400 2925
rect 29354 2737 29360 2913
rect 29394 2737 29400 2913
rect 29354 2725 29400 2737
rect 29472 2913 29518 2925
rect 29472 2737 29478 2913
rect 29512 2737 29518 2913
rect 29472 2725 29518 2737
rect 29590 2913 29636 2925
rect 29590 2737 29596 2913
rect 29630 2737 29636 2913
rect 29590 2725 29636 2737
rect 28651 2631 28687 2725
rect 28887 2631 28923 2725
rect 29123 2632 29159 2725
rect 29285 2677 29351 2684
rect 29285 2643 29301 2677
rect 29335 2643 29351 2677
rect 29285 2632 29351 2643
rect 29123 2631 29351 2632
rect 28651 2602 29351 2631
rect 28651 2601 29233 2602
rect 28771 2488 28805 2601
rect 29167 2560 29233 2601
rect 29167 2526 29183 2560
rect 29217 2526 29233 2560
rect 29167 2519 29233 2526
rect 29595 2492 29630 2725
rect 29882 2492 30023 4451
rect 30472 4038 30506 4822
rect 31185 4760 31219 4822
rect 30774 4722 31516 4760
rect 30584 4551 30594 4619
rect 30649 4551 30659 4619
rect 30774 4598 30808 4722
rect 31010 4598 31044 4722
rect 31246 4598 31280 4722
rect 31482 4598 31516 4722
rect 30768 4586 30814 4598
rect 30768 4210 30774 4586
rect 30808 4210 30814 4586
rect 30768 4198 30814 4210
rect 30886 4586 30932 4598
rect 30886 4210 30892 4586
rect 30926 4210 30932 4586
rect 30886 4198 30932 4210
rect 31004 4586 31050 4598
rect 31004 4210 31010 4586
rect 31044 4210 31050 4586
rect 31004 4198 31050 4210
rect 31122 4586 31168 4598
rect 31122 4210 31128 4586
rect 31162 4210 31168 4586
rect 31122 4198 31168 4210
rect 31240 4586 31286 4598
rect 31240 4210 31246 4586
rect 31280 4210 31286 4586
rect 31240 4198 31286 4210
rect 31358 4586 31404 4598
rect 31358 4210 31364 4586
rect 31398 4210 31404 4586
rect 31358 4198 31404 4210
rect 31476 4586 31522 4598
rect 31476 4210 31482 4586
rect 31516 4210 31522 4586
rect 31642 4381 31716 4393
rect 31638 4290 31648 4381
rect 31710 4290 31720 4381
rect 31642 4278 31716 4290
rect 31476 4198 31522 4210
rect 31888 4039 31922 4822
rect 32257 4794 32293 4888
rect 32493 4794 32529 4888
rect 32729 4795 32765 4888
rect 32891 4840 32957 4847
rect 32891 4806 32907 4840
rect 32941 4806 32957 4840
rect 32891 4795 32957 4806
rect 32729 4794 32957 4795
rect 32257 4765 32957 4794
rect 32257 4764 32839 4765
rect 31983 4732 32059 4737
rect 31980 4676 31990 4732
rect 32043 4731 32059 4732
rect 32043 4676 32309 4731
rect 31983 4671 32309 4676
rect 32104 4629 32195 4634
rect 32104 4540 32114 4629
rect 32187 4540 32195 4629
rect 32104 4528 32195 4540
rect 32141 4134 32195 4528
rect 32255 4219 32309 4671
rect 32377 4651 32411 4764
rect 32773 4723 32839 4764
rect 32773 4689 32789 4723
rect 32823 4689 32839 4723
rect 32773 4682 32839 4689
rect 33201 4655 33236 4888
rect 32847 4651 33236 4655
rect 32371 4639 32417 4651
rect 32371 4263 32377 4639
rect 32411 4263 32417 4639
rect 32371 4251 32417 4263
rect 32489 4639 32535 4651
rect 32489 4263 32495 4639
rect 32529 4263 32535 4639
rect 32489 4251 32535 4263
rect 32607 4639 32653 4651
rect 32607 4263 32613 4639
rect 32647 4290 32653 4639
rect 32724 4639 32770 4651
rect 32724 4463 32730 4639
rect 32764 4463 32770 4639
rect 32724 4456 32770 4463
rect 32842 4639 33236 4651
rect 32842 4463 32848 4639
rect 32882 4626 33236 4639
rect 32882 4463 32888 4626
rect 33061 4624 33236 4626
rect 33061 4566 33103 4624
rect 33215 4566 33236 4624
rect 33061 4537 33236 4566
rect 32724 4451 32773 4456
rect 32842 4451 32888 4463
rect 32730 4290 32773 4451
rect 32647 4263 32773 4290
rect 32871 4376 33778 4392
rect 32871 4295 32887 4376
rect 32995 4295 33778 4376
rect 32871 4278 33778 4295
rect 32607 4251 32773 4263
rect 32613 4247 32773 4251
rect 32255 4213 32486 4219
rect 32255 4179 32436 4213
rect 32470 4179 32486 4213
rect 32255 4163 32486 4179
rect 32538 4213 32604 4219
rect 32538 4179 32554 4213
rect 32588 4179 32604 4213
rect 32538 4134 32604 4179
rect 32141 4126 32604 4134
rect 32141 4094 32605 4126
rect 32697 4110 32773 4247
rect 32693 4050 32703 4110
rect 32765 4050 32775 4110
rect 31615 4038 31922 4039
rect 30472 4033 30788 4038
rect 31502 4033 31922 4038
rect 30472 4022 30855 4033
rect 30472 3995 30804 4022
rect 30472 3866 30506 3995
rect 30788 3988 30804 3995
rect 30838 3988 30855 4022
rect 30788 3982 30855 3988
rect 31435 4022 31922 4033
rect 32701 4024 32771 4050
rect 31435 3988 31452 4022
rect 31486 3995 31922 4022
rect 31486 3988 31502 3995
rect 31615 3994 31922 3995
rect 31435 3982 31502 3988
rect 30613 3955 30669 3967
rect 30613 3921 30619 3955
rect 30653 3954 30669 3955
rect 31726 3954 31782 3966
rect 30653 3938 31120 3954
rect 30653 3921 31070 3938
rect 30613 3905 31070 3921
rect 31054 3904 31070 3905
rect 31104 3904 31120 3938
rect 31054 3897 31120 3904
rect 31172 3939 31742 3954
rect 31172 3905 31188 3939
rect 31222 3920 31742 3939
rect 31776 3920 31782 3954
rect 31222 3905 31782 3920
rect 31172 3895 31239 3905
rect 31726 3904 31782 3905
rect 31888 3866 31922 3994
rect 30466 3854 30512 3866
rect 30466 3678 30472 3854
rect 30506 3678 30512 3854
rect 30466 3666 30512 3678
rect 30584 3854 30630 3866
rect 30584 3678 30590 3854
rect 30624 3678 30630 3854
rect 30584 3666 30630 3678
rect 30886 3854 30932 3866
rect 30589 3372 30623 3666
rect 30886 3478 30892 3854
rect 30926 3478 30932 3854
rect 30886 3466 30932 3478
rect 31004 3854 31050 3866
rect 31004 3478 31010 3854
rect 31044 3478 31050 3854
rect 31004 3466 31050 3478
rect 31122 3854 31168 3866
rect 31122 3478 31128 3854
rect 31162 3478 31168 3854
rect 31122 3466 31168 3478
rect 31240 3854 31286 3866
rect 31240 3478 31246 3854
rect 31280 3478 31286 3854
rect 31240 3466 31286 3478
rect 31358 3854 31404 3866
rect 31358 3478 31364 3854
rect 31398 3478 31404 3854
rect 31764 3854 31810 3866
rect 31764 3678 31770 3854
rect 31804 3678 31810 3854
rect 31764 3666 31810 3678
rect 31882 3854 31928 3866
rect 31882 3678 31888 3854
rect 31922 3678 31928 3854
rect 31882 3666 31928 3678
rect 31358 3466 31404 3478
rect 31246 3372 31280 3466
rect 31770 3372 31803 3666
rect 30589 3340 31803 3372
rect 30955 3316 31361 3340
rect 30955 3193 31067 3316
rect 31241 3193 31361 3316
rect 30955 3149 31361 3193
rect 29241 2488 30023 2492
rect 28765 2476 28811 2488
rect 28370 2251 28703 2348
rect 28513 2208 28613 2220
rect 28513 2127 28524 2208
rect 28606 2127 28616 2208
rect 28513 2120 28613 2127
rect 28535 1971 28589 2120
rect 28649 2056 28703 2251
rect 28765 2100 28771 2476
rect 28805 2100 28811 2476
rect 28765 2088 28811 2100
rect 28883 2476 28929 2488
rect 28883 2100 28889 2476
rect 28923 2100 28929 2476
rect 28883 2088 28929 2100
rect 29001 2476 29047 2488
rect 29001 2100 29007 2476
rect 29041 2127 29047 2476
rect 29118 2476 29164 2488
rect 29118 2300 29124 2476
rect 29158 2300 29164 2476
rect 29118 2293 29164 2300
rect 29236 2476 30023 2488
rect 29236 2300 29242 2476
rect 29276 2463 30023 2476
rect 29276 2300 29282 2463
rect 29526 2381 30023 2463
rect 29118 2288 29167 2293
rect 29236 2288 29282 2300
rect 29124 2127 29167 2288
rect 29041 2100 29167 2127
rect 29001 2088 29167 2100
rect 29007 2084 29167 2088
rect 28649 2050 28880 2056
rect 28649 2016 28830 2050
rect 28864 2016 28880 2050
rect 28649 2000 28880 2016
rect 28932 2050 28998 2056
rect 28932 2016 28948 2050
rect 28982 2016 28998 2050
rect 28932 1971 28998 2016
rect 28535 1963 28998 1971
rect 28535 1931 28999 1963
rect 29091 1947 29167 2084
rect 29087 1887 29097 1947
rect 29159 1887 29169 1947
rect 30971 1726 31416 1732
rect 30971 1526 30983 1726
rect 31404 1526 31416 1726
rect 30971 1520 31139 1526
rect 31129 1452 31139 1520
rect 31271 1520 31416 1526
rect 31271 1452 31281 1520
rect 31139 1412 31271 1452
rect 31138 1346 31271 1412
rect 30467 1303 31940 1346
rect 30467 1000 30501 1303
rect 30833 1200 30867 1303
rect 31069 1200 31103 1303
rect 31305 1200 31339 1303
rect 31541 1200 31575 1303
rect 30827 1188 30873 1200
rect 30343 988 30389 1000
rect 30343 812 30349 988
rect 30383 812 30389 988
rect 30343 800 30389 812
rect 30461 988 30507 1000
rect 30461 812 30467 988
rect 30501 812 30507 988
rect 30461 800 30507 812
rect 30579 988 30625 1000
rect 30579 812 30585 988
rect 30619 812 30625 988
rect 30579 800 30625 812
rect 30697 988 30743 1000
rect 30827 988 30833 1188
rect 30697 812 30703 988
rect 30737 812 30833 988
rect 30867 812 30873 1188
rect 30697 800 30743 812
rect 30827 800 30873 812
rect 30945 1188 30991 1200
rect 30945 812 30951 1188
rect 30985 812 30991 1188
rect 30945 800 30991 812
rect 31063 1188 31109 1200
rect 31063 812 31069 1188
rect 31103 812 31109 1188
rect 31063 800 31109 812
rect 31181 1188 31227 1200
rect 31181 812 31187 1188
rect 31221 812 31227 1188
rect 31181 800 31227 812
rect 31299 1188 31345 1200
rect 31299 812 31305 1188
rect 31339 812 31345 1188
rect 31299 800 31345 812
rect 31417 1188 31463 1200
rect 31417 812 31423 1188
rect 31457 812 31463 1188
rect 31417 800 31463 812
rect 31535 1188 31581 1200
rect 31535 812 31541 1188
rect 31575 988 31581 1188
rect 31906 1000 31940 1303
rect 32447 1223 32583 1243
rect 32447 1161 32483 1223
rect 32543 1161 32583 1223
rect 32447 1133 32583 1161
rect 32143 1103 33120 1133
rect 31664 988 31710 1000
rect 31575 812 31670 988
rect 31704 812 31710 988
rect 31535 800 31581 812
rect 31664 800 31710 812
rect 31782 988 31828 1000
rect 31782 812 31788 988
rect 31822 812 31828 988
rect 31782 800 31828 812
rect 31900 988 31946 1000
rect 31900 812 31906 988
rect 31940 812 31946 988
rect 31900 800 31946 812
rect 32018 988 32064 1000
rect 32143 997 32175 1103
rect 32379 997 32411 1103
rect 32615 997 32647 1103
rect 32851 997 32883 1103
rect 33086 997 33120 1103
rect 32018 812 32024 988
rect 32058 812 32064 988
rect 32018 800 32064 812
rect 32136 985 32182 997
rect 32136 809 32142 985
rect 32176 809 32182 985
rect 30349 766 30383 800
rect 30951 766 30985 800
rect 31187 766 31221 800
rect 30349 731 30508 766
rect 30951 731 31221 766
rect 31788 766 31822 800
rect 32024 766 32058 800
rect 32136 797 32182 809
rect 32254 985 32300 997
rect 32254 809 32260 985
rect 32294 809 32300 985
rect 32254 797 32300 809
rect 32372 985 32418 997
rect 32372 809 32378 985
rect 32412 809 32418 985
rect 32372 797 32418 809
rect 32490 985 32536 997
rect 32490 809 32496 985
rect 32530 809 32536 985
rect 32490 797 32536 809
rect 32608 985 32654 997
rect 32608 809 32614 985
rect 32648 809 32654 985
rect 32608 797 32654 809
rect 32726 985 32772 997
rect 32726 809 32732 985
rect 32766 809 32772 985
rect 32726 797 32772 809
rect 32844 985 32890 997
rect 32844 809 32850 985
rect 32884 809 32890 985
rect 32844 797 32890 809
rect 32962 985 33008 997
rect 32962 809 32968 985
rect 33002 809 33008 985
rect 32962 797 33008 809
rect 33080 985 33126 997
rect 33080 809 33086 985
rect 33120 809 33126 985
rect 33080 797 33126 809
rect 33198 985 33244 997
rect 33198 809 33204 985
rect 33238 809 33244 985
rect 33198 797 33244 809
rect 31788 731 32058 766
rect 29718 583 30336 646
rect 30403 583 30413 646
rect 29718 582 30372 583
rect 28839 118 28975 138
rect 28839 56 28875 118
rect 28935 56 28975 118
rect 28839 28 28975 56
rect 28535 -2 29512 28
rect 28535 -108 28567 -2
rect 28771 -108 28803 -2
rect 29007 -108 29039 -2
rect 29243 -108 29275 -2
rect 29478 -108 29512 -2
rect 28528 -120 28574 -108
rect 28528 -296 28534 -120
rect 28568 -296 28574 -120
rect 28528 -308 28574 -296
rect 28646 -120 28692 -108
rect 28646 -296 28652 -120
rect 28686 -296 28692 -120
rect 28646 -308 28692 -296
rect 28764 -120 28810 -108
rect 28764 -296 28770 -120
rect 28804 -296 28810 -120
rect 28764 -308 28810 -296
rect 28882 -120 28928 -108
rect 28882 -296 28888 -120
rect 28922 -296 28928 -120
rect 28882 -308 28928 -296
rect 29000 -120 29046 -108
rect 29000 -296 29006 -120
rect 29040 -296 29046 -120
rect 29000 -308 29046 -296
rect 29118 -120 29164 -108
rect 29118 -296 29124 -120
rect 29158 -296 29164 -120
rect 29118 -308 29164 -296
rect 29236 -120 29282 -108
rect 29236 -296 29242 -120
rect 29276 -296 29282 -120
rect 29236 -308 29282 -296
rect 29354 -120 29400 -108
rect 29354 -296 29360 -120
rect 29394 -296 29400 -120
rect 29354 -308 29400 -296
rect 29472 -120 29518 -108
rect 29472 -296 29478 -120
rect 29512 -296 29518 -120
rect 29472 -308 29518 -296
rect 29590 -120 29636 -108
rect 29590 -296 29596 -120
rect 29630 -296 29636 -120
rect 29590 -308 29636 -296
rect 28651 -402 28687 -308
rect 28887 -402 28923 -308
rect 29123 -401 29159 -308
rect 29285 -356 29351 -349
rect 29285 -390 29301 -356
rect 29335 -390 29351 -356
rect 29285 -401 29351 -390
rect 29123 -402 29351 -401
rect 28651 -431 29351 -402
rect 28651 -432 29233 -431
rect 28771 -545 28805 -432
rect 29167 -473 29233 -432
rect 29167 -507 29183 -473
rect 29217 -507 29233 -473
rect 29167 -514 29233 -507
rect 29595 -541 29630 -308
rect 29718 -541 29809 582
rect 29241 -545 29809 -541
rect 28765 -557 28811 -545
rect 28625 -693 28725 -685
rect 28619 -780 28629 -693
rect 28718 -780 28728 -693
rect 28625 -785 28725 -780
rect 28220 -913 28589 -813
rect 22375 -1108 22385 -994
rect 22508 -1108 22518 -994
rect 28535 -1062 28589 -913
rect 28649 -977 28703 -785
rect 28765 -933 28771 -557
rect 28805 -933 28811 -557
rect 28765 -945 28811 -933
rect 28883 -557 28929 -545
rect 28883 -933 28889 -557
rect 28923 -933 28929 -557
rect 28883 -945 28929 -933
rect 29001 -557 29047 -545
rect 29001 -933 29007 -557
rect 29041 -906 29047 -557
rect 29118 -557 29164 -545
rect 29118 -733 29124 -557
rect 29158 -733 29164 -557
rect 29118 -740 29164 -733
rect 29236 -557 29809 -545
rect 29236 -733 29242 -557
rect 29276 -570 29809 -557
rect 29276 -733 29282 -570
rect 29526 -650 29809 -570
rect 29898 457 30336 520
rect 30403 457 30413 520
rect 29118 -745 29167 -740
rect 29236 -745 29282 -733
rect 29124 -906 29167 -745
rect 29041 -933 29167 -906
rect 29001 -945 29167 -933
rect 29007 -949 29167 -945
rect 28649 -983 28880 -977
rect 28649 -1017 28830 -983
rect 28864 -1017 28880 -983
rect 28649 -1033 28880 -1017
rect 28932 -983 28998 -977
rect 28932 -1017 28948 -983
rect 28982 -1017 28998 -983
rect 28932 -1062 28998 -1017
rect 28535 -1070 28998 -1062
rect 28535 -1102 28999 -1070
rect 29091 -1086 29167 -949
rect 29087 -1146 29097 -1086
rect 29159 -1146 29169 -1086
rect 28910 -1802 29046 -1782
rect 25675 -1853 25754 -1841
rect 23196 -1901 23275 -1889
rect 23196 -1998 23202 -1901
rect 23126 -2018 23202 -1998
rect 23269 -1998 23275 -1901
rect 25675 -1964 25681 -1853
rect 25748 -1964 25754 -1853
rect 26823 -1847 26902 -1835
rect 26823 -1964 26829 -1847
rect 26896 -1964 26902 -1847
rect 28910 -1864 28946 -1802
rect 29006 -1864 29046 -1802
rect 28910 -1892 29046 -1864
rect 28606 -1922 29583 -1892
rect 23269 -2018 23346 -1998
rect 23126 -2126 23170 -2018
rect 23302 -2126 23346 -2018
rect 24923 -2060 24979 -2052
rect 23126 -2168 23346 -2126
rect 23997 -2068 24979 -2060
rect 23997 -2102 24939 -2068
rect 24973 -2102 24979 -2068
rect 25642 -2072 25652 -1964
rect 25784 -2027 25794 -1964
rect 25784 -2038 25796 -2027
rect 25784 -2072 25797 -2038
rect 26053 -2048 26109 -2046
rect 23997 -2118 24979 -2102
rect 25652 -2110 25797 -2072
rect 23997 -2119 24976 -2118
rect 22730 -2198 23707 -2168
rect 22730 -2304 22762 -2198
rect 22966 -2304 22998 -2198
rect 23202 -2304 23234 -2198
rect 23438 -2304 23470 -2198
rect 23673 -2304 23707 -2198
rect 22723 -2316 22769 -2304
rect 22723 -2492 22729 -2316
rect 22763 -2492 22769 -2316
rect 22723 -2504 22769 -2492
rect 22841 -2316 22887 -2304
rect 22841 -2492 22847 -2316
rect 22881 -2492 22887 -2316
rect 22841 -2504 22887 -2492
rect 22959 -2316 23005 -2304
rect 22959 -2492 22965 -2316
rect 22999 -2492 23005 -2316
rect 22959 -2504 23005 -2492
rect 23077 -2316 23123 -2304
rect 23077 -2492 23083 -2316
rect 23117 -2492 23123 -2316
rect 23077 -2504 23123 -2492
rect 23195 -2316 23241 -2304
rect 23195 -2492 23201 -2316
rect 23235 -2492 23241 -2316
rect 23195 -2504 23241 -2492
rect 23313 -2316 23359 -2304
rect 23313 -2492 23319 -2316
rect 23353 -2492 23359 -2316
rect 23313 -2504 23359 -2492
rect 23431 -2316 23477 -2304
rect 23431 -2492 23437 -2316
rect 23471 -2492 23477 -2316
rect 23431 -2504 23477 -2492
rect 23549 -2316 23595 -2304
rect 23549 -2492 23555 -2316
rect 23589 -2492 23595 -2316
rect 23549 -2504 23595 -2492
rect 23667 -2316 23713 -2304
rect 23667 -2492 23673 -2316
rect 23707 -2492 23713 -2316
rect 23667 -2504 23713 -2492
rect 23785 -2316 23831 -2304
rect 23785 -2492 23791 -2316
rect 23825 -2492 23831 -2316
rect 23785 -2504 23831 -2492
rect 22846 -2598 22882 -2504
rect 23082 -2598 23118 -2504
rect 23318 -2597 23354 -2504
rect 23480 -2552 23546 -2545
rect 23480 -2586 23496 -2552
rect 23530 -2586 23546 -2552
rect 23480 -2597 23546 -2586
rect 23318 -2598 23546 -2597
rect 22846 -2627 23546 -2598
rect 22846 -2628 23428 -2627
rect 21497 -2798 21650 -2660
rect 22966 -2741 23000 -2628
rect 23362 -2669 23428 -2628
rect 23362 -2703 23378 -2669
rect 23412 -2703 23428 -2669
rect 23362 -2710 23428 -2703
rect 23790 -2709 23825 -2504
rect 23997 -2709 24064 -2119
rect 25756 -2142 25797 -2110
rect 26043 -2114 26053 -2048
rect 26109 -2114 26119 -2048
rect 26789 -2072 26799 -1964
rect 26931 -2027 26941 -1964
rect 26931 -2038 26943 -2027
rect 28606 -2028 28638 -1922
rect 28842 -2028 28874 -1922
rect 29078 -2028 29110 -1922
rect 29314 -2028 29346 -1922
rect 29549 -2028 29583 -1922
rect 26931 -2072 26944 -2038
rect 26799 -2110 26944 -2072
rect 26903 -2138 26944 -2110
rect 25172 -2170 25442 -2142
rect 24913 -2236 24923 -2170
rect 24989 -2236 24999 -2170
rect 25172 -2232 25206 -2170
rect 25408 -2232 25442 -2170
rect 25526 -2170 25797 -2142
rect 26314 -2166 26584 -2138
rect 25526 -2232 25560 -2170
rect 25762 -2232 25797 -2170
rect 25938 -2182 26109 -2166
rect 25938 -2216 26069 -2182
rect 26103 -2216 26109 -2182
rect 25938 -2232 26109 -2216
rect 26314 -2228 26348 -2166
rect 26550 -2228 26584 -2166
rect 26668 -2166 26944 -2138
rect 26668 -2228 26702 -2166
rect 26904 -2228 26944 -2166
rect 28599 -2040 28645 -2028
rect 28599 -2216 28605 -2040
rect 28639 -2216 28645 -2040
rect 28599 -2228 28645 -2216
rect 28717 -2040 28763 -2028
rect 28717 -2216 28723 -2040
rect 28757 -2216 28763 -2040
rect 28717 -2228 28763 -2216
rect 28835 -2040 28881 -2028
rect 28835 -2216 28841 -2040
rect 28875 -2216 28881 -2040
rect 28835 -2228 28881 -2216
rect 28953 -2040 28999 -2028
rect 28953 -2216 28959 -2040
rect 28993 -2216 28999 -2040
rect 28953 -2228 28999 -2216
rect 29071 -2040 29117 -2028
rect 29071 -2216 29077 -2040
rect 29111 -2216 29117 -2040
rect 29071 -2228 29117 -2216
rect 29189 -2040 29235 -2028
rect 29189 -2216 29195 -2040
rect 29229 -2216 29235 -2040
rect 29189 -2228 29235 -2216
rect 29307 -2040 29353 -2028
rect 29307 -2216 29313 -2040
rect 29347 -2216 29353 -2040
rect 29307 -2228 29353 -2216
rect 29425 -2040 29471 -2028
rect 29425 -2216 29431 -2040
rect 29465 -2216 29471 -2040
rect 29425 -2228 29471 -2216
rect 29543 -2040 29589 -2028
rect 29543 -2216 29549 -2040
rect 29583 -2216 29589 -2040
rect 29543 -2228 29589 -2216
rect 29661 -2040 29707 -2028
rect 29661 -2216 29667 -2040
rect 29701 -2216 29707 -2040
rect 29661 -2228 29707 -2216
rect 25048 -2244 25094 -2232
rect 25048 -2620 25054 -2244
rect 25088 -2620 25094 -2244
rect 25048 -2632 25094 -2620
rect 25166 -2244 25212 -2232
rect 25166 -2620 25172 -2244
rect 25206 -2620 25212 -2244
rect 25166 -2632 25212 -2620
rect 25284 -2244 25330 -2232
rect 25284 -2620 25290 -2244
rect 25324 -2620 25330 -2244
rect 25284 -2632 25330 -2620
rect 25402 -2244 25448 -2232
rect 25402 -2620 25408 -2244
rect 25442 -2620 25448 -2244
rect 25402 -2632 25448 -2620
rect 25520 -2244 25566 -2232
rect 25520 -2620 25526 -2244
rect 25560 -2620 25566 -2244
rect 25520 -2632 25566 -2620
rect 25638 -2244 25684 -2232
rect 25638 -2620 25644 -2244
rect 25678 -2620 25684 -2244
rect 25638 -2632 25684 -2620
rect 25756 -2244 25802 -2232
rect 25756 -2620 25762 -2244
rect 25796 -2620 25802 -2244
rect 25756 -2632 25802 -2620
rect 23790 -2737 24064 -2709
rect 23436 -2741 24064 -2737
rect 20282 -2866 20391 -2812
rect 19602 -2905 19829 -2869
rect 19602 -3012 19637 -2905
rect 19763 -2939 19829 -2905
rect 19763 -2973 19779 -2939
rect 19813 -2973 19829 -2939
rect 20110 -2881 20207 -2866
rect 20110 -2948 20167 -2881
rect 19763 -2979 19829 -2973
rect 20004 -2984 20273 -2948
rect 20004 -3012 20037 -2984
rect 20240 -3012 20273 -2984
rect 20357 -3012 20391 -2866
rect 21208 -2873 21218 -2798
rect 21286 -2873 21650 -2798
rect 21235 -2874 21650 -2873
rect 22960 -2753 23006 -2741
rect 19478 -3024 19524 -3012
rect 19478 -3200 19484 -3024
rect 19518 -3200 19524 -3024
rect 19478 -3212 19524 -3200
rect 19596 -3024 19642 -3012
rect 19596 -3200 19602 -3024
rect 19636 -3200 19642 -3024
rect 19596 -3212 19642 -3200
rect 19714 -3024 19760 -3012
rect 19714 -3200 19720 -3024
rect 19754 -3200 19760 -3024
rect 19714 -3212 19760 -3200
rect 19832 -3024 19878 -3012
rect 19832 -3200 19838 -3024
rect 19872 -3079 19878 -3024
rect 19997 -3024 20043 -3012
rect 19997 -3079 20003 -3024
rect 19872 -3167 20003 -3079
rect 19872 -3200 19878 -3167
rect 19832 -3212 19878 -3200
rect 19997 -3200 20003 -3167
rect 20037 -3200 20043 -3024
rect 19997 -3212 20043 -3200
rect 20115 -3024 20161 -3012
rect 20115 -3200 20121 -3024
rect 20155 -3200 20161 -3024
rect 20115 -3212 20161 -3200
rect 20233 -3024 20279 -3012
rect 20233 -3200 20239 -3024
rect 20273 -3200 20279 -3024
rect 20233 -3212 20279 -3200
rect 20351 -3024 20397 -3012
rect 20351 -3200 20357 -3024
rect 20391 -3200 20397 -3024
rect 22960 -3129 22966 -2753
rect 23000 -3129 23006 -2753
rect 22960 -3141 23006 -3129
rect 23078 -2753 23124 -2741
rect 23078 -3129 23084 -2753
rect 23118 -3129 23124 -2753
rect 23078 -3141 23124 -3129
rect 23196 -2753 23242 -2741
rect 23196 -3129 23202 -2753
rect 23236 -3105 23242 -2753
rect 23313 -2753 23359 -2741
rect 23313 -2929 23319 -2753
rect 23353 -2929 23359 -2753
rect 23313 -2941 23359 -2929
rect 23431 -2753 24064 -2741
rect 23431 -2929 23437 -2753
rect 23471 -2766 24064 -2753
rect 25054 -2674 25088 -2632
rect 25290 -2674 25324 -2632
rect 25054 -2702 25324 -2674
rect 25408 -2673 25442 -2632
rect 25644 -2673 25678 -2632
rect 25408 -2702 25678 -2673
rect 25054 -2750 25088 -2702
rect 23471 -2929 23477 -2766
rect 25054 -2780 25117 -2750
rect 23431 -2941 23477 -2929
rect 25082 -2872 25117 -2780
rect 25082 -2908 25309 -2872
rect 25579 -2883 25589 -2786
rect 25688 -2883 25698 -2786
rect 25762 -2815 25796 -2632
rect 25762 -2869 25871 -2815
rect 23319 -3057 23354 -2941
rect 25082 -3015 25117 -2908
rect 25243 -2942 25309 -2908
rect 25243 -2976 25259 -2942
rect 25293 -2976 25309 -2942
rect 25590 -2884 25687 -2883
rect 25590 -2951 25647 -2884
rect 25243 -2982 25309 -2976
rect 25484 -2987 25753 -2951
rect 25484 -3015 25517 -2987
rect 25720 -3015 25753 -2987
rect 25837 -3015 25871 -2869
rect 24958 -3027 25004 -3015
rect 23450 -3057 23558 -3047
rect 23319 -3105 23450 -3057
rect 23558 -3089 23703 -3083
rect 23236 -3129 23450 -3105
rect 23196 -3141 23450 -3129
rect 23202 -3145 23450 -3141
rect 20351 -3212 20397 -3200
rect 21267 -3146 22113 -3145
rect 21267 -3173 22838 -3146
rect 21267 -3179 23075 -3173
rect 19484 -3251 19518 -3212
rect 19720 -3251 19754 -3212
rect 19484 -3287 19754 -3251
rect 20121 -3250 20154 -3212
rect 20357 -3250 20390 -3212
rect 20121 -3286 20390 -3250
rect 21267 -3213 23025 -3179
rect 23059 -3213 23075 -3179
rect 21267 -3229 23075 -3213
rect 23127 -3179 23193 -3173
rect 23127 -3213 23143 -3179
rect 23177 -3213 23193 -3179
rect 23376 -3189 23450 -3145
rect 23691 -3156 23703 -3089
rect 23558 -3162 23703 -3156
rect 23450 -3199 23558 -3189
rect 21267 -3245 22838 -3229
rect 21267 -3246 22775 -3245
rect 21267 -3249 22310 -3246
rect 19484 -3288 19650 -3287
rect 19518 -3367 19650 -3288
rect 19508 -3475 19518 -3367
rect 19650 -3475 19660 -3367
rect 19542 -3603 19548 -3475
rect 19615 -3603 19621 -3475
rect 19542 -3615 19621 -3603
rect 16122 -3849 17099 -3819
rect 19316 -3821 19379 -3804
rect 19241 -3825 19379 -3821
rect 16122 -3955 16154 -3849
rect 16358 -3955 16390 -3849
rect 16594 -3955 16626 -3849
rect 16830 -3955 16862 -3849
rect 17065 -3955 17099 -3849
rect 17409 -3859 19379 -3825
rect 17407 -3888 19379 -3859
rect 17407 -3904 17453 -3888
rect 19241 -3890 19379 -3888
rect 16115 -3967 16161 -3955
rect 16115 -4143 16121 -3967
rect 16155 -4143 16161 -3967
rect 16115 -4155 16161 -4143
rect 16233 -3967 16279 -3955
rect 16233 -4143 16239 -3967
rect 16273 -4143 16279 -3967
rect 16233 -4155 16279 -4143
rect 16351 -3967 16397 -3955
rect 16351 -4143 16357 -3967
rect 16391 -4143 16397 -3967
rect 16351 -4155 16397 -4143
rect 16469 -3967 16515 -3955
rect 16469 -4143 16475 -3967
rect 16509 -4143 16515 -3967
rect 16469 -4155 16515 -4143
rect 16587 -3967 16633 -3955
rect 16587 -4143 16593 -3967
rect 16627 -4143 16633 -3967
rect 16587 -4155 16633 -4143
rect 16705 -3967 16751 -3955
rect 16705 -4143 16711 -3967
rect 16745 -4143 16751 -3967
rect 16705 -4155 16751 -4143
rect 16823 -3967 16869 -3955
rect 16823 -4143 16829 -3967
rect 16863 -4143 16869 -3967
rect 16823 -4155 16869 -4143
rect 16941 -3967 16987 -3955
rect 16941 -4143 16947 -3967
rect 16981 -4143 16987 -3967
rect 16941 -4155 16987 -4143
rect 17059 -3967 17105 -3955
rect 17059 -4143 17065 -3967
rect 17099 -4143 17105 -3967
rect 17059 -4155 17105 -4143
rect 17177 -3967 17223 -3955
rect 17177 -4143 17183 -3967
rect 17217 -4143 17223 -3967
rect 17177 -4155 17223 -4143
rect 16238 -4249 16274 -4155
rect 16474 -4249 16510 -4155
rect 16710 -4248 16746 -4155
rect 16872 -4203 16938 -4196
rect 16872 -4237 16888 -4203
rect 16922 -4237 16938 -4203
rect 16872 -4248 16938 -4237
rect 16710 -4249 16938 -4248
rect 16238 -4278 16938 -4249
rect 16238 -4279 16820 -4278
rect 16358 -4392 16392 -4279
rect 16754 -4320 16820 -4279
rect 16754 -4354 16770 -4320
rect 16804 -4354 16820 -4320
rect 16754 -4361 16820 -4354
rect 17182 -4373 17217 -4155
rect 17406 -4356 17453 -3904
rect 20303 -3894 20382 -3882
rect 20303 -4012 20309 -3894
rect 20376 -4012 20382 -3894
rect 18365 -4120 18375 -4012
rect 18507 -4120 18517 -4012
rect 20263 -4120 20273 -4012
rect 20405 -4120 20415 -4012
rect 18375 -4160 18507 -4120
rect 20273 -4160 20405 -4120
rect 18374 -4226 18507 -4160
rect 20272 -4226 20405 -4160
rect 17703 -4269 19176 -4226
rect 17406 -4372 17452 -4356
rect 17371 -4373 17452 -4372
rect 17182 -4388 17452 -4373
rect 16828 -4392 17452 -4388
rect 16352 -4404 16398 -4392
rect 16087 -4882 16097 -4764
rect 16215 -4796 16225 -4764
rect 16352 -4780 16358 -4404
rect 16392 -4780 16398 -4404
rect 16352 -4792 16398 -4780
rect 16470 -4404 16516 -4392
rect 16470 -4780 16476 -4404
rect 16510 -4780 16516 -4404
rect 16470 -4792 16516 -4780
rect 16588 -4404 16634 -4392
rect 16588 -4780 16594 -4404
rect 16628 -4756 16634 -4404
rect 16705 -4404 16751 -4392
rect 16705 -4580 16711 -4404
rect 16745 -4580 16751 -4404
rect 16705 -4592 16751 -4580
rect 16823 -4404 17452 -4392
rect 16823 -4580 16829 -4404
rect 16863 -4416 17452 -4404
rect 16863 -4417 17105 -4416
rect 16863 -4580 16869 -4417
rect 17371 -4418 17452 -4416
rect 17703 -4572 17737 -4269
rect 18069 -4372 18103 -4269
rect 18305 -4372 18339 -4269
rect 18541 -4372 18575 -4269
rect 18777 -4372 18811 -4269
rect 18063 -4384 18109 -4372
rect 16823 -4592 16869 -4580
rect 17579 -4584 17625 -4572
rect 16711 -4708 16746 -4592
rect 16842 -4708 16950 -4698
rect 16711 -4756 16842 -4708
rect 16950 -4745 17098 -4739
rect 16628 -4780 16842 -4756
rect 16588 -4792 16842 -4780
rect 16594 -4796 16842 -4792
rect 16215 -4824 16230 -4796
rect 16215 -4830 16467 -4824
rect 16215 -4864 16417 -4830
rect 16451 -4864 16467 -4830
rect 16215 -4880 16467 -4864
rect 16519 -4830 16585 -4824
rect 16519 -4864 16535 -4830
rect 16569 -4864 16585 -4830
rect 16768 -4840 16842 -4796
rect 17086 -4812 17098 -4745
rect 17579 -4760 17585 -4584
rect 17619 -4760 17625 -4584
rect 17579 -4772 17625 -4760
rect 17697 -4584 17743 -4572
rect 17697 -4760 17703 -4584
rect 17737 -4760 17743 -4584
rect 17697 -4772 17743 -4760
rect 17815 -4584 17861 -4572
rect 17815 -4760 17821 -4584
rect 17855 -4760 17861 -4584
rect 17815 -4772 17861 -4760
rect 17933 -4584 17979 -4572
rect 18063 -4584 18069 -4384
rect 17933 -4760 17939 -4584
rect 17973 -4760 18069 -4584
rect 18103 -4760 18109 -4384
rect 17933 -4772 17979 -4760
rect 18063 -4772 18109 -4760
rect 18181 -4384 18227 -4372
rect 18181 -4760 18187 -4384
rect 18221 -4760 18227 -4384
rect 18181 -4772 18227 -4760
rect 18299 -4384 18345 -4372
rect 18299 -4760 18305 -4384
rect 18339 -4760 18345 -4384
rect 18299 -4772 18345 -4760
rect 18417 -4384 18463 -4372
rect 18417 -4760 18423 -4384
rect 18457 -4760 18463 -4384
rect 18417 -4772 18463 -4760
rect 18535 -4384 18581 -4372
rect 18535 -4760 18541 -4384
rect 18575 -4760 18581 -4384
rect 18535 -4772 18581 -4760
rect 18653 -4384 18699 -4372
rect 18653 -4760 18659 -4384
rect 18693 -4760 18699 -4384
rect 18653 -4772 18699 -4760
rect 18771 -4384 18817 -4372
rect 18771 -4760 18777 -4384
rect 18811 -4584 18817 -4384
rect 19142 -4572 19176 -4269
rect 19601 -4269 21074 -4226
rect 19601 -4572 19635 -4269
rect 19967 -4372 20001 -4269
rect 20203 -4372 20237 -4269
rect 20439 -4372 20473 -4269
rect 20675 -4372 20709 -4269
rect 19961 -4384 20007 -4372
rect 18900 -4584 18946 -4572
rect 18811 -4760 18906 -4584
rect 18940 -4760 18946 -4584
rect 18771 -4772 18817 -4760
rect 18900 -4772 18946 -4760
rect 19018 -4584 19064 -4572
rect 19018 -4760 19024 -4584
rect 19058 -4760 19064 -4584
rect 19018 -4772 19064 -4760
rect 19136 -4584 19182 -4572
rect 19136 -4760 19142 -4584
rect 19176 -4760 19182 -4584
rect 19136 -4772 19182 -4760
rect 19254 -4584 19300 -4572
rect 19254 -4760 19260 -4584
rect 19294 -4760 19300 -4584
rect 19254 -4772 19300 -4760
rect 19477 -4584 19523 -4572
rect 19477 -4760 19483 -4584
rect 19517 -4760 19523 -4584
rect 19477 -4772 19523 -4760
rect 19595 -4584 19641 -4572
rect 19595 -4760 19601 -4584
rect 19635 -4760 19641 -4584
rect 19595 -4772 19641 -4760
rect 19713 -4584 19759 -4572
rect 19713 -4760 19719 -4584
rect 19753 -4760 19759 -4584
rect 19713 -4772 19759 -4760
rect 19831 -4584 19877 -4572
rect 19961 -4584 19967 -4384
rect 19831 -4760 19837 -4584
rect 19871 -4760 19967 -4584
rect 20001 -4760 20007 -4384
rect 19831 -4772 19877 -4760
rect 19961 -4772 20007 -4760
rect 20079 -4384 20125 -4372
rect 20079 -4760 20085 -4384
rect 20119 -4760 20125 -4384
rect 20079 -4772 20125 -4760
rect 20197 -4384 20243 -4372
rect 20197 -4760 20203 -4384
rect 20237 -4760 20243 -4384
rect 20197 -4772 20243 -4760
rect 20315 -4384 20361 -4372
rect 20315 -4760 20321 -4384
rect 20355 -4760 20361 -4384
rect 20315 -4772 20361 -4760
rect 20433 -4384 20479 -4372
rect 20433 -4760 20439 -4384
rect 20473 -4760 20479 -4384
rect 20433 -4772 20479 -4760
rect 20551 -4384 20597 -4372
rect 20551 -4760 20557 -4384
rect 20591 -4760 20597 -4384
rect 20551 -4772 20597 -4760
rect 20669 -4384 20715 -4372
rect 20669 -4760 20675 -4384
rect 20709 -4584 20715 -4384
rect 21040 -4572 21074 -4269
rect 20798 -4584 20844 -4572
rect 20709 -4760 20804 -4584
rect 20838 -4760 20844 -4584
rect 20669 -4772 20715 -4760
rect 20798 -4772 20844 -4760
rect 20916 -4584 20962 -4572
rect 20916 -4760 20922 -4584
rect 20956 -4760 20962 -4584
rect 20916 -4772 20962 -4760
rect 21034 -4584 21080 -4572
rect 21034 -4760 21040 -4584
rect 21074 -4760 21080 -4584
rect 21034 -4772 21080 -4760
rect 21152 -4584 21198 -4572
rect 21152 -4760 21158 -4584
rect 21192 -4760 21198 -4584
rect 21152 -4772 21198 -4760
rect 16950 -4818 17098 -4812
rect 17585 -4806 17619 -4772
rect 18187 -4806 18221 -4772
rect 18423 -4806 18457 -4772
rect 16842 -4850 16950 -4840
rect 17585 -4841 17744 -4806
rect 18187 -4841 18457 -4806
rect 19024 -4806 19058 -4772
rect 19260 -4806 19294 -4772
rect 19024 -4841 19294 -4806
rect 19483 -4806 19517 -4772
rect 20085 -4806 20119 -4772
rect 20321 -4806 20355 -4772
rect 19483 -4841 19642 -4806
rect 20085 -4841 20355 -4806
rect 20922 -4806 20956 -4772
rect 21158 -4806 21192 -4772
rect 20922 -4841 21192 -4806
rect 16215 -4882 16230 -4880
rect 16130 -4896 16230 -4882
rect 16130 -4939 16230 -4938
rect 15751 -4960 16230 -4939
rect 16519 -4960 16585 -4864
rect 15751 -5008 16585 -4960
rect 15751 -5037 16230 -5008
rect 15751 -5039 15856 -5037
rect 16130 -5038 16230 -5037
rect 15584 -5224 15594 -5145
rect 15687 -5224 15697 -5145
rect 16587 -5160 16666 -5148
rect 15595 -6398 15688 -5224
rect 16587 -5253 16593 -5160
rect 16513 -5273 16593 -5253
rect 16660 -5253 16666 -5160
rect 16660 -5273 16733 -5253
rect 16513 -5381 16557 -5273
rect 16689 -5381 16733 -5273
rect 16513 -5423 16733 -5381
rect 16117 -5453 17094 -5423
rect 16117 -5559 16149 -5453
rect 16353 -5559 16385 -5453
rect 16589 -5559 16621 -5453
rect 16825 -5559 16857 -5453
rect 17060 -5559 17094 -5453
rect 16110 -5571 16156 -5559
rect 16110 -5747 16116 -5571
rect 16150 -5747 16156 -5571
rect 16110 -5759 16156 -5747
rect 16228 -5571 16274 -5559
rect 16228 -5747 16234 -5571
rect 16268 -5747 16274 -5571
rect 16228 -5759 16274 -5747
rect 16346 -5571 16392 -5559
rect 16346 -5747 16352 -5571
rect 16386 -5747 16392 -5571
rect 16346 -5759 16392 -5747
rect 16464 -5571 16510 -5559
rect 16464 -5747 16470 -5571
rect 16504 -5747 16510 -5571
rect 16464 -5759 16510 -5747
rect 16582 -5571 16628 -5559
rect 16582 -5747 16588 -5571
rect 16622 -5747 16628 -5571
rect 16582 -5759 16628 -5747
rect 16700 -5571 16746 -5559
rect 16700 -5747 16706 -5571
rect 16740 -5747 16746 -5571
rect 16700 -5759 16746 -5747
rect 16818 -5571 16864 -5559
rect 16818 -5747 16824 -5571
rect 16858 -5747 16864 -5571
rect 16818 -5759 16864 -5747
rect 16936 -5571 16982 -5559
rect 16936 -5747 16942 -5571
rect 16976 -5747 16982 -5571
rect 16936 -5759 16982 -5747
rect 17054 -5571 17100 -5559
rect 17054 -5747 17060 -5571
rect 17094 -5747 17100 -5571
rect 17054 -5759 17100 -5747
rect 17172 -5571 17218 -5559
rect 17172 -5747 17178 -5571
rect 17212 -5747 17218 -5571
rect 17172 -5759 17218 -5747
rect 17710 -5625 17744 -4841
rect 18423 -4903 18457 -4841
rect 18012 -4941 18754 -4903
rect 18012 -5065 18046 -4941
rect 18248 -5065 18282 -4941
rect 18484 -5065 18518 -4941
rect 18720 -5065 18754 -4941
rect 19010 -5048 19020 -4982
rect 19083 -5048 19093 -4982
rect 18006 -5077 18052 -5065
rect 18006 -5453 18012 -5077
rect 18046 -5453 18052 -5077
rect 18006 -5465 18052 -5453
rect 18124 -5077 18170 -5065
rect 18124 -5453 18130 -5077
rect 18164 -5453 18170 -5077
rect 18124 -5465 18170 -5453
rect 18242 -5077 18288 -5065
rect 18242 -5453 18248 -5077
rect 18282 -5453 18288 -5077
rect 18242 -5465 18288 -5453
rect 18360 -5077 18406 -5065
rect 18360 -5453 18366 -5077
rect 18400 -5453 18406 -5077
rect 18360 -5465 18406 -5453
rect 18478 -5077 18524 -5065
rect 18478 -5453 18484 -5077
rect 18518 -5453 18524 -5077
rect 18478 -5465 18524 -5453
rect 18596 -5077 18642 -5065
rect 18596 -5453 18602 -5077
rect 18636 -5453 18642 -5077
rect 18596 -5465 18642 -5453
rect 18714 -5077 18760 -5065
rect 18714 -5453 18720 -5077
rect 18754 -5453 18760 -5077
rect 18714 -5465 18760 -5453
rect 19126 -5624 19160 -4841
rect 18853 -5625 19160 -5624
rect 17710 -5630 18026 -5625
rect 18740 -5630 19160 -5625
rect 17710 -5641 18093 -5630
rect 17710 -5668 18042 -5641
rect 16233 -5853 16269 -5759
rect 16469 -5853 16505 -5759
rect 16705 -5852 16741 -5759
rect 16867 -5807 16933 -5800
rect 16867 -5841 16883 -5807
rect 16917 -5841 16933 -5807
rect 16867 -5852 16933 -5841
rect 16705 -5853 16933 -5852
rect 16233 -5882 16933 -5853
rect 16233 -5883 16815 -5882
rect 16353 -5996 16387 -5883
rect 16749 -5924 16815 -5883
rect 16749 -5958 16765 -5924
rect 16799 -5958 16815 -5924
rect 16749 -5965 16815 -5958
rect 17177 -5992 17212 -5759
rect 17710 -5797 17744 -5668
rect 18026 -5675 18042 -5668
rect 18076 -5675 18093 -5641
rect 18026 -5681 18093 -5675
rect 18673 -5641 19160 -5630
rect 18673 -5675 18690 -5641
rect 18724 -5668 19160 -5641
rect 18724 -5675 18740 -5668
rect 18853 -5669 19160 -5668
rect 18673 -5681 18740 -5675
rect 17851 -5708 17907 -5696
rect 17851 -5742 17857 -5708
rect 17891 -5709 17907 -5708
rect 18964 -5709 19020 -5697
rect 17891 -5725 18358 -5709
rect 17891 -5742 18308 -5725
rect 17851 -5758 18308 -5742
rect 18292 -5759 18308 -5758
rect 18342 -5759 18358 -5725
rect 18292 -5766 18358 -5759
rect 18410 -5724 18980 -5709
rect 18410 -5758 18426 -5724
rect 18460 -5743 18980 -5724
rect 19014 -5743 19020 -5709
rect 18460 -5758 19020 -5743
rect 18410 -5768 18477 -5758
rect 18964 -5759 19020 -5758
rect 19126 -5797 19160 -5669
rect 19608 -5625 19642 -4841
rect 20321 -4903 20355 -4841
rect 19910 -4941 20652 -4903
rect 19910 -5065 19944 -4941
rect 20146 -5065 20180 -4941
rect 20382 -5065 20416 -4941
rect 20618 -5065 20652 -4941
rect 19904 -5077 19950 -5065
rect 19904 -5453 19910 -5077
rect 19944 -5453 19950 -5077
rect 19904 -5465 19950 -5453
rect 20022 -5077 20068 -5065
rect 20022 -5453 20028 -5077
rect 20062 -5453 20068 -5077
rect 20022 -5465 20068 -5453
rect 20140 -5077 20186 -5065
rect 20140 -5453 20146 -5077
rect 20180 -5453 20186 -5077
rect 20140 -5465 20186 -5453
rect 20258 -5077 20304 -5065
rect 20258 -5453 20264 -5077
rect 20298 -5453 20304 -5077
rect 20258 -5465 20304 -5453
rect 20376 -5077 20422 -5065
rect 20376 -5453 20382 -5077
rect 20416 -5453 20422 -5077
rect 20376 -5465 20422 -5453
rect 20494 -5077 20540 -5065
rect 20494 -5453 20500 -5077
rect 20534 -5453 20540 -5077
rect 20494 -5465 20540 -5453
rect 20612 -5077 20658 -5065
rect 20612 -5453 20618 -5077
rect 20652 -5453 20658 -5077
rect 20612 -5465 20658 -5453
rect 21024 -5624 21058 -4841
rect 20636 -5625 20705 -5624
rect 20751 -5625 21058 -5624
rect 19608 -5630 19924 -5625
rect 20636 -5629 21058 -5625
rect 19608 -5641 19991 -5630
rect 19608 -5668 19940 -5641
rect 19608 -5797 19642 -5668
rect 19924 -5675 19940 -5668
rect 19974 -5675 19991 -5641
rect 19924 -5681 19991 -5675
rect 20569 -5640 21058 -5629
rect 20569 -5674 20586 -5640
rect 20620 -5668 21058 -5640
rect 20620 -5674 20636 -5668
rect 20751 -5669 21058 -5668
rect 20569 -5680 20636 -5674
rect 19749 -5708 19805 -5696
rect 19749 -5742 19755 -5708
rect 19789 -5709 19805 -5708
rect 20862 -5709 20918 -5697
rect 19789 -5725 20256 -5709
rect 19789 -5742 20206 -5725
rect 19749 -5758 20206 -5742
rect 20190 -5759 20206 -5758
rect 20240 -5759 20256 -5725
rect 20190 -5766 20256 -5759
rect 20308 -5724 20878 -5709
rect 20308 -5758 20324 -5724
rect 20358 -5743 20878 -5724
rect 20912 -5743 20918 -5709
rect 20358 -5758 20918 -5743
rect 20308 -5768 20375 -5758
rect 20862 -5759 20918 -5758
rect 21024 -5797 21058 -5669
rect 21139 -5019 21206 -4995
rect 21139 -5053 21156 -5019
rect 21190 -5053 21206 -5019
rect 16823 -5996 17212 -5992
rect 16347 -6008 16393 -5996
rect 16347 -6384 16353 -6008
rect 16387 -6384 16393 -6008
rect 16347 -6396 16393 -6384
rect 16465 -6008 16511 -5996
rect 16465 -6384 16471 -6008
rect 16505 -6384 16511 -6008
rect 16465 -6396 16511 -6384
rect 16583 -6008 16629 -5996
rect 16583 -6384 16589 -6008
rect 16623 -6360 16629 -6008
rect 16700 -6008 16746 -5996
rect 16700 -6184 16706 -6008
rect 16740 -6184 16746 -6008
rect 16700 -6196 16746 -6184
rect 16818 -6008 17212 -5996
rect 17704 -5809 17750 -5797
rect 17704 -5985 17710 -5809
rect 17744 -5985 17750 -5809
rect 17704 -5997 17750 -5985
rect 17822 -5809 17868 -5797
rect 17822 -5985 17828 -5809
rect 17862 -5985 17868 -5809
rect 17822 -5997 17868 -5985
rect 18124 -5809 18170 -5797
rect 16818 -6184 16824 -6008
rect 16858 -6021 17212 -6008
rect 16858 -6184 16864 -6021
rect 17134 -6024 17212 -6021
rect 17134 -6076 17144 -6024
rect 17207 -6076 17217 -6024
rect 17139 -6082 17212 -6076
rect 16818 -6196 16864 -6184
rect 16706 -6312 16741 -6196
rect 17827 -6291 17861 -5997
rect 18124 -6185 18130 -5809
rect 18164 -6185 18170 -5809
rect 18124 -6197 18170 -6185
rect 18242 -5809 18288 -5797
rect 18242 -6185 18248 -5809
rect 18282 -6185 18288 -5809
rect 18242 -6197 18288 -6185
rect 18360 -5809 18406 -5797
rect 18360 -6185 18366 -5809
rect 18400 -6185 18406 -5809
rect 18360 -6197 18406 -6185
rect 18478 -5809 18524 -5797
rect 18478 -6185 18484 -5809
rect 18518 -6185 18524 -5809
rect 18478 -6197 18524 -6185
rect 18596 -5809 18642 -5797
rect 18596 -6185 18602 -5809
rect 18636 -6185 18642 -5809
rect 19002 -5809 19048 -5797
rect 19002 -5985 19008 -5809
rect 19042 -5985 19048 -5809
rect 19002 -5997 19048 -5985
rect 19120 -5809 19166 -5797
rect 19120 -5985 19126 -5809
rect 19160 -5985 19166 -5809
rect 19120 -5997 19166 -5985
rect 19602 -5809 19648 -5797
rect 19602 -5985 19608 -5809
rect 19642 -5985 19648 -5809
rect 19602 -5997 19648 -5985
rect 19720 -5809 19766 -5797
rect 19720 -5985 19726 -5809
rect 19760 -5985 19766 -5809
rect 19720 -5997 19766 -5985
rect 20022 -5809 20068 -5797
rect 18596 -6197 18642 -6185
rect 18484 -6291 18518 -6197
rect 19008 -6291 19041 -5997
rect 16837 -6312 16945 -6302
rect 16706 -6360 16837 -6312
rect 17827 -6323 19041 -6291
rect 19725 -6291 19759 -5997
rect 20022 -6185 20028 -5809
rect 20062 -6185 20068 -5809
rect 20022 -6197 20068 -6185
rect 20140 -5809 20186 -5797
rect 20140 -6185 20146 -5809
rect 20180 -6185 20186 -5809
rect 20140 -6197 20186 -6185
rect 20258 -5809 20304 -5797
rect 20258 -6185 20264 -5809
rect 20298 -6185 20304 -5809
rect 20258 -6197 20304 -6185
rect 20376 -5809 20422 -5797
rect 20376 -6185 20382 -5809
rect 20416 -6185 20422 -5809
rect 20376 -6197 20422 -6185
rect 20494 -5809 20540 -5797
rect 20494 -6185 20500 -5809
rect 20534 -6185 20540 -5809
rect 20900 -5809 20946 -5797
rect 20900 -5985 20906 -5809
rect 20940 -5985 20946 -5809
rect 20900 -5997 20946 -5985
rect 21018 -5809 21064 -5797
rect 21018 -5985 21024 -5809
rect 21058 -5985 21064 -5809
rect 21018 -5997 21064 -5985
rect 20494 -6197 20540 -6185
rect 20382 -6291 20416 -6197
rect 20906 -6291 20939 -5997
rect 19725 -6323 20939 -6291
rect 16945 -6354 17101 -6348
rect 16623 -6384 16837 -6360
rect 16583 -6396 16837 -6384
rect 15595 -6400 16180 -6398
rect 16589 -6400 16837 -6396
rect 15595 -6428 16225 -6400
rect 15595 -6434 16462 -6428
rect 15595 -6468 16412 -6434
rect 16446 -6468 16462 -6434
rect 15595 -6484 16462 -6468
rect 16514 -6434 16580 -6428
rect 16514 -6468 16530 -6434
rect 16564 -6468 16580 -6434
rect 16763 -6444 16837 -6400
rect 17089 -6421 17101 -6354
rect 18320 -6408 18452 -6323
rect 20218 -6408 20350 -6323
rect 16945 -6427 17101 -6421
rect 16837 -6454 16945 -6444
rect 15595 -6500 16225 -6484
rect 15595 -6504 16180 -6500
rect 15595 -6505 15696 -6504
rect 16125 -6553 16225 -6542
rect 15255 -6591 15423 -6572
rect 15255 -6678 15282 -6591
rect 15384 -6678 15423 -6591
rect 16089 -6659 16099 -6553
rect 16211 -6564 16225 -6553
rect 16514 -6564 16580 -6468
rect 18310 -6516 18320 -6408
rect 18452 -6516 18462 -6408
rect 20208 -6516 20218 -6408
rect 20350 -6516 20360 -6408
rect 21139 -6436 21206 -5053
rect 21267 -5482 21423 -3249
rect 22108 -3250 22310 -3249
rect 21267 -5580 21279 -5482
rect 21411 -5580 21423 -5482
rect 21267 -5586 21423 -5580
rect 21550 -3661 22094 -3634
rect 21550 -3767 21942 -3661
rect 22054 -3674 22094 -3661
rect 22054 -3767 22096 -3674
rect 21550 -3778 22096 -3767
rect 21550 -3779 22094 -3778
rect 16211 -6612 16580 -6564
rect 16211 -6642 16225 -6612
rect 16211 -6659 16221 -6642
rect 15255 -6684 15423 -6678
rect 16513 -6715 16579 -6612
rect 18336 -6656 18342 -6516
rect 18409 -6656 18415 -6516
rect 18336 -6668 18415 -6656
rect 21139 -6715 21205 -6436
rect 16511 -6795 21205 -6715
rect 19922 -7306 20386 -7274
rect 20474 -7290 20484 -7230
rect 20546 -7290 20556 -7230
rect 19922 -7314 20385 -7306
rect 19922 -7462 19976 -7314
rect 14264 -7794 15027 -7714
rect 14014 -7807 15027 -7794
rect 13974 -7819 15027 -7807
rect 13509 -7932 13543 -7819
rect 13979 -7823 15027 -7819
rect 14329 -7824 15027 -7823
rect 19611 -7563 19976 -7462
rect 20036 -7359 20267 -7343
rect 20036 -7393 20217 -7359
rect 20251 -7393 20267 -7359
rect 20036 -7399 20267 -7393
rect 20319 -7359 20385 -7314
rect 20319 -7393 20335 -7359
rect 20369 -7393 20385 -7359
rect 20319 -7399 20385 -7393
rect 13905 -7857 13971 -7850
rect 13905 -7891 13921 -7857
rect 13955 -7891 13971 -7857
rect 13905 -7932 13971 -7891
rect 13389 -7933 13971 -7932
rect 13389 -7962 14089 -7933
rect 13389 -8056 13425 -7962
rect 13625 -8056 13661 -7962
rect 13861 -7963 14089 -7962
rect 13861 -8056 13897 -7963
rect 14023 -7974 14089 -7963
rect 14023 -8008 14039 -7974
rect 14073 -8008 14089 -7974
rect 14023 -8015 14089 -8008
rect 14333 -8056 14368 -7824
rect 13266 -8068 13312 -8056
rect 13266 -8244 13272 -8068
rect 13306 -8244 13312 -8068
rect 13266 -8256 13312 -8244
rect 13384 -8068 13430 -8056
rect 13384 -8244 13390 -8068
rect 13424 -8244 13430 -8068
rect 13384 -8256 13430 -8244
rect 13502 -8068 13548 -8056
rect 13502 -8244 13508 -8068
rect 13542 -8244 13548 -8068
rect 13502 -8256 13548 -8244
rect 13620 -8068 13666 -8056
rect 13620 -8244 13626 -8068
rect 13660 -8244 13666 -8068
rect 13620 -8256 13666 -8244
rect 13738 -8068 13784 -8056
rect 13738 -8244 13744 -8068
rect 13778 -8244 13784 -8068
rect 13738 -8256 13784 -8244
rect 13856 -8068 13902 -8056
rect 13856 -8244 13862 -8068
rect 13896 -8244 13902 -8068
rect 13856 -8256 13902 -8244
rect 13974 -8068 14020 -8056
rect 13974 -8244 13980 -8068
rect 14014 -8244 14020 -8068
rect 13974 -8256 14020 -8244
rect 14092 -8068 14138 -8056
rect 14092 -8244 14098 -8068
rect 14132 -8244 14138 -8068
rect 14092 -8256 14138 -8244
rect 14210 -8068 14256 -8056
rect 14210 -8244 14216 -8068
rect 14250 -8244 14256 -8068
rect 14210 -8256 14256 -8244
rect 14328 -8068 14374 -8056
rect 14328 -8244 14334 -8068
rect 14368 -8244 14374 -8068
rect 14328 -8256 14374 -8244
rect 13273 -8362 13305 -8256
rect 13509 -8362 13541 -8256
rect 13745 -8362 13777 -8256
rect 13981 -8362 14013 -8256
rect 14216 -8362 14250 -8256
rect 13273 -8392 14250 -8362
rect 13577 -8420 13713 -8392
rect 13577 -8482 13613 -8420
rect 13673 -8482 13713 -8420
rect 13577 -8502 13713 -8482
rect 19611 -8592 19697 -7563
rect 20036 -7591 20090 -7399
rect 20478 -7427 20554 -7290
rect 20394 -7431 20554 -7427
rect 19765 -7598 20090 -7591
rect 19760 -7687 19770 -7598
rect 19839 -7687 20090 -7598
rect 19765 -7691 20090 -7687
rect 20152 -7443 20198 -7431
rect 20152 -7819 20158 -7443
rect 20192 -7819 20198 -7443
rect 20152 -7831 20198 -7819
rect 20270 -7443 20316 -7431
rect 20270 -7819 20276 -7443
rect 20310 -7819 20316 -7443
rect 20270 -7831 20316 -7819
rect 20388 -7443 20554 -7431
rect 20388 -7819 20394 -7443
rect 20428 -7470 20554 -7443
rect 20428 -7819 20434 -7470
rect 20511 -7631 20554 -7470
rect 20388 -7831 20434 -7819
rect 20505 -7636 20554 -7631
rect 20505 -7643 20551 -7636
rect 20505 -7819 20511 -7643
rect 20545 -7819 20551 -7643
rect 20505 -7831 20551 -7819
rect 20623 -7643 20669 -7631
rect 20623 -7819 20629 -7643
rect 20663 -7806 20669 -7643
rect 21550 -7726 21706 -3779
rect 21806 -4773 22093 -4744
rect 21806 -4879 21941 -4773
rect 22053 -4775 22093 -4773
rect 22059 -4786 22093 -4775
rect 21806 -4881 21947 -4879
rect 22059 -4881 22094 -4786
rect 21806 -4890 22094 -4881
rect 21806 -4891 22093 -4890
rect 21806 -4892 22061 -4891
rect 21809 -7229 21961 -4892
rect 22217 -5144 22310 -3250
rect 22373 -3309 22839 -3287
rect 23127 -3309 23193 -3213
rect 24958 -3203 24964 -3027
rect 24998 -3203 25004 -3027
rect 24958 -3215 25004 -3203
rect 25076 -3027 25122 -3015
rect 25076 -3203 25082 -3027
rect 25116 -3203 25122 -3027
rect 25076 -3215 25122 -3203
rect 25194 -3027 25240 -3015
rect 25194 -3203 25200 -3027
rect 25234 -3203 25240 -3027
rect 25194 -3215 25240 -3203
rect 25312 -3027 25358 -3015
rect 25312 -3203 25318 -3027
rect 25352 -3082 25358 -3027
rect 25477 -3027 25523 -3015
rect 25477 -3082 25483 -3027
rect 25352 -3170 25483 -3082
rect 25352 -3203 25358 -3170
rect 25312 -3215 25358 -3203
rect 25477 -3203 25483 -3170
rect 25517 -3203 25523 -3027
rect 25477 -3215 25523 -3203
rect 25595 -3027 25641 -3015
rect 25595 -3203 25601 -3027
rect 25635 -3203 25641 -3027
rect 25595 -3215 25641 -3203
rect 25713 -3027 25759 -3015
rect 25713 -3203 25719 -3027
rect 25753 -3203 25759 -3027
rect 25713 -3215 25759 -3203
rect 25831 -3027 25877 -3015
rect 25831 -3203 25837 -3027
rect 25871 -3203 25877 -3027
rect 25831 -3215 25877 -3203
rect 24964 -3254 24998 -3215
rect 25200 -3254 25234 -3215
rect 24964 -3289 25234 -3254
rect 25601 -3253 25634 -3215
rect 25837 -3253 25870 -3215
rect 25601 -3289 25870 -3253
rect 22373 -3357 23193 -3309
rect 24998 -3290 25234 -3289
rect 22373 -3388 22839 -3357
rect 24998 -3364 25130 -3290
rect 22373 -3644 22478 -3388
rect 24988 -3472 24998 -3364
rect 25130 -3472 25140 -3364
rect 23211 -3551 23290 -3539
rect 22373 -3750 22436 -3644
rect 22548 -3750 22558 -3644
rect 23211 -3648 23217 -3551
rect 23140 -3668 23217 -3648
rect 23284 -3648 23290 -3551
rect 25027 -3602 25033 -3472
rect 25100 -3602 25106 -3472
rect 25027 -3614 25106 -3602
rect 23284 -3668 23360 -3648
rect 22373 -3761 22522 -3750
rect 22373 -4938 22478 -3761
rect 23140 -3776 23184 -3668
rect 23316 -3776 23360 -3668
rect 23140 -3818 23360 -3776
rect 25938 -3803 26000 -2232
rect 26190 -2240 26236 -2228
rect 26190 -2616 26196 -2240
rect 26230 -2616 26236 -2240
rect 26190 -2628 26236 -2616
rect 26308 -2240 26354 -2228
rect 26308 -2616 26314 -2240
rect 26348 -2616 26354 -2240
rect 26308 -2628 26354 -2616
rect 26426 -2240 26472 -2228
rect 26426 -2616 26432 -2240
rect 26466 -2616 26472 -2240
rect 26426 -2628 26472 -2616
rect 26544 -2240 26590 -2228
rect 26544 -2616 26550 -2240
rect 26584 -2616 26590 -2240
rect 26544 -2628 26590 -2616
rect 26662 -2240 26708 -2228
rect 26662 -2616 26668 -2240
rect 26702 -2616 26708 -2240
rect 26662 -2628 26708 -2616
rect 26780 -2240 26826 -2228
rect 26780 -2616 26786 -2240
rect 26820 -2616 26826 -2240
rect 26780 -2628 26826 -2616
rect 26898 -2240 26944 -2228
rect 26898 -2616 26904 -2240
rect 26938 -2616 26944 -2240
rect 28722 -2322 28758 -2228
rect 28958 -2322 28994 -2228
rect 29194 -2321 29230 -2228
rect 29356 -2276 29422 -2269
rect 29356 -2310 29372 -2276
rect 29406 -2310 29422 -2276
rect 29356 -2321 29422 -2310
rect 29194 -2322 29422 -2321
rect 28722 -2351 29422 -2322
rect 28722 -2352 29304 -2351
rect 28842 -2465 28876 -2352
rect 29238 -2393 29304 -2352
rect 29238 -2427 29254 -2393
rect 29288 -2427 29304 -2393
rect 29238 -2434 29304 -2427
rect 29666 -2461 29701 -2228
rect 29312 -2462 29701 -2461
rect 29898 -2462 29989 457
rect 30474 -53 30508 731
rect 31187 669 31221 731
rect 30776 631 31518 669
rect 30586 460 30596 528
rect 30651 460 30661 528
rect 30776 507 30810 631
rect 31012 507 31046 631
rect 31248 507 31282 631
rect 31484 507 31518 631
rect 30770 495 30816 507
rect 30770 119 30776 495
rect 30810 119 30816 495
rect 30770 107 30816 119
rect 30888 495 30934 507
rect 30888 119 30894 495
rect 30928 119 30934 495
rect 30888 107 30934 119
rect 31006 495 31052 507
rect 31006 119 31012 495
rect 31046 119 31052 495
rect 31006 107 31052 119
rect 31124 495 31170 507
rect 31124 119 31130 495
rect 31164 119 31170 495
rect 31124 107 31170 119
rect 31242 495 31288 507
rect 31242 119 31248 495
rect 31282 119 31288 495
rect 31242 107 31288 119
rect 31360 495 31406 507
rect 31360 119 31366 495
rect 31400 119 31406 495
rect 31360 107 31406 119
rect 31478 495 31524 507
rect 31478 119 31484 495
rect 31518 119 31524 495
rect 31644 290 31718 302
rect 31640 199 31650 290
rect 31712 199 31722 290
rect 31644 187 31718 199
rect 31478 107 31524 119
rect 31890 -52 31924 731
rect 32259 703 32295 797
rect 32495 703 32531 797
rect 32731 704 32767 797
rect 32893 749 32959 756
rect 32893 715 32909 749
rect 32943 715 32959 749
rect 32893 704 32959 715
rect 32731 703 32959 704
rect 32259 674 32959 703
rect 32259 673 32841 674
rect 31985 641 32061 646
rect 31982 585 31992 641
rect 32045 640 32061 641
rect 32045 585 32311 640
rect 31985 580 32311 585
rect 32106 538 32197 543
rect 32106 449 32116 538
rect 32189 449 32197 538
rect 32106 437 32197 449
rect 32143 43 32197 437
rect 32257 128 32311 580
rect 32379 560 32413 673
rect 32775 632 32841 673
rect 32775 598 32791 632
rect 32825 598 32841 632
rect 32775 591 32841 598
rect 33203 564 33238 797
rect 32849 560 33238 564
rect 32373 548 32419 560
rect 32373 172 32379 548
rect 32413 172 32419 548
rect 32373 160 32419 172
rect 32491 548 32537 560
rect 32491 172 32497 548
rect 32531 172 32537 548
rect 32491 160 32537 172
rect 32609 548 32655 560
rect 32609 172 32615 548
rect 32649 199 32655 548
rect 32726 548 32772 560
rect 32726 372 32732 548
rect 32766 372 32772 548
rect 32726 365 32772 372
rect 32844 548 33238 560
rect 32844 372 32850 548
rect 32884 538 33238 548
rect 32884 535 33097 538
rect 32884 372 32890 535
rect 33063 467 33097 535
rect 33224 467 33238 538
rect 33063 446 33238 467
rect 32726 360 32775 365
rect 32844 360 32890 372
rect 32732 199 32775 360
rect 32649 172 32775 199
rect 32916 289 33779 301
rect 32916 198 32932 289
rect 33056 198 33779 289
rect 32916 188 33779 198
rect 32609 160 32775 172
rect 32615 156 32775 160
rect 32257 122 32488 128
rect 32257 88 32438 122
rect 32472 88 32488 122
rect 32257 72 32488 88
rect 32540 122 32606 128
rect 32540 88 32556 122
rect 32590 88 32606 122
rect 32540 43 32606 88
rect 32143 35 32606 43
rect 32143 3 32607 35
rect 32699 19 32775 156
rect 32695 -41 32705 19
rect 32767 -41 32777 19
rect 31617 -53 31924 -52
rect 30474 -58 30790 -53
rect 31504 -58 31924 -53
rect 30474 -69 30857 -58
rect 30474 -96 30806 -69
rect 30474 -225 30508 -96
rect 30790 -103 30806 -96
rect 30840 -103 30857 -69
rect 30790 -109 30857 -103
rect 31437 -69 31924 -58
rect 32703 -67 32773 -41
rect 31437 -103 31454 -69
rect 31488 -96 31924 -69
rect 31488 -103 31504 -96
rect 31617 -97 31924 -96
rect 31437 -109 31504 -103
rect 30615 -136 30671 -124
rect 30615 -170 30621 -136
rect 30655 -137 30671 -136
rect 31728 -137 31784 -125
rect 30655 -153 31122 -137
rect 30655 -170 31072 -153
rect 30615 -186 31072 -170
rect 31056 -187 31072 -186
rect 31106 -187 31122 -153
rect 31056 -194 31122 -187
rect 31174 -152 31744 -137
rect 31174 -186 31190 -152
rect 31224 -171 31744 -152
rect 31778 -171 31784 -137
rect 31224 -186 31784 -171
rect 31174 -196 31241 -186
rect 31728 -187 31784 -186
rect 31890 -225 31924 -97
rect 30468 -237 30514 -225
rect 30468 -413 30474 -237
rect 30508 -413 30514 -237
rect 30468 -425 30514 -413
rect 30586 -237 30632 -225
rect 30586 -413 30592 -237
rect 30626 -413 30632 -237
rect 30586 -425 30632 -413
rect 30888 -237 30934 -225
rect 30591 -719 30625 -425
rect 30888 -613 30894 -237
rect 30928 -613 30934 -237
rect 30888 -625 30934 -613
rect 31006 -237 31052 -225
rect 31006 -613 31012 -237
rect 31046 -613 31052 -237
rect 31006 -625 31052 -613
rect 31124 -237 31170 -225
rect 31124 -613 31130 -237
rect 31164 -613 31170 -237
rect 31124 -625 31170 -613
rect 31242 -237 31288 -225
rect 31242 -613 31248 -237
rect 31282 -613 31288 -237
rect 31242 -625 31288 -613
rect 31360 -237 31406 -225
rect 31360 -613 31366 -237
rect 31400 -613 31406 -237
rect 31766 -237 31812 -225
rect 31766 -413 31772 -237
rect 31806 -413 31812 -237
rect 31766 -425 31812 -413
rect 31884 -237 31930 -225
rect 31884 -413 31890 -237
rect 31924 -413 31930 -237
rect 31884 -425 31930 -413
rect 31360 -625 31406 -613
rect 31248 -719 31282 -625
rect 31772 -719 31805 -425
rect 30591 -751 31805 -719
rect 30957 -775 31363 -751
rect 30957 -898 31069 -775
rect 31243 -898 31363 -775
rect 30957 -942 31363 -898
rect 30971 -1769 31416 -1763
rect 30971 -1969 30983 -1769
rect 31404 -1969 31416 -1769
rect 30971 -1975 31139 -1969
rect 31129 -2043 31139 -1975
rect 31271 -1975 31416 -1969
rect 31271 -2043 31281 -1975
rect 31139 -2083 31271 -2043
rect 31138 -2149 31271 -2083
rect 29312 -2465 29989 -2462
rect 26898 -2628 26944 -2616
rect 28836 -2477 28882 -2465
rect 26196 -2670 26230 -2628
rect 26432 -2670 26466 -2628
rect 26196 -2698 26466 -2670
rect 26550 -2669 26584 -2628
rect 26786 -2669 26820 -2628
rect 26550 -2698 26820 -2669
rect 26196 -2746 26230 -2698
rect 26196 -2776 26259 -2746
rect 26224 -2868 26259 -2776
rect 26731 -2806 26831 -2785
rect 26731 -2860 26745 -2806
rect 26810 -2860 26831 -2806
rect 26731 -2865 26831 -2860
rect 26904 -2811 26938 -2628
rect 26904 -2865 27013 -2811
rect 26224 -2904 26451 -2868
rect 26224 -3011 26259 -2904
rect 26385 -2938 26451 -2904
rect 26385 -2972 26401 -2938
rect 26435 -2972 26451 -2938
rect 26732 -2880 26829 -2865
rect 26732 -2947 26789 -2880
rect 26385 -2978 26451 -2972
rect 26626 -2983 26895 -2947
rect 26626 -3011 26659 -2983
rect 26862 -3011 26895 -2983
rect 26979 -3011 27013 -2865
rect 28671 -2814 28775 -2806
rect 28671 -2915 28681 -2814
rect 28767 -2897 28777 -2814
rect 28836 -2853 28842 -2477
rect 28876 -2853 28882 -2477
rect 28836 -2865 28882 -2853
rect 28954 -2477 29000 -2465
rect 28954 -2853 28960 -2477
rect 28994 -2853 29000 -2477
rect 28954 -2865 29000 -2853
rect 29072 -2477 29118 -2465
rect 29072 -2853 29078 -2477
rect 29112 -2826 29118 -2477
rect 29189 -2477 29235 -2465
rect 29189 -2653 29195 -2477
rect 29229 -2653 29235 -2477
rect 29189 -2660 29235 -2653
rect 29307 -2477 29989 -2465
rect 29307 -2653 29313 -2477
rect 29347 -2490 29989 -2477
rect 29347 -2653 29353 -2490
rect 29597 -2570 29989 -2490
rect 30467 -2192 31940 -2149
rect 30467 -2495 30501 -2192
rect 30833 -2295 30867 -2192
rect 31069 -2295 31103 -2192
rect 31305 -2295 31339 -2192
rect 31541 -2295 31575 -2192
rect 30827 -2307 30873 -2295
rect 30343 -2507 30389 -2495
rect 29189 -2665 29238 -2660
rect 29307 -2665 29353 -2653
rect 29195 -2826 29238 -2665
rect 30343 -2683 30349 -2507
rect 30383 -2683 30389 -2507
rect 30343 -2695 30389 -2683
rect 30461 -2507 30507 -2495
rect 30461 -2683 30467 -2507
rect 30501 -2683 30507 -2507
rect 30461 -2695 30507 -2683
rect 30579 -2507 30625 -2495
rect 30579 -2683 30585 -2507
rect 30619 -2683 30625 -2507
rect 30579 -2695 30625 -2683
rect 30697 -2507 30743 -2495
rect 30827 -2507 30833 -2307
rect 30697 -2683 30703 -2507
rect 30737 -2683 30833 -2507
rect 30867 -2683 30873 -2307
rect 30697 -2695 30743 -2683
rect 30827 -2695 30873 -2683
rect 30945 -2307 30991 -2295
rect 30945 -2683 30951 -2307
rect 30985 -2683 30991 -2307
rect 30945 -2695 30991 -2683
rect 31063 -2307 31109 -2295
rect 31063 -2683 31069 -2307
rect 31103 -2683 31109 -2307
rect 31063 -2695 31109 -2683
rect 31181 -2307 31227 -2295
rect 31181 -2683 31187 -2307
rect 31221 -2683 31227 -2307
rect 31181 -2695 31227 -2683
rect 31299 -2307 31345 -2295
rect 31299 -2683 31305 -2307
rect 31339 -2683 31345 -2307
rect 31299 -2695 31345 -2683
rect 31417 -2307 31463 -2295
rect 31417 -2683 31423 -2307
rect 31457 -2683 31463 -2307
rect 31417 -2695 31463 -2683
rect 31535 -2307 31581 -2295
rect 31535 -2683 31541 -2307
rect 31575 -2507 31581 -2307
rect 31906 -2495 31940 -2192
rect 32447 -2272 32583 -2252
rect 32447 -2334 32483 -2272
rect 32543 -2334 32583 -2272
rect 32447 -2362 32583 -2334
rect 32143 -2392 33120 -2362
rect 31664 -2507 31710 -2495
rect 31575 -2683 31670 -2507
rect 31704 -2683 31710 -2507
rect 31535 -2695 31581 -2683
rect 31664 -2695 31710 -2683
rect 31782 -2507 31828 -2495
rect 31782 -2683 31788 -2507
rect 31822 -2683 31828 -2507
rect 31782 -2695 31828 -2683
rect 31900 -2507 31946 -2495
rect 31900 -2683 31906 -2507
rect 31940 -2683 31946 -2507
rect 31900 -2695 31946 -2683
rect 32018 -2507 32064 -2495
rect 32143 -2498 32175 -2392
rect 32379 -2498 32411 -2392
rect 32615 -2498 32647 -2392
rect 32851 -2498 32883 -2392
rect 33086 -2498 33120 -2392
rect 32018 -2683 32024 -2507
rect 32058 -2683 32064 -2507
rect 32018 -2695 32064 -2683
rect 32136 -2510 32182 -2498
rect 32136 -2686 32142 -2510
rect 32176 -2686 32182 -2510
rect 30349 -2729 30383 -2695
rect 30951 -2729 30985 -2695
rect 31187 -2729 31221 -2695
rect 30349 -2764 30508 -2729
rect 30951 -2764 31221 -2729
rect 31788 -2729 31822 -2695
rect 32024 -2729 32058 -2695
rect 32136 -2698 32182 -2686
rect 32254 -2510 32300 -2498
rect 32254 -2686 32260 -2510
rect 32294 -2686 32300 -2510
rect 32254 -2698 32300 -2686
rect 32372 -2510 32418 -2498
rect 32372 -2686 32378 -2510
rect 32412 -2686 32418 -2510
rect 32372 -2698 32418 -2686
rect 32490 -2510 32536 -2498
rect 32490 -2686 32496 -2510
rect 32530 -2686 32536 -2510
rect 32490 -2698 32536 -2686
rect 32608 -2510 32654 -2498
rect 32608 -2686 32614 -2510
rect 32648 -2686 32654 -2510
rect 32608 -2698 32654 -2686
rect 32726 -2510 32772 -2498
rect 32726 -2686 32732 -2510
rect 32766 -2686 32772 -2510
rect 32726 -2698 32772 -2686
rect 32844 -2510 32890 -2498
rect 32844 -2686 32850 -2510
rect 32884 -2686 32890 -2510
rect 32844 -2698 32890 -2686
rect 32962 -2510 33008 -2498
rect 32962 -2686 32968 -2510
rect 33002 -2686 33008 -2510
rect 32962 -2698 33008 -2686
rect 33080 -2510 33126 -2498
rect 33080 -2686 33086 -2510
rect 33120 -2686 33126 -2510
rect 33080 -2698 33126 -2686
rect 33198 -2510 33244 -2498
rect 33198 -2686 33204 -2510
rect 33238 -2686 33244 -2510
rect 33198 -2698 33244 -2686
rect 31788 -2764 32058 -2729
rect 29112 -2853 29238 -2826
rect 29072 -2865 29238 -2853
rect 29078 -2869 29238 -2865
rect 28767 -2903 28951 -2897
rect 28767 -2915 28901 -2903
rect 28671 -2937 28901 -2915
rect 28935 -2937 28951 -2903
rect 28671 -2953 28951 -2937
rect 29003 -2903 29069 -2897
rect 29003 -2937 29019 -2903
rect 29053 -2937 29069 -2903
rect 29003 -2982 29069 -2937
rect 28448 -2988 29069 -2982
rect 26100 -3023 26146 -3011
rect 26100 -3199 26106 -3023
rect 26140 -3199 26146 -3023
rect 26100 -3211 26146 -3199
rect 26218 -3023 26264 -3011
rect 26218 -3199 26224 -3023
rect 26258 -3199 26264 -3023
rect 26218 -3211 26264 -3199
rect 26336 -3023 26382 -3011
rect 26336 -3199 26342 -3023
rect 26376 -3199 26382 -3023
rect 26336 -3211 26382 -3199
rect 26454 -3023 26500 -3011
rect 26454 -3199 26460 -3023
rect 26494 -3078 26500 -3023
rect 26619 -3023 26665 -3011
rect 26619 -3078 26625 -3023
rect 26494 -3166 26625 -3078
rect 26494 -3199 26500 -3166
rect 26454 -3211 26500 -3199
rect 26619 -3199 26625 -3166
rect 26659 -3199 26665 -3023
rect 26619 -3211 26665 -3199
rect 26737 -3023 26783 -3011
rect 26737 -3199 26743 -3023
rect 26777 -3199 26783 -3023
rect 26737 -3211 26783 -3199
rect 26855 -3023 26901 -3011
rect 26855 -3199 26861 -3023
rect 26895 -3199 26901 -3023
rect 26855 -3211 26901 -3199
rect 26973 -3023 27019 -3011
rect 26973 -3199 26979 -3023
rect 27013 -3199 27019 -3023
rect 28443 -3048 28453 -2988
rect 28538 -2990 29069 -2988
rect 28538 -3022 29070 -2990
rect 29162 -3006 29238 -2869
rect 28538 -3048 28548 -3022
rect 28448 -3055 28543 -3048
rect 29158 -3066 29168 -3006
rect 29230 -3066 29240 -3006
rect 29895 -3038 30336 -2975
rect 30403 -3038 30413 -2975
rect 26973 -3211 27019 -3199
rect 26106 -3250 26140 -3211
rect 26342 -3250 26376 -3211
rect 26106 -3286 26376 -3250
rect 26743 -3249 26776 -3211
rect 26979 -3249 27012 -3211
rect 26743 -3285 27012 -3249
rect 26106 -3287 26272 -3286
rect 26140 -3366 26272 -3287
rect 26130 -3474 26140 -3366
rect 26272 -3474 26282 -3366
rect 26161 -3611 26167 -3474
rect 26234 -3611 26240 -3474
rect 26161 -3623 26240 -3611
rect 22744 -3848 23721 -3818
rect 25938 -3820 26001 -3803
rect 25863 -3824 26001 -3820
rect 22744 -3954 22776 -3848
rect 22980 -3954 23012 -3848
rect 23216 -3954 23248 -3848
rect 23452 -3954 23484 -3848
rect 23687 -3954 23721 -3848
rect 24031 -3858 26001 -3824
rect 24029 -3887 26001 -3858
rect 24029 -3903 24075 -3887
rect 25863 -3889 26001 -3887
rect 22737 -3966 22783 -3954
rect 22737 -4142 22743 -3966
rect 22777 -4142 22783 -3966
rect 22737 -4154 22783 -4142
rect 22855 -3966 22901 -3954
rect 22855 -4142 22861 -3966
rect 22895 -4142 22901 -3966
rect 22855 -4154 22901 -4142
rect 22973 -3966 23019 -3954
rect 22973 -4142 22979 -3966
rect 23013 -4142 23019 -3966
rect 22973 -4154 23019 -4142
rect 23091 -3966 23137 -3954
rect 23091 -4142 23097 -3966
rect 23131 -4142 23137 -3966
rect 23091 -4154 23137 -4142
rect 23209 -3966 23255 -3954
rect 23209 -4142 23215 -3966
rect 23249 -4142 23255 -3966
rect 23209 -4154 23255 -4142
rect 23327 -3966 23373 -3954
rect 23327 -4142 23333 -3966
rect 23367 -4142 23373 -3966
rect 23327 -4154 23373 -4142
rect 23445 -3966 23491 -3954
rect 23445 -4142 23451 -3966
rect 23485 -4142 23491 -3966
rect 23445 -4154 23491 -4142
rect 23563 -3966 23609 -3954
rect 23563 -4142 23569 -3966
rect 23603 -4142 23609 -3966
rect 23563 -4154 23609 -4142
rect 23681 -3966 23727 -3954
rect 23681 -4142 23687 -3966
rect 23721 -4142 23727 -3966
rect 23681 -4154 23727 -4142
rect 23799 -3966 23845 -3954
rect 23799 -4142 23805 -3966
rect 23839 -4142 23845 -3966
rect 23799 -4154 23845 -4142
rect 22860 -4248 22896 -4154
rect 23096 -4248 23132 -4154
rect 23332 -4247 23368 -4154
rect 23494 -4202 23560 -4195
rect 23494 -4236 23510 -4202
rect 23544 -4236 23560 -4202
rect 23494 -4247 23560 -4236
rect 23332 -4248 23560 -4247
rect 22860 -4277 23560 -4248
rect 22860 -4278 23442 -4277
rect 22980 -4391 23014 -4278
rect 23376 -4319 23442 -4278
rect 23376 -4353 23392 -4319
rect 23426 -4353 23442 -4319
rect 23376 -4360 23442 -4353
rect 23804 -4372 23839 -4154
rect 24028 -4355 24075 -3903
rect 26924 -3896 27003 -3884
rect 26924 -4011 26930 -3896
rect 26997 -4011 27003 -3896
rect 24987 -4119 24997 -4011
rect 25129 -4119 25139 -4011
rect 26885 -4119 26895 -4011
rect 27027 -4119 27037 -4011
rect 24997 -4159 25129 -4119
rect 26895 -4159 27027 -4119
rect 24996 -4225 25129 -4159
rect 26894 -4225 27027 -4159
rect 24325 -4268 25798 -4225
rect 24028 -4371 24074 -4355
rect 23993 -4372 24074 -4371
rect 23804 -4387 24074 -4372
rect 23450 -4391 24074 -4387
rect 22974 -4403 23020 -4391
rect 22709 -4881 22719 -4763
rect 22837 -4795 22847 -4763
rect 22974 -4779 22980 -4403
rect 23014 -4779 23020 -4403
rect 22974 -4791 23020 -4779
rect 23092 -4403 23138 -4391
rect 23092 -4779 23098 -4403
rect 23132 -4779 23138 -4403
rect 23092 -4791 23138 -4779
rect 23210 -4403 23256 -4391
rect 23210 -4779 23216 -4403
rect 23250 -4755 23256 -4403
rect 23327 -4403 23373 -4391
rect 23327 -4579 23333 -4403
rect 23367 -4579 23373 -4403
rect 23327 -4591 23373 -4579
rect 23445 -4403 24074 -4391
rect 23445 -4579 23451 -4403
rect 23485 -4415 24074 -4403
rect 23485 -4416 23727 -4415
rect 23485 -4579 23491 -4416
rect 23993 -4417 24074 -4415
rect 24325 -4571 24359 -4268
rect 24691 -4371 24725 -4268
rect 24927 -4371 24961 -4268
rect 25163 -4371 25197 -4268
rect 25399 -4371 25433 -4268
rect 24685 -4383 24731 -4371
rect 23445 -4591 23491 -4579
rect 24201 -4583 24247 -4571
rect 23333 -4707 23368 -4591
rect 23464 -4707 23572 -4697
rect 23333 -4755 23464 -4707
rect 23572 -4738 23721 -4732
rect 23250 -4779 23464 -4755
rect 23210 -4791 23464 -4779
rect 23216 -4795 23464 -4791
rect 22837 -4823 22852 -4795
rect 22837 -4829 23089 -4823
rect 22837 -4863 23039 -4829
rect 23073 -4863 23089 -4829
rect 22837 -4879 23089 -4863
rect 23141 -4829 23207 -4823
rect 23141 -4863 23157 -4829
rect 23191 -4863 23207 -4829
rect 23390 -4839 23464 -4795
rect 23709 -4805 23721 -4738
rect 24201 -4759 24207 -4583
rect 24241 -4759 24247 -4583
rect 24201 -4771 24247 -4759
rect 24319 -4583 24365 -4571
rect 24319 -4759 24325 -4583
rect 24359 -4759 24365 -4583
rect 24319 -4771 24365 -4759
rect 24437 -4583 24483 -4571
rect 24437 -4759 24443 -4583
rect 24477 -4759 24483 -4583
rect 24437 -4771 24483 -4759
rect 24555 -4583 24601 -4571
rect 24685 -4583 24691 -4383
rect 24555 -4759 24561 -4583
rect 24595 -4759 24691 -4583
rect 24725 -4759 24731 -4383
rect 24555 -4771 24601 -4759
rect 24685 -4771 24731 -4759
rect 24803 -4383 24849 -4371
rect 24803 -4759 24809 -4383
rect 24843 -4759 24849 -4383
rect 24803 -4771 24849 -4759
rect 24921 -4383 24967 -4371
rect 24921 -4759 24927 -4383
rect 24961 -4759 24967 -4383
rect 24921 -4771 24967 -4759
rect 25039 -4383 25085 -4371
rect 25039 -4759 25045 -4383
rect 25079 -4759 25085 -4383
rect 25039 -4771 25085 -4759
rect 25157 -4383 25203 -4371
rect 25157 -4759 25163 -4383
rect 25197 -4759 25203 -4383
rect 25157 -4771 25203 -4759
rect 25275 -4383 25321 -4371
rect 25275 -4759 25281 -4383
rect 25315 -4759 25321 -4383
rect 25275 -4771 25321 -4759
rect 25393 -4383 25439 -4371
rect 25393 -4759 25399 -4383
rect 25433 -4583 25439 -4383
rect 25764 -4571 25798 -4268
rect 26223 -4268 27696 -4225
rect 26223 -4571 26257 -4268
rect 26589 -4371 26623 -4268
rect 26825 -4371 26859 -4268
rect 27061 -4371 27095 -4268
rect 27297 -4371 27331 -4268
rect 26583 -4383 26629 -4371
rect 25522 -4583 25568 -4571
rect 25433 -4759 25528 -4583
rect 25562 -4759 25568 -4583
rect 25393 -4771 25439 -4759
rect 25522 -4771 25568 -4759
rect 25640 -4583 25686 -4571
rect 25640 -4759 25646 -4583
rect 25680 -4759 25686 -4583
rect 25640 -4771 25686 -4759
rect 25758 -4583 25804 -4571
rect 25758 -4759 25764 -4583
rect 25798 -4759 25804 -4583
rect 25758 -4771 25804 -4759
rect 25876 -4583 25922 -4571
rect 25876 -4759 25882 -4583
rect 25916 -4759 25922 -4583
rect 25876 -4771 25922 -4759
rect 26099 -4583 26145 -4571
rect 26099 -4759 26105 -4583
rect 26139 -4759 26145 -4583
rect 26099 -4771 26145 -4759
rect 26217 -4583 26263 -4571
rect 26217 -4759 26223 -4583
rect 26257 -4759 26263 -4583
rect 26217 -4771 26263 -4759
rect 26335 -4583 26381 -4571
rect 26335 -4759 26341 -4583
rect 26375 -4759 26381 -4583
rect 26335 -4771 26381 -4759
rect 26453 -4583 26499 -4571
rect 26583 -4583 26589 -4383
rect 26453 -4759 26459 -4583
rect 26493 -4759 26589 -4583
rect 26623 -4759 26629 -4383
rect 26453 -4771 26499 -4759
rect 26583 -4771 26629 -4759
rect 26701 -4383 26747 -4371
rect 26701 -4759 26707 -4383
rect 26741 -4759 26747 -4383
rect 26701 -4771 26747 -4759
rect 26819 -4383 26865 -4371
rect 26819 -4759 26825 -4383
rect 26859 -4759 26865 -4383
rect 26819 -4771 26865 -4759
rect 26937 -4383 26983 -4371
rect 26937 -4759 26943 -4383
rect 26977 -4759 26983 -4383
rect 26937 -4771 26983 -4759
rect 27055 -4383 27101 -4371
rect 27055 -4759 27061 -4383
rect 27095 -4759 27101 -4383
rect 27055 -4771 27101 -4759
rect 27173 -4383 27219 -4371
rect 27173 -4759 27179 -4383
rect 27213 -4759 27219 -4383
rect 27173 -4771 27219 -4759
rect 27291 -4383 27337 -4371
rect 27291 -4759 27297 -4383
rect 27331 -4583 27337 -4383
rect 27662 -4571 27696 -4268
rect 27420 -4583 27466 -4571
rect 27331 -4759 27426 -4583
rect 27460 -4759 27466 -4583
rect 27291 -4771 27337 -4759
rect 27420 -4771 27466 -4759
rect 27538 -4583 27584 -4571
rect 27538 -4759 27544 -4583
rect 27578 -4759 27584 -4583
rect 27538 -4771 27584 -4759
rect 27656 -4583 27702 -4571
rect 27656 -4759 27662 -4583
rect 27696 -4759 27702 -4583
rect 27656 -4771 27702 -4759
rect 27774 -4583 27820 -4571
rect 27774 -4759 27780 -4583
rect 27814 -4759 27820 -4583
rect 27774 -4771 27820 -4759
rect 23572 -4811 23721 -4805
rect 24207 -4805 24241 -4771
rect 24809 -4805 24843 -4771
rect 25045 -4805 25079 -4771
rect 23464 -4849 23572 -4839
rect 24207 -4840 24366 -4805
rect 24809 -4840 25079 -4805
rect 25646 -4805 25680 -4771
rect 25882 -4805 25916 -4771
rect 25646 -4840 25916 -4805
rect 26105 -4805 26139 -4771
rect 26707 -4805 26741 -4771
rect 26943 -4805 26977 -4771
rect 26105 -4840 26264 -4805
rect 26707 -4840 26977 -4805
rect 27544 -4805 27578 -4771
rect 27780 -4805 27814 -4771
rect 27544 -4840 27814 -4805
rect 22837 -4881 22852 -4879
rect 22752 -4895 22852 -4881
rect 22752 -4938 22852 -4937
rect 22373 -4959 22852 -4938
rect 23141 -4959 23207 -4863
rect 22373 -5007 23207 -4959
rect 22373 -5036 22852 -5007
rect 22373 -5038 22478 -5036
rect 22752 -5037 22852 -5036
rect 22206 -5223 22216 -5144
rect 22309 -5223 22319 -5144
rect 23208 -5160 23287 -5148
rect 22217 -6397 22310 -5223
rect 23208 -5252 23214 -5160
rect 23135 -5272 23214 -5252
rect 23281 -5252 23287 -5160
rect 23281 -5272 23355 -5252
rect 23135 -5380 23179 -5272
rect 23311 -5380 23355 -5272
rect 23135 -5422 23355 -5380
rect 22739 -5452 23716 -5422
rect 22739 -5558 22771 -5452
rect 22975 -5558 23007 -5452
rect 23211 -5558 23243 -5452
rect 23447 -5558 23479 -5452
rect 23682 -5558 23716 -5452
rect 22732 -5570 22778 -5558
rect 22732 -5746 22738 -5570
rect 22772 -5746 22778 -5570
rect 22732 -5758 22778 -5746
rect 22850 -5570 22896 -5558
rect 22850 -5746 22856 -5570
rect 22890 -5746 22896 -5570
rect 22850 -5758 22896 -5746
rect 22968 -5570 23014 -5558
rect 22968 -5746 22974 -5570
rect 23008 -5746 23014 -5570
rect 22968 -5758 23014 -5746
rect 23086 -5570 23132 -5558
rect 23086 -5746 23092 -5570
rect 23126 -5746 23132 -5570
rect 23086 -5758 23132 -5746
rect 23204 -5570 23250 -5558
rect 23204 -5746 23210 -5570
rect 23244 -5746 23250 -5570
rect 23204 -5758 23250 -5746
rect 23322 -5570 23368 -5558
rect 23322 -5746 23328 -5570
rect 23362 -5746 23368 -5570
rect 23322 -5758 23368 -5746
rect 23440 -5570 23486 -5558
rect 23440 -5746 23446 -5570
rect 23480 -5746 23486 -5570
rect 23440 -5758 23486 -5746
rect 23558 -5570 23604 -5558
rect 23558 -5746 23564 -5570
rect 23598 -5746 23604 -5570
rect 23558 -5758 23604 -5746
rect 23676 -5570 23722 -5558
rect 23676 -5746 23682 -5570
rect 23716 -5746 23722 -5570
rect 23676 -5758 23722 -5746
rect 23794 -5570 23840 -5558
rect 23794 -5746 23800 -5570
rect 23834 -5746 23840 -5570
rect 23794 -5758 23840 -5746
rect 24332 -5624 24366 -4840
rect 25045 -4902 25079 -4840
rect 24634 -4940 25376 -4902
rect 24634 -5064 24668 -4940
rect 24870 -5064 24904 -4940
rect 25106 -5064 25140 -4940
rect 25342 -5064 25376 -4940
rect 25632 -5047 25642 -4981
rect 25705 -5047 25715 -4981
rect 24628 -5076 24674 -5064
rect 24628 -5452 24634 -5076
rect 24668 -5452 24674 -5076
rect 24628 -5464 24674 -5452
rect 24746 -5076 24792 -5064
rect 24746 -5452 24752 -5076
rect 24786 -5452 24792 -5076
rect 24746 -5464 24792 -5452
rect 24864 -5076 24910 -5064
rect 24864 -5452 24870 -5076
rect 24904 -5452 24910 -5076
rect 24864 -5464 24910 -5452
rect 24982 -5076 25028 -5064
rect 24982 -5452 24988 -5076
rect 25022 -5452 25028 -5076
rect 24982 -5464 25028 -5452
rect 25100 -5076 25146 -5064
rect 25100 -5452 25106 -5076
rect 25140 -5452 25146 -5076
rect 25100 -5464 25146 -5452
rect 25218 -5076 25264 -5064
rect 25218 -5452 25224 -5076
rect 25258 -5452 25264 -5076
rect 25218 -5464 25264 -5452
rect 25336 -5076 25382 -5064
rect 25336 -5452 25342 -5076
rect 25376 -5452 25382 -5076
rect 25336 -5464 25382 -5452
rect 25748 -5623 25782 -4840
rect 25475 -5624 25782 -5623
rect 24332 -5629 24648 -5624
rect 25362 -5629 25782 -5624
rect 24332 -5640 24715 -5629
rect 24332 -5667 24664 -5640
rect 22855 -5852 22891 -5758
rect 23091 -5852 23127 -5758
rect 23327 -5851 23363 -5758
rect 23489 -5806 23555 -5799
rect 23489 -5840 23505 -5806
rect 23539 -5840 23555 -5806
rect 23489 -5851 23555 -5840
rect 23327 -5852 23555 -5851
rect 22855 -5881 23555 -5852
rect 22855 -5882 23437 -5881
rect 22975 -5995 23009 -5882
rect 23371 -5923 23437 -5882
rect 23371 -5957 23387 -5923
rect 23421 -5957 23437 -5923
rect 23371 -5964 23437 -5957
rect 23799 -5991 23834 -5758
rect 24332 -5796 24366 -5667
rect 24648 -5674 24664 -5667
rect 24698 -5674 24715 -5640
rect 24648 -5680 24715 -5674
rect 25295 -5640 25782 -5629
rect 25295 -5674 25312 -5640
rect 25346 -5667 25782 -5640
rect 25346 -5674 25362 -5667
rect 25475 -5668 25782 -5667
rect 25295 -5680 25362 -5674
rect 24473 -5707 24529 -5695
rect 24473 -5741 24479 -5707
rect 24513 -5708 24529 -5707
rect 25586 -5708 25642 -5696
rect 24513 -5724 24980 -5708
rect 24513 -5741 24930 -5724
rect 24473 -5757 24930 -5741
rect 24914 -5758 24930 -5757
rect 24964 -5758 24980 -5724
rect 24914 -5765 24980 -5758
rect 25032 -5723 25602 -5708
rect 25032 -5757 25048 -5723
rect 25082 -5742 25602 -5723
rect 25636 -5742 25642 -5708
rect 25082 -5757 25642 -5742
rect 25032 -5767 25099 -5757
rect 25586 -5758 25642 -5757
rect 25748 -5796 25782 -5668
rect 26230 -5624 26264 -4840
rect 26943 -4902 26977 -4840
rect 26532 -4940 27274 -4902
rect 26532 -5064 26566 -4940
rect 26768 -5064 26802 -4940
rect 27004 -5064 27038 -4940
rect 27240 -5064 27274 -4940
rect 26526 -5076 26572 -5064
rect 26526 -5452 26532 -5076
rect 26566 -5452 26572 -5076
rect 26526 -5464 26572 -5452
rect 26644 -5076 26690 -5064
rect 26644 -5452 26650 -5076
rect 26684 -5452 26690 -5076
rect 26644 -5464 26690 -5452
rect 26762 -5076 26808 -5064
rect 26762 -5452 26768 -5076
rect 26802 -5452 26808 -5076
rect 26762 -5464 26808 -5452
rect 26880 -5076 26926 -5064
rect 26880 -5452 26886 -5076
rect 26920 -5452 26926 -5076
rect 26880 -5464 26926 -5452
rect 26998 -5076 27044 -5064
rect 26998 -5452 27004 -5076
rect 27038 -5452 27044 -5076
rect 26998 -5464 27044 -5452
rect 27116 -5076 27162 -5064
rect 27116 -5452 27122 -5076
rect 27156 -5452 27162 -5076
rect 27116 -5464 27162 -5452
rect 27234 -5076 27280 -5064
rect 27234 -5452 27240 -5076
rect 27274 -5452 27280 -5076
rect 27234 -5464 27280 -5452
rect 27646 -5623 27680 -4840
rect 28907 -4872 29043 -4852
rect 28907 -4934 28943 -4872
rect 29003 -4934 29043 -4872
rect 28907 -4962 29043 -4934
rect 28603 -4992 29580 -4962
rect 27258 -5624 27327 -5623
rect 27373 -5624 27680 -5623
rect 26230 -5629 26546 -5624
rect 27258 -5628 27680 -5624
rect 26230 -5640 26613 -5629
rect 26230 -5667 26562 -5640
rect 26230 -5796 26264 -5667
rect 26546 -5674 26562 -5667
rect 26596 -5674 26613 -5640
rect 26546 -5680 26613 -5674
rect 27191 -5639 27680 -5628
rect 27191 -5673 27208 -5639
rect 27242 -5667 27680 -5639
rect 27242 -5673 27258 -5667
rect 27373 -5668 27680 -5667
rect 27191 -5679 27258 -5673
rect 26371 -5707 26427 -5695
rect 26371 -5741 26377 -5707
rect 26411 -5708 26427 -5707
rect 27484 -5708 27540 -5696
rect 26411 -5724 26878 -5708
rect 26411 -5741 26828 -5724
rect 26371 -5757 26828 -5741
rect 26812 -5758 26828 -5757
rect 26862 -5758 26878 -5724
rect 26812 -5765 26878 -5758
rect 26930 -5723 27500 -5708
rect 26930 -5757 26946 -5723
rect 26980 -5742 27500 -5723
rect 27534 -5742 27540 -5708
rect 26980 -5757 27540 -5742
rect 26930 -5767 26997 -5757
rect 27484 -5758 27540 -5757
rect 27646 -5796 27680 -5668
rect 27761 -5018 27828 -4994
rect 27761 -5052 27778 -5018
rect 27812 -5052 27828 -5018
rect 23445 -5995 23834 -5991
rect 22969 -6007 23015 -5995
rect 22969 -6383 22975 -6007
rect 23009 -6383 23015 -6007
rect 22969 -6395 23015 -6383
rect 23087 -6007 23133 -5995
rect 23087 -6383 23093 -6007
rect 23127 -6383 23133 -6007
rect 23087 -6395 23133 -6383
rect 23205 -6007 23251 -5995
rect 23205 -6383 23211 -6007
rect 23245 -6359 23251 -6007
rect 23322 -6007 23368 -5995
rect 23322 -6183 23328 -6007
rect 23362 -6183 23368 -6007
rect 23322 -6195 23368 -6183
rect 23440 -6007 23834 -5995
rect 24326 -5808 24372 -5796
rect 24326 -5984 24332 -5808
rect 24366 -5984 24372 -5808
rect 24326 -5996 24372 -5984
rect 24444 -5808 24490 -5796
rect 24444 -5984 24450 -5808
rect 24484 -5984 24490 -5808
rect 24444 -5996 24490 -5984
rect 24746 -5808 24792 -5796
rect 23440 -6183 23446 -6007
rect 23480 -6020 23834 -6007
rect 23480 -6183 23486 -6020
rect 23756 -6023 23834 -6020
rect 23756 -6075 23766 -6023
rect 23829 -6075 23839 -6023
rect 23761 -6081 23834 -6075
rect 23440 -6195 23486 -6183
rect 23328 -6311 23363 -6195
rect 24449 -6290 24483 -5996
rect 24746 -6184 24752 -5808
rect 24786 -6184 24792 -5808
rect 24746 -6196 24792 -6184
rect 24864 -5808 24910 -5796
rect 24864 -6184 24870 -5808
rect 24904 -6184 24910 -5808
rect 24864 -6196 24910 -6184
rect 24982 -5808 25028 -5796
rect 24982 -6184 24988 -5808
rect 25022 -6184 25028 -5808
rect 24982 -6196 25028 -6184
rect 25100 -5808 25146 -5796
rect 25100 -6184 25106 -5808
rect 25140 -6184 25146 -5808
rect 25100 -6196 25146 -6184
rect 25218 -5808 25264 -5796
rect 25218 -6184 25224 -5808
rect 25258 -6184 25264 -5808
rect 25624 -5808 25670 -5796
rect 25624 -5984 25630 -5808
rect 25664 -5984 25670 -5808
rect 25624 -5996 25670 -5984
rect 25742 -5808 25788 -5796
rect 25742 -5984 25748 -5808
rect 25782 -5984 25788 -5808
rect 25742 -5996 25788 -5984
rect 26224 -5808 26270 -5796
rect 26224 -5984 26230 -5808
rect 26264 -5984 26270 -5808
rect 26224 -5996 26270 -5984
rect 26342 -5808 26388 -5796
rect 26342 -5984 26348 -5808
rect 26382 -5984 26388 -5808
rect 26342 -5996 26388 -5984
rect 26644 -5808 26690 -5796
rect 25218 -6196 25264 -6184
rect 25106 -6290 25140 -6196
rect 25630 -6290 25663 -5996
rect 23459 -6311 23567 -6301
rect 23328 -6359 23459 -6311
rect 24449 -6322 25663 -6290
rect 26347 -6290 26381 -5996
rect 26644 -6184 26650 -5808
rect 26684 -6184 26690 -5808
rect 26644 -6196 26690 -6184
rect 26762 -5808 26808 -5796
rect 26762 -6184 26768 -5808
rect 26802 -6184 26808 -5808
rect 26762 -6196 26808 -6184
rect 26880 -5808 26926 -5796
rect 26880 -6184 26886 -5808
rect 26920 -6184 26926 -5808
rect 26880 -6196 26926 -6184
rect 26998 -5808 27044 -5796
rect 26998 -6184 27004 -5808
rect 27038 -6184 27044 -5808
rect 26998 -6196 27044 -6184
rect 27116 -5808 27162 -5796
rect 27116 -6184 27122 -5808
rect 27156 -6184 27162 -5808
rect 27522 -5808 27568 -5796
rect 27522 -5984 27528 -5808
rect 27562 -5984 27568 -5808
rect 27522 -5996 27568 -5984
rect 27640 -5808 27686 -5796
rect 27640 -5984 27646 -5808
rect 27680 -5984 27686 -5808
rect 27640 -5996 27686 -5984
rect 27116 -6196 27162 -6184
rect 27004 -6290 27038 -6196
rect 27528 -6290 27561 -5996
rect 26347 -6322 27561 -6290
rect 23567 -6355 23712 -6349
rect 23245 -6383 23459 -6359
rect 23205 -6395 23459 -6383
rect 22217 -6399 22802 -6397
rect 23211 -6399 23459 -6395
rect 22217 -6427 22847 -6399
rect 22217 -6433 23084 -6427
rect 22217 -6467 23034 -6433
rect 23068 -6467 23084 -6433
rect 22217 -6483 23084 -6467
rect 23136 -6433 23202 -6427
rect 23136 -6467 23152 -6433
rect 23186 -6467 23202 -6433
rect 23385 -6443 23459 -6399
rect 23700 -6422 23712 -6355
rect 24942 -6407 25074 -6322
rect 26840 -6407 26972 -6322
rect 23567 -6428 23712 -6422
rect 23459 -6453 23567 -6443
rect 22217 -6499 22847 -6483
rect 22217 -6503 22802 -6499
rect 22217 -6504 22318 -6503
rect 22747 -6552 22847 -6541
rect 22711 -6658 22721 -6552
rect 22833 -6563 22847 -6552
rect 23136 -6563 23202 -6467
rect 24932 -6515 24942 -6407
rect 25074 -6515 25084 -6407
rect 26830 -6515 26840 -6407
rect 26972 -6515 26982 -6407
rect 27761 -6435 27828 -5052
rect 28603 -5098 28635 -4992
rect 28839 -5098 28871 -4992
rect 29075 -5098 29107 -4992
rect 29311 -5098 29343 -4992
rect 29546 -5098 29580 -4992
rect 28596 -5110 28642 -5098
rect 28596 -5286 28602 -5110
rect 28636 -5286 28642 -5110
rect 28596 -5298 28642 -5286
rect 28714 -5110 28760 -5098
rect 28714 -5286 28720 -5110
rect 28754 -5286 28760 -5110
rect 28714 -5298 28760 -5286
rect 28832 -5110 28878 -5098
rect 28832 -5286 28838 -5110
rect 28872 -5286 28878 -5110
rect 28832 -5298 28878 -5286
rect 28950 -5110 28996 -5098
rect 28950 -5286 28956 -5110
rect 28990 -5286 28996 -5110
rect 28950 -5298 28996 -5286
rect 29068 -5110 29114 -5098
rect 29068 -5286 29074 -5110
rect 29108 -5286 29114 -5110
rect 29068 -5298 29114 -5286
rect 29186 -5110 29232 -5098
rect 29186 -5286 29192 -5110
rect 29226 -5286 29232 -5110
rect 29186 -5298 29232 -5286
rect 29304 -5110 29350 -5098
rect 29304 -5286 29310 -5110
rect 29344 -5286 29350 -5110
rect 29304 -5298 29350 -5286
rect 29422 -5110 29468 -5098
rect 29422 -5286 29428 -5110
rect 29462 -5286 29468 -5110
rect 29422 -5298 29468 -5286
rect 29540 -5110 29586 -5098
rect 29540 -5286 29546 -5110
rect 29580 -5286 29586 -5110
rect 29540 -5298 29586 -5286
rect 29658 -5110 29704 -5098
rect 29658 -5286 29664 -5110
rect 29698 -5286 29704 -5110
rect 29658 -5298 29704 -5286
rect 28719 -5392 28755 -5298
rect 28955 -5392 28991 -5298
rect 29191 -5391 29227 -5298
rect 29353 -5346 29419 -5339
rect 29353 -5380 29369 -5346
rect 29403 -5380 29419 -5346
rect 29353 -5391 29419 -5380
rect 29191 -5392 29419 -5391
rect 28719 -5421 29419 -5392
rect 28719 -5422 29301 -5421
rect 27889 -5481 28045 -5475
rect 27889 -5579 27901 -5481
rect 28033 -5579 28045 -5481
rect 28839 -5535 28873 -5422
rect 29235 -5463 29301 -5422
rect 29235 -5497 29251 -5463
rect 29285 -5497 29301 -5463
rect 29235 -5504 29301 -5497
rect 29663 -5531 29698 -5298
rect 29309 -5532 29844 -5531
rect 29895 -5532 29990 -3038
rect 30474 -3548 30508 -2764
rect 31187 -2826 31221 -2764
rect 30776 -2864 31518 -2826
rect 30586 -3035 30596 -2967
rect 30651 -3035 30661 -2967
rect 30776 -2988 30810 -2864
rect 31012 -2988 31046 -2864
rect 31248 -2988 31282 -2864
rect 31484 -2988 31518 -2864
rect 30770 -3000 30816 -2988
rect 30770 -3376 30776 -3000
rect 30810 -3376 30816 -3000
rect 30770 -3388 30816 -3376
rect 30888 -3000 30934 -2988
rect 30888 -3376 30894 -3000
rect 30928 -3376 30934 -3000
rect 30888 -3388 30934 -3376
rect 31006 -3000 31052 -2988
rect 31006 -3376 31012 -3000
rect 31046 -3376 31052 -3000
rect 31006 -3388 31052 -3376
rect 31124 -3000 31170 -2988
rect 31124 -3376 31130 -3000
rect 31164 -3376 31170 -3000
rect 31124 -3388 31170 -3376
rect 31242 -3000 31288 -2988
rect 31242 -3376 31248 -3000
rect 31282 -3376 31288 -3000
rect 31242 -3388 31288 -3376
rect 31360 -3000 31406 -2988
rect 31360 -3376 31366 -3000
rect 31400 -3376 31406 -3000
rect 31360 -3388 31406 -3376
rect 31478 -3000 31524 -2988
rect 31478 -3376 31484 -3000
rect 31518 -3376 31524 -3000
rect 31644 -3205 31718 -3193
rect 31640 -3296 31650 -3205
rect 31712 -3296 31722 -3205
rect 31644 -3308 31718 -3296
rect 31478 -3388 31524 -3376
rect 31890 -3547 31924 -2764
rect 32259 -2792 32295 -2698
rect 32495 -2792 32531 -2698
rect 32731 -2791 32767 -2698
rect 32893 -2746 32959 -2739
rect 32893 -2780 32909 -2746
rect 32943 -2780 32959 -2746
rect 32893 -2791 32959 -2780
rect 32731 -2792 32959 -2791
rect 32259 -2821 32959 -2792
rect 32259 -2822 32841 -2821
rect 31985 -2854 32061 -2849
rect 31982 -2910 31992 -2854
rect 32045 -2855 32061 -2854
rect 32045 -2910 32311 -2855
rect 31985 -2915 32311 -2910
rect 32106 -2957 32197 -2952
rect 32106 -3046 32116 -2957
rect 32189 -3046 32197 -2957
rect 32106 -3058 32197 -3046
rect 32143 -3452 32197 -3058
rect 32257 -3367 32311 -2915
rect 32379 -2935 32413 -2822
rect 32775 -2863 32841 -2822
rect 32775 -2897 32791 -2863
rect 32825 -2897 32841 -2863
rect 32775 -2904 32841 -2897
rect 33203 -2931 33238 -2698
rect 32849 -2935 33238 -2931
rect 32373 -2947 32419 -2935
rect 32373 -3323 32379 -2947
rect 32413 -3323 32419 -2947
rect 32373 -3335 32419 -3323
rect 32491 -2947 32537 -2935
rect 32491 -3323 32497 -2947
rect 32531 -3323 32537 -2947
rect 32491 -3335 32537 -3323
rect 32609 -2947 32655 -2935
rect 32609 -3323 32615 -2947
rect 32649 -3296 32655 -2947
rect 32726 -2947 32772 -2935
rect 32726 -3123 32732 -2947
rect 32766 -3123 32772 -2947
rect 32726 -3130 32772 -3123
rect 32844 -2947 33238 -2935
rect 32844 -3123 32850 -2947
rect 32884 -2960 33238 -2947
rect 32884 -3123 32890 -2960
rect 33063 -3049 33238 -2960
rect 33107 -3050 33238 -3049
rect 32726 -3135 32775 -3130
rect 32844 -3135 32890 -3123
rect 32732 -3296 32775 -3135
rect 32649 -3323 32775 -3296
rect 32609 -3335 32775 -3323
rect 32615 -3339 32775 -3335
rect 32257 -3373 32488 -3367
rect 32257 -3407 32438 -3373
rect 32472 -3407 32488 -3373
rect 32257 -3423 32488 -3407
rect 32540 -3373 32606 -3367
rect 32540 -3407 32556 -3373
rect 32590 -3407 32606 -3373
rect 32540 -3452 32606 -3407
rect 32143 -3460 32606 -3452
rect 32143 -3492 32607 -3460
rect 32699 -3476 32775 -3339
rect 32695 -3536 32705 -3476
rect 32767 -3536 32777 -3476
rect 31617 -3548 31924 -3547
rect 30474 -3553 30790 -3548
rect 31504 -3553 31924 -3548
rect 30474 -3564 30857 -3553
rect 30474 -3591 30806 -3564
rect 30474 -3720 30508 -3591
rect 30790 -3598 30806 -3591
rect 30840 -3598 30857 -3564
rect 30790 -3604 30857 -3598
rect 31437 -3564 31924 -3553
rect 32703 -3562 32773 -3536
rect 31437 -3598 31454 -3564
rect 31488 -3591 31924 -3564
rect 31488 -3598 31504 -3591
rect 31617 -3592 31924 -3591
rect 31437 -3604 31504 -3598
rect 30615 -3631 30671 -3619
rect 30615 -3665 30621 -3631
rect 30655 -3632 30671 -3631
rect 31728 -3632 31784 -3620
rect 30655 -3648 31122 -3632
rect 30655 -3665 31072 -3648
rect 30615 -3681 31072 -3665
rect 31056 -3682 31072 -3681
rect 31106 -3682 31122 -3648
rect 31056 -3689 31122 -3682
rect 31174 -3647 31744 -3632
rect 31174 -3681 31190 -3647
rect 31224 -3666 31744 -3647
rect 31778 -3666 31784 -3632
rect 31224 -3681 31784 -3666
rect 31174 -3691 31241 -3681
rect 31728 -3682 31784 -3681
rect 31890 -3720 31924 -3592
rect 30468 -3732 30514 -3720
rect 30468 -3908 30474 -3732
rect 30508 -3908 30514 -3732
rect 30468 -3920 30514 -3908
rect 30586 -3732 30632 -3720
rect 30586 -3908 30592 -3732
rect 30626 -3908 30632 -3732
rect 30586 -3920 30632 -3908
rect 30888 -3732 30934 -3720
rect 30591 -4214 30625 -3920
rect 30888 -4108 30894 -3732
rect 30928 -4108 30934 -3732
rect 30888 -4120 30934 -4108
rect 31006 -3732 31052 -3720
rect 31006 -4108 31012 -3732
rect 31046 -4108 31052 -3732
rect 31006 -4120 31052 -4108
rect 31124 -3732 31170 -3720
rect 31124 -4108 31130 -3732
rect 31164 -4108 31170 -3732
rect 31124 -4120 31170 -4108
rect 31242 -3732 31288 -3720
rect 31242 -4108 31248 -3732
rect 31282 -4108 31288 -3732
rect 31242 -4120 31288 -4108
rect 31360 -3732 31406 -3720
rect 31360 -4108 31366 -3732
rect 31400 -4108 31406 -3732
rect 31766 -3732 31812 -3720
rect 31766 -3908 31772 -3732
rect 31806 -3908 31812 -3732
rect 31766 -3920 31812 -3908
rect 31884 -3732 31930 -3720
rect 31884 -3908 31890 -3732
rect 31924 -3908 31930 -3732
rect 31884 -3920 31930 -3908
rect 31360 -4120 31406 -4108
rect 31248 -4214 31282 -4120
rect 31772 -4214 31805 -3920
rect 30591 -4246 31805 -4214
rect 30957 -4270 31363 -4246
rect 30957 -4393 31069 -4270
rect 31243 -4393 31363 -4270
rect 30957 -4437 31363 -4393
rect 29309 -5535 29990 -5532
rect 27889 -5585 28045 -5579
rect 28833 -5547 28879 -5535
rect 28281 -5802 28391 -5801
rect 28279 -5803 28657 -5802
rect 28279 -5808 28658 -5803
rect 28273 -5898 28283 -5808
rect 28367 -5898 28658 -5808
rect 28279 -5902 28658 -5898
rect 28281 -5903 28391 -5902
rect 28581 -5903 28658 -5902
rect 28603 -6052 28657 -5903
rect 28833 -5923 28839 -5547
rect 28873 -5923 28879 -5547
rect 28833 -5935 28879 -5923
rect 28951 -5547 28997 -5535
rect 28951 -5923 28957 -5547
rect 28991 -5923 28997 -5547
rect 28951 -5935 28997 -5923
rect 29069 -5547 29115 -5535
rect 29069 -5923 29075 -5547
rect 29109 -5896 29115 -5547
rect 29186 -5547 29232 -5535
rect 29186 -5723 29192 -5547
rect 29226 -5723 29232 -5547
rect 29186 -5730 29232 -5723
rect 29304 -5547 29990 -5535
rect 29304 -5723 29310 -5547
rect 29344 -5560 29990 -5547
rect 29344 -5723 29350 -5560
rect 29594 -5640 29990 -5560
rect 29186 -5735 29235 -5730
rect 29304 -5735 29350 -5723
rect 29192 -5896 29235 -5735
rect 33125 -5758 33238 -3050
rect 33284 -3206 33781 -3193
rect 33284 -3297 33299 -3206
rect 33409 -3297 33781 -3206
rect 33284 -3306 33781 -3297
rect 29562 -5762 33238 -5758
rect 29109 -5923 29235 -5896
rect 29069 -5935 29235 -5923
rect 29075 -5939 29235 -5935
rect 28713 -5955 28786 -5950
rect 28707 -6019 28717 -5955
rect 28783 -5967 28793 -5955
rect 28783 -5973 28948 -5967
rect 28783 -6007 28898 -5973
rect 28932 -6007 28948 -5973
rect 28783 -6019 28948 -6007
rect 28713 -6023 28948 -6019
rect 29000 -5973 29066 -5967
rect 29000 -6007 29016 -5973
rect 29050 -6007 29066 -5973
rect 29000 -6052 29066 -6007
rect 28603 -6060 29066 -6052
rect 28603 -6092 29067 -6060
rect 29159 -6076 29235 -5939
rect 29559 -5876 33238 -5762
rect 29155 -6136 29165 -6076
rect 29227 -6136 29237 -6076
rect 22833 -6611 23202 -6563
rect 22833 -6641 22847 -6611
rect 22833 -6658 22843 -6641
rect 23135 -6714 23201 -6611
rect 24964 -6650 24970 -6515
rect 25037 -6650 25043 -6515
rect 24964 -6662 25043 -6650
rect 27761 -6714 27827 -6435
rect 23133 -6794 27827 -6714
rect 29559 -7229 29724 -5876
rect 30971 -6117 31416 -6111
rect 30971 -6317 30983 -6117
rect 31404 -6317 31416 -6117
rect 30971 -6323 31139 -6317
rect 31129 -6391 31139 -6323
rect 31271 -6323 31416 -6317
rect 31271 -6391 31281 -6323
rect 31139 -6431 31271 -6391
rect 31138 -6497 31271 -6431
rect 30467 -6540 31940 -6497
rect 30467 -6843 30501 -6540
rect 30833 -6643 30867 -6540
rect 31069 -6643 31103 -6540
rect 31305 -6643 31339 -6540
rect 31541 -6643 31575 -6540
rect 30827 -6655 30873 -6643
rect 30343 -6855 30389 -6843
rect 30343 -7031 30349 -6855
rect 30383 -7031 30389 -6855
rect 30343 -7043 30389 -7031
rect 30461 -6855 30507 -6843
rect 30461 -7031 30467 -6855
rect 30501 -7031 30507 -6855
rect 30461 -7043 30507 -7031
rect 30579 -6855 30625 -6843
rect 30579 -7031 30585 -6855
rect 30619 -7031 30625 -6855
rect 30579 -7043 30625 -7031
rect 30697 -6855 30743 -6843
rect 30827 -6855 30833 -6655
rect 30697 -7031 30703 -6855
rect 30737 -7031 30833 -6855
rect 30867 -7031 30873 -6655
rect 30697 -7043 30743 -7031
rect 30827 -7043 30873 -7031
rect 30945 -6655 30991 -6643
rect 30945 -7031 30951 -6655
rect 30985 -7031 30991 -6655
rect 30945 -7043 30991 -7031
rect 31063 -6655 31109 -6643
rect 31063 -7031 31069 -6655
rect 31103 -7031 31109 -6655
rect 31063 -7043 31109 -7031
rect 31181 -6655 31227 -6643
rect 31181 -7031 31187 -6655
rect 31221 -7031 31227 -6655
rect 31181 -7043 31227 -7031
rect 31299 -6655 31345 -6643
rect 31299 -7031 31305 -6655
rect 31339 -7031 31345 -6655
rect 31299 -7043 31345 -7031
rect 31417 -6655 31463 -6643
rect 31417 -7031 31423 -6655
rect 31457 -7031 31463 -6655
rect 31417 -7043 31463 -7031
rect 31535 -6655 31581 -6643
rect 31535 -7031 31541 -6655
rect 31575 -6855 31581 -6655
rect 31906 -6843 31940 -6540
rect 32447 -6620 32583 -6600
rect 32447 -6682 32483 -6620
rect 32543 -6682 32583 -6620
rect 32447 -6710 32583 -6682
rect 32143 -6740 33120 -6710
rect 31664 -6855 31710 -6843
rect 31575 -7031 31670 -6855
rect 31704 -7031 31710 -6855
rect 31535 -7043 31581 -7031
rect 31664 -7043 31710 -7031
rect 31782 -6855 31828 -6843
rect 31782 -7031 31788 -6855
rect 31822 -7031 31828 -6855
rect 31782 -7043 31828 -7031
rect 31900 -6855 31946 -6843
rect 31900 -7031 31906 -6855
rect 31940 -7031 31946 -6855
rect 31900 -7043 31946 -7031
rect 32018 -6855 32064 -6843
rect 32143 -6846 32175 -6740
rect 32379 -6846 32411 -6740
rect 32615 -6846 32647 -6740
rect 32851 -6846 32883 -6740
rect 33086 -6846 33120 -6740
rect 32018 -7031 32024 -6855
rect 32058 -7031 32064 -6855
rect 32018 -7043 32064 -7031
rect 32136 -6858 32182 -6846
rect 32136 -7034 32142 -6858
rect 32176 -7034 32182 -6858
rect 30349 -7077 30383 -7043
rect 30951 -7077 30985 -7043
rect 31187 -7077 31221 -7043
rect 30349 -7112 30508 -7077
rect 30951 -7112 31221 -7077
rect 31788 -7077 31822 -7043
rect 32024 -7077 32058 -7043
rect 32136 -7046 32182 -7034
rect 32254 -6858 32300 -6846
rect 32254 -7034 32260 -6858
rect 32294 -7034 32300 -6858
rect 32254 -7046 32300 -7034
rect 32372 -6858 32418 -6846
rect 32372 -7034 32378 -6858
rect 32412 -7034 32418 -6858
rect 32372 -7046 32418 -7034
rect 32490 -6858 32536 -6846
rect 32490 -7034 32496 -6858
rect 32530 -7034 32536 -6858
rect 32490 -7046 32536 -7034
rect 32608 -6858 32654 -6846
rect 32608 -7034 32614 -6858
rect 32648 -7034 32654 -6858
rect 32608 -7046 32654 -7034
rect 32726 -6858 32772 -6846
rect 32726 -7034 32732 -6858
rect 32766 -7034 32772 -6858
rect 32726 -7046 32772 -7034
rect 32844 -6858 32890 -6846
rect 32844 -7034 32850 -6858
rect 32884 -7034 32890 -6858
rect 32844 -7046 32890 -7034
rect 32962 -6858 33008 -6846
rect 32962 -7034 32968 -6858
rect 33002 -7034 33008 -6858
rect 32962 -7046 33008 -7034
rect 33080 -6858 33126 -6846
rect 33080 -7034 33086 -6858
rect 33120 -7034 33126 -6858
rect 33080 -7046 33126 -7034
rect 33198 -6858 33244 -6846
rect 33198 -7034 33204 -6858
rect 33238 -7034 33244 -6858
rect 33198 -7046 33244 -7034
rect 31788 -7112 32058 -7077
rect 21809 -7380 29724 -7229
rect 30317 -7193 30414 -7187
rect 30317 -7264 30329 -7193
rect 30402 -7197 30414 -7193
rect 30403 -7260 30414 -7197
rect 30402 -7264 30414 -7260
rect 30317 -7270 30414 -7264
rect 21888 -7382 29724 -7380
rect 29895 -7323 30359 -7322
rect 29895 -7386 30336 -7323
rect 30403 -7386 30413 -7323
rect 29895 -7389 30359 -7386
rect 27381 -7458 28669 -7457
rect 20913 -7806 21706 -7726
rect 20663 -7819 21706 -7806
rect 20623 -7831 21706 -7819
rect 20158 -7944 20192 -7831
rect 20628 -7835 21706 -7831
rect 24307 -7459 28793 -7458
rect 24307 -7468 28794 -7459
rect 24307 -7558 28697 -7468
rect 28781 -7558 28794 -7468
rect 24307 -7564 28794 -7558
rect 24307 -7565 28793 -7564
rect 20554 -7869 20620 -7862
rect 20554 -7903 20570 -7869
rect 20604 -7903 20620 -7869
rect 20554 -7944 20620 -7903
rect 20038 -7945 20620 -7944
rect 20038 -7974 20738 -7945
rect 20038 -8068 20074 -7974
rect 20274 -8068 20310 -7974
rect 20510 -7975 20738 -7974
rect 20510 -8068 20546 -7975
rect 20672 -7986 20738 -7975
rect 20672 -8020 20688 -7986
rect 20722 -8020 20738 -7986
rect 20672 -8027 20738 -8020
rect 20982 -8068 21017 -7835
rect 19915 -8080 19961 -8068
rect 19915 -8256 19921 -8080
rect 19955 -8256 19961 -8080
rect 19915 -8268 19961 -8256
rect 20033 -8080 20079 -8068
rect 20033 -8256 20039 -8080
rect 20073 -8256 20079 -8080
rect 20033 -8268 20079 -8256
rect 20151 -8080 20197 -8068
rect 20151 -8256 20157 -8080
rect 20191 -8256 20197 -8080
rect 20151 -8268 20197 -8256
rect 20269 -8080 20315 -8068
rect 20269 -8256 20275 -8080
rect 20309 -8256 20315 -8080
rect 20269 -8268 20315 -8256
rect 20387 -8080 20433 -8068
rect 20387 -8256 20393 -8080
rect 20427 -8256 20433 -8080
rect 20387 -8268 20433 -8256
rect 20505 -8080 20551 -8068
rect 20505 -8256 20511 -8080
rect 20545 -8256 20551 -8080
rect 20505 -8268 20551 -8256
rect 20623 -8080 20669 -8068
rect 20623 -8256 20629 -8080
rect 20663 -8256 20669 -8080
rect 20623 -8268 20669 -8256
rect 20741 -8080 20787 -8068
rect 20741 -8256 20747 -8080
rect 20781 -8256 20787 -8080
rect 20741 -8268 20787 -8256
rect 20859 -8080 20905 -8068
rect 20859 -8256 20865 -8080
rect 20899 -8256 20905 -8080
rect 20859 -8268 20905 -8256
rect 20977 -8080 21023 -8068
rect 20977 -8256 20983 -8080
rect 21017 -8256 21023 -8080
rect 20977 -8268 21023 -8256
rect 19922 -8374 19954 -8268
rect 20158 -8374 20190 -8268
rect 20394 -8374 20426 -8268
rect 20630 -8374 20662 -8268
rect 20865 -8374 20899 -8268
rect 19922 -8404 20899 -8374
rect 20226 -8432 20362 -8404
rect 20226 -8494 20262 -8432
rect 20322 -8494 20362 -8432
rect 20226 -8514 20362 -8494
rect -1124 -8696 416 -8695
rect 12795 -8696 13219 -8695
rect -1124 -8701 13219 -8696
rect -1124 -8705 6527 -8701
rect -1124 -8774 1487 -8705
rect 1583 -8774 6527 -8705
rect -1124 -8775 6527 -8774
rect 6627 -8775 13219 -8701
rect -1124 -8780 13219 -8775
rect 13733 -8667 19697 -8592
rect -258 -8781 12841 -8780
rect -638 -8811 12908 -8809
rect 13733 -8811 13814 -8667
rect 24307 -8706 24463 -7565
rect 28914 -7717 29050 -7697
rect 28914 -7779 28950 -7717
rect 29010 -7779 29050 -7717
rect 28914 -7807 29050 -7779
rect 28610 -7837 29587 -7807
rect 28610 -7943 28642 -7837
rect 28846 -7943 28878 -7837
rect 29082 -7943 29114 -7837
rect 29318 -7943 29350 -7837
rect 29553 -7943 29587 -7837
rect 28603 -7955 28649 -7943
rect 28603 -8131 28609 -7955
rect 28643 -8131 28649 -7955
rect 28603 -8143 28649 -8131
rect 28721 -7955 28767 -7943
rect 28721 -8131 28727 -7955
rect 28761 -8131 28767 -7955
rect 28721 -8143 28767 -8131
rect 28839 -7955 28885 -7943
rect 28839 -8131 28845 -7955
rect 28879 -8131 28885 -7955
rect 28839 -8143 28885 -8131
rect 28957 -7955 29003 -7943
rect 28957 -8131 28963 -7955
rect 28997 -8131 29003 -7955
rect 28957 -8143 29003 -8131
rect 29075 -7955 29121 -7943
rect 29075 -8131 29081 -7955
rect 29115 -8131 29121 -7955
rect 29075 -8143 29121 -8131
rect 29193 -7955 29239 -7943
rect 29193 -8131 29199 -7955
rect 29233 -8131 29239 -7955
rect 29193 -8143 29239 -8131
rect 29311 -7955 29357 -7943
rect 29311 -8131 29317 -7955
rect 29351 -8131 29357 -7955
rect 29311 -8143 29357 -8131
rect 29429 -7955 29475 -7943
rect 29429 -8131 29435 -7955
rect 29469 -8131 29475 -7955
rect 29429 -8143 29475 -8131
rect 29547 -7955 29593 -7943
rect 29547 -8131 29553 -7955
rect 29587 -8131 29593 -7955
rect 29547 -8143 29593 -8131
rect 29665 -7955 29711 -7943
rect 29665 -8131 29671 -7955
rect 29705 -8131 29711 -7955
rect 29665 -8143 29711 -8131
rect 27624 -8202 28208 -8201
rect -638 -8817 13814 -8811
rect -638 -8903 -627 -8817
rect -528 -8903 13814 -8817
rect -638 -8911 13814 -8903
rect -258 -8912 13814 -8911
rect 13842 -8787 24463 -8706
rect 24501 -8211 28209 -8202
rect 24501 -8301 28112 -8211
rect 28196 -8301 28209 -8211
rect 28726 -8237 28762 -8143
rect 28962 -8237 28998 -8143
rect 29198 -8236 29234 -8143
rect 29360 -8191 29426 -8184
rect 29360 -8225 29376 -8191
rect 29410 -8225 29426 -8191
rect 29360 -8236 29426 -8225
rect 29198 -8237 29426 -8236
rect 28726 -8266 29426 -8237
rect 28726 -8267 29308 -8266
rect 24501 -8307 28209 -8301
rect 24501 -8308 28208 -8307
rect 24501 -8309 26686 -8308
rect 13842 -8788 19532 -8787
rect -535 -8951 416 -8950
rect -535 -8952 12857 -8951
rect 13842 -8952 13926 -8788
rect 24501 -8829 24657 -8309
rect 28846 -8380 28880 -8267
rect 29242 -8308 29308 -8267
rect 29242 -8342 29258 -8308
rect 29292 -8342 29308 -8308
rect 29242 -8349 29308 -8342
rect 29670 -8376 29705 -8143
rect 29895 -8376 29990 -7389
rect 30474 -7896 30508 -7112
rect 31187 -7174 31221 -7112
rect 30776 -7212 31518 -7174
rect 30586 -7383 30596 -7315
rect 30651 -7383 30661 -7315
rect 30776 -7336 30810 -7212
rect 31012 -7336 31046 -7212
rect 31248 -7336 31282 -7212
rect 31484 -7336 31518 -7212
rect 30770 -7348 30816 -7336
rect 30770 -7724 30776 -7348
rect 30810 -7724 30816 -7348
rect 30770 -7736 30816 -7724
rect 30888 -7348 30934 -7336
rect 30888 -7724 30894 -7348
rect 30928 -7724 30934 -7348
rect 30888 -7736 30934 -7724
rect 31006 -7348 31052 -7336
rect 31006 -7724 31012 -7348
rect 31046 -7724 31052 -7348
rect 31006 -7736 31052 -7724
rect 31124 -7348 31170 -7336
rect 31124 -7724 31130 -7348
rect 31164 -7724 31170 -7348
rect 31124 -7736 31170 -7724
rect 31242 -7348 31288 -7336
rect 31242 -7724 31248 -7348
rect 31282 -7724 31288 -7348
rect 31242 -7736 31288 -7724
rect 31360 -7348 31406 -7336
rect 31360 -7724 31366 -7348
rect 31400 -7724 31406 -7348
rect 31360 -7736 31406 -7724
rect 31478 -7348 31524 -7336
rect 31478 -7724 31484 -7348
rect 31518 -7724 31524 -7348
rect 31644 -7553 31718 -7541
rect 31640 -7644 31650 -7553
rect 31712 -7644 31722 -7553
rect 31644 -7656 31718 -7644
rect 31478 -7736 31524 -7724
rect 31890 -7895 31924 -7112
rect 32259 -7140 32295 -7046
rect 32495 -7140 32531 -7046
rect 32731 -7139 32767 -7046
rect 32893 -7094 32959 -7087
rect 32893 -7128 32909 -7094
rect 32943 -7128 32959 -7094
rect 32893 -7139 32959 -7128
rect 32731 -7140 32959 -7139
rect 32259 -7169 32959 -7140
rect 32259 -7170 32841 -7169
rect 31985 -7202 32061 -7197
rect 31982 -7258 31992 -7202
rect 32045 -7203 32061 -7202
rect 32045 -7258 32311 -7203
rect 31985 -7263 32311 -7258
rect 32106 -7305 32197 -7300
rect 32106 -7394 32116 -7305
rect 32189 -7394 32197 -7305
rect 32106 -7406 32197 -7394
rect 32143 -7800 32197 -7406
rect 32257 -7715 32311 -7263
rect 32379 -7283 32413 -7170
rect 32775 -7211 32841 -7170
rect 32775 -7245 32791 -7211
rect 32825 -7245 32841 -7211
rect 32775 -7252 32841 -7245
rect 33203 -7279 33238 -7046
rect 32849 -7283 33238 -7279
rect 32373 -7295 32419 -7283
rect 32373 -7671 32379 -7295
rect 32413 -7671 32419 -7295
rect 32373 -7683 32419 -7671
rect 32491 -7295 32537 -7283
rect 32491 -7671 32497 -7295
rect 32531 -7671 32537 -7295
rect 32491 -7683 32537 -7671
rect 32609 -7295 32655 -7283
rect 32609 -7671 32615 -7295
rect 32649 -7644 32655 -7295
rect 32726 -7295 32772 -7283
rect 32726 -7471 32732 -7295
rect 32766 -7471 32772 -7295
rect 32726 -7478 32772 -7471
rect 32844 -7294 33238 -7283
rect 32844 -7295 33081 -7294
rect 32844 -7471 32850 -7295
rect 32884 -7308 33081 -7295
rect 32884 -7471 32890 -7308
rect 33063 -7382 33081 -7308
rect 33223 -7382 33238 -7294
rect 33063 -7397 33238 -7382
rect 32726 -7483 32775 -7478
rect 32844 -7483 32890 -7471
rect 32732 -7644 32775 -7483
rect 32649 -7671 32775 -7644
rect 33069 -7553 33781 -7535
rect 33069 -7645 33079 -7553
rect 33223 -7645 33781 -7553
rect 33069 -7656 33781 -7645
rect 32609 -7683 32775 -7671
rect 32615 -7687 32775 -7683
rect 32257 -7721 32488 -7715
rect 32257 -7755 32438 -7721
rect 32472 -7755 32488 -7721
rect 32257 -7771 32488 -7755
rect 32540 -7721 32606 -7715
rect 32540 -7755 32556 -7721
rect 32590 -7755 32606 -7721
rect 32540 -7800 32606 -7755
rect 32143 -7808 32606 -7800
rect 32143 -7840 32607 -7808
rect 32699 -7824 32775 -7687
rect 32695 -7884 32705 -7824
rect 32767 -7884 32777 -7824
rect 31617 -7896 31924 -7895
rect 30474 -7901 30790 -7896
rect 31504 -7901 31924 -7896
rect 30474 -7912 30857 -7901
rect 30474 -7939 30806 -7912
rect 30474 -8068 30508 -7939
rect 30790 -7946 30806 -7939
rect 30840 -7946 30857 -7912
rect 30790 -7952 30857 -7946
rect 31437 -7912 31924 -7901
rect 32703 -7910 32773 -7884
rect 31437 -7946 31454 -7912
rect 31488 -7939 31924 -7912
rect 31488 -7946 31504 -7939
rect 31617 -7940 31924 -7939
rect 31437 -7952 31504 -7946
rect 30615 -7979 30671 -7967
rect 30615 -8013 30621 -7979
rect 30655 -7980 30671 -7979
rect 31728 -7980 31784 -7968
rect 30655 -7996 31122 -7980
rect 30655 -8013 31072 -7996
rect 30615 -8029 31072 -8013
rect 31056 -8030 31072 -8029
rect 31106 -8030 31122 -7996
rect 31056 -8037 31122 -8030
rect 31174 -7995 31744 -7980
rect 31174 -8029 31190 -7995
rect 31224 -8014 31744 -7995
rect 31778 -8014 31784 -7980
rect 31224 -8029 31784 -8014
rect 31174 -8039 31241 -8029
rect 31728 -8030 31784 -8029
rect 31890 -8068 31924 -7940
rect 30468 -8080 30514 -8068
rect 30468 -8256 30474 -8080
rect 30508 -8256 30514 -8080
rect 30468 -8268 30514 -8256
rect 30586 -8080 30632 -8068
rect 30586 -8256 30592 -8080
rect 30626 -8256 30632 -8080
rect 30586 -8268 30632 -8256
rect 30888 -8080 30934 -8068
rect 29316 -8380 29990 -8376
rect 28840 -8392 28886 -8380
rect -535 -8954 13926 -8952
rect -535 -8960 6335 -8954
rect -535 -9026 -510 -8960
rect -366 -9026 6335 -8960
rect 6427 -9026 13926 -8954
rect -535 -9035 13926 -9026
rect -258 -9036 13926 -9035
rect 12834 -9037 13926 -9036
rect 13954 -8911 24657 -8829
rect -938 -9085 416 -9084
rect 13954 -9085 14032 -8911
rect 24501 -8912 24657 -8911
rect 24706 -8518 25111 -8516
rect 24706 -8520 28404 -8518
rect 24706 -8527 28778 -8520
rect 24706 -8617 28281 -8527
rect 28365 -8617 28778 -8527
rect 24706 -8622 28778 -8617
rect 24706 -8623 28404 -8622
rect 24706 -8624 25111 -8623
rect 24706 -8952 24862 -8624
rect 28724 -8812 28778 -8622
rect 28840 -8768 28846 -8392
rect 28880 -8768 28886 -8392
rect 28840 -8780 28886 -8768
rect 28958 -8392 29004 -8380
rect 28958 -8768 28964 -8392
rect 28998 -8768 29004 -8392
rect 28958 -8780 29004 -8768
rect 29076 -8392 29122 -8380
rect 29076 -8768 29082 -8392
rect 29116 -8741 29122 -8392
rect 29193 -8392 29239 -8380
rect 29193 -8568 29199 -8392
rect 29233 -8568 29239 -8392
rect 29193 -8575 29239 -8568
rect 29311 -8392 29990 -8380
rect 29311 -8568 29317 -8392
rect 29351 -8405 29990 -8392
rect 29351 -8568 29357 -8405
rect 29601 -8485 29990 -8405
rect 29193 -8580 29242 -8575
rect 29311 -8580 29357 -8568
rect 30591 -8562 30625 -8268
rect 30888 -8456 30894 -8080
rect 30928 -8456 30934 -8080
rect 30888 -8468 30934 -8456
rect 31006 -8080 31052 -8068
rect 31006 -8456 31012 -8080
rect 31046 -8456 31052 -8080
rect 31006 -8468 31052 -8456
rect 31124 -8080 31170 -8068
rect 31124 -8456 31130 -8080
rect 31164 -8456 31170 -8080
rect 31124 -8468 31170 -8456
rect 31242 -8080 31288 -8068
rect 31242 -8456 31248 -8080
rect 31282 -8456 31288 -8080
rect 31242 -8468 31288 -8456
rect 31360 -8080 31406 -8068
rect 31360 -8456 31366 -8080
rect 31400 -8456 31406 -8080
rect 31766 -8080 31812 -8068
rect 31766 -8256 31772 -8080
rect 31806 -8256 31812 -8080
rect 31766 -8268 31812 -8256
rect 31884 -8080 31930 -8068
rect 31884 -8256 31890 -8080
rect 31924 -8256 31930 -8080
rect 31884 -8268 31930 -8256
rect 31360 -8468 31406 -8456
rect 31248 -8562 31282 -8468
rect 31772 -8562 31805 -8268
rect 29199 -8741 29242 -8580
rect 30591 -8594 31805 -8562
rect 29116 -8768 29242 -8741
rect 29076 -8780 29242 -8768
rect 29082 -8784 29242 -8780
rect 28724 -8818 28955 -8812
rect 28724 -8852 28905 -8818
rect 28939 -8852 28955 -8818
rect 28724 -8868 28955 -8852
rect 29007 -8818 29073 -8812
rect 29007 -8852 29023 -8818
rect 29057 -8852 29073 -8818
rect -938 -9100 14032 -9085
rect -938 -9171 -925 -9100
rect -811 -9171 14032 -9100
rect -938 -9186 14032 -9171
rect 14060 -8961 24862 -8952
rect 14060 -9029 19767 -8961
rect 19836 -9029 24862 -8961
rect 14060 -9036 24862 -9029
rect 24909 -8873 25065 -8871
rect 28593 -8873 28656 -8872
rect 24909 -8876 28668 -8873
rect 24909 -8951 28594 -8876
rect 28655 -8897 28668 -8876
rect 29007 -8897 29073 -8852
rect 28655 -8905 29073 -8897
rect 28655 -8937 29074 -8905
rect 29166 -8921 29242 -8784
rect 30957 -8618 31363 -8594
rect 30957 -8741 31069 -8618
rect 31243 -8741 31363 -8618
rect 30957 -8785 31363 -8741
rect 28655 -8951 28668 -8937
rect 24909 -8961 28668 -8951
rect -938 -9187 12916 -9186
rect -258 -9188 12916 -9187
rect -1123 -9223 -983 -9222
rect -1123 -9224 416 -9223
rect 1588 -9224 1794 -9222
rect 14060 -9224 14155 -9036
rect -1123 -9238 14155 -9224
rect -1123 -9304 1619 -9238
rect 1763 -9304 14155 -9238
rect -1123 -9325 14155 -9304
rect 14183 -9086 19039 -9085
rect 24909 -9086 25065 -8961
rect 29162 -8981 29172 -8921
rect 29234 -8981 29244 -8921
rect 14183 -9186 25065 -9086
rect -1123 -9326 -983 -9325
rect -258 -9326 12685 -9325
rect 14183 -9363 14273 -9186
rect 1325 -9383 14273 -9363
rect 1325 -9437 1333 -9383
rect 1428 -9437 14273 -9383
rect 1325 -9444 14273 -9437
rect 27889 -9274 28045 -9260
rect 27889 -9355 27908 -9274
rect 28025 -9355 28045 -9274
rect 27889 -9593 28045 -9355
<< via1 >>
rect 7024 5807 7084 5869
rect 13573 5806 13633 5868
rect 20227 5827 20287 5889
rect 7246 4657 7308 4665
rect 7246 4611 7252 4657
rect 7252 4611 7304 4657
rect 7304 4611 7308 4657
rect 7246 4605 7308 4611
rect -994 4273 -910 4331
rect -756 3943 -688 3946
rect -756 3898 -749 3943
rect -749 3898 -692 3943
rect -692 3898 -688 3943
rect -756 3894 -688 3898
rect 360 3907 420 3969
rect 3350 3730 3384 3762
rect 3384 3730 3451 3762
rect 3451 3730 3482 3762
rect 3350 3654 3482 3730
rect 5832 3780 5866 3816
rect 5866 3780 5933 3816
rect 5933 3780 5964 3816
rect 5832 3708 5964 3780
rect 582 2757 644 2765
rect 582 2711 588 2757
rect 588 2711 640 2757
rect 640 2711 644 2757
rect 582 2705 644 2711
rect 6233 3718 6289 3732
rect 6233 3684 6249 3718
rect 6249 3684 6283 3718
rect 6283 3684 6289 3718
rect 6233 3666 6289 3684
rect 6979 3782 7008 3816
rect 7008 3782 7075 3816
rect 7075 3782 7111 3816
rect 6979 3708 7111 3782
rect 5103 3594 5169 3610
rect 5103 3560 5119 3594
rect 5119 3560 5153 3594
rect 5153 3560 5169 3594
rect 5103 3544 5169 3560
rect 5769 2897 5868 2994
rect 3630 2690 3738 2723
rect 3630 2623 3725 2690
rect 3725 2623 3738 2690
rect 3630 2591 3738 2623
rect 2122 2013 2234 2119
rect 352 1322 412 1384
rect 2121 1005 2233 1007
rect 2121 901 2239 1005
rect 2127 899 2239 901
rect 5178 2319 5310 2416
rect 5178 2308 5211 2319
rect 5211 2308 5278 2319
rect 5278 2308 5310 2319
rect 2616 2030 2728 2136
rect 3364 2079 3396 2112
rect 3396 2079 3463 2112
rect 3463 2079 3496 2112
rect 3364 2004 3496 2079
rect 6925 2920 6990 2974
rect 13795 4656 13857 4664
rect 13795 4610 13801 4656
rect 13801 4610 13853 4656
rect 13853 4610 13857 4656
rect 13795 4604 13857 4610
rect 13229 4175 13286 4229
rect 20449 4677 20511 4685
rect 20449 4631 20455 4677
rect 20455 4631 20507 4677
rect 20507 4631 20511 4677
rect 20449 4625 20511 4631
rect 9899 3818 9933 3850
rect 9933 3818 10000 3850
rect 10000 3818 10031 3850
rect 9899 3742 10031 3818
rect 12381 3869 12416 3904
rect 12416 3869 12483 3904
rect 12483 3869 12513 3904
rect 12381 3796 12513 3869
rect 12782 3806 12838 3820
rect 12782 3772 12798 3806
rect 12798 3772 12832 3806
rect 12832 3772 12838 3806
rect 12782 3754 12838 3772
rect 13528 3871 13560 3904
rect 13560 3871 13627 3904
rect 13627 3871 13660 3904
rect 13528 3796 13660 3871
rect 11652 3682 11718 3698
rect 11652 3648 11668 3682
rect 11668 3648 11702 3682
rect 11702 3648 11718 3682
rect 11652 3632 11718 3648
rect 12318 2985 12417 3082
rect 10179 2772 10287 2811
rect 10179 2705 10271 2772
rect 10271 2705 10287 2772
rect 10179 2679 10287 2705
rect 6320 2321 6452 2414
rect 6320 2306 6349 2321
rect 6349 2306 6416 2321
rect 6416 2306 6452 2321
rect 8671 2101 8783 2207
rect 5177 1661 5309 1769
rect 7075 1737 7108 1769
rect 7108 1737 7175 1769
rect 7175 1737 7207 1769
rect 7075 1661 7207 1737
rect 2899 899 3017 1017
rect 3644 1040 3752 1073
rect 3644 973 3740 1040
rect 3740 973 3752 1040
rect 3644 941 3752 973
rect 2396 557 2489 636
rect -955 91 -868 195
rect -158 94 -81 190
rect 574 172 636 180
rect 574 126 580 172
rect 580 126 632 172
rect 632 126 636 172
rect 574 120 636 126
rect 3359 473 3394 508
rect 3394 473 3461 508
rect 3461 473 3491 508
rect 3359 400 3491 473
rect 5822 783 5885 799
rect 5822 749 5851 783
rect 5851 749 5885 783
rect 5822 733 5885 749
rect 3946 -295 4009 -243
rect 3639 -568 3747 -531
rect 3639 -635 3738 -568
rect 3738 -635 3747 -568
rect 3639 -663 3747 -635
rect 2901 -878 3013 -772
rect 5122 -721 5254 -627
rect 5122 -735 5151 -721
rect 5151 -735 5218 -721
rect 5218 -735 5254 -721
rect 7020 -735 7152 -627
rect 333 -1956 393 -1894
rect 3342 -2050 3372 -2018
rect 3372 -2050 3439 -2018
rect 3439 -2050 3474 -2018
rect 3342 -2126 3474 -2050
rect 5824 -1995 5852 -1964
rect 5852 -1995 5919 -1964
rect 5919 -1995 5956 -1964
rect 5824 -2072 5956 -1995
rect 6225 -2062 6281 -2048
rect 6225 -2096 6241 -2062
rect 6241 -2096 6275 -2062
rect 6275 -2096 6281 -2062
rect 6225 -2114 6281 -2096
rect 6971 -1998 7008 -1964
rect 7008 -1998 7075 -1964
rect 7075 -1998 7103 -1964
rect 6971 -2072 7103 -1998
rect 5095 -2186 5161 -2170
rect 5095 -2220 5111 -2186
rect 5111 -2220 5145 -2186
rect 5145 -2220 5161 -2186
rect 5095 -2236 5161 -2220
rect 555 -3106 617 -3098
rect 555 -3152 561 -3106
rect 561 -3152 613 -3106
rect 613 -3152 617 -3106
rect 555 -3158 617 -3152
rect 5761 -2883 5860 -2786
rect 3622 -3097 3730 -3057
rect 3622 -3164 3715 -3097
rect 3715 -3164 3730 -3097
rect 3622 -3189 3730 -3164
rect 2114 -3767 2226 -3661
rect 349 -4716 409 -4654
rect 5170 -3458 5302 -3364
rect 5170 -3472 5192 -3458
rect 5192 -3472 5259 -3458
rect 5259 -3472 5302 -3458
rect 2608 -3750 2720 -3644
rect 3356 -3703 3393 -3668
rect 3393 -3703 3460 -3668
rect 3460 -3703 3488 -3668
rect 3356 -3776 3488 -3703
rect 6917 -2860 6982 -2806
rect 11727 2415 11859 2504
rect 11727 2396 11756 2415
rect 11756 2396 11823 2415
rect 11823 2396 11859 2415
rect 9165 2118 9277 2224
rect 9913 2166 9947 2200
rect 9947 2166 10014 2200
rect 10014 2166 10045 2200
rect 9913 2092 10045 2166
rect 13474 3008 13539 3062
rect 14569 2996 14637 3071
rect 12869 2407 13001 2502
rect 12869 2394 12895 2407
rect 12895 2394 12962 2407
rect 12962 2394 13001 2407
rect 11726 1749 11858 1857
rect 13624 1824 13662 1857
rect 13662 1824 13729 1857
rect 13729 1824 13756 1857
rect 13624 1749 13756 1824
rect 9448 987 9566 1105
rect 10193 1122 10301 1161
rect 10193 1055 10289 1122
rect 10289 1055 10301 1122
rect 10193 1029 10301 1055
rect 8945 645 9038 724
rect 9908 566 9939 596
rect 9939 566 10006 596
rect 10006 566 10040 596
rect 9908 488 10040 566
rect 12371 871 12434 887
rect 12371 837 12400 871
rect 12400 837 12434 871
rect 12371 821 12434 837
rect 10495 -207 10558 -155
rect 10188 -479 10296 -443
rect 10188 -546 10286 -479
rect 10286 -546 10296 -479
rect 10188 -575 10296 -546
rect 9450 -790 9562 -684
rect 11671 -636 11803 -539
rect 11671 -647 11700 -636
rect 11700 -647 11767 -636
rect 11767 -647 11803 -636
rect 13569 -647 13701 -539
rect 14638 295 14758 384
rect 9893 -2052 9927 -2020
rect 9927 -2052 9994 -2020
rect 9994 -2052 10025 -2020
rect 9893 -2128 10025 -2052
rect 12375 -1999 12408 -1966
rect 12408 -1999 12475 -1966
rect 12475 -1999 12507 -1966
rect 12375 -2074 12507 -1999
rect 12776 -2064 12832 -2050
rect 12776 -2098 12792 -2064
rect 12792 -2098 12826 -2064
rect 12826 -2098 12832 -2064
rect 12776 -2116 12832 -2098
rect 13522 -1999 13556 -1966
rect 13556 -1999 13623 -1966
rect 13623 -1999 13654 -1966
rect 13522 -2074 13654 -1999
rect 11646 -2188 11712 -2172
rect 11646 -2222 11662 -2188
rect 11662 -2222 11696 -2188
rect 11696 -2222 11712 -2188
rect 11646 -2238 11712 -2222
rect 8012 -2872 8080 -2797
rect 12312 -2885 12411 -2788
rect 10173 -3103 10281 -3059
rect 10173 -3170 10265 -3103
rect 10265 -3170 10281 -3103
rect 10173 -3191 10281 -3170
rect 6312 -3463 6444 -3366
rect 6312 -3474 6345 -3463
rect 6345 -3474 6412 -3463
rect 6412 -3474 6444 -3463
rect 5169 -4119 5301 -4011
rect 7067 -4044 7099 -4011
rect 7099 -4044 7166 -4011
rect 7166 -4044 7199 -4011
rect 7067 -4119 7199 -4044
rect 2891 -4881 3009 -4763
rect 3636 -4747 3744 -4707
rect 3636 -4814 3723 -4747
rect 3723 -4814 3744 -4747
rect 3636 -4839 3744 -4814
rect 2388 -5223 2481 -5144
rect -760 -5537 -679 -5474
rect 571 -5866 633 -5858
rect 571 -5912 577 -5866
rect 577 -5912 629 -5866
rect 629 -5912 633 -5866
rect 571 -5918 633 -5912
rect 3351 -5302 3382 -5272
rect 3382 -5302 3449 -5272
rect 3449 -5302 3483 -5272
rect 3351 -5380 3483 -5302
rect 5814 -4997 5877 -4981
rect 5814 -5031 5843 -4997
rect 5843 -5031 5877 -4997
rect 5814 -5047 5877 -5031
rect 3938 -6075 4001 -6023
rect 3631 -6339 3739 -6311
rect 3631 -6406 3723 -6339
rect 3723 -6406 3739 -6339
rect 3631 -6443 3739 -6406
rect 2893 -6658 3005 -6552
rect 5114 -6507 5246 -6407
rect 5114 -6515 5144 -6507
rect 5144 -6515 5211 -6507
rect 5211 -6515 5246 -6507
rect 7012 -6515 7144 -6407
rect 8665 -3769 8777 -3663
rect 7281 -7229 7343 -7223
rect 7281 -7275 7287 -7229
rect 7287 -7275 7339 -7229
rect 7339 -7275 7343 -7229
rect 7281 -7283 7343 -7275
rect 6342 -7548 6418 -7462
rect 6573 -7680 6702 -7589
rect 11721 -3461 11853 -3366
rect 11721 -3474 11750 -3461
rect 11750 -3474 11817 -3461
rect 11817 -3474 11853 -3461
rect 9159 -3752 9271 -3646
rect 9907 -3696 9938 -3670
rect 9938 -3696 10005 -3670
rect 10005 -3696 10039 -3670
rect 9907 -3778 10039 -3696
rect 13468 -2862 13533 -2808
rect 16553 3748 16586 3782
rect 16586 3748 16653 3782
rect 16653 3748 16685 3782
rect 16553 3674 16685 3748
rect 19035 3804 19067 3836
rect 19067 3804 19134 3836
rect 19134 3804 19167 3836
rect 19035 3728 19167 3804
rect 19436 3738 19492 3752
rect 19436 3704 19452 3738
rect 19452 3704 19486 3738
rect 19486 3704 19492 3738
rect 19436 3686 19492 3704
rect 20182 3803 20214 3836
rect 20214 3803 20281 3836
rect 20281 3803 20314 3836
rect 20182 3728 20314 3803
rect 18306 3614 18372 3630
rect 18306 3580 18322 3614
rect 18322 3580 18356 3614
rect 18356 3580 18372 3614
rect 18306 3564 18372 3580
rect 18972 2917 19071 3014
rect 16833 2706 16941 2743
rect 16833 2639 16921 2706
rect 16921 2639 16941 2706
rect 16833 2611 16941 2639
rect 15324 1025 15436 1027
rect 15324 921 15442 1025
rect 15330 920 15442 921
rect 15330 919 15442 920
rect 18381 2343 18513 2436
rect 18381 2328 18409 2343
rect 18409 2328 18476 2343
rect 18476 2328 18513 2343
rect 15819 2050 15931 2156
rect 16567 2100 16601 2132
rect 16601 2100 16668 2132
rect 16668 2100 16699 2132
rect 16567 2024 16699 2100
rect 20128 2940 20193 2994
rect 23178 3817 23206 3850
rect 23206 3817 23273 3850
rect 23273 3817 23310 3850
rect 23178 3742 23310 3817
rect 25660 3869 25690 3904
rect 25690 3869 25757 3904
rect 25757 3869 25792 3904
rect 25660 3796 25792 3869
rect 26061 3806 26117 3820
rect 26061 3772 26077 3806
rect 26077 3772 26111 3806
rect 26111 3772 26117 3806
rect 26061 3754 26117 3772
rect 26807 3875 26839 3904
rect 26839 3875 26906 3904
rect 26906 3875 26939 3904
rect 26807 3796 26939 3875
rect 24931 3682 24997 3698
rect 24931 3648 24947 3682
rect 24947 3648 24981 3682
rect 24981 3648 24997 3682
rect 24931 3632 24997 3648
rect 25597 2985 25696 3082
rect 23458 2782 23566 2811
rect 23458 2715 23553 2782
rect 23553 2715 23566 2782
rect 23458 2679 23566 2715
rect 19523 2346 19655 2434
rect 19523 2326 19555 2346
rect 19555 2326 19622 2346
rect 19622 2326 19655 2346
rect 21950 2101 22062 2207
rect 18380 1681 18512 1789
rect 20278 1752 20308 1789
rect 20308 1752 20375 1789
rect 20375 1752 20410 1789
rect 20278 1681 20410 1752
rect 16102 919 16220 1037
rect 16847 1055 16955 1093
rect 16847 988 16938 1055
rect 16938 988 16955 1055
rect 16847 961 16955 988
rect 15599 577 15692 656
rect 16562 497 16596 528
rect 16596 497 16663 528
rect 16663 497 16694 528
rect 16562 420 16694 497
rect 19025 803 19088 819
rect 19025 769 19054 803
rect 19054 769 19088 803
rect 19025 753 19088 769
rect 17149 -275 17212 -223
rect 16842 -550 16950 -511
rect 16842 -617 16940 -550
rect 16940 -617 16950 -550
rect 16842 -643 16950 -617
rect 16104 -858 16216 -752
rect 18325 -702 18457 -607
rect 18325 -715 18349 -702
rect 18349 -715 18416 -702
rect 18416 -715 18457 -702
rect 20223 -715 20355 -607
rect 21276 -1003 21399 -994
rect 21276 -1102 21285 -1003
rect 21285 -1102 21391 -1003
rect 21391 -1102 21399 -1003
rect 21276 -1108 21399 -1102
rect 16548 -2055 16578 -2019
rect 16578 -2055 16645 -2019
rect 16645 -2055 16680 -2019
rect 16548 -2127 16680 -2055
rect 19030 -1995 19063 -1965
rect 19063 -1995 19130 -1965
rect 19130 -1995 19162 -1965
rect 19030 -2073 19162 -1995
rect 19431 -2063 19487 -2049
rect 19431 -2097 19447 -2063
rect 19447 -2097 19481 -2063
rect 19481 -2097 19487 -2063
rect 19431 -2115 19487 -2097
rect 20177 -1998 20212 -1965
rect 20212 -1998 20279 -1965
rect 20279 -1998 20309 -1965
rect 20177 -2073 20309 -1998
rect 18301 -2187 18367 -2171
rect 18301 -2221 18317 -2187
rect 18317 -2221 18351 -2187
rect 18351 -2221 18367 -2187
rect 18301 -2237 18367 -2221
rect 18967 -2884 19066 -2787
rect 16828 -3094 16936 -3058
rect 16828 -3161 16926 -3094
rect 16926 -3161 16936 -3094
rect 16828 -3190 16936 -3161
rect 12863 -3472 12995 -3368
rect 12863 -3476 12891 -3472
rect 12891 -3476 12958 -3472
rect 12958 -3476 12995 -3472
rect 15253 -3770 15457 -3657
rect 15405 -3771 15457 -3770
rect 11720 -4121 11852 -4013
rect 13618 -4045 13655 -4013
rect 13655 -4045 13722 -4013
rect 13722 -4045 13750 -4013
rect 13618 -4121 13750 -4045
rect 9442 -4883 9560 -4765
rect 10187 -4748 10295 -4709
rect 10187 -4815 10281 -4748
rect 10281 -4815 10295 -4748
rect 10187 -4841 10295 -4815
rect 8939 -5225 9032 -5146
rect 9902 -5307 9938 -5274
rect 9938 -5307 10005 -5274
rect 10005 -5307 10034 -5274
rect 9902 -5382 10034 -5307
rect 12365 -4999 12428 -4983
rect 12365 -5033 12394 -4999
rect 12394 -5033 12428 -4999
rect 12365 -5049 12428 -5033
rect 10489 -6077 10552 -6025
rect 10182 -6348 10290 -6313
rect 10182 -6415 10270 -6348
rect 10270 -6415 10290 -6348
rect 10182 -6445 10290 -6415
rect 9444 -6660 9556 -6554
rect 11665 -6508 11797 -6409
rect 11665 -6517 11692 -6508
rect 11692 -6517 11759 -6508
rect 11759 -6517 11797 -6508
rect 13563 -6517 13695 -6409
rect 13835 -7224 13897 -7218
rect 13835 -7270 13841 -7224
rect 13841 -7270 13893 -7224
rect 13893 -7270 13897 -7224
rect 13835 -7278 13897 -7270
rect 7059 -8487 7119 -8425
rect 18376 -3457 18508 -3365
rect 18376 -3473 18402 -3457
rect 18402 -3473 18469 -3457
rect 18469 -3473 18508 -3457
rect 15814 -3751 15926 -3645
rect 16562 -3701 16598 -3669
rect 16598 -3701 16665 -3669
rect 16665 -3701 16694 -3669
rect 16562 -3777 16694 -3701
rect 20123 -2861 20188 -2807
rect 25006 2402 25138 2504
rect 25006 2396 25030 2402
rect 25030 2396 25097 2402
rect 25097 2396 25138 2402
rect 22444 2118 22556 2224
rect 23192 2166 23229 2200
rect 23229 2166 23296 2200
rect 23296 2166 23324 2200
rect 23192 2092 23324 2166
rect 26753 3008 26818 3062
rect 27731 2996 27799 3071
rect 26148 2404 26280 2502
rect 26148 2394 26173 2404
rect 26173 2394 26240 2404
rect 26240 2394 26280 2404
rect 25005 1749 25137 1857
rect 26903 1821 26936 1857
rect 26936 1821 27003 1857
rect 27003 1821 27035 1857
rect 26903 1749 27035 1821
rect 22727 987 22845 1105
rect 23472 1121 23580 1161
rect 23472 1054 23558 1121
rect 23558 1054 23580 1121
rect 23472 1029 23580 1054
rect 22224 645 22317 724
rect 21745 218 21841 318
rect 23187 558 23221 596
rect 23221 558 23288 596
rect 23288 558 23319 596
rect 23187 488 23319 558
rect 25650 871 25713 887
rect 25650 837 25679 871
rect 25679 837 25713 871
rect 25650 821 25713 837
rect 23774 -207 23837 -155
rect 23467 -484 23575 -443
rect 23467 -551 23564 -484
rect 23564 -551 23575 -484
rect 23467 -575 23575 -551
rect 22729 -790 22841 -684
rect 24950 -636 25082 -539
rect 24950 -647 24980 -636
rect 24980 -647 25047 -636
rect 25047 -647 25082 -636
rect 26848 -647 26980 -539
rect 28880 5660 28940 5722
rect 31137 5617 31269 5651
rect 31137 5543 31269 5617
rect 32481 5252 32541 5314
rect 28225 4575 28304 4649
rect 28377 4439 28458 4535
rect 30334 4674 30401 4737
rect 29102 4510 29164 4518
rect 29102 4464 29108 4510
rect 29108 4464 29160 4510
rect 29160 4464 29164 4510
rect 29102 4458 29164 4464
rect 30334 4548 30401 4611
rect 28875 3089 28935 3151
rect 30594 4602 30649 4619
rect 30594 4568 30599 4602
rect 30599 4568 30633 4602
rect 30633 4568 30649 4602
rect 30594 4551 30649 4568
rect 31648 4290 31710 4381
rect 31990 4721 32043 4732
rect 31990 4687 31999 4721
rect 31999 4687 32033 4721
rect 32033 4687 32043 4721
rect 31990 4676 32043 4687
rect 32114 4540 32187 4629
rect 33103 4566 33215 4624
rect 32887 4295 32995 4376
rect 32703 4102 32765 4110
rect 32703 4056 32709 4102
rect 32709 4056 32761 4102
rect 32761 4056 32765 4102
rect 32703 4050 32765 4056
rect 31067 3307 31241 3316
rect 31067 3205 31086 3307
rect 31086 3205 31221 3307
rect 31221 3205 31241 3307
rect 31067 3193 31241 3205
rect 28524 2127 28606 2208
rect 29097 1939 29159 1947
rect 29097 1893 29103 1939
rect 29103 1893 29155 1939
rect 29155 1893 29159 1939
rect 29097 1887 29159 1893
rect 31139 1526 31271 1560
rect 31139 1452 31271 1526
rect 32483 1161 32543 1223
rect 30336 583 30403 646
rect 28875 56 28935 118
rect 28629 -780 28718 -693
rect 22385 -1003 22508 -994
rect 22385 -1102 22394 -1003
rect 22394 -1102 22500 -1003
rect 22500 -1102 22508 -1003
rect 22385 -1108 22508 -1102
rect 30336 457 30403 520
rect 29097 -1094 29159 -1086
rect 29097 -1140 29103 -1094
rect 29103 -1140 29155 -1094
rect 29155 -1140 29159 -1094
rect 29097 -1146 29159 -1140
rect 28946 -1864 29006 -1802
rect 23170 -2050 23202 -2018
rect 23202 -2050 23269 -2018
rect 23269 -2050 23302 -2018
rect 23170 -2126 23302 -2050
rect 25652 -2002 25681 -1964
rect 25681 -2002 25748 -1964
rect 25748 -2002 25784 -1964
rect 25652 -2072 25784 -2002
rect 26053 -2062 26109 -2048
rect 26053 -2096 26069 -2062
rect 26069 -2096 26103 -2062
rect 26103 -2096 26109 -2062
rect 26053 -2114 26109 -2096
rect 26799 -1996 26829 -1964
rect 26829 -1996 26896 -1964
rect 26896 -1996 26931 -1964
rect 26799 -2072 26931 -1996
rect 24923 -2186 24989 -2170
rect 24923 -2220 24939 -2186
rect 24939 -2220 24973 -2186
rect 24973 -2220 24989 -2186
rect 24923 -2236 24989 -2220
rect 21218 -2873 21286 -2798
rect 25589 -2883 25688 -2786
rect 23450 -3089 23558 -3057
rect 23450 -3156 23542 -3089
rect 23542 -3156 23558 -3089
rect 23450 -3189 23558 -3156
rect 19518 -3454 19650 -3367
rect 19518 -3475 19548 -3454
rect 19548 -3475 19615 -3454
rect 19615 -3475 19650 -3454
rect 18375 -4120 18507 -4012
rect 20273 -4043 20309 -4012
rect 20309 -4043 20376 -4012
rect 20376 -4043 20405 -4012
rect 20273 -4120 20405 -4043
rect 16097 -4882 16215 -4764
rect 16842 -4745 16950 -4708
rect 16842 -4812 16937 -4745
rect 16937 -4812 16950 -4745
rect 16842 -4840 16950 -4812
rect 15594 -5224 15687 -5145
rect 16557 -5309 16593 -5273
rect 16593 -5309 16660 -5273
rect 16660 -5309 16689 -5273
rect 16557 -5381 16689 -5309
rect 19020 -4998 19083 -4982
rect 19020 -5032 19049 -4998
rect 19049 -5032 19083 -4998
rect 19020 -5048 19083 -5032
rect 17144 -6076 17207 -6024
rect 16837 -6354 16945 -6312
rect 16837 -6421 16940 -6354
rect 16940 -6421 16945 -6354
rect 16837 -6444 16945 -6421
rect 15282 -6603 15384 -6591
rect 15282 -6671 15301 -6603
rect 15301 -6671 15371 -6603
rect 15371 -6671 15384 -6603
rect 15282 -6678 15384 -6671
rect 16099 -6659 16211 -6553
rect 18320 -6507 18452 -6408
rect 18320 -6516 18342 -6507
rect 18342 -6516 18409 -6507
rect 18409 -6516 18452 -6507
rect 20218 -6516 20350 -6408
rect 21942 -3767 22054 -3661
rect 20484 -7236 20546 -7230
rect 20484 -7282 20490 -7236
rect 20490 -7282 20542 -7236
rect 20542 -7282 20546 -7236
rect 20484 -7290 20546 -7282
rect 13613 -8482 13673 -8420
rect 19770 -7687 19839 -7598
rect 21941 -4775 22053 -4773
rect 21941 -4879 22059 -4775
rect 21947 -4881 22059 -4879
rect 24998 -3453 25130 -3364
rect 24998 -3472 25033 -3453
rect 25033 -3472 25100 -3453
rect 25100 -3472 25130 -3453
rect 22436 -3750 22548 -3644
rect 23184 -3700 23217 -3668
rect 23217 -3700 23284 -3668
rect 23284 -3700 23316 -3668
rect 23184 -3776 23316 -3700
rect 30596 511 30651 528
rect 30596 477 30601 511
rect 30601 477 30635 511
rect 30635 477 30651 511
rect 30596 460 30651 477
rect 31650 199 31712 290
rect 31992 630 32045 641
rect 31992 596 32001 630
rect 32001 596 32035 630
rect 32035 596 32045 630
rect 31992 585 32045 596
rect 32116 449 32189 538
rect 32932 198 33056 289
rect 32705 11 32767 19
rect 32705 -35 32711 11
rect 32711 -35 32763 11
rect 32763 -35 32767 11
rect 32705 -41 32767 -35
rect 31069 -784 31243 -775
rect 31069 -886 31088 -784
rect 31088 -886 31223 -784
rect 31223 -886 31243 -784
rect 31069 -898 31243 -886
rect 31139 -1969 31271 -1935
rect 31139 -2043 31271 -1969
rect 26745 -2860 26810 -2806
rect 28681 -2915 28767 -2814
rect 32483 -2334 32543 -2272
rect 28453 -3048 28538 -2988
rect 29168 -3014 29230 -3006
rect 29168 -3060 29174 -3014
rect 29174 -3060 29226 -3014
rect 29226 -3060 29230 -3014
rect 29168 -3066 29230 -3060
rect 30336 -3038 30403 -2975
rect 26140 -3462 26272 -3366
rect 26140 -3474 26167 -3462
rect 26167 -3474 26234 -3462
rect 26234 -3474 26272 -3462
rect 24997 -4119 25129 -4011
rect 26895 -4045 26930 -4011
rect 26930 -4045 26997 -4011
rect 26997 -4045 27027 -4011
rect 26895 -4119 27027 -4045
rect 22719 -4881 22837 -4763
rect 23464 -4738 23572 -4707
rect 23464 -4805 23560 -4738
rect 23560 -4805 23572 -4738
rect 23464 -4839 23572 -4805
rect 22216 -5223 22309 -5144
rect 23179 -5309 23214 -5272
rect 23214 -5309 23281 -5272
rect 23281 -5309 23311 -5272
rect 23179 -5380 23311 -5309
rect 25642 -4997 25705 -4981
rect 25642 -5031 25671 -4997
rect 25671 -5031 25705 -4997
rect 25642 -5047 25705 -5031
rect 28943 -4934 29003 -4872
rect 23766 -6075 23829 -6023
rect 23459 -6355 23567 -6311
rect 23459 -6422 23551 -6355
rect 23551 -6422 23567 -6355
rect 23459 -6443 23567 -6422
rect 22721 -6658 22833 -6552
rect 24942 -6501 25074 -6407
rect 24942 -6515 24970 -6501
rect 24970 -6515 25037 -6501
rect 25037 -6515 25074 -6501
rect 26840 -6515 26972 -6407
rect 27908 -5570 28025 -5489
rect 30596 -2984 30651 -2967
rect 30596 -3018 30601 -2984
rect 30601 -3018 30635 -2984
rect 30635 -3018 30651 -2984
rect 30596 -3035 30651 -3018
rect 31650 -3296 31712 -3205
rect 31992 -2865 32045 -2854
rect 31992 -2899 32001 -2865
rect 32001 -2899 32035 -2865
rect 32035 -2899 32045 -2865
rect 31992 -2910 32045 -2899
rect 32116 -3046 32189 -2957
rect 32705 -3484 32767 -3476
rect 32705 -3530 32711 -3484
rect 32711 -3530 32763 -3484
rect 32763 -3530 32767 -3484
rect 32705 -3536 32767 -3530
rect 31069 -4279 31243 -4270
rect 31069 -4381 31088 -4279
rect 31088 -4381 31223 -4279
rect 31223 -4381 31243 -4279
rect 31069 -4393 31243 -4381
rect 28283 -5898 28367 -5808
rect 33299 -3297 33409 -3206
rect 28717 -6019 28783 -5955
rect 29165 -6084 29227 -6076
rect 29165 -6130 29171 -6084
rect 29171 -6130 29223 -6084
rect 29223 -6130 29227 -6084
rect 29165 -6136 29227 -6130
rect 31139 -6317 31271 -6283
rect 31139 -6391 31271 -6317
rect 32483 -6682 32543 -6620
rect 30336 -7260 30402 -7197
rect 30402 -7260 30403 -7197
rect 30336 -7386 30403 -7323
rect 28697 -7558 28781 -7468
rect 20262 -8494 20322 -8432
rect 1487 -8774 1583 -8705
rect 6527 -8775 6627 -8701
rect 28950 -7779 29010 -7717
rect -627 -8903 -528 -8817
rect 28112 -8301 28196 -8211
rect 30596 -7332 30651 -7315
rect 30596 -7366 30601 -7332
rect 30601 -7366 30635 -7332
rect 30635 -7366 30651 -7332
rect 30596 -7383 30651 -7366
rect 31650 -7644 31712 -7553
rect 31992 -7213 32045 -7202
rect 31992 -7247 32001 -7213
rect 32001 -7247 32035 -7213
rect 32035 -7247 32045 -7213
rect 31992 -7258 32045 -7247
rect 32116 -7394 32189 -7305
rect 33081 -7382 33223 -7294
rect 33079 -7645 33223 -7553
rect 32705 -7832 32767 -7824
rect 32705 -7878 32711 -7832
rect 32711 -7878 32763 -7832
rect 32763 -7878 32767 -7832
rect 32705 -7884 32767 -7878
rect 6335 -9026 6427 -8954
rect 28281 -8617 28365 -8527
rect 19767 -9029 19836 -8961
rect 28594 -8951 28655 -8876
rect 31069 -8627 31243 -8618
rect 31069 -8729 31088 -8627
rect 31088 -8729 31223 -8627
rect 31223 -8729 31243 -8627
rect 31069 -8741 31243 -8729
rect 29172 -8929 29234 -8921
rect 29172 -8975 29178 -8929
rect 29178 -8975 29230 -8929
rect 29230 -8975 29234 -8929
rect 29172 -8981 29234 -8975
rect 1333 -9437 1428 -9383
rect 27908 -9355 28025 -9274
<< metal2 >>
rect 20227 5889 20287 5899
rect 7024 5869 7084 5879
rect 7024 5797 7084 5807
rect 13573 5868 13633 5878
rect 20227 5817 20287 5827
rect 13573 5796 13633 5806
rect 28880 5722 28940 5732
rect 28880 5650 28940 5660
rect 31126 5662 31279 5672
rect 31126 5523 31279 5533
rect 32481 5314 32541 5324
rect 32481 5242 32541 5252
rect 30334 4742 30401 4747
rect 30327 4737 32043 4742
rect 20449 4693 20511 4695
rect 20449 4685 20513 4693
rect 20511 4683 20513 4685
rect 7246 4673 7308 4675
rect 7246 4665 7310 4673
rect 7308 4663 7310 4665
rect 7246 4591 7310 4601
rect 13795 4672 13857 4674
rect 13795 4664 13859 4672
rect 13857 4662 13859 4664
rect 30327 4674 30334 4737
rect 30401 4732 32043 4737
rect 30401 4676 31990 4732
rect 30401 4674 32043 4676
rect 30327 4666 32043 4674
rect 30334 4664 30401 4666
rect 28225 4650 28304 4659
rect 20449 4611 20513 4621
rect 24276 4649 28304 4650
rect 13795 4590 13859 4600
rect 24276 4575 28225 4649
rect 32114 4629 32187 4639
rect 30334 4620 30401 4621
rect 30594 4620 32114 4629
rect 24276 4574 28304 4575
rect -780 4445 -664 4455
rect -790 4389 -780 4435
rect -664 4434 16113 4435
rect 24276 4434 24345 4574
rect 28225 4565 28304 4574
rect 30326 4619 32114 4620
rect 30326 4611 30594 4619
rect 30326 4548 30334 4611
rect 30401 4551 30594 4611
rect 30649 4551 32114 4619
rect 30401 4548 32114 4551
rect 28377 4535 28458 4545
rect 30326 4541 32114 4548
rect 30327 4540 30416 4541
rect 33090 4636 33228 4646
rect 33090 4544 33228 4554
rect 30334 4538 30401 4540
rect -664 4389 24345 4434
rect -790 4375 24345 4389
rect 24399 4527 24473 4528
rect 24399 4526 26733 4527
rect 24399 4445 28377 4526
rect 24399 4347 24473 4445
rect 26547 4444 28377 4445
rect 32114 4530 32187 4540
rect 29102 4526 29164 4528
rect 29102 4518 29166 4526
rect 29164 4516 29166 4518
rect 29102 4444 29166 4454
rect 28377 4429 28458 4439
rect -1000 4331 24473 4347
rect -1000 4273 -994 4331
rect -910 4281 24473 4331
rect 31648 4381 33005 4391
rect 31710 4376 33005 4381
rect 31710 4295 32887 4376
rect 32995 4295 33005 4376
rect 31710 4290 33005 4295
rect -910 4273 -899 4281
rect -1000 4262 -899 4273
rect 360 3969 420 3979
rect -756 3950 -688 3956
rect -767 3946 -676 3950
rect -767 3894 -756 3946
rect -688 3894 -676 3946
rect 360 3897 420 3907
rect -955 201 -868 205
rect -767 201 -676 3894
rect 582 2773 644 2775
rect 582 2765 646 2773
rect 644 2763 646 2765
rect 582 2691 646 2701
rect 352 1384 412 1394
rect 352 1312 412 1322
rect -964 195 -80 201
rect -964 91 -955 195
rect -868 190 -80 195
rect -868 94 -158 190
rect -81 94 -80 190
rect 574 188 636 190
rect 574 180 638 188
rect 636 178 638 180
rect 574 106 638 116
rect -868 91 -80 94
rect -964 84 -80 91
rect -955 81 -868 84
rect -773 -5466 -670 -5456
rect -773 -5555 -670 -5545
rect -637 -8817 -519 84
rect 333 -1894 393 -1884
rect 333 -1966 393 -1956
rect 555 -3090 617 -3088
rect 555 -3098 619 -3090
rect 617 -3100 619 -3098
rect 555 -3172 619 -3162
rect 349 -4654 409 -4644
rect 349 -4726 409 -4716
rect 571 -5850 633 -5848
rect 571 -5858 635 -5850
rect 633 -5860 635 -5858
rect 571 -5932 635 -5922
rect -637 -8903 -627 -8817
rect -528 -8903 -519 -8817
rect -637 -8911 -519 -8903
rect -627 -8913 -528 -8911
rect 1326 -9383 1433 4281
rect 31648 4280 33005 4290
rect 1474 4249 17633 4251
rect 28107 4249 28168 4250
rect 1474 4229 28199 4249
rect 1474 4175 13229 4229
rect 13286 4175 28199 4229
rect 1474 4156 28199 4175
rect 1474 4155 24458 4156
rect 1475 -8705 1593 4155
rect 28107 4029 28199 4156
rect 32703 4118 32765 4120
rect 32703 4110 32767 4118
rect 32765 4108 32767 4110
rect 32703 4036 32767 4046
rect 12370 3915 12523 3925
rect 9888 3861 10041 3871
rect 5821 3827 5974 3837
rect 3339 3773 3492 3783
rect 6968 3827 7121 3837
rect 6233 3732 6289 3742
rect 5821 3688 5974 3698
rect 3339 3634 3492 3644
rect 6108 3666 6233 3728
rect 6289 3666 6290 3728
rect 13517 3915 13670 3925
rect 12782 3820 12838 3830
rect 12370 3776 12523 3786
rect 9888 3722 10041 3732
rect 12657 3754 12782 3816
rect 12838 3754 12839 3816
rect 25649 3915 25802 3925
rect 23167 3861 23320 3871
rect 19024 3847 19177 3857
rect 13517 3776 13670 3786
rect 16542 3793 16695 3803
rect 11652 3705 11718 3708
rect 6968 3688 7121 3698
rect 10726 3698 11718 3705
rect 5103 3617 5169 3620
rect 4177 3610 5169 3617
rect 4177 3544 5103 3610
rect 3610 2581 3620 2734
rect 3749 2581 3759 2734
rect 2110 2146 2277 2147
rect 2617 2146 2733 2147
rect 2110 2136 2733 2146
rect 2110 2119 2616 2136
rect 2110 2013 2122 2119
rect 2234 2030 2616 2119
rect 2728 2030 2733 2136
rect 2234 2013 2733 2030
rect 2110 2004 2733 2013
rect 3353 2123 3506 2133
rect 3353 1984 3506 1994
rect 2109 1025 2274 1035
rect 2109 1024 2277 1025
rect 2899 1024 3017 1027
rect 2109 1017 3017 1024
rect 2109 1007 2899 1017
rect 2109 901 2121 1007
rect 2233 1005 2899 1007
rect 2109 899 2127 901
rect 2239 899 2899 1005
rect 3624 931 3634 1084
rect 3763 931 3773 1084
rect 2109 892 3017 899
rect 2115 890 3017 892
rect 2152 889 3017 890
rect 2386 645 2501 655
rect 2386 538 2501 548
rect 2896 -762 3012 889
rect 3348 519 3501 529
rect 3348 380 3501 390
rect 3946 -239 4009 -233
rect 4177 -239 4245 3544
rect 5103 3534 5169 3544
rect 6108 3005 6168 3666
rect 6233 3656 6289 3666
rect 6030 3004 6168 3005
rect 5768 2994 6168 3004
rect 5768 2897 5769 2994
rect 5868 2897 6168 2994
rect 10726 3632 11652 3698
rect 6925 2983 6990 2984
rect 8020 2983 8234 2993
rect 6924 2974 8058 2983
rect 6924 2920 6925 2974
rect 6990 2920 8058 2974
rect 6924 2909 8058 2920
rect 5768 2889 6168 2897
rect 8020 2908 8058 2909
rect 8203 2908 8234 2983
rect 8020 2895 8234 2908
rect 5768 2885 6077 2889
rect 10159 2669 10169 2822
rect 10298 2669 10308 2822
rect 5168 2426 5321 2436
rect 5168 2287 5321 2297
rect 6310 2424 6463 2434
rect 6310 2285 6463 2295
rect 8659 2234 8826 2235
rect 9166 2234 9282 2235
rect 8659 2224 9282 2234
rect 8659 2207 9165 2224
rect 8659 2101 8671 2207
rect 8783 2118 9165 2207
rect 9277 2118 9282 2224
rect 8783 2101 9282 2118
rect 8659 2092 9282 2101
rect 9902 2211 10055 2221
rect 9902 2072 10055 2082
rect 5166 1780 5319 1790
rect 5166 1641 5319 1651
rect 7064 1780 7217 1790
rect 7064 1641 7217 1651
rect 9448 1112 9566 1115
rect 8656 1105 9566 1112
rect 8656 987 9448 1105
rect 10173 1019 10183 1172
rect 10312 1019 10322 1172
rect 8656 977 9566 987
rect 5807 809 5885 819
rect 5807 713 5885 723
rect 3941 -243 4245 -239
rect 3941 -295 3946 -243
rect 4009 -295 4245 -243
rect 3941 -301 4245 -295
rect 3946 -305 4009 -301
rect 3619 -673 3629 -520
rect 3758 -673 3768 -520
rect 5112 -617 5265 -607
rect 5112 -756 5265 -746
rect 7010 -617 7163 -607
rect 7010 -756 7163 -746
rect 2896 -772 3013 -762
rect 2896 -878 2901 -772
rect 2896 -888 3013 -878
rect 2896 -889 3012 -888
rect 8656 -1207 8822 977
rect 8935 733 9050 743
rect 8935 626 9050 636
rect 9445 -674 9561 977
rect 9897 607 10050 617
rect 9897 468 10050 478
rect 10495 -151 10558 -145
rect 10726 -151 10794 3632
rect 11652 3622 11718 3632
rect 12657 3093 12717 3754
rect 12782 3744 12838 3754
rect 20171 3847 20324 3857
rect 19436 3752 19492 3762
rect 19024 3708 19177 3718
rect 16542 3654 16695 3664
rect 19311 3686 19436 3748
rect 19492 3686 19493 3748
rect 26796 3915 26949 3925
rect 26061 3820 26117 3830
rect 25649 3776 25802 3786
rect 23167 3722 23320 3732
rect 25936 3754 26061 3816
rect 26117 3754 26118 3816
rect 26796 3776 26949 3786
rect 20171 3708 20324 3718
rect 24931 3705 24997 3708
rect 24005 3698 24997 3705
rect 18306 3637 18372 3640
rect 12579 3092 12717 3093
rect 12317 3082 12717 3092
rect 12317 2985 12318 3082
rect 12417 2985 12717 3082
rect 17380 3630 18372 3637
rect 17380 3564 18306 3630
rect 13474 3071 13539 3072
rect 14569 3071 14637 3081
rect 13473 3062 14569 3071
rect 13473 3008 13474 3062
rect 13539 3008 14569 3062
rect 13473 2997 14569 3008
rect 14569 2986 14637 2996
rect 12317 2977 12717 2985
rect 12317 2973 12626 2977
rect 16813 2601 16823 2754
rect 16952 2601 16962 2754
rect 11717 2514 11870 2524
rect 11717 2375 11870 2385
rect 12859 2512 13012 2522
rect 12859 2373 13012 2383
rect 14638 2166 15582 2169
rect 15820 2166 15936 2167
rect 14638 2156 15936 2166
rect 14638 2050 15819 2156
rect 15931 2050 15936 2156
rect 14638 2024 15936 2050
rect 16556 2143 16709 2153
rect 11715 1868 11868 1878
rect 11715 1729 11868 1739
rect 13613 1868 13766 1878
rect 13613 1729 13766 1739
rect 12356 897 12434 907
rect 12356 801 12434 811
rect 14638 384 14758 2024
rect 16556 2004 16709 2014
rect 15312 1045 15477 1055
rect 15312 1044 15480 1045
rect 16102 1044 16220 1047
rect 15312 1037 16220 1044
rect 15312 1027 16102 1037
rect 15312 921 15324 1027
rect 15436 1025 16102 1027
rect 15312 919 15330 921
rect 15442 919 16102 1025
rect 16827 951 16837 1104
rect 16966 951 16976 1104
rect 15312 912 16220 919
rect 15318 910 16220 912
rect 15355 909 16220 910
rect 15589 665 15704 675
rect 15589 558 15704 568
rect 14638 285 14758 295
rect 10490 -155 10794 -151
rect 10490 -207 10495 -155
rect 10558 -207 10794 -155
rect 10490 -213 10794 -207
rect 10495 -217 10558 -213
rect 10168 -585 10178 -432
rect 10307 -585 10317 -432
rect 11661 -529 11814 -519
rect 11661 -668 11814 -658
rect 13559 -529 13712 -519
rect 13559 -668 13712 -658
rect 9445 -684 9562 -674
rect 9445 -790 9450 -684
rect 9445 -800 9562 -790
rect 16099 -742 16215 909
rect 16551 539 16704 549
rect 16551 400 16704 410
rect 17149 -219 17212 -213
rect 17380 -219 17448 3564
rect 18306 3554 18372 3564
rect 19311 3025 19371 3686
rect 19436 3676 19492 3686
rect 19233 3024 19371 3025
rect 18971 3014 19371 3024
rect 18971 2917 18972 3014
rect 19071 2917 19371 3014
rect 24005 3632 24931 3698
rect 20128 3003 20193 3004
rect 21192 3003 21289 3013
rect 20127 2994 21192 3003
rect 20127 2940 20128 2994
rect 20193 2940 21192 2994
rect 20127 2929 21192 2940
rect 21289 2929 21290 3003
rect 21192 2919 21289 2929
rect 18971 2909 19371 2917
rect 18971 2905 19280 2909
rect 23438 2669 23448 2822
rect 23577 2669 23587 2822
rect 18371 2446 18524 2456
rect 18371 2307 18524 2317
rect 19513 2444 19666 2454
rect 19513 2305 19666 2315
rect 21938 2234 22105 2235
rect 22445 2234 22561 2235
rect 21938 2224 22561 2234
rect 21938 2207 22444 2224
rect 21938 2101 21950 2207
rect 22062 2118 22444 2207
rect 22556 2118 22561 2224
rect 22062 2101 22561 2118
rect 21938 2092 22561 2101
rect 23181 2211 23334 2221
rect 23181 2072 23334 2082
rect 18369 1800 18522 1810
rect 18369 1661 18522 1671
rect 20267 1800 20420 1810
rect 20267 1661 20420 1671
rect 22727 1112 22845 1115
rect 21964 1105 22845 1112
rect 21964 987 22727 1105
rect 23452 1019 23462 1172
rect 23591 1019 23601 1172
rect 21964 978 22845 987
rect 19010 829 19088 839
rect 19010 733 19088 743
rect 21745 318 21841 328
rect 21745 208 21841 218
rect 17144 -223 17448 -219
rect 17144 -275 17149 -223
rect 17212 -275 17448 -223
rect 17144 -281 17448 -275
rect 17149 -285 17212 -281
rect 16822 -653 16832 -500
rect 16961 -653 16971 -500
rect 18315 -597 18468 -587
rect 18315 -736 18468 -726
rect 20213 -597 20366 -587
rect 20213 -736 20366 -726
rect 16099 -752 16216 -742
rect 9445 -801 9561 -800
rect 16099 -858 16104 -752
rect 16099 -868 16216 -858
rect 16099 -869 16215 -868
rect 21265 -986 21407 -976
rect 21265 -1129 21407 -1120
rect 8656 -1353 14570 -1207
rect 8745 -1358 14570 -1353
rect 21965 -1229 22075 978
rect 22106 977 22845 978
rect 22214 733 22329 743
rect 22214 626 22329 636
rect 22724 -674 22840 977
rect 23176 607 23329 617
rect 23176 468 23329 478
rect 23774 -151 23837 -145
rect 24005 -151 24073 3632
rect 24931 3622 24997 3632
rect 25936 3093 25996 3754
rect 26061 3744 26117 3754
rect 25858 3092 25996 3093
rect 25596 3082 25996 3092
rect 25596 2985 25597 3082
rect 25696 2985 25996 3082
rect 26753 3071 26818 3072
rect 27731 3071 27799 3081
rect 26752 3062 27731 3071
rect 26752 3008 26753 3062
rect 26818 3008 27731 3062
rect 26752 2997 27731 3008
rect 27731 2986 27799 2996
rect 25596 2977 25996 2985
rect 25596 2973 25905 2977
rect 24996 2514 25149 2524
rect 24996 2375 25149 2385
rect 26138 2512 26291 2522
rect 26138 2373 26291 2383
rect 28107 2219 28198 4029
rect 31048 3332 31259 3342
rect 31048 3165 31259 3175
rect 28875 3151 28935 3161
rect 28875 3079 28935 3089
rect 28107 2208 28606 2219
rect 28107 2127 28524 2208
rect 28107 2118 28606 2127
rect 28524 2117 28606 2118
rect 29097 1955 29159 1957
rect 29097 1947 29161 1955
rect 29159 1945 29161 1947
rect 24994 1868 25147 1878
rect 24994 1729 25147 1739
rect 26892 1868 27045 1878
rect 29097 1873 29161 1883
rect 26892 1729 27045 1739
rect 31128 1571 31281 1581
rect 31128 1432 31281 1442
rect 32483 1223 32543 1233
rect 32483 1151 32543 1161
rect 25635 897 25713 907
rect 25635 801 25713 811
rect 30336 651 30403 656
rect 30329 646 32045 651
rect 30329 583 30336 646
rect 30403 641 32045 646
rect 30403 585 31992 641
rect 30403 583 32045 585
rect 30329 575 32045 583
rect 30336 573 30403 575
rect 32116 538 32189 548
rect 30336 529 30403 530
rect 30596 529 32116 538
rect 30328 528 32116 529
rect 30328 520 30596 528
rect 30328 457 30336 520
rect 30403 460 30596 520
rect 30651 460 32116 528
rect 30403 457 32116 460
rect 30328 450 32116 457
rect 30329 449 30418 450
rect 30336 447 30403 449
rect 32116 439 32189 449
rect 31650 290 33069 300
rect 31712 289 33069 290
rect 31712 199 32932 289
rect 31650 198 32932 199
rect 33056 198 33069 289
rect 31650 189 33069 198
rect 32932 188 33056 189
rect 28875 118 28935 128
rect 28875 46 28935 56
rect 32705 27 32767 29
rect 32705 19 32769 27
rect 32767 17 32769 19
rect 32705 -55 32769 -45
rect 23769 -155 24073 -151
rect 23769 -207 23774 -155
rect 23837 -207 24073 -155
rect 23769 -213 24073 -207
rect 23774 -217 23837 -213
rect 23447 -585 23457 -432
rect 23586 -585 23596 -432
rect 24940 -529 25093 -519
rect 24940 -668 25093 -658
rect 26838 -529 26991 -519
rect 26838 -668 26991 -658
rect 22724 -684 22841 -674
rect 22724 -790 22729 -684
rect 28629 -692 28718 -683
rect 22724 -800 22841 -790
rect 28113 -693 28718 -692
rect 28113 -780 28629 -693
rect 28113 -784 28718 -780
rect 22724 -801 22840 -800
rect 22374 -986 22516 -976
rect 22374 -1130 22516 -1120
rect 5813 -1953 5966 -1943
rect 3331 -2007 3484 -1997
rect 6960 -1953 7113 -1943
rect 6225 -2048 6281 -2038
rect 5813 -2092 5966 -2082
rect 3331 -2146 3484 -2136
rect 6100 -2114 6225 -2052
rect 6281 -2114 6282 -2052
rect 12364 -1955 12517 -1945
rect 6960 -2092 7113 -2082
rect 9882 -2009 10035 -1999
rect 5095 -2163 5161 -2160
rect 4169 -2170 5161 -2163
rect 4169 -2236 5095 -2170
rect 3602 -3199 3612 -3046
rect 3741 -3199 3751 -3046
rect 2102 -3634 2269 -3633
rect 2609 -3634 2725 -3633
rect 2102 -3644 2725 -3634
rect 2102 -3661 2608 -3644
rect 2102 -3767 2114 -3661
rect 2226 -3750 2608 -3661
rect 2720 -3750 2725 -3644
rect 2226 -3767 2725 -3750
rect 2102 -3776 2725 -3767
rect 3345 -3657 3498 -3647
rect 3345 -3796 3498 -3786
rect 1998 -4745 2232 -4740
rect 1998 -4750 2266 -4745
rect 2232 -4755 2266 -4750
rect 2232 -4756 2269 -4755
rect 2891 -4756 3009 -4753
rect 2232 -4763 3009 -4756
rect 2232 -4881 2891 -4763
rect 3616 -4849 3626 -4696
rect 3755 -4849 3765 -4696
rect 2232 -4887 3009 -4881
rect 1998 -4891 3009 -4887
rect 1998 -4897 2232 -4891
rect 2378 -5135 2493 -5125
rect 2378 -5242 2493 -5232
rect 2888 -6542 3004 -4891
rect 3340 -5261 3493 -5251
rect 3340 -5400 3493 -5390
rect 3938 -6019 4001 -6013
rect 4169 -6019 4237 -2236
rect 5095 -2246 5161 -2236
rect 6100 -2775 6160 -2114
rect 6225 -2124 6281 -2114
rect 13511 -1955 13664 -1945
rect 12776 -2050 12832 -2040
rect 12364 -2094 12517 -2084
rect 9882 -2148 10035 -2138
rect 12651 -2116 12776 -2054
rect 12832 -2116 12833 -2054
rect 13511 -2094 13664 -2084
rect 11646 -2165 11712 -2162
rect 6022 -2776 6160 -2775
rect 5760 -2786 6160 -2776
rect 5760 -2883 5761 -2786
rect 5860 -2883 6160 -2786
rect 10720 -2172 11712 -2165
rect 10720 -2238 11646 -2172
rect 6917 -2797 6982 -2796
rect 8012 -2797 8080 -2787
rect 6916 -2806 8012 -2797
rect 6916 -2860 6917 -2806
rect 6982 -2860 8012 -2806
rect 6916 -2871 8012 -2860
rect 8012 -2882 8080 -2872
rect 5760 -2891 6160 -2883
rect 5760 -2895 6069 -2891
rect 10153 -3201 10163 -3048
rect 10292 -3201 10302 -3048
rect 5160 -3354 5313 -3344
rect 5160 -3493 5313 -3483
rect 6302 -3356 6455 -3346
rect 6302 -3495 6455 -3485
rect 9160 -3636 9276 -3635
rect 8899 -3639 9276 -3636
rect 8653 -3646 9276 -3639
rect 8653 -3663 9159 -3646
rect 8653 -3769 8665 -3663
rect 8777 -3752 9159 -3663
rect 9271 -3752 9276 -3646
rect 8777 -3769 9276 -3752
rect 8653 -3778 9276 -3769
rect 9896 -3659 10049 -3649
rect 9896 -3798 10049 -3788
rect 5158 -4000 5311 -3990
rect 5158 -4139 5311 -4129
rect 7056 -4000 7209 -3990
rect 7056 -4139 7209 -4129
rect 8633 -4757 8856 -4747
rect 9442 -4758 9560 -4755
rect 8856 -4765 9560 -4758
rect 8856 -4883 9442 -4765
rect 10167 -4851 10177 -4698
rect 10306 -4851 10316 -4698
rect 8856 -4893 9560 -4883
rect 8633 -4903 8856 -4893
rect 5799 -4971 5877 -4961
rect 5799 -5067 5877 -5057
rect 8929 -5137 9044 -5127
rect 8929 -5244 9044 -5234
rect 3933 -6023 4237 -6019
rect 3933 -6075 3938 -6023
rect 4001 -6075 4237 -6023
rect 3933 -6081 4237 -6075
rect 3938 -6085 4001 -6081
rect 3611 -6453 3621 -6300
rect 3750 -6453 3760 -6300
rect 5104 -6397 5257 -6387
rect 5104 -6536 5257 -6526
rect 7002 -6397 7155 -6387
rect 7002 -6536 7155 -6526
rect 2888 -6552 3005 -6542
rect 2888 -6658 2893 -6552
rect 2888 -6668 3005 -6658
rect 9439 -6544 9555 -4893
rect 9891 -5263 10044 -5253
rect 9891 -5402 10044 -5392
rect 10489 -6021 10552 -6015
rect 10720 -6021 10788 -2238
rect 11646 -2248 11712 -2238
rect 12651 -2777 12711 -2116
rect 12776 -2126 12832 -2116
rect 12573 -2778 12711 -2777
rect 12311 -2788 12711 -2778
rect 12311 -2885 12312 -2788
rect 12411 -2885 12711 -2788
rect 13468 -2799 13533 -2798
rect 14436 -2799 14566 -1358
rect 21965 -1361 27874 -1229
rect 21965 -1362 22069 -1361
rect 27745 -1385 27874 -1361
rect 27745 -1474 27875 -1385
rect 19019 -1954 19172 -1944
rect 16537 -2008 16690 -1998
rect 20166 -1954 20319 -1944
rect 19431 -2049 19487 -2039
rect 19019 -2093 19172 -2083
rect 16537 -2147 16690 -2137
rect 19306 -2115 19431 -2053
rect 19487 -2115 19488 -2053
rect 25641 -1953 25794 -1943
rect 20166 -2093 20319 -2083
rect 23159 -2007 23312 -1997
rect 18301 -2164 18367 -2161
rect 13467 -2808 14566 -2799
rect 13467 -2862 13468 -2808
rect 13533 -2862 14566 -2808
rect 13467 -2873 14566 -2862
rect 14436 -2876 14566 -2873
rect 17375 -2171 18367 -2164
rect 17375 -2237 18301 -2171
rect 12311 -2893 12711 -2885
rect 12311 -2897 12620 -2893
rect 16808 -3200 16818 -3047
rect 16947 -3200 16957 -3047
rect 11711 -3356 11864 -3346
rect 11711 -3495 11864 -3485
rect 12853 -3358 13006 -3348
rect 12853 -3497 13006 -3487
rect 15241 -3634 15407 -3632
rect 15241 -3635 15475 -3634
rect 15815 -3635 15931 -3634
rect 15241 -3645 15931 -3635
rect 15241 -3657 15814 -3645
rect 15241 -3770 15253 -3657
rect 15457 -3751 15814 -3657
rect 15926 -3751 15931 -3645
rect 15241 -3771 15405 -3770
rect 15457 -3771 15931 -3751
rect 15241 -3777 15931 -3771
rect 16551 -3658 16704 -3648
rect 15241 -3778 15465 -3777
rect 16551 -3797 16704 -3787
rect 11709 -4002 11862 -3992
rect 11709 -4141 11862 -4131
rect 13607 -4002 13760 -3992
rect 13607 -4141 13760 -4131
rect 15307 -4756 15472 -4746
rect 15307 -4757 15475 -4756
rect 16097 -4757 16215 -4754
rect 15307 -4764 16215 -4757
rect 15307 -4772 16097 -4764
rect 15307 -4884 15314 -4772
rect 15458 -4882 16097 -4772
rect 16822 -4850 16832 -4697
rect 16961 -4850 16971 -4697
rect 15458 -4884 16215 -4882
rect 15307 -4889 16215 -4884
rect 15313 -4891 16215 -4889
rect 15314 -4892 16215 -4891
rect 15314 -4894 15458 -4892
rect 12350 -4973 12428 -4963
rect 12350 -5069 12428 -5059
rect 15584 -5136 15699 -5126
rect 15584 -5243 15699 -5233
rect 10484 -6025 10788 -6021
rect 10484 -6077 10489 -6025
rect 10552 -6077 10788 -6025
rect 10484 -6083 10788 -6077
rect 10489 -6087 10552 -6083
rect 10162 -6455 10172 -6302
rect 10301 -6455 10311 -6302
rect 11655 -6399 11808 -6389
rect 11655 -6538 11808 -6528
rect 13553 -6399 13706 -6389
rect 13553 -6538 13706 -6528
rect 16094 -6543 16210 -4892
rect 16546 -5262 16699 -5252
rect 16546 -5401 16699 -5391
rect 17144 -6020 17207 -6014
rect 17375 -6020 17443 -2237
rect 18301 -2247 18367 -2237
rect 19306 -2776 19366 -2115
rect 19431 -2125 19487 -2115
rect 26788 -1953 26941 -1943
rect 26053 -2048 26109 -2038
rect 25641 -2092 25794 -2082
rect 23159 -2146 23312 -2136
rect 25928 -2114 26053 -2052
rect 26109 -2114 26110 -2052
rect 26788 -2092 26941 -2082
rect 24923 -2163 24989 -2160
rect 19228 -2777 19366 -2776
rect 18966 -2787 19366 -2777
rect 18966 -2884 18967 -2787
rect 19066 -2884 19366 -2787
rect 23997 -2170 24989 -2163
rect 23997 -2236 24923 -2170
rect 20123 -2798 20188 -2797
rect 21218 -2798 21286 -2788
rect 20122 -2807 21218 -2798
rect 20122 -2861 20123 -2807
rect 20188 -2861 21218 -2807
rect 20122 -2872 21218 -2861
rect 21218 -2883 21286 -2873
rect 18966 -2892 19366 -2884
rect 18966 -2896 19275 -2892
rect 23430 -3199 23440 -3046
rect 23569 -3199 23579 -3046
rect 18366 -3355 18519 -3345
rect 18366 -3494 18519 -3484
rect 19508 -3357 19661 -3347
rect 19508 -3496 19661 -3486
rect 22437 -3634 22553 -3633
rect 21930 -3644 22553 -3634
rect 21930 -3661 22436 -3644
rect 21930 -3767 21942 -3661
rect 22054 -3750 22436 -3661
rect 22548 -3750 22553 -3644
rect 22054 -3767 22553 -3750
rect 21930 -3776 22553 -3767
rect 23173 -3657 23326 -3647
rect 23173 -3796 23326 -3786
rect 18364 -4001 18517 -3991
rect 18364 -4140 18517 -4130
rect 20262 -4001 20415 -3991
rect 20262 -4140 20415 -4130
rect 21929 -4755 22094 -4745
rect 21929 -4756 22097 -4755
rect 22719 -4756 22837 -4753
rect 21929 -4763 22837 -4756
rect 21929 -4773 22719 -4763
rect 21929 -4879 21941 -4773
rect 22053 -4775 22719 -4773
rect 21929 -4881 21947 -4879
rect 22059 -4881 22719 -4775
rect 23444 -4849 23454 -4696
rect 23583 -4849 23593 -4696
rect 21929 -4888 22837 -4881
rect 21935 -4890 22837 -4888
rect 21972 -4891 22837 -4890
rect 19005 -4972 19083 -4962
rect 19005 -5068 19083 -5058
rect 22206 -5135 22321 -5125
rect 22206 -5242 22321 -5232
rect 17139 -6024 17443 -6020
rect 17139 -6076 17144 -6024
rect 17207 -6076 17443 -6024
rect 17139 -6082 17443 -6076
rect 17144 -6086 17207 -6082
rect 16817 -6454 16827 -6301
rect 16956 -6454 16966 -6301
rect 18310 -6398 18463 -6388
rect 18310 -6537 18463 -6527
rect 20208 -6398 20361 -6388
rect 20208 -6537 20361 -6527
rect 22716 -6542 22832 -4891
rect 23168 -5261 23321 -5251
rect 23168 -5400 23321 -5390
rect 23766 -6019 23829 -6013
rect 23997 -6019 24065 -2236
rect 24923 -2246 24989 -2236
rect 25928 -2775 25988 -2114
rect 26053 -2124 26109 -2114
rect 25850 -2776 25988 -2775
rect 25588 -2786 25988 -2776
rect 25588 -2883 25589 -2786
rect 25688 -2883 25988 -2786
rect 26745 -2797 26810 -2796
rect 27745 -2797 27876 -1474
rect 26744 -2806 27876 -2797
rect 26744 -2860 26745 -2806
rect 26810 -2860 27876 -2806
rect 26744 -2871 27876 -2860
rect 27745 -2873 27876 -2871
rect 27840 -2874 27876 -2873
rect 25588 -2891 25988 -2883
rect 25588 -2895 25897 -2891
rect 24988 -3354 25141 -3344
rect 24988 -3493 25141 -3483
rect 26130 -3356 26283 -3346
rect 26130 -3495 26283 -3485
rect 24986 -4000 25139 -3990
rect 24986 -4139 25139 -4129
rect 26884 -4000 27037 -3990
rect 26884 -4139 27037 -4129
rect 25627 -4971 25705 -4961
rect 25627 -5067 25705 -5057
rect 27900 -5483 28032 -5473
rect 27900 -5589 28032 -5579
rect 23761 -6023 24065 -6019
rect 23761 -6075 23766 -6023
rect 23829 -6075 24065 -6023
rect 28113 -5942 28210 -784
rect 28629 -790 28718 -784
rect 31050 -759 31261 -749
rect 31050 -926 31261 -916
rect 29097 -1078 29159 -1076
rect 29097 -1086 29161 -1078
rect 29159 -1088 29161 -1086
rect 29097 -1160 29161 -1150
rect 28946 -1802 29006 -1792
rect 28946 -1874 29006 -1864
rect 31128 -1924 31281 -1914
rect 31128 -2063 31281 -2053
rect 32483 -2272 32543 -2262
rect 32483 -2344 32543 -2334
rect 28681 -2814 28767 -2804
rect 30329 -2837 30422 -2833
rect 28681 -2925 28767 -2915
rect 30299 -2843 30436 -2837
rect 30299 -2920 30329 -2843
rect 30422 -2844 30436 -2843
rect 30422 -2854 32045 -2844
rect 30422 -2910 31992 -2854
rect 30422 -2920 32045 -2910
rect 30299 -2927 30436 -2920
rect 30329 -2930 30422 -2927
rect 32116 -2957 32189 -2947
rect 30336 -2966 30403 -2965
rect 30596 -2966 32116 -2957
rect 30328 -2967 32116 -2966
rect 30328 -2975 30596 -2967
rect 28453 -2988 28538 -2978
rect 28453 -3058 28538 -3048
rect 29168 -2998 29230 -2996
rect 29168 -3006 29232 -2998
rect 29230 -3008 29232 -3006
rect 30328 -3038 30336 -2975
rect 30403 -3035 30596 -2975
rect 30651 -3035 32116 -2967
rect 30403 -3038 32116 -3035
rect 30328 -3045 32116 -3038
rect 30329 -3046 30418 -3045
rect 30336 -3048 30403 -3046
rect 32116 -3056 32189 -3046
rect 29168 -3080 29232 -3070
rect 32943 -3195 33425 -3194
rect 31650 -3205 33425 -3195
rect 31712 -3206 33425 -3205
rect 31712 -3296 33299 -3206
rect 31650 -3297 33299 -3296
rect 33409 -3297 33425 -3206
rect 31650 -3306 33425 -3297
rect 33299 -3307 33409 -3306
rect 32705 -3468 32767 -3466
rect 32705 -3476 32769 -3468
rect 32767 -3478 32769 -3476
rect 32705 -3550 32769 -3540
rect 31050 -4254 31261 -4244
rect 31050 -4421 31261 -4411
rect 28943 -4872 29003 -4862
rect 28943 -4944 29003 -4934
rect 28283 -5808 28367 -5798
rect 28283 -5907 28367 -5898
rect 28113 -5944 28751 -5942
rect 28113 -5945 28776 -5944
rect 28113 -5955 28783 -5945
rect 28113 -6019 28717 -5955
rect 28113 -6029 28783 -6019
rect 29894 -5972 33430 -5884
rect 28113 -6031 28708 -6029
rect 23761 -6081 24065 -6075
rect 29165 -6068 29227 -6066
rect 29165 -6076 29229 -6068
rect 29227 -6078 29229 -6076
rect 23766 -6085 23829 -6081
rect 29165 -6150 29229 -6140
rect 23439 -6453 23449 -6300
rect 23578 -6453 23588 -6300
rect 24932 -6397 25085 -6387
rect 24932 -6536 25085 -6526
rect 26830 -6397 26983 -6387
rect 26830 -6536 26983 -6526
rect 9439 -6554 9556 -6544
rect 9439 -6660 9444 -6554
rect 16094 -6553 16211 -6543
rect 2888 -6669 3004 -6668
rect 9439 -6670 9556 -6660
rect 15255 -6591 15423 -6581
rect 9439 -6671 9555 -6670
rect 15255 -6678 15282 -6591
rect 15384 -6678 15423 -6591
rect 16094 -6659 16099 -6553
rect 16094 -6669 16211 -6659
rect 22716 -6552 22833 -6542
rect 22716 -6658 22721 -6552
rect 22716 -6668 22833 -6658
rect 22716 -6669 22832 -6668
rect 16094 -6670 16210 -6669
rect 15255 -6926 15423 -6678
rect 29894 -6926 29988 -5972
rect 31128 -6272 31281 -6262
rect 31128 -6411 31281 -6401
rect 32483 -6620 32543 -6610
rect 32483 -6692 32543 -6682
rect 15255 -7100 29988 -6926
rect 15354 -7101 29988 -7100
rect 30336 -7192 30403 -7187
rect 30329 -7197 32045 -7192
rect 7281 -7219 7345 -7209
rect 7343 -7283 7345 -7281
rect 7281 -7291 7345 -7283
rect 13835 -7214 13899 -7204
rect 13897 -7278 13899 -7276
rect 13835 -7286 13899 -7278
rect 20484 -7226 20548 -7216
rect 13835 -7288 13897 -7286
rect 30329 -7260 30336 -7197
rect 30403 -7202 32045 -7197
rect 30403 -7258 31992 -7202
rect 30403 -7260 32045 -7258
rect 30329 -7268 32045 -7260
rect 30336 -7270 30403 -7268
rect 33081 -7285 33223 -7284
rect 33316 -7285 33430 -5972
rect 20546 -7290 20548 -7288
rect 7281 -7293 7343 -7291
rect 20484 -7298 20548 -7290
rect 33068 -7294 33430 -7285
rect 20484 -7300 20546 -7298
rect 32116 -7305 32189 -7295
rect 30336 -7314 30403 -7313
rect 30596 -7314 32116 -7305
rect 30328 -7315 32116 -7314
rect 30328 -7323 30596 -7315
rect 30328 -7386 30336 -7323
rect 30403 -7383 30596 -7323
rect 30651 -7383 32116 -7315
rect 30403 -7386 32116 -7383
rect 30328 -7393 32116 -7386
rect 30329 -7394 30418 -7393
rect 33068 -7382 33081 -7294
rect 33223 -7382 33430 -7294
rect 33068 -7393 33430 -7382
rect 30336 -7396 30403 -7394
rect 32116 -7404 32189 -7394
rect 6342 -7454 6418 -7452
rect 1475 -8774 1487 -8705
rect 1583 -8774 1593 -8705
rect 1475 -8780 1593 -8774
rect 6335 -7462 6427 -7454
rect 6335 -7548 6342 -7462
rect 6418 -7548 6427 -7462
rect 1487 -8784 1583 -8780
rect 6335 -8954 6427 -7548
rect 28697 -7468 28781 -7458
rect 28697 -7568 28781 -7558
rect 31650 -7553 33223 -7543
rect 6522 -7589 6702 -7579
rect 6522 -7680 6573 -7589
rect 19770 -7598 19839 -7588
rect 6522 -7690 6702 -7680
rect 19762 -7687 19770 -7598
rect 19839 -7687 19840 -7598
rect 31712 -7644 33079 -7553
rect 31650 -7645 33079 -7644
rect 31650 -7654 33223 -7645
rect 33079 -7655 33223 -7654
rect 6522 -8701 6631 -7690
rect 7059 -8425 7119 -8415
rect 7059 -8497 7119 -8487
rect 13613 -8420 13673 -8410
rect 13613 -8492 13673 -8482
rect 6522 -8775 6527 -8701
rect 6627 -8775 6631 -8701
rect 6522 -8781 6631 -8775
rect 6527 -8785 6627 -8781
rect 6335 -9036 6427 -9026
rect 19762 -8846 19840 -7687
rect 28950 -7717 29010 -7707
rect 28950 -7789 29010 -7779
rect 32705 -7816 32767 -7814
rect 32705 -7824 32769 -7816
rect 32767 -7826 32769 -7824
rect 32705 -7898 32769 -7888
rect 28112 -8211 28196 -8201
rect 28112 -8311 28196 -8301
rect 20262 -8432 20322 -8422
rect 20262 -8504 20322 -8494
rect 28281 -8527 28365 -8517
rect 28281 -8627 28365 -8617
rect 31050 -8602 31261 -8592
rect 31050 -8769 31261 -8759
rect 19762 -8961 19841 -8846
rect 28594 -8876 28655 -8866
rect 28594 -8961 28655 -8951
rect 29172 -8913 29234 -8911
rect 29172 -8921 29236 -8913
rect 29234 -8923 29236 -8921
rect 19762 -9029 19767 -8961
rect 19836 -9029 19841 -8961
rect 29172 -8995 29236 -8985
rect 19762 -9032 19841 -9029
rect 19767 -9039 19836 -9032
rect 27900 -9268 28032 -9258
rect 27900 -9374 28032 -9364
rect 1326 -9437 1333 -9383
rect 1428 -9389 1433 -9383
rect 1428 -9437 1432 -9389
rect 1326 -9448 1432 -9437
<< via2 >>
rect 7024 5807 7084 5869
rect 13573 5806 13633 5868
rect 20227 5827 20287 5889
rect 28880 5660 28940 5722
rect 31126 5651 31279 5662
rect 31126 5543 31137 5651
rect 31137 5543 31269 5651
rect 31269 5543 31279 5651
rect 31126 5533 31279 5543
rect 32481 5252 32541 5314
rect 7246 4605 7308 4663
rect 7308 4605 7310 4663
rect 7246 4601 7310 4605
rect 13795 4604 13857 4662
rect 13857 4604 13859 4662
rect 20449 4625 20511 4683
rect 20511 4625 20513 4683
rect 20449 4621 20513 4625
rect 13795 4600 13859 4604
rect -780 4389 -664 4445
rect 33090 4624 33228 4636
rect 33090 4566 33103 4624
rect 33103 4566 33215 4624
rect 33215 4566 33228 4624
rect 33090 4554 33228 4566
rect 29102 4458 29164 4516
rect 29164 4458 29166 4516
rect 29102 4454 29166 4458
rect 360 3907 420 3969
rect 582 2705 644 2763
rect 644 2705 646 2763
rect 582 2701 646 2705
rect 352 1322 412 1384
rect 574 120 636 178
rect 636 120 638 178
rect 574 116 638 120
rect -773 -5474 -670 -5466
rect -773 -5537 -760 -5474
rect -760 -5537 -679 -5474
rect -679 -5537 -670 -5474
rect -773 -5545 -670 -5537
rect 333 -1956 393 -1894
rect 555 -3158 617 -3100
rect 617 -3158 619 -3100
rect 555 -3162 619 -3158
rect 349 -4716 409 -4654
rect 571 -5918 633 -5860
rect 633 -5918 635 -5860
rect 571 -5922 635 -5918
rect 32703 4050 32765 4108
rect 32765 4050 32767 4108
rect 32703 4046 32767 4050
rect 12370 3904 12523 3915
rect 9888 3850 10041 3861
rect 5821 3816 5974 3827
rect 3339 3762 3492 3773
rect 3339 3654 3350 3762
rect 3350 3654 3482 3762
rect 3482 3654 3492 3762
rect 5821 3708 5832 3816
rect 5832 3708 5964 3816
rect 5964 3708 5974 3816
rect 6968 3816 7121 3827
rect 5821 3698 5974 3708
rect 3339 3644 3492 3654
rect 6968 3708 6979 3816
rect 6979 3708 7111 3816
rect 7111 3708 7121 3816
rect 9888 3742 9899 3850
rect 9899 3742 10031 3850
rect 10031 3742 10041 3850
rect 12370 3796 12381 3904
rect 12381 3796 12513 3904
rect 12513 3796 12523 3904
rect 13517 3904 13670 3915
rect 12370 3786 12523 3796
rect 9888 3732 10041 3742
rect 13517 3796 13528 3904
rect 13528 3796 13660 3904
rect 13660 3796 13670 3904
rect 25649 3904 25802 3915
rect 19024 3836 19177 3847
rect 13517 3786 13670 3796
rect 16542 3782 16695 3793
rect 6968 3698 7121 3708
rect 3620 2723 3749 2734
rect 3620 2591 3630 2723
rect 3630 2591 3738 2723
rect 3738 2591 3749 2723
rect 3620 2581 3749 2591
rect 3353 2112 3506 2123
rect 3353 2004 3364 2112
rect 3364 2004 3496 2112
rect 3496 2004 3506 2112
rect 3353 1994 3506 2004
rect 3634 1073 3763 1084
rect 3634 941 3644 1073
rect 3644 941 3752 1073
rect 3752 941 3763 1073
rect 3634 931 3763 941
rect 2386 636 2501 645
rect 2386 557 2396 636
rect 2396 557 2489 636
rect 2489 557 2501 636
rect 2386 548 2501 557
rect 3348 508 3501 519
rect 3348 400 3359 508
rect 3359 400 3491 508
rect 3491 400 3501 508
rect 3348 390 3501 400
rect 8058 2908 8203 2983
rect 10169 2811 10298 2822
rect 10169 2679 10179 2811
rect 10179 2679 10287 2811
rect 10287 2679 10298 2811
rect 10169 2669 10298 2679
rect 5168 2416 5321 2426
rect 5168 2308 5178 2416
rect 5178 2308 5310 2416
rect 5310 2308 5321 2416
rect 5168 2297 5321 2308
rect 6310 2414 6463 2424
rect 6310 2306 6320 2414
rect 6320 2306 6452 2414
rect 6452 2306 6463 2414
rect 6310 2295 6463 2306
rect 9902 2200 10055 2211
rect 9902 2092 9913 2200
rect 9913 2092 10045 2200
rect 10045 2092 10055 2200
rect 9902 2082 10055 2092
rect 5166 1769 5319 1780
rect 5166 1661 5177 1769
rect 5177 1661 5309 1769
rect 5309 1661 5319 1769
rect 5166 1651 5319 1661
rect 7064 1769 7217 1780
rect 7064 1661 7075 1769
rect 7075 1661 7207 1769
rect 7207 1661 7217 1769
rect 7064 1651 7217 1661
rect 10183 1161 10312 1172
rect 10183 1029 10193 1161
rect 10193 1029 10301 1161
rect 10301 1029 10312 1161
rect 10183 1019 10312 1029
rect 5807 799 5885 809
rect 5807 733 5822 799
rect 5822 733 5885 799
rect 5807 723 5885 733
rect 3629 -531 3758 -520
rect 3629 -663 3639 -531
rect 3639 -663 3747 -531
rect 3747 -663 3758 -531
rect 3629 -673 3758 -663
rect 5112 -627 5265 -617
rect 5112 -735 5122 -627
rect 5122 -735 5254 -627
rect 5254 -735 5265 -627
rect 5112 -746 5265 -735
rect 7010 -627 7163 -617
rect 7010 -735 7020 -627
rect 7020 -735 7152 -627
rect 7152 -735 7163 -627
rect 7010 -746 7163 -735
rect 8935 724 9050 733
rect 8935 645 8945 724
rect 8945 645 9038 724
rect 9038 645 9050 724
rect 8935 636 9050 645
rect 9897 596 10050 607
rect 9897 488 9908 596
rect 9908 488 10040 596
rect 10040 488 10050 596
rect 9897 478 10050 488
rect 16542 3674 16553 3782
rect 16553 3674 16685 3782
rect 16685 3674 16695 3782
rect 19024 3728 19035 3836
rect 19035 3728 19167 3836
rect 19167 3728 19177 3836
rect 20171 3836 20324 3847
rect 19024 3718 19177 3728
rect 16542 3664 16695 3674
rect 20171 3728 20182 3836
rect 20182 3728 20314 3836
rect 20314 3728 20324 3836
rect 20171 3718 20324 3728
rect 23167 3850 23320 3861
rect 23167 3742 23178 3850
rect 23178 3742 23310 3850
rect 23310 3742 23320 3850
rect 25649 3796 25660 3904
rect 25660 3796 25792 3904
rect 25792 3796 25802 3904
rect 26796 3904 26949 3915
rect 25649 3786 25802 3796
rect 23167 3732 23320 3742
rect 26796 3796 26807 3904
rect 26807 3796 26939 3904
rect 26939 3796 26949 3904
rect 26796 3786 26949 3796
rect 16823 2743 16952 2754
rect 16823 2611 16833 2743
rect 16833 2611 16941 2743
rect 16941 2611 16952 2743
rect 16823 2601 16952 2611
rect 11717 2504 11870 2514
rect 11717 2396 11727 2504
rect 11727 2396 11859 2504
rect 11859 2396 11870 2504
rect 11717 2385 11870 2396
rect 12859 2502 13012 2512
rect 12859 2394 12869 2502
rect 12869 2394 13001 2502
rect 13001 2394 13012 2502
rect 12859 2383 13012 2394
rect 16556 2132 16709 2143
rect 16556 2024 16567 2132
rect 16567 2024 16699 2132
rect 16699 2024 16709 2132
rect 11715 1857 11868 1868
rect 11715 1749 11726 1857
rect 11726 1749 11858 1857
rect 11858 1749 11868 1857
rect 11715 1739 11868 1749
rect 13613 1857 13766 1868
rect 13613 1749 13624 1857
rect 13624 1749 13756 1857
rect 13756 1749 13766 1857
rect 13613 1739 13766 1749
rect 12356 887 12434 897
rect 12356 821 12371 887
rect 12371 821 12434 887
rect 12356 811 12434 821
rect 16556 2014 16709 2024
rect 16837 1093 16966 1104
rect 16837 961 16847 1093
rect 16847 961 16955 1093
rect 16955 961 16966 1093
rect 16837 951 16966 961
rect 15589 656 15704 665
rect 15589 577 15599 656
rect 15599 577 15692 656
rect 15692 577 15704 656
rect 15589 568 15704 577
rect 10178 -443 10307 -432
rect 10178 -575 10188 -443
rect 10188 -575 10296 -443
rect 10296 -575 10307 -443
rect 10178 -585 10307 -575
rect 11661 -539 11814 -529
rect 11661 -647 11671 -539
rect 11671 -647 11803 -539
rect 11803 -647 11814 -539
rect 11661 -658 11814 -647
rect 13559 -539 13712 -529
rect 13559 -647 13569 -539
rect 13569 -647 13701 -539
rect 13701 -647 13712 -539
rect 13559 -658 13712 -647
rect 16551 528 16704 539
rect 16551 420 16562 528
rect 16562 420 16694 528
rect 16694 420 16704 528
rect 16551 410 16704 420
rect 21192 2929 21289 3003
rect 23448 2811 23577 2822
rect 23448 2679 23458 2811
rect 23458 2679 23566 2811
rect 23566 2679 23577 2811
rect 23448 2669 23577 2679
rect 18371 2436 18524 2446
rect 18371 2328 18381 2436
rect 18381 2328 18513 2436
rect 18513 2328 18524 2436
rect 18371 2317 18524 2328
rect 19513 2434 19666 2444
rect 19513 2326 19523 2434
rect 19523 2326 19655 2434
rect 19655 2326 19666 2434
rect 19513 2315 19666 2326
rect 23181 2200 23334 2211
rect 23181 2092 23192 2200
rect 23192 2092 23324 2200
rect 23324 2092 23334 2200
rect 23181 2082 23334 2092
rect 18369 1789 18522 1800
rect 18369 1681 18380 1789
rect 18380 1681 18512 1789
rect 18512 1681 18522 1789
rect 18369 1671 18522 1681
rect 20267 1789 20420 1800
rect 20267 1681 20278 1789
rect 20278 1681 20410 1789
rect 20410 1681 20420 1789
rect 20267 1671 20420 1681
rect 23462 1161 23591 1172
rect 23462 1029 23472 1161
rect 23472 1029 23580 1161
rect 23580 1029 23591 1161
rect 23462 1019 23591 1029
rect 19010 819 19088 829
rect 19010 753 19025 819
rect 19025 753 19088 819
rect 19010 743 19088 753
rect 21745 218 21841 318
rect 16832 -511 16961 -500
rect 16832 -643 16842 -511
rect 16842 -643 16950 -511
rect 16950 -643 16961 -511
rect 16832 -653 16961 -643
rect 18315 -607 18468 -597
rect 18315 -715 18325 -607
rect 18325 -715 18457 -607
rect 18457 -715 18468 -607
rect 18315 -726 18468 -715
rect 20213 -607 20366 -597
rect 20213 -715 20223 -607
rect 20223 -715 20355 -607
rect 20355 -715 20366 -607
rect 20213 -726 20366 -715
rect 21265 -994 21407 -986
rect 21265 -1108 21276 -994
rect 21276 -1108 21399 -994
rect 21399 -1108 21407 -994
rect 21265 -1120 21407 -1108
rect 22214 724 22329 733
rect 22214 645 22224 724
rect 22224 645 22317 724
rect 22317 645 22329 724
rect 22214 636 22329 645
rect 23176 596 23329 607
rect 23176 488 23187 596
rect 23187 488 23319 596
rect 23319 488 23329 596
rect 23176 478 23329 488
rect 24996 2504 25149 2514
rect 24996 2396 25006 2504
rect 25006 2396 25138 2504
rect 25138 2396 25149 2504
rect 24996 2385 25149 2396
rect 26138 2502 26291 2512
rect 26138 2394 26148 2502
rect 26148 2394 26280 2502
rect 26280 2394 26291 2502
rect 26138 2383 26291 2394
rect 31048 3316 31259 3332
rect 31048 3193 31067 3316
rect 31067 3193 31241 3316
rect 31241 3193 31259 3316
rect 31048 3175 31259 3193
rect 28875 3089 28935 3151
rect 29097 1887 29159 1945
rect 29159 1887 29161 1945
rect 29097 1883 29161 1887
rect 24994 1857 25147 1868
rect 24994 1749 25005 1857
rect 25005 1749 25137 1857
rect 25137 1749 25147 1857
rect 24994 1739 25147 1749
rect 26892 1857 27045 1868
rect 26892 1749 26903 1857
rect 26903 1749 27035 1857
rect 27035 1749 27045 1857
rect 26892 1739 27045 1749
rect 31128 1560 31281 1571
rect 31128 1452 31139 1560
rect 31139 1452 31271 1560
rect 31271 1452 31281 1560
rect 31128 1442 31281 1452
rect 32483 1161 32543 1223
rect 25635 887 25713 897
rect 25635 821 25650 887
rect 25650 821 25713 887
rect 25635 811 25713 821
rect 28875 56 28935 118
rect 32705 -41 32767 17
rect 32767 -41 32769 17
rect 32705 -45 32769 -41
rect 23457 -443 23586 -432
rect 23457 -575 23467 -443
rect 23467 -575 23575 -443
rect 23575 -575 23586 -443
rect 23457 -585 23586 -575
rect 24940 -539 25093 -529
rect 24940 -647 24950 -539
rect 24950 -647 25082 -539
rect 25082 -647 25093 -539
rect 24940 -658 25093 -647
rect 26838 -539 26991 -529
rect 26838 -647 26848 -539
rect 26848 -647 26980 -539
rect 26980 -647 26991 -539
rect 26838 -658 26991 -647
rect 22374 -994 22516 -986
rect 22374 -1108 22385 -994
rect 22385 -1108 22508 -994
rect 22508 -1108 22516 -994
rect 22374 -1120 22516 -1108
rect 5813 -1964 5966 -1953
rect 3331 -2018 3484 -2007
rect 3331 -2126 3342 -2018
rect 3342 -2126 3474 -2018
rect 3474 -2126 3484 -2018
rect 5813 -2072 5824 -1964
rect 5824 -2072 5956 -1964
rect 5956 -2072 5966 -1964
rect 6960 -1964 7113 -1953
rect 5813 -2082 5966 -2072
rect 3331 -2136 3484 -2126
rect 6960 -2072 6971 -1964
rect 6971 -2072 7103 -1964
rect 7103 -2072 7113 -1964
rect 12364 -1966 12517 -1955
rect 6960 -2082 7113 -2072
rect 9882 -2020 10035 -2009
rect 3612 -3057 3741 -3046
rect 3612 -3189 3622 -3057
rect 3622 -3189 3730 -3057
rect 3730 -3189 3741 -3057
rect 3612 -3199 3741 -3189
rect 3345 -3668 3498 -3657
rect 3345 -3776 3356 -3668
rect 3356 -3776 3488 -3668
rect 3488 -3776 3498 -3668
rect 3345 -3786 3498 -3776
rect 1998 -4887 2232 -4750
rect 3626 -4707 3755 -4696
rect 3626 -4839 3636 -4707
rect 3636 -4839 3744 -4707
rect 3744 -4839 3755 -4707
rect 3626 -4849 3755 -4839
rect 2378 -5144 2493 -5135
rect 2378 -5223 2388 -5144
rect 2388 -5223 2481 -5144
rect 2481 -5223 2493 -5144
rect 2378 -5232 2493 -5223
rect 3340 -5272 3493 -5261
rect 3340 -5380 3351 -5272
rect 3351 -5380 3483 -5272
rect 3483 -5380 3493 -5272
rect 3340 -5390 3493 -5380
rect 9882 -2128 9893 -2020
rect 9893 -2128 10025 -2020
rect 10025 -2128 10035 -2020
rect 12364 -2074 12375 -1966
rect 12375 -2074 12507 -1966
rect 12507 -2074 12517 -1966
rect 13511 -1966 13664 -1955
rect 12364 -2084 12517 -2074
rect 9882 -2138 10035 -2128
rect 13511 -2074 13522 -1966
rect 13522 -2074 13654 -1966
rect 13654 -2074 13664 -1966
rect 13511 -2084 13664 -2074
rect 10163 -3059 10292 -3048
rect 10163 -3191 10173 -3059
rect 10173 -3191 10281 -3059
rect 10281 -3191 10292 -3059
rect 10163 -3201 10292 -3191
rect 5160 -3364 5313 -3354
rect 5160 -3472 5170 -3364
rect 5170 -3472 5302 -3364
rect 5302 -3472 5313 -3364
rect 5160 -3483 5313 -3472
rect 6302 -3366 6455 -3356
rect 6302 -3474 6312 -3366
rect 6312 -3474 6444 -3366
rect 6444 -3474 6455 -3366
rect 6302 -3485 6455 -3474
rect 9896 -3670 10049 -3659
rect 9896 -3778 9907 -3670
rect 9907 -3778 10039 -3670
rect 10039 -3778 10049 -3670
rect 9896 -3788 10049 -3778
rect 5158 -4011 5311 -4000
rect 5158 -4119 5169 -4011
rect 5169 -4119 5301 -4011
rect 5301 -4119 5311 -4011
rect 5158 -4129 5311 -4119
rect 7056 -4011 7209 -4000
rect 7056 -4119 7067 -4011
rect 7067 -4119 7199 -4011
rect 7199 -4119 7209 -4011
rect 7056 -4129 7209 -4119
rect 8633 -4893 8856 -4757
rect 10177 -4709 10306 -4698
rect 10177 -4841 10187 -4709
rect 10187 -4841 10295 -4709
rect 10295 -4841 10306 -4709
rect 10177 -4851 10306 -4841
rect 5799 -4981 5877 -4971
rect 5799 -5047 5814 -4981
rect 5814 -5047 5877 -4981
rect 5799 -5057 5877 -5047
rect 8929 -5146 9044 -5137
rect 8929 -5225 8939 -5146
rect 8939 -5225 9032 -5146
rect 9032 -5225 9044 -5146
rect 8929 -5234 9044 -5225
rect 3621 -6311 3750 -6300
rect 3621 -6443 3631 -6311
rect 3631 -6443 3739 -6311
rect 3739 -6443 3750 -6311
rect 3621 -6453 3750 -6443
rect 5104 -6407 5257 -6397
rect 5104 -6515 5114 -6407
rect 5114 -6515 5246 -6407
rect 5246 -6515 5257 -6407
rect 5104 -6526 5257 -6515
rect 7002 -6407 7155 -6397
rect 7002 -6515 7012 -6407
rect 7012 -6515 7144 -6407
rect 7144 -6515 7155 -6407
rect 7002 -6526 7155 -6515
rect 9891 -5274 10044 -5263
rect 9891 -5382 9902 -5274
rect 9902 -5382 10034 -5274
rect 10034 -5382 10044 -5274
rect 9891 -5392 10044 -5382
rect 19019 -1965 19172 -1954
rect 16537 -2019 16690 -2008
rect 16537 -2127 16548 -2019
rect 16548 -2127 16680 -2019
rect 16680 -2127 16690 -2019
rect 19019 -2073 19030 -1965
rect 19030 -2073 19162 -1965
rect 19162 -2073 19172 -1965
rect 20166 -1965 20319 -1954
rect 19019 -2083 19172 -2073
rect 16537 -2137 16690 -2127
rect 20166 -2073 20177 -1965
rect 20177 -2073 20309 -1965
rect 20309 -2073 20319 -1965
rect 25641 -1964 25794 -1953
rect 20166 -2083 20319 -2073
rect 23159 -2018 23312 -2007
rect 16818 -3058 16947 -3047
rect 16818 -3190 16828 -3058
rect 16828 -3190 16936 -3058
rect 16936 -3190 16947 -3058
rect 16818 -3200 16947 -3190
rect 11711 -3366 11864 -3356
rect 11711 -3474 11721 -3366
rect 11721 -3474 11853 -3366
rect 11853 -3474 11864 -3366
rect 11711 -3485 11864 -3474
rect 12853 -3368 13006 -3358
rect 12853 -3476 12863 -3368
rect 12863 -3476 12995 -3368
rect 12995 -3476 13006 -3368
rect 12853 -3487 13006 -3476
rect 16551 -3669 16704 -3658
rect 16551 -3777 16562 -3669
rect 16562 -3777 16694 -3669
rect 16694 -3777 16704 -3669
rect 16551 -3787 16704 -3777
rect 11709 -4013 11862 -4002
rect 11709 -4121 11720 -4013
rect 11720 -4121 11852 -4013
rect 11852 -4121 11862 -4013
rect 11709 -4131 11862 -4121
rect 13607 -4013 13760 -4002
rect 13607 -4121 13618 -4013
rect 13618 -4121 13750 -4013
rect 13750 -4121 13760 -4013
rect 13607 -4131 13760 -4121
rect 15314 -4884 15458 -4772
rect 16832 -4708 16961 -4697
rect 16832 -4840 16842 -4708
rect 16842 -4840 16950 -4708
rect 16950 -4840 16961 -4708
rect 16832 -4850 16961 -4840
rect 12350 -4983 12428 -4973
rect 12350 -5049 12365 -4983
rect 12365 -5049 12428 -4983
rect 12350 -5059 12428 -5049
rect 15584 -5145 15699 -5136
rect 15584 -5224 15594 -5145
rect 15594 -5224 15687 -5145
rect 15687 -5224 15699 -5145
rect 15584 -5233 15699 -5224
rect 10172 -6313 10301 -6302
rect 10172 -6445 10182 -6313
rect 10182 -6445 10290 -6313
rect 10290 -6445 10301 -6313
rect 10172 -6455 10301 -6445
rect 11655 -6409 11808 -6399
rect 11655 -6517 11665 -6409
rect 11665 -6517 11797 -6409
rect 11797 -6517 11808 -6409
rect 11655 -6528 11808 -6517
rect 13553 -6409 13706 -6399
rect 13553 -6517 13563 -6409
rect 13563 -6517 13695 -6409
rect 13695 -6517 13706 -6409
rect 13553 -6528 13706 -6517
rect 16546 -5273 16699 -5262
rect 16546 -5381 16557 -5273
rect 16557 -5381 16689 -5273
rect 16689 -5381 16699 -5273
rect 16546 -5391 16699 -5381
rect 23159 -2126 23170 -2018
rect 23170 -2126 23302 -2018
rect 23302 -2126 23312 -2018
rect 25641 -2072 25652 -1964
rect 25652 -2072 25784 -1964
rect 25784 -2072 25794 -1964
rect 26788 -1964 26941 -1953
rect 25641 -2082 25794 -2072
rect 23159 -2136 23312 -2126
rect 26788 -2072 26799 -1964
rect 26799 -2072 26931 -1964
rect 26931 -2072 26941 -1964
rect 26788 -2082 26941 -2072
rect 23440 -3057 23569 -3046
rect 23440 -3189 23450 -3057
rect 23450 -3189 23558 -3057
rect 23558 -3189 23569 -3057
rect 23440 -3199 23569 -3189
rect 18366 -3365 18519 -3355
rect 18366 -3473 18376 -3365
rect 18376 -3473 18508 -3365
rect 18508 -3473 18519 -3365
rect 18366 -3484 18519 -3473
rect 19508 -3367 19661 -3357
rect 19508 -3475 19518 -3367
rect 19518 -3475 19650 -3367
rect 19650 -3475 19661 -3367
rect 19508 -3486 19661 -3475
rect 23173 -3668 23326 -3657
rect 23173 -3776 23184 -3668
rect 23184 -3776 23316 -3668
rect 23316 -3776 23326 -3668
rect 23173 -3786 23326 -3776
rect 18364 -4012 18517 -4001
rect 18364 -4120 18375 -4012
rect 18375 -4120 18507 -4012
rect 18507 -4120 18517 -4012
rect 18364 -4130 18517 -4120
rect 20262 -4012 20415 -4001
rect 20262 -4120 20273 -4012
rect 20273 -4120 20405 -4012
rect 20405 -4120 20415 -4012
rect 20262 -4130 20415 -4120
rect 23454 -4707 23583 -4696
rect 23454 -4839 23464 -4707
rect 23464 -4839 23572 -4707
rect 23572 -4839 23583 -4707
rect 23454 -4849 23583 -4839
rect 19005 -4982 19083 -4972
rect 19005 -5048 19020 -4982
rect 19020 -5048 19083 -4982
rect 19005 -5058 19083 -5048
rect 22206 -5144 22321 -5135
rect 22206 -5223 22216 -5144
rect 22216 -5223 22309 -5144
rect 22309 -5223 22321 -5144
rect 22206 -5232 22321 -5223
rect 16827 -6312 16956 -6301
rect 16827 -6444 16837 -6312
rect 16837 -6444 16945 -6312
rect 16945 -6444 16956 -6312
rect 16827 -6454 16956 -6444
rect 18310 -6408 18463 -6398
rect 18310 -6516 18320 -6408
rect 18320 -6516 18452 -6408
rect 18452 -6516 18463 -6408
rect 18310 -6527 18463 -6516
rect 20208 -6408 20361 -6398
rect 20208 -6516 20218 -6408
rect 20218 -6516 20350 -6408
rect 20350 -6516 20361 -6408
rect 20208 -6527 20361 -6516
rect 23168 -5272 23321 -5261
rect 23168 -5380 23179 -5272
rect 23179 -5380 23311 -5272
rect 23311 -5380 23321 -5272
rect 23168 -5390 23321 -5380
rect 24988 -3364 25141 -3354
rect 24988 -3472 24998 -3364
rect 24998 -3472 25130 -3364
rect 25130 -3472 25141 -3364
rect 24988 -3483 25141 -3472
rect 26130 -3366 26283 -3356
rect 26130 -3474 26140 -3366
rect 26140 -3474 26272 -3366
rect 26272 -3474 26283 -3366
rect 26130 -3485 26283 -3474
rect 24986 -4011 25139 -4000
rect 24986 -4119 24997 -4011
rect 24997 -4119 25129 -4011
rect 25129 -4119 25139 -4011
rect 24986 -4129 25139 -4119
rect 26884 -4011 27037 -4000
rect 26884 -4119 26895 -4011
rect 26895 -4119 27027 -4011
rect 27027 -4119 27037 -4011
rect 26884 -4129 27037 -4119
rect 25627 -4981 25705 -4971
rect 25627 -5047 25642 -4981
rect 25642 -5047 25705 -4981
rect 25627 -5057 25705 -5047
rect 27900 -5489 28032 -5483
rect 27900 -5570 27908 -5489
rect 27908 -5570 28025 -5489
rect 28025 -5570 28032 -5489
rect 27900 -5579 28032 -5570
rect 31050 -775 31261 -759
rect 31050 -898 31069 -775
rect 31069 -898 31243 -775
rect 31243 -898 31261 -775
rect 31050 -916 31261 -898
rect 29097 -1146 29159 -1088
rect 29159 -1146 29161 -1088
rect 29097 -1150 29161 -1146
rect 28946 -1864 29006 -1802
rect 31128 -1935 31281 -1924
rect 31128 -2043 31139 -1935
rect 31139 -2043 31271 -1935
rect 31271 -2043 31281 -1935
rect 31128 -2053 31281 -2043
rect 32483 -2334 32543 -2272
rect 28681 -2915 28767 -2814
rect 30329 -2920 30422 -2843
rect 28453 -3048 28538 -2988
rect 29168 -3066 29230 -3008
rect 29230 -3066 29232 -3008
rect 29168 -3070 29232 -3066
rect 32705 -3536 32767 -3478
rect 32767 -3536 32769 -3478
rect 32705 -3540 32769 -3536
rect 31050 -4270 31261 -4254
rect 31050 -4393 31069 -4270
rect 31069 -4393 31243 -4270
rect 31243 -4393 31261 -4270
rect 31050 -4411 31261 -4393
rect 28943 -4934 29003 -4872
rect 28283 -5898 28367 -5808
rect 28717 -6019 28783 -5955
rect 29165 -6136 29227 -6078
rect 29227 -6136 29229 -6078
rect 29165 -6140 29229 -6136
rect 23449 -6311 23578 -6300
rect 23449 -6443 23459 -6311
rect 23459 -6443 23567 -6311
rect 23567 -6443 23578 -6311
rect 23449 -6453 23578 -6443
rect 24932 -6407 25085 -6397
rect 24932 -6515 24942 -6407
rect 24942 -6515 25074 -6407
rect 25074 -6515 25085 -6407
rect 24932 -6526 25085 -6515
rect 26830 -6407 26983 -6397
rect 26830 -6515 26840 -6407
rect 26840 -6515 26972 -6407
rect 26972 -6515 26983 -6407
rect 26830 -6526 26983 -6515
rect 31128 -6283 31281 -6272
rect 31128 -6391 31139 -6283
rect 31139 -6391 31271 -6283
rect 31271 -6391 31281 -6283
rect 31128 -6401 31281 -6391
rect 32483 -6682 32543 -6620
rect 7281 -7223 7345 -7219
rect 7281 -7281 7343 -7223
rect 7343 -7281 7345 -7223
rect 13835 -7218 13899 -7214
rect 13835 -7276 13897 -7218
rect 13897 -7276 13899 -7218
rect 20484 -7230 20548 -7226
rect 20484 -7288 20546 -7230
rect 20546 -7288 20548 -7230
rect 28697 -7558 28781 -7468
rect 7059 -8487 7119 -8425
rect 13613 -8482 13673 -8420
rect 28950 -7779 29010 -7717
rect 32705 -7884 32767 -7826
rect 32767 -7884 32769 -7826
rect 32705 -7888 32769 -7884
rect 28114 -8301 28196 -8211
rect 20262 -8494 20322 -8432
rect 28281 -8617 28365 -8527
rect 31050 -8618 31261 -8602
rect 31050 -8741 31069 -8618
rect 31069 -8741 31243 -8618
rect 31243 -8741 31261 -8618
rect 31050 -8759 31261 -8741
rect 28594 -8951 28655 -8876
rect 29172 -8981 29234 -8923
rect 29234 -8981 29236 -8923
rect 29172 -8985 29236 -8981
rect 27900 -9274 28032 -9268
rect 27900 -9355 27908 -9274
rect 27908 -9355 28025 -9274
rect 28025 -9355 28032 -9274
rect 27900 -9364 28032 -9355
<< metal3 >>
rect 20211 5893 20309 5911
rect 7008 5873 7106 5891
rect 7008 5801 7018 5873
rect 7088 5801 7106 5873
rect 7008 5793 7106 5801
rect 13557 5872 13655 5890
rect 13557 5800 13567 5872
rect 13637 5800 13655 5872
rect 20211 5821 20221 5893
rect 20291 5821 20309 5893
rect 20211 5813 20309 5821
rect 13557 5792 13655 5800
rect 28864 5726 28962 5744
rect 28864 5654 28874 5726
rect 28944 5654 28962 5726
rect 28864 5646 28962 5654
rect 31094 5514 31104 5693
rect 31303 5514 31313 5693
rect 32465 5318 32563 5336
rect 32465 5246 32475 5318
rect 32545 5246 32563 5318
rect 32465 5238 32563 5246
rect 20429 4689 20531 4705
rect 7226 4669 7328 4685
rect 7226 4601 7240 4669
rect 7314 4601 7328 4669
rect 7226 4587 7328 4601
rect 13775 4668 13877 4684
rect 13775 4600 13789 4668
rect 13863 4600 13877 4668
rect 20429 4621 20443 4689
rect 20517 4621 20531 4689
rect 20429 4607 20531 4621
rect 33080 4644 33439 4645
rect 33080 4636 33535 4644
rect 13775 4586 13877 4600
rect 33080 4554 33090 4636
rect 33228 4554 33535 4636
rect 33080 4545 33535 4554
rect 29082 4522 29184 4538
rect 29082 4454 29096 4522
rect 29170 4454 29184 4522
rect -790 4445 -654 4450
rect -790 4389 -780 4445
rect -664 4389 -654 4445
rect 29082 4440 29184 4454
rect -790 4384 -654 4389
rect -783 -5466 -660 4384
rect 33361 4215 33535 4545
rect 32560 4024 32570 4140
rect 32908 4024 32918 4140
rect 344 3973 442 3991
rect 344 3901 354 3973
rect 424 3901 442 3973
rect 344 3893 442 3901
rect 3307 3625 3317 3804
rect 3516 3625 3526 3804
rect 5789 3679 5799 3858
rect 5998 3679 6008 3858
rect 6936 3679 6946 3858
rect 7145 3679 7155 3858
rect 9856 3713 9866 3892
rect 10065 3713 10075 3892
rect 12338 3767 12348 3946
rect 12547 3767 12557 3946
rect 13485 3767 13495 3946
rect 13694 3767 13704 3946
rect 16510 3645 16520 3824
rect 16719 3645 16729 3824
rect 18992 3699 19002 3878
rect 19201 3699 19211 3878
rect 20139 3699 20149 3878
rect 20348 3699 20358 3878
rect 23135 3713 23145 3892
rect 23344 3713 23354 3892
rect 25617 3767 25627 3946
rect 25826 3767 25836 3946
rect 26764 3767 26774 3946
rect 26973 3767 26983 3946
rect 28859 3155 28957 3173
rect 28859 3083 28869 3155
rect 28939 3083 28957 3155
rect 31015 3153 31025 3348
rect 31291 3153 31301 3348
rect 28859 3075 28957 3083
rect 21390 3008 21647 3009
rect 21182 3003 21647 3008
rect 8048 2985 8213 2988
rect 8048 2983 8412 2985
rect 8048 2908 8058 2983
rect 8203 2908 8412 2983
rect 21182 2929 21192 3003
rect 21289 2929 21647 3003
rect 21182 2924 21647 2929
rect 8048 2903 8412 2908
rect 562 2769 664 2785
rect 562 2701 576 2769
rect 650 2701 664 2769
rect 562 2687 664 2701
rect 3601 2756 3780 2766
rect 3601 2548 3780 2557
rect 5135 2266 5144 2445
rect 5343 2266 5353 2445
rect 6277 2264 6286 2443
rect 6485 2264 6495 2443
rect 3321 1975 3331 2154
rect 3530 1975 3540 2154
rect 5134 1632 5144 1811
rect 5343 1632 5353 1811
rect 7032 1632 7042 1811
rect 7241 1632 7251 1811
rect 336 1388 434 1406
rect 336 1316 346 1388
rect 416 1316 434 1388
rect 336 1308 434 1316
rect 3615 1106 3794 1116
rect 3615 898 3794 907
rect 2397 813 2489 814
rect 5795 813 5899 815
rect 2397 809 5899 813
rect 2397 723 5807 809
rect 5885 723 5899 809
rect 2397 710 5899 723
rect 2397 650 2489 710
rect 2376 645 2511 650
rect 2376 548 2386 645
rect 2501 548 2511 645
rect 2376 543 2511 548
rect 3316 371 3326 550
rect 3525 371 3535 550
rect 554 184 656 200
rect 554 116 568 184
rect 642 116 656 184
rect 554 102 656 116
rect 3610 -498 3789 -488
rect 3610 -706 3789 -697
rect 5078 -777 5088 -598
rect 5287 -777 5297 -598
rect 6976 -777 6986 -598
rect 7185 -777 7195 -598
rect 1634 -1500 1835 -1499
rect 8268 -1500 8412 2903
rect 10150 2844 10329 2854
rect 10150 2636 10329 2645
rect 16804 2776 16983 2786
rect 16804 2568 16983 2577
rect 11684 2354 11693 2533
rect 11892 2354 11902 2533
rect 12826 2352 12835 2531
rect 13034 2352 13044 2531
rect 18338 2286 18347 2465
rect 18546 2286 18556 2465
rect 19480 2284 19489 2463
rect 19688 2284 19698 2463
rect 9870 2063 9880 2242
rect 10079 2063 10089 2242
rect 16524 1995 16534 2174
rect 16733 1995 16743 2174
rect 11683 1720 11693 1899
rect 11892 1720 11902 1899
rect 13581 1720 13591 1899
rect 13790 1720 13800 1899
rect 18337 1652 18347 1831
rect 18546 1652 18556 1831
rect 20235 1652 20245 1831
rect 20444 1652 20454 1831
rect 10164 1194 10343 1204
rect 10164 986 10343 995
rect 16818 1126 16997 1136
rect 16818 918 16997 927
rect 8946 901 9038 902
rect 12344 901 12448 903
rect 8946 897 12448 901
rect 8946 811 12356 897
rect 12434 811 12448 897
rect 8946 798 12448 811
rect 15600 833 15692 834
rect 18998 833 19102 835
rect 15600 829 19102 833
rect 8946 738 9038 798
rect 15600 743 19010 829
rect 19088 743 19102 829
rect 8925 733 9060 738
rect 8925 636 8935 733
rect 9050 636 9060 733
rect 15600 730 19102 743
rect 15600 670 15692 730
rect 15579 665 15714 670
rect 8925 631 9060 636
rect 9865 459 9875 638
rect 10074 459 10084 638
rect 15579 568 15589 665
rect 15704 568 15714 665
rect 15579 563 15714 568
rect 16519 391 16529 570
rect 16728 391 16738 570
rect 10159 -410 10338 -400
rect 16813 -478 16992 -468
rect 10159 -618 10338 -609
rect 11627 -689 11637 -510
rect 11836 -689 11846 -510
rect 13525 -689 13535 -510
rect 13734 -689 13744 -510
rect 16813 -686 16992 -677
rect 18281 -757 18291 -578
rect 18490 -757 18500 -578
rect 20179 -757 20189 -578
rect 20388 -757 20398 -578
rect 21254 -986 21421 -976
rect 21254 -1120 21265 -986
rect 21407 -1120 21421 -986
rect 21254 -1246 21421 -1120
rect 9521 -1247 21421 -1246
rect 1634 -1672 8412 -1500
rect 8633 -1418 21421 -1247
rect 8633 -1419 20532 -1418
rect 317 -1890 415 -1872
rect 317 -1962 327 -1890
rect 397 -1962 415 -1890
rect 317 -1970 415 -1962
rect 535 -3094 637 -3078
rect 535 -3162 549 -3094
rect 623 -3162 637 -3094
rect 535 -3176 637 -3162
rect 333 -4650 431 -4632
rect 333 -4722 343 -4650
rect 413 -4722 431 -4650
rect 333 -4730 431 -4722
rect 1634 -4745 1835 -1672
rect 3299 -2155 3309 -1976
rect 3508 -2155 3518 -1976
rect 5781 -2101 5791 -1922
rect 5990 -2101 6000 -1922
rect 6928 -2101 6938 -1922
rect 7137 -2101 7147 -1922
rect 3593 -3024 3772 -3014
rect 3593 -3232 3772 -3223
rect 5127 -3514 5136 -3335
rect 5335 -3514 5345 -3335
rect 6269 -3516 6278 -3337
rect 6477 -3516 6487 -3337
rect 3313 -3805 3323 -3626
rect 3522 -3805 3532 -3626
rect 5126 -4148 5136 -3969
rect 5335 -4148 5345 -3969
rect 7024 -4148 7034 -3969
rect 7233 -4148 7243 -3969
rect 8633 -4578 8819 -1419
rect 21498 -1500 21647 2924
rect 23429 2844 23608 2854
rect 23429 2636 23608 2645
rect 24963 2354 24972 2533
rect 25171 2354 25181 2533
rect 26105 2352 26114 2531
rect 26313 2352 26323 2531
rect 23149 2063 23159 2242
rect 23358 2063 23368 2242
rect 29077 1951 29179 1967
rect 24962 1720 24972 1899
rect 25171 1720 25181 1899
rect 26860 1720 26870 1899
rect 27069 1720 27079 1899
rect 29077 1883 29091 1951
rect 29165 1883 29179 1951
rect 29077 1869 29179 1883
rect 31096 1423 31106 1602
rect 31305 1423 31315 1602
rect 32467 1227 32565 1245
rect 23443 1194 23622 1204
rect 32467 1155 32477 1227
rect 32547 1155 32565 1227
rect 32467 1147 32565 1155
rect 23443 986 23622 995
rect 22225 901 22317 902
rect 25623 901 25727 903
rect 22225 897 25727 901
rect 22225 811 25635 897
rect 25713 811 25727 897
rect 22225 798 25727 811
rect 22225 738 22317 798
rect 22204 733 22339 738
rect 22204 636 22214 733
rect 22329 636 22339 733
rect 22204 631 22339 636
rect 23144 459 23154 638
rect 23353 459 23363 638
rect 21735 318 22077 323
rect 21735 218 21745 318
rect 21841 218 22077 318
rect 21735 213 22077 218
rect 21736 210 22077 213
rect 15038 -1687 21647 -1500
rect 21927 -1496 22077 210
rect 28859 122 28957 140
rect 28859 50 28869 122
rect 28939 50 28957 122
rect 28859 42 28957 50
rect 32562 -67 32572 49
rect 32910 -67 32920 49
rect 23438 -410 23617 -400
rect 23438 -618 23617 -609
rect 24906 -689 24916 -510
rect 25115 -689 25125 -510
rect 26804 -689 26814 -510
rect 27013 -689 27023 -510
rect 31017 -938 31027 -743
rect 31293 -938 31303 -743
rect 22363 -986 22530 -976
rect 22363 -1120 22374 -986
rect 22516 -1120 22530 -986
rect 22363 -1248 22530 -1120
rect 29077 -1082 29179 -1066
rect 29077 -1150 29091 -1082
rect 29165 -1150 29179 -1082
rect 29077 -1164 29179 -1150
rect 33361 -1248 33534 4215
rect 22363 -1334 33534 -1248
rect 22364 -1418 33534 -1334
rect 33361 -1421 33534 -1418
rect 30076 -1496 30195 -1494
rect 9850 -2157 9860 -1978
rect 10059 -2157 10069 -1978
rect 12332 -2103 12342 -1924
rect 12541 -2103 12551 -1924
rect 13479 -2103 13489 -1924
rect 13688 -2103 13698 -1924
rect 10144 -3026 10323 -3016
rect 10144 -3234 10323 -3225
rect 11678 -3516 11687 -3337
rect 11886 -3516 11896 -3337
rect 12820 -3518 12829 -3339
rect 13028 -3518 13038 -3339
rect 9864 -3807 9874 -3628
rect 10073 -3807 10083 -3628
rect 11677 -4150 11687 -3971
rect 11886 -4150 11896 -3971
rect 13575 -4150 13585 -3971
rect 13784 -4150 13794 -3971
rect 3607 -4674 3786 -4664
rect 1633 -4750 2245 -4745
rect 1633 -4887 1998 -4750
rect 2232 -4887 2245 -4750
rect 8632 -4703 8820 -4578
rect 10158 -4676 10337 -4666
rect 8622 -4757 8866 -4703
rect 8622 -4798 8633 -4757
rect 3607 -4882 3786 -4873
rect 1633 -4891 2245 -4887
rect 1988 -4892 2242 -4891
rect 8623 -4893 8633 -4798
rect 8856 -4893 8866 -4757
rect 15038 -4741 15239 -1687
rect 21927 -1691 30195 -1496
rect 28930 -1798 29028 -1780
rect 28930 -1870 28940 -1798
rect 29010 -1870 29028 -1798
rect 28930 -1878 29028 -1870
rect 16505 -2156 16515 -1977
rect 16714 -2156 16724 -1977
rect 18987 -2102 18997 -1923
rect 19196 -2102 19206 -1923
rect 20134 -2102 20144 -1923
rect 20343 -2102 20353 -1923
rect 23127 -2155 23137 -1976
rect 23336 -2155 23346 -1976
rect 25609 -2101 25619 -1922
rect 25818 -2101 25828 -1922
rect 26756 -2101 26766 -1922
rect 26965 -2101 26975 -1922
rect 28109 -2811 28777 -2809
rect 28108 -2814 28777 -2811
rect 28108 -2915 28681 -2814
rect 28767 -2915 28777 -2814
rect 28108 -2920 28777 -2915
rect 30076 -2838 30195 -1691
rect 31096 -2072 31106 -1893
rect 31305 -2072 31315 -1893
rect 32467 -2268 32565 -2250
rect 32467 -2340 32477 -2268
rect 32547 -2340 32565 -2268
rect 32467 -2348 32565 -2340
rect 30076 -2843 30432 -2838
rect 30076 -2920 30329 -2843
rect 30422 -2920 30432 -2843
rect 16799 -3025 16978 -3015
rect 16799 -3233 16978 -3224
rect 23421 -3024 23600 -3014
rect 23421 -3232 23600 -3223
rect 18333 -3515 18342 -3336
rect 18541 -3515 18551 -3336
rect 19475 -3517 19484 -3338
rect 19683 -3517 19693 -3338
rect 24955 -3514 24964 -3335
rect 25163 -3514 25173 -3335
rect 26097 -3516 26106 -3337
rect 26305 -3516 26315 -3337
rect 16519 -3806 16529 -3627
rect 16728 -3806 16738 -3627
rect 23141 -3805 23151 -3626
rect 23350 -3805 23360 -3626
rect 18332 -4149 18342 -3970
rect 18541 -4149 18551 -3970
rect 20230 -4149 20240 -3970
rect 20439 -4149 20449 -3970
rect 24954 -4148 24964 -3969
rect 25163 -4148 25173 -3969
rect 26852 -4148 26862 -3969
rect 27061 -4148 27071 -3969
rect 16813 -4675 16992 -4665
rect 15038 -4772 15486 -4741
rect 15038 -4794 15314 -4772
rect 10158 -4884 10337 -4875
rect 15039 -4884 15314 -4794
rect 15458 -4884 15486 -4772
rect 16813 -4883 16992 -4874
rect 23435 -4674 23614 -4664
rect 23435 -4882 23614 -4873
rect 8623 -4898 8866 -4893
rect 15039 -4902 15486 -4884
rect 2389 -4967 2481 -4966
rect 5787 -4967 5891 -4965
rect 2389 -4971 5891 -4967
rect 2389 -5057 5799 -4971
rect 5877 -5057 5891 -4971
rect 2389 -5070 5891 -5057
rect 8940 -4969 9032 -4968
rect 12338 -4969 12442 -4967
rect 8940 -4973 12442 -4969
rect 8940 -5059 12350 -4973
rect 12428 -5059 12442 -4973
rect 2389 -5130 2481 -5070
rect 8940 -5072 12442 -5059
rect 15595 -4968 15687 -4967
rect 18993 -4968 19097 -4966
rect 15595 -4972 19097 -4968
rect 15595 -5058 19005 -4972
rect 19083 -5058 19097 -4972
rect 15595 -5071 19097 -5058
rect 22217 -4967 22309 -4966
rect 25615 -4967 25719 -4965
rect 22217 -4971 25719 -4967
rect 22217 -5057 25627 -4971
rect 25705 -5057 25719 -4971
rect 22217 -5070 25719 -5057
rect 2368 -5135 2503 -5130
rect 8940 -5132 9032 -5072
rect 15595 -5131 15687 -5071
rect 22217 -5130 22309 -5070
rect 2368 -5232 2378 -5135
rect 2493 -5232 2503 -5135
rect 8919 -5137 9054 -5132
rect 2368 -5237 2503 -5232
rect 3308 -5409 3318 -5230
rect 3517 -5409 3527 -5230
rect 8919 -5234 8929 -5137
rect 9044 -5234 9054 -5137
rect 15574 -5136 15709 -5131
rect 8919 -5239 9054 -5234
rect 9859 -5411 9869 -5232
rect 10068 -5411 10078 -5232
rect 15574 -5233 15584 -5136
rect 15699 -5233 15709 -5136
rect 22196 -5135 22331 -5130
rect 15574 -5238 15709 -5233
rect 16514 -5410 16524 -5231
rect 16723 -5410 16733 -5231
rect 22196 -5232 22206 -5135
rect 22321 -5232 22331 -5135
rect 22196 -5237 22331 -5232
rect 23136 -5409 23146 -5230
rect 23345 -5409 23355 -5230
rect -783 -5545 -773 -5466
rect -670 -5545 -660 -5466
rect -783 -5550 -660 -5545
rect 27887 -5483 28047 -5477
rect 27887 -5579 27900 -5483
rect 28032 -5579 28047 -5483
rect 551 -5854 653 -5838
rect 551 -5922 565 -5854
rect 639 -5922 653 -5854
rect 551 -5936 653 -5922
rect 3602 -6278 3781 -6268
rect 10153 -6280 10332 -6270
rect 3602 -6486 3781 -6477
rect 5070 -6557 5080 -6378
rect 5279 -6557 5289 -6378
rect 6968 -6557 6978 -6378
rect 7177 -6557 7187 -6378
rect 16808 -6279 16987 -6269
rect 10153 -6488 10332 -6479
rect 11621 -6559 11631 -6380
rect 11830 -6559 11840 -6380
rect 13519 -6559 13529 -6380
rect 13728 -6559 13738 -6380
rect 23430 -6278 23609 -6268
rect 16808 -6487 16987 -6478
rect 18276 -6558 18286 -6379
rect 18485 -6558 18495 -6379
rect 20174 -6558 20184 -6379
rect 20383 -6558 20393 -6379
rect 23430 -6486 23609 -6477
rect 24898 -6557 24908 -6378
rect 25107 -6557 25117 -6378
rect 26796 -6557 26806 -6378
rect 27005 -6557 27015 -6378
rect 7261 -7219 7363 -7205
rect 7261 -7287 7275 -7219
rect 7349 -7287 7363 -7219
rect 7261 -7303 7363 -7287
rect 13815 -7214 13917 -7200
rect 13815 -7282 13829 -7214
rect 13903 -7282 13917 -7214
rect 13815 -7298 13917 -7282
rect 20464 -7226 20566 -7212
rect 20464 -7294 20478 -7226
rect 20552 -7294 20566 -7226
rect 20464 -7310 20566 -7294
rect 7043 -8419 7141 -8411
rect 7043 -8491 7053 -8419
rect 7123 -8491 7141 -8419
rect 7043 -8509 7141 -8491
rect 13597 -8414 13695 -8406
rect 13597 -8486 13607 -8414
rect 13677 -8486 13695 -8414
rect 13597 -8504 13695 -8486
rect 20246 -8426 20344 -8418
rect 20246 -8498 20256 -8426
rect 20326 -8498 20344 -8426
rect 20246 -8516 20344 -8498
rect 27887 -9268 28047 -5579
rect 28108 -5587 28208 -2920
rect 30076 -2925 30432 -2920
rect 30076 -2927 30395 -2925
rect 28443 -2988 28548 -2983
rect 28443 -3048 28453 -2988
rect 28538 -3048 28548 -2988
rect 28443 -3085 28548 -3048
rect 29148 -3002 29250 -2986
rect 29148 -3070 29162 -3002
rect 29236 -3070 29250 -3002
rect 29148 -3084 29250 -3070
rect 28108 -8211 28209 -5587
rect 28277 -5803 28379 -5794
rect 28273 -5808 28379 -5803
rect 28273 -5898 28283 -5808
rect 28367 -5898 28379 -5808
rect 28273 -5903 28379 -5898
rect 28108 -8301 28114 -8211
rect 28196 -8301 28209 -8211
rect 28108 -8311 28209 -8301
rect 28277 -5905 28379 -5903
rect 28277 -8522 28377 -5905
rect 28271 -8527 28377 -8522
rect 28271 -8617 28281 -8527
rect 28365 -8617 28377 -8527
rect 28271 -8622 28377 -8617
rect 28277 -8624 28377 -8622
rect 28454 -8871 28531 -3085
rect 32562 -3562 32572 -3446
rect 32910 -3562 32920 -3446
rect 31017 -4433 31027 -4238
rect 31293 -4433 31303 -4238
rect 28927 -4868 29025 -4850
rect 28927 -4940 28937 -4868
rect 29007 -4940 29025 -4868
rect 28927 -4948 29025 -4940
rect 28707 -5955 28793 -5950
rect 28707 -6019 28717 -5955
rect 28783 -6019 28793 -5955
rect 28707 -7453 28793 -6019
rect 29145 -6072 29247 -6056
rect 29145 -6140 29159 -6072
rect 29233 -6140 29247 -6072
rect 29145 -6154 29247 -6140
rect 31096 -6420 31106 -6241
rect 31305 -6420 31315 -6241
rect 32467 -6616 32565 -6598
rect 32467 -6688 32477 -6616
rect 32547 -6688 32565 -6616
rect 32467 -6696 32565 -6688
rect 28692 -7468 28793 -7453
rect 28692 -7558 28697 -7468
rect 28781 -7558 28793 -7468
rect 28692 -7567 28793 -7558
rect 28934 -7713 29032 -7695
rect 28934 -7785 28944 -7713
rect 29014 -7785 29032 -7713
rect 28934 -7793 29032 -7785
rect 32562 -7910 32572 -7794
rect 32910 -7910 32920 -7794
rect 31017 -8781 31027 -8586
rect 31293 -8781 31303 -8586
rect 28454 -8876 28665 -8871
rect 28454 -8951 28594 -8876
rect 28655 -8951 28665 -8876
rect 28454 -8956 28665 -8951
rect 29152 -8917 29254 -8901
rect 29152 -8985 29166 -8917
rect 29240 -8985 29254 -8917
rect 29152 -8999 29254 -8985
rect 27887 -9364 27900 -9268
rect 28032 -9364 28047 -9268
rect 27887 -9390 28047 -9364
<< via3 >>
rect 7018 5869 7088 5873
rect 7018 5807 7024 5869
rect 7024 5807 7084 5869
rect 7084 5807 7088 5869
rect 7018 5801 7088 5807
rect 13567 5868 13637 5872
rect 13567 5806 13573 5868
rect 13573 5806 13633 5868
rect 13633 5806 13637 5868
rect 13567 5800 13637 5806
rect 20221 5889 20291 5893
rect 20221 5827 20227 5889
rect 20227 5827 20287 5889
rect 20287 5827 20291 5889
rect 20221 5821 20291 5827
rect 28874 5722 28944 5726
rect 28874 5660 28880 5722
rect 28880 5660 28940 5722
rect 28940 5660 28944 5722
rect 28874 5654 28944 5660
rect 31104 5662 31303 5693
rect 31104 5533 31126 5662
rect 31126 5533 31279 5662
rect 31279 5533 31303 5662
rect 31104 5514 31303 5533
rect 32475 5314 32545 5318
rect 32475 5252 32481 5314
rect 32481 5252 32541 5314
rect 32541 5252 32545 5314
rect 32475 5246 32545 5252
rect 7240 4663 7314 4669
rect 7240 4601 7246 4663
rect 7246 4601 7310 4663
rect 7310 4601 7314 4663
rect 13789 4662 13863 4668
rect 13789 4600 13795 4662
rect 13795 4600 13859 4662
rect 13859 4600 13863 4662
rect 20443 4683 20517 4689
rect 20443 4621 20449 4683
rect 20449 4621 20513 4683
rect 20513 4621 20517 4683
rect 29096 4516 29170 4522
rect 29096 4454 29102 4516
rect 29102 4454 29166 4516
rect 29166 4454 29170 4516
rect 32570 4108 32908 4140
rect 32570 4046 32703 4108
rect 32703 4046 32767 4108
rect 32767 4046 32908 4108
rect 32570 4024 32908 4046
rect 354 3969 424 3973
rect 354 3907 360 3969
rect 360 3907 420 3969
rect 420 3907 424 3969
rect 354 3901 424 3907
rect 3317 3773 3516 3804
rect 3317 3644 3339 3773
rect 3339 3644 3492 3773
rect 3492 3644 3516 3773
rect 3317 3625 3516 3644
rect 5799 3827 5998 3858
rect 5799 3698 5821 3827
rect 5821 3698 5974 3827
rect 5974 3698 5998 3827
rect 5799 3679 5998 3698
rect 6946 3827 7145 3858
rect 6946 3698 6968 3827
rect 6968 3698 7121 3827
rect 7121 3698 7145 3827
rect 6946 3679 7145 3698
rect 9866 3861 10065 3892
rect 9866 3732 9888 3861
rect 9888 3732 10041 3861
rect 10041 3732 10065 3861
rect 9866 3713 10065 3732
rect 12348 3915 12547 3946
rect 12348 3786 12370 3915
rect 12370 3786 12523 3915
rect 12523 3786 12547 3915
rect 12348 3767 12547 3786
rect 13495 3915 13694 3946
rect 13495 3786 13517 3915
rect 13517 3786 13670 3915
rect 13670 3786 13694 3915
rect 13495 3767 13694 3786
rect 16520 3793 16719 3824
rect 16520 3664 16542 3793
rect 16542 3664 16695 3793
rect 16695 3664 16719 3793
rect 16520 3645 16719 3664
rect 19002 3847 19201 3878
rect 19002 3718 19024 3847
rect 19024 3718 19177 3847
rect 19177 3718 19201 3847
rect 19002 3699 19201 3718
rect 20149 3847 20348 3878
rect 20149 3718 20171 3847
rect 20171 3718 20324 3847
rect 20324 3718 20348 3847
rect 20149 3699 20348 3718
rect 23145 3861 23344 3892
rect 23145 3732 23167 3861
rect 23167 3732 23320 3861
rect 23320 3732 23344 3861
rect 23145 3713 23344 3732
rect 25627 3915 25826 3946
rect 25627 3786 25649 3915
rect 25649 3786 25802 3915
rect 25802 3786 25826 3915
rect 25627 3767 25826 3786
rect 26774 3915 26973 3946
rect 26774 3786 26796 3915
rect 26796 3786 26949 3915
rect 26949 3786 26973 3915
rect 26774 3767 26973 3786
rect 28869 3151 28939 3155
rect 28869 3089 28875 3151
rect 28875 3089 28935 3151
rect 28935 3089 28939 3151
rect 28869 3083 28939 3089
rect 31025 3332 31291 3348
rect 31025 3175 31048 3332
rect 31048 3175 31259 3332
rect 31259 3175 31291 3332
rect 31025 3153 31291 3175
rect 576 2763 650 2769
rect 576 2701 582 2763
rect 582 2701 646 2763
rect 646 2701 650 2763
rect 3601 2734 3780 2756
rect 3601 2581 3620 2734
rect 3620 2581 3749 2734
rect 3749 2581 3780 2734
rect 3601 2557 3780 2581
rect 5144 2426 5343 2445
rect 5144 2297 5168 2426
rect 5168 2297 5321 2426
rect 5321 2297 5343 2426
rect 5144 2266 5343 2297
rect 6286 2424 6485 2443
rect 6286 2295 6310 2424
rect 6310 2295 6463 2424
rect 6463 2295 6485 2424
rect 6286 2264 6485 2295
rect 3331 2123 3530 2154
rect 3331 1994 3353 2123
rect 3353 1994 3506 2123
rect 3506 1994 3530 2123
rect 3331 1975 3530 1994
rect 5144 1780 5343 1811
rect 5144 1651 5166 1780
rect 5166 1651 5319 1780
rect 5319 1651 5343 1780
rect 5144 1632 5343 1651
rect 7042 1780 7241 1811
rect 7042 1651 7064 1780
rect 7064 1651 7217 1780
rect 7217 1651 7241 1780
rect 7042 1632 7241 1651
rect 346 1384 416 1388
rect 346 1322 352 1384
rect 352 1322 412 1384
rect 412 1322 416 1384
rect 346 1316 416 1322
rect 3615 1084 3794 1106
rect 3615 931 3634 1084
rect 3634 931 3763 1084
rect 3763 931 3794 1084
rect 3615 907 3794 931
rect 3326 519 3525 550
rect 3326 390 3348 519
rect 3348 390 3501 519
rect 3501 390 3525 519
rect 3326 371 3525 390
rect 568 178 642 184
rect 568 116 574 178
rect 574 116 638 178
rect 638 116 642 178
rect 3610 -520 3789 -498
rect 3610 -673 3629 -520
rect 3629 -673 3758 -520
rect 3758 -673 3789 -520
rect 3610 -697 3789 -673
rect 5088 -617 5287 -598
rect 5088 -746 5112 -617
rect 5112 -746 5265 -617
rect 5265 -746 5287 -617
rect 5088 -777 5287 -746
rect 6986 -617 7185 -598
rect 6986 -746 7010 -617
rect 7010 -746 7163 -617
rect 7163 -746 7185 -617
rect 6986 -777 7185 -746
rect 10150 2822 10329 2844
rect 10150 2669 10169 2822
rect 10169 2669 10298 2822
rect 10298 2669 10329 2822
rect 10150 2645 10329 2669
rect 16804 2754 16983 2776
rect 16804 2601 16823 2754
rect 16823 2601 16952 2754
rect 16952 2601 16983 2754
rect 16804 2577 16983 2601
rect 11693 2514 11892 2533
rect 11693 2385 11717 2514
rect 11717 2385 11870 2514
rect 11870 2385 11892 2514
rect 11693 2354 11892 2385
rect 12835 2512 13034 2531
rect 12835 2383 12859 2512
rect 12859 2383 13012 2512
rect 13012 2383 13034 2512
rect 12835 2352 13034 2383
rect 18347 2446 18546 2465
rect 18347 2317 18371 2446
rect 18371 2317 18524 2446
rect 18524 2317 18546 2446
rect 18347 2286 18546 2317
rect 19489 2444 19688 2463
rect 19489 2315 19513 2444
rect 19513 2315 19666 2444
rect 19666 2315 19688 2444
rect 19489 2284 19688 2315
rect 9880 2211 10079 2242
rect 9880 2082 9902 2211
rect 9902 2082 10055 2211
rect 10055 2082 10079 2211
rect 9880 2063 10079 2082
rect 16534 2143 16733 2174
rect 16534 2014 16556 2143
rect 16556 2014 16709 2143
rect 16709 2014 16733 2143
rect 16534 1995 16733 2014
rect 11693 1868 11892 1899
rect 11693 1739 11715 1868
rect 11715 1739 11868 1868
rect 11868 1739 11892 1868
rect 11693 1720 11892 1739
rect 13591 1868 13790 1899
rect 13591 1739 13613 1868
rect 13613 1739 13766 1868
rect 13766 1739 13790 1868
rect 13591 1720 13790 1739
rect 18347 1800 18546 1831
rect 18347 1671 18369 1800
rect 18369 1671 18522 1800
rect 18522 1671 18546 1800
rect 18347 1652 18546 1671
rect 20245 1800 20444 1831
rect 20245 1671 20267 1800
rect 20267 1671 20420 1800
rect 20420 1671 20444 1800
rect 20245 1652 20444 1671
rect 10164 1172 10343 1194
rect 10164 1019 10183 1172
rect 10183 1019 10312 1172
rect 10312 1019 10343 1172
rect 10164 995 10343 1019
rect 16818 1104 16997 1126
rect 16818 951 16837 1104
rect 16837 951 16966 1104
rect 16966 951 16997 1104
rect 16818 927 16997 951
rect 9875 607 10074 638
rect 9875 478 9897 607
rect 9897 478 10050 607
rect 10050 478 10074 607
rect 9875 459 10074 478
rect 16529 539 16728 570
rect 16529 410 16551 539
rect 16551 410 16704 539
rect 16704 410 16728 539
rect 16529 391 16728 410
rect 10159 -432 10338 -410
rect 10159 -585 10178 -432
rect 10178 -585 10307 -432
rect 10307 -585 10338 -432
rect 16813 -500 16992 -478
rect 10159 -609 10338 -585
rect 11637 -529 11836 -510
rect 11637 -658 11661 -529
rect 11661 -658 11814 -529
rect 11814 -658 11836 -529
rect 11637 -689 11836 -658
rect 13535 -529 13734 -510
rect 13535 -658 13559 -529
rect 13559 -658 13712 -529
rect 13712 -658 13734 -529
rect 13535 -689 13734 -658
rect 16813 -653 16832 -500
rect 16832 -653 16961 -500
rect 16961 -653 16992 -500
rect 16813 -677 16992 -653
rect 18291 -597 18490 -578
rect 18291 -726 18315 -597
rect 18315 -726 18468 -597
rect 18468 -726 18490 -597
rect 18291 -757 18490 -726
rect 20189 -597 20388 -578
rect 20189 -726 20213 -597
rect 20213 -726 20366 -597
rect 20366 -726 20388 -597
rect 20189 -757 20388 -726
rect 327 -1894 397 -1890
rect 327 -1956 333 -1894
rect 333 -1956 393 -1894
rect 393 -1956 397 -1894
rect 327 -1962 397 -1956
rect 549 -3100 623 -3094
rect 549 -3162 555 -3100
rect 555 -3162 619 -3100
rect 619 -3162 623 -3100
rect 343 -4654 413 -4650
rect 343 -4716 349 -4654
rect 349 -4716 409 -4654
rect 409 -4716 413 -4654
rect 343 -4722 413 -4716
rect 3309 -2007 3508 -1976
rect 3309 -2136 3331 -2007
rect 3331 -2136 3484 -2007
rect 3484 -2136 3508 -2007
rect 3309 -2155 3508 -2136
rect 5791 -1953 5990 -1922
rect 5791 -2082 5813 -1953
rect 5813 -2082 5966 -1953
rect 5966 -2082 5990 -1953
rect 5791 -2101 5990 -2082
rect 6938 -1953 7137 -1922
rect 6938 -2082 6960 -1953
rect 6960 -2082 7113 -1953
rect 7113 -2082 7137 -1953
rect 6938 -2101 7137 -2082
rect 3593 -3046 3772 -3024
rect 3593 -3199 3612 -3046
rect 3612 -3199 3741 -3046
rect 3741 -3199 3772 -3046
rect 3593 -3223 3772 -3199
rect 5136 -3354 5335 -3335
rect 5136 -3483 5160 -3354
rect 5160 -3483 5313 -3354
rect 5313 -3483 5335 -3354
rect 5136 -3514 5335 -3483
rect 6278 -3356 6477 -3337
rect 6278 -3485 6302 -3356
rect 6302 -3485 6455 -3356
rect 6455 -3485 6477 -3356
rect 6278 -3516 6477 -3485
rect 3323 -3657 3522 -3626
rect 3323 -3786 3345 -3657
rect 3345 -3786 3498 -3657
rect 3498 -3786 3522 -3657
rect 3323 -3805 3522 -3786
rect 5136 -4000 5335 -3969
rect 5136 -4129 5158 -4000
rect 5158 -4129 5311 -4000
rect 5311 -4129 5335 -4000
rect 5136 -4148 5335 -4129
rect 7034 -4000 7233 -3969
rect 7034 -4129 7056 -4000
rect 7056 -4129 7209 -4000
rect 7209 -4129 7233 -4000
rect 7034 -4148 7233 -4129
rect 23429 2822 23608 2844
rect 23429 2669 23448 2822
rect 23448 2669 23577 2822
rect 23577 2669 23608 2822
rect 23429 2645 23608 2669
rect 24972 2514 25171 2533
rect 24972 2385 24996 2514
rect 24996 2385 25149 2514
rect 25149 2385 25171 2514
rect 24972 2354 25171 2385
rect 26114 2512 26313 2531
rect 26114 2383 26138 2512
rect 26138 2383 26291 2512
rect 26291 2383 26313 2512
rect 26114 2352 26313 2383
rect 23159 2211 23358 2242
rect 23159 2082 23181 2211
rect 23181 2082 23334 2211
rect 23334 2082 23358 2211
rect 23159 2063 23358 2082
rect 24972 1868 25171 1899
rect 24972 1739 24994 1868
rect 24994 1739 25147 1868
rect 25147 1739 25171 1868
rect 24972 1720 25171 1739
rect 26870 1868 27069 1899
rect 26870 1739 26892 1868
rect 26892 1739 27045 1868
rect 27045 1739 27069 1868
rect 26870 1720 27069 1739
rect 29091 1945 29165 1951
rect 29091 1883 29097 1945
rect 29097 1883 29161 1945
rect 29161 1883 29165 1945
rect 31106 1571 31305 1602
rect 31106 1442 31128 1571
rect 31128 1442 31281 1571
rect 31281 1442 31305 1571
rect 31106 1423 31305 1442
rect 23443 1172 23622 1194
rect 23443 1019 23462 1172
rect 23462 1019 23591 1172
rect 23591 1019 23622 1172
rect 32477 1223 32547 1227
rect 32477 1161 32483 1223
rect 32483 1161 32543 1223
rect 32543 1161 32547 1223
rect 32477 1155 32547 1161
rect 23443 995 23622 1019
rect 23154 607 23353 638
rect 23154 478 23176 607
rect 23176 478 23329 607
rect 23329 478 23353 607
rect 23154 459 23353 478
rect 28869 118 28939 122
rect 28869 56 28875 118
rect 28875 56 28935 118
rect 28935 56 28939 118
rect 28869 50 28939 56
rect 32572 17 32910 49
rect 32572 -45 32705 17
rect 32705 -45 32769 17
rect 32769 -45 32910 17
rect 32572 -67 32910 -45
rect 23438 -432 23617 -410
rect 23438 -585 23457 -432
rect 23457 -585 23586 -432
rect 23586 -585 23617 -432
rect 23438 -609 23617 -585
rect 24916 -529 25115 -510
rect 24916 -658 24940 -529
rect 24940 -658 25093 -529
rect 25093 -658 25115 -529
rect 24916 -689 25115 -658
rect 26814 -529 27013 -510
rect 26814 -658 26838 -529
rect 26838 -658 26991 -529
rect 26991 -658 27013 -529
rect 26814 -689 27013 -658
rect 31027 -759 31293 -743
rect 31027 -916 31050 -759
rect 31050 -916 31261 -759
rect 31261 -916 31293 -759
rect 31027 -938 31293 -916
rect 29091 -1088 29165 -1082
rect 29091 -1150 29097 -1088
rect 29097 -1150 29161 -1088
rect 29161 -1150 29165 -1088
rect 9860 -2009 10059 -1978
rect 9860 -2138 9882 -2009
rect 9882 -2138 10035 -2009
rect 10035 -2138 10059 -2009
rect 9860 -2157 10059 -2138
rect 12342 -1955 12541 -1924
rect 12342 -2084 12364 -1955
rect 12364 -2084 12517 -1955
rect 12517 -2084 12541 -1955
rect 12342 -2103 12541 -2084
rect 13489 -1955 13688 -1924
rect 13489 -2084 13511 -1955
rect 13511 -2084 13664 -1955
rect 13664 -2084 13688 -1955
rect 13489 -2103 13688 -2084
rect 10144 -3048 10323 -3026
rect 10144 -3201 10163 -3048
rect 10163 -3201 10292 -3048
rect 10292 -3201 10323 -3048
rect 10144 -3225 10323 -3201
rect 11687 -3356 11886 -3337
rect 11687 -3485 11711 -3356
rect 11711 -3485 11864 -3356
rect 11864 -3485 11886 -3356
rect 11687 -3516 11886 -3485
rect 12829 -3358 13028 -3339
rect 12829 -3487 12853 -3358
rect 12853 -3487 13006 -3358
rect 13006 -3487 13028 -3358
rect 12829 -3518 13028 -3487
rect 9874 -3659 10073 -3628
rect 9874 -3788 9896 -3659
rect 9896 -3788 10049 -3659
rect 10049 -3788 10073 -3659
rect 9874 -3807 10073 -3788
rect 11687 -4002 11886 -3971
rect 11687 -4131 11709 -4002
rect 11709 -4131 11862 -4002
rect 11862 -4131 11886 -4002
rect 11687 -4150 11886 -4131
rect 13585 -4002 13784 -3971
rect 13585 -4131 13607 -4002
rect 13607 -4131 13760 -4002
rect 13760 -4131 13784 -4002
rect 13585 -4150 13784 -4131
rect 3607 -4696 3786 -4674
rect 3607 -4849 3626 -4696
rect 3626 -4849 3755 -4696
rect 3755 -4849 3786 -4696
rect 10158 -4698 10337 -4676
rect 3607 -4873 3786 -4849
rect 10158 -4851 10177 -4698
rect 10177 -4851 10306 -4698
rect 10306 -4851 10337 -4698
rect 28940 -1802 29010 -1798
rect 28940 -1864 28946 -1802
rect 28946 -1864 29006 -1802
rect 29006 -1864 29010 -1802
rect 28940 -1870 29010 -1864
rect 16515 -2008 16714 -1977
rect 16515 -2137 16537 -2008
rect 16537 -2137 16690 -2008
rect 16690 -2137 16714 -2008
rect 16515 -2156 16714 -2137
rect 18997 -1954 19196 -1923
rect 18997 -2083 19019 -1954
rect 19019 -2083 19172 -1954
rect 19172 -2083 19196 -1954
rect 18997 -2102 19196 -2083
rect 20144 -1954 20343 -1923
rect 20144 -2083 20166 -1954
rect 20166 -2083 20319 -1954
rect 20319 -2083 20343 -1954
rect 20144 -2102 20343 -2083
rect 23137 -2007 23336 -1976
rect 23137 -2136 23159 -2007
rect 23159 -2136 23312 -2007
rect 23312 -2136 23336 -2007
rect 23137 -2155 23336 -2136
rect 25619 -1953 25818 -1922
rect 25619 -2082 25641 -1953
rect 25641 -2082 25794 -1953
rect 25794 -2082 25818 -1953
rect 25619 -2101 25818 -2082
rect 26766 -1953 26965 -1922
rect 26766 -2082 26788 -1953
rect 26788 -2082 26941 -1953
rect 26941 -2082 26965 -1953
rect 26766 -2101 26965 -2082
rect 31106 -1924 31305 -1893
rect 31106 -2053 31128 -1924
rect 31128 -2053 31281 -1924
rect 31281 -2053 31305 -1924
rect 31106 -2072 31305 -2053
rect 32477 -2272 32547 -2268
rect 32477 -2334 32483 -2272
rect 32483 -2334 32543 -2272
rect 32543 -2334 32547 -2272
rect 32477 -2340 32547 -2334
rect 16799 -3047 16978 -3025
rect 16799 -3200 16818 -3047
rect 16818 -3200 16947 -3047
rect 16947 -3200 16978 -3047
rect 16799 -3224 16978 -3200
rect 23421 -3046 23600 -3024
rect 23421 -3199 23440 -3046
rect 23440 -3199 23569 -3046
rect 23569 -3199 23600 -3046
rect 23421 -3223 23600 -3199
rect 18342 -3355 18541 -3336
rect 18342 -3484 18366 -3355
rect 18366 -3484 18519 -3355
rect 18519 -3484 18541 -3355
rect 18342 -3515 18541 -3484
rect 19484 -3357 19683 -3338
rect 19484 -3486 19508 -3357
rect 19508 -3486 19661 -3357
rect 19661 -3486 19683 -3357
rect 19484 -3517 19683 -3486
rect 24964 -3354 25163 -3335
rect 24964 -3483 24988 -3354
rect 24988 -3483 25141 -3354
rect 25141 -3483 25163 -3354
rect 24964 -3514 25163 -3483
rect 26106 -3356 26305 -3337
rect 26106 -3485 26130 -3356
rect 26130 -3485 26283 -3356
rect 26283 -3485 26305 -3356
rect 26106 -3516 26305 -3485
rect 16529 -3658 16728 -3627
rect 16529 -3787 16551 -3658
rect 16551 -3787 16704 -3658
rect 16704 -3787 16728 -3658
rect 16529 -3806 16728 -3787
rect 23151 -3657 23350 -3626
rect 23151 -3786 23173 -3657
rect 23173 -3786 23326 -3657
rect 23326 -3786 23350 -3657
rect 23151 -3805 23350 -3786
rect 18342 -4001 18541 -3970
rect 18342 -4130 18364 -4001
rect 18364 -4130 18517 -4001
rect 18517 -4130 18541 -4001
rect 18342 -4149 18541 -4130
rect 20240 -4001 20439 -3970
rect 20240 -4130 20262 -4001
rect 20262 -4130 20415 -4001
rect 20415 -4130 20439 -4001
rect 20240 -4149 20439 -4130
rect 24964 -4000 25163 -3969
rect 24964 -4129 24986 -4000
rect 24986 -4129 25139 -4000
rect 25139 -4129 25163 -4000
rect 24964 -4148 25163 -4129
rect 26862 -4000 27061 -3969
rect 26862 -4129 26884 -4000
rect 26884 -4129 27037 -4000
rect 27037 -4129 27061 -4000
rect 26862 -4148 27061 -4129
rect 16813 -4697 16992 -4675
rect 10158 -4875 10337 -4851
rect 16813 -4850 16832 -4697
rect 16832 -4850 16961 -4697
rect 16961 -4850 16992 -4697
rect 16813 -4874 16992 -4850
rect 23435 -4696 23614 -4674
rect 23435 -4849 23454 -4696
rect 23454 -4849 23583 -4696
rect 23583 -4849 23614 -4696
rect 23435 -4873 23614 -4849
rect 3318 -5261 3517 -5230
rect 3318 -5390 3340 -5261
rect 3340 -5390 3493 -5261
rect 3493 -5390 3517 -5261
rect 3318 -5409 3517 -5390
rect 9869 -5263 10068 -5232
rect 9869 -5392 9891 -5263
rect 9891 -5392 10044 -5263
rect 10044 -5392 10068 -5263
rect 9869 -5411 10068 -5392
rect 16524 -5262 16723 -5231
rect 16524 -5391 16546 -5262
rect 16546 -5391 16699 -5262
rect 16699 -5391 16723 -5262
rect 16524 -5410 16723 -5391
rect 23146 -5261 23345 -5230
rect 23146 -5390 23168 -5261
rect 23168 -5390 23321 -5261
rect 23321 -5390 23345 -5261
rect 23146 -5409 23345 -5390
rect 565 -5860 639 -5854
rect 565 -5922 571 -5860
rect 571 -5922 635 -5860
rect 635 -5922 639 -5860
rect 3602 -6300 3781 -6278
rect 3602 -6453 3621 -6300
rect 3621 -6453 3750 -6300
rect 3750 -6453 3781 -6300
rect 10153 -6302 10332 -6280
rect 3602 -6477 3781 -6453
rect 5080 -6397 5279 -6378
rect 5080 -6526 5104 -6397
rect 5104 -6526 5257 -6397
rect 5257 -6526 5279 -6397
rect 5080 -6557 5279 -6526
rect 6978 -6397 7177 -6378
rect 6978 -6526 7002 -6397
rect 7002 -6526 7155 -6397
rect 7155 -6526 7177 -6397
rect 6978 -6557 7177 -6526
rect 10153 -6455 10172 -6302
rect 10172 -6455 10301 -6302
rect 10301 -6455 10332 -6302
rect 16808 -6301 16987 -6279
rect 10153 -6479 10332 -6455
rect 11631 -6399 11830 -6380
rect 11631 -6528 11655 -6399
rect 11655 -6528 11808 -6399
rect 11808 -6528 11830 -6399
rect 11631 -6559 11830 -6528
rect 13529 -6399 13728 -6380
rect 13529 -6528 13553 -6399
rect 13553 -6528 13706 -6399
rect 13706 -6528 13728 -6399
rect 13529 -6559 13728 -6528
rect 16808 -6454 16827 -6301
rect 16827 -6454 16956 -6301
rect 16956 -6454 16987 -6301
rect 23430 -6300 23609 -6278
rect 16808 -6478 16987 -6454
rect 18286 -6398 18485 -6379
rect 18286 -6527 18310 -6398
rect 18310 -6527 18463 -6398
rect 18463 -6527 18485 -6398
rect 18286 -6558 18485 -6527
rect 20184 -6398 20383 -6379
rect 20184 -6527 20208 -6398
rect 20208 -6527 20361 -6398
rect 20361 -6527 20383 -6398
rect 20184 -6558 20383 -6527
rect 23430 -6453 23449 -6300
rect 23449 -6453 23578 -6300
rect 23578 -6453 23609 -6300
rect 23430 -6477 23609 -6453
rect 24908 -6397 25107 -6378
rect 24908 -6526 24932 -6397
rect 24932 -6526 25085 -6397
rect 25085 -6526 25107 -6397
rect 24908 -6557 25107 -6526
rect 26806 -6397 27005 -6378
rect 26806 -6526 26830 -6397
rect 26830 -6526 26983 -6397
rect 26983 -6526 27005 -6397
rect 26806 -6557 27005 -6526
rect 7275 -7281 7281 -7219
rect 7281 -7281 7345 -7219
rect 7345 -7281 7349 -7219
rect 7275 -7287 7349 -7281
rect 13829 -7276 13835 -7214
rect 13835 -7276 13899 -7214
rect 13899 -7276 13903 -7214
rect 13829 -7282 13903 -7276
rect 20478 -7288 20484 -7226
rect 20484 -7288 20548 -7226
rect 20548 -7288 20552 -7226
rect 20478 -7294 20552 -7288
rect 7053 -8425 7123 -8419
rect 7053 -8487 7059 -8425
rect 7059 -8487 7119 -8425
rect 7119 -8487 7123 -8425
rect 7053 -8491 7123 -8487
rect 13607 -8420 13677 -8414
rect 13607 -8482 13613 -8420
rect 13613 -8482 13673 -8420
rect 13673 -8482 13677 -8420
rect 13607 -8486 13677 -8482
rect 20256 -8432 20326 -8426
rect 20256 -8494 20262 -8432
rect 20262 -8494 20322 -8432
rect 20322 -8494 20326 -8432
rect 20256 -8498 20326 -8494
rect 29162 -3008 29236 -3002
rect 29162 -3070 29168 -3008
rect 29168 -3070 29232 -3008
rect 29232 -3070 29236 -3008
rect 32572 -3478 32910 -3446
rect 32572 -3540 32705 -3478
rect 32705 -3540 32769 -3478
rect 32769 -3540 32910 -3478
rect 32572 -3562 32910 -3540
rect 31027 -4254 31293 -4238
rect 31027 -4411 31050 -4254
rect 31050 -4411 31261 -4254
rect 31261 -4411 31293 -4254
rect 31027 -4433 31293 -4411
rect 28937 -4872 29007 -4868
rect 28937 -4934 28943 -4872
rect 28943 -4934 29003 -4872
rect 29003 -4934 29007 -4872
rect 28937 -4940 29007 -4934
rect 29159 -6078 29233 -6072
rect 29159 -6140 29165 -6078
rect 29165 -6140 29229 -6078
rect 29229 -6140 29233 -6078
rect 31106 -6272 31305 -6241
rect 31106 -6401 31128 -6272
rect 31128 -6401 31281 -6272
rect 31281 -6401 31305 -6272
rect 31106 -6420 31305 -6401
rect 32477 -6620 32547 -6616
rect 32477 -6682 32483 -6620
rect 32483 -6682 32543 -6620
rect 32543 -6682 32547 -6620
rect 32477 -6688 32547 -6682
rect 28944 -7717 29014 -7713
rect 28944 -7779 28950 -7717
rect 28950 -7779 29010 -7717
rect 29010 -7779 29014 -7717
rect 28944 -7785 29014 -7779
rect 32572 -7826 32910 -7794
rect 32572 -7888 32705 -7826
rect 32705 -7888 32769 -7826
rect 32769 -7888 32910 -7826
rect 32572 -7910 32910 -7888
rect 31027 -8602 31293 -8586
rect 31027 -8759 31050 -8602
rect 31050 -8759 31261 -8602
rect 31261 -8759 31293 -8602
rect 31027 -8781 31293 -8759
rect 29166 -8923 29240 -8917
rect 29166 -8985 29172 -8923
rect 29172 -8985 29236 -8923
rect 29236 -8985 29240 -8923
<< metal4 >>
rect 31555 6061 33576 6062
rect 28152 6060 33576 6061
rect 1234 6053 6886 6054
rect 13285 6053 33576 6060
rect 1234 5893 33576 6053
rect 1234 5873 20221 5893
rect 1234 5801 7018 5873
rect 7088 5872 20221 5873
rect 7088 5801 13567 5872
rect 1234 5800 13567 5801
rect 13637 5821 20221 5872
rect 20291 5821 33576 5893
rect 13637 5800 33576 5821
rect 1234 5762 33576 5800
rect 1234 5755 21786 5762
rect 1234 5754 6886 5755
rect 1234 4133 1640 5754
rect 27939 5726 33576 5762
rect 27939 5654 28874 5726
rect 28944 5693 33576 5726
rect 28944 5654 31104 5693
rect 27939 5602 31104 5654
rect 7552 4568 7553 4776
rect 13584 4752 14094 4753
rect 13584 4571 13585 4752
rect 20251 4560 20252 4736
rect 7547 4134 11104 4166
rect 13860 4139 17417 4166
rect 20695 4139 24252 4166
rect 27939 4146 28406 5602
rect 30962 5599 31104 5602
rect 31082 5514 31104 5599
rect 31303 5600 33576 5693
rect 31303 5599 31431 5600
rect 31303 5514 31327 5599
rect 31082 5511 31327 5514
rect 32315 5318 32701 5600
rect 32315 5277 32475 5318
rect 32317 5246 32475 5277
rect 32545 5277 32701 5318
rect 32545 5246 32699 5277
rect 32317 5224 32699 5246
rect 29313 4392 29314 4563
rect 27314 4139 28406 4146
rect 32569 4141 32625 4142
rect 13860 4134 28406 4139
rect 118 4129 4275 4133
rect 7547 4129 28406 4134
rect 118 3973 28406 4129
rect 118 3901 354 3973
rect 424 3946 28406 3973
rect 424 3901 12348 3946
rect 118 3892 12348 3901
rect 118 3879 9866 3892
rect 1239 3858 9866 3879
rect 1239 3804 5799 3858
rect 1239 3625 3317 3804
rect 3516 3679 5799 3804
rect 5998 3679 6946 3858
rect 7145 3713 9866 3858
rect 10065 3767 12348 3892
rect 12547 3767 13495 3946
rect 13694 3892 25627 3946
rect 13694 3878 23145 3892
rect 13694 3824 19002 3878
rect 13694 3767 16520 3824
rect 10065 3713 16520 3767
rect 7145 3679 16520 3713
rect 3516 3645 16520 3679
rect 16719 3699 19002 3824
rect 19201 3699 20149 3878
rect 20348 3713 23145 3878
rect 23344 3767 25627 3892
rect 25826 3767 26774 3946
rect 26973 3767 28406 3946
rect 32565 4140 32625 4141
rect 32862 4141 32901 4142
rect 32862 4140 32916 4141
rect 32565 4024 32570 4140
rect 32908 4024 32916 4140
rect 32565 3883 32625 4024
rect 23344 3713 28406 3767
rect 32862 3883 32916 4024
rect 20348 3699 28406 3713
rect 16719 3645 28406 3699
rect 3516 3625 28406 3645
rect 1239 3507 28406 3625
rect 1239 3506 11104 3507
rect 13657 3506 24252 3507
rect 1239 3419 7724 3506
rect 1239 3404 5133 3419
rect 1239 1535 1917 3404
rect 105 1388 1917 1535
rect 105 1316 346 1388
rect 416 1316 1917 1388
rect 105 1294 1917 1316
rect 1239 -1720 1917 1294
rect 2776 2154 3671 2368
rect 2776 1975 3331 2154
rect 3530 1986 3671 2154
rect 3530 1981 4016 1986
rect 5894 1981 6241 1984
rect 7108 1981 7724 3419
rect 3530 1975 7724 1981
rect 2776 1811 7724 1975
rect 2776 1632 5144 1811
rect 5343 1632 7042 1811
rect 7241 1632 7724 1811
rect 2776 1476 7724 1632
rect 2776 746 2946 1476
rect 7108 1471 7724 1476
rect 9325 2242 10220 2456
rect 9325 2063 9880 2242
rect 10079 2074 10220 2242
rect 10079 2069 10565 2074
rect 12443 2069 12790 2072
rect 13657 2069 14273 3506
rect 16499 3439 20927 3506
rect 10079 2063 14273 2069
rect 9325 1899 14273 2063
rect 9325 1720 11693 1899
rect 11892 1720 13591 1899
rect 13790 1720 14273 1899
rect 9325 1564 14273 1720
rect 9325 834 9495 1564
rect 13657 1559 14273 1564
rect 15979 2174 16874 2388
rect 15979 1995 16534 2174
rect 16733 2006 16874 2174
rect 16733 2001 17219 2006
rect 19097 2001 19444 2004
rect 20311 2001 20927 3439
rect 26936 3484 28406 3507
rect 16733 1995 20927 2001
rect 15979 1831 20927 1995
rect 15979 1652 18347 1831
rect 18546 1652 20245 1831
rect 20444 1652 20927 1831
rect 15979 1496 20927 1652
rect 2776 550 4044 746
rect 2776 371 3326 550
rect 3525 371 4044 550
rect 2776 102 4044 371
rect 9325 638 10593 834
rect 9325 459 9875 638
rect 10074 459 10593 638
rect 9325 190 10593 459
rect 15979 766 16149 1496
rect 20311 1491 20927 1496
rect 22604 2242 23499 2456
rect 22604 2063 23159 2242
rect 23358 2074 23499 2242
rect 23358 2069 23844 2074
rect 25722 2069 26069 2072
rect 26936 2069 27552 3484
rect 23358 2063 27552 2069
rect 22604 1899 27552 2063
rect 22604 1720 24972 1899
rect 25171 1720 26870 1899
rect 27069 1720 27552 1899
rect 22604 1564 27552 1720
rect 22604 834 22774 1564
rect 26936 1559 27552 1564
rect 27939 3253 28406 3484
rect 27939 3155 29421 3253
rect 27939 3083 28869 3155
rect 28939 3083 29421 3155
rect 27939 3015 29421 3083
rect 15979 570 17247 766
rect 15979 391 16529 570
rect 16728 391 17247 570
rect 15979 122 17247 391
rect 22604 638 23872 834
rect 22604 459 23154 638
rect 23353 459 23872 638
rect 22604 190 23872 459
rect 27939 237 28406 3015
rect 28959 2000 29318 2002
rect 30847 1767 32200 1778
rect 33044 1767 33576 5600
rect 30847 1602 33576 1767
rect 30847 1508 31106 1602
rect 31084 1423 31106 1508
rect 31305 1508 33576 1602
rect 31305 1423 31329 1508
rect 32002 1506 33576 1508
rect 31084 1420 31329 1423
rect 32317 1227 32703 1506
rect 32317 1186 32477 1227
rect 32319 1155 32477 1186
rect 32547 1186 32703 1227
rect 32547 1155 32701 1186
rect 32319 1133 32701 1155
rect 27939 122 29424 237
rect 27939 50 28869 122
rect 28939 50 29424 122
rect 32571 50 32627 51
rect 27939 -1 29424 50
rect 32567 49 32627 50
rect 32864 50 32903 51
rect 32864 49 32918 50
rect 5064 -598 5309 -595
rect 5064 -616 5088 -598
rect 5287 -616 5309 -598
rect 6962 -598 7207 -595
rect 6962 -616 6986 -598
rect 7185 -616 7207 -598
rect 11613 -510 11858 -507
rect 11613 -528 11637 -510
rect 11836 -528 11858 -510
rect 13511 -510 13756 -507
rect 13511 -528 13535 -510
rect 13734 -528 13756 -510
rect 4960 -920 4984 -683
rect 5494 -920 6830 -734
rect 11509 -832 11533 -595
rect 12043 -832 13379 -646
rect 18267 -578 18512 -575
rect 18267 -596 18291 -578
rect 18490 -596 18512 -578
rect 20165 -578 20410 -575
rect 20165 -596 20189 -578
rect 20388 -596 20410 -578
rect 11509 -837 13876 -832
rect 11897 -839 13568 -837
rect 18163 -900 18187 -663
rect 18697 -900 20033 -714
rect 24892 -510 25137 -507
rect 24892 -528 24916 -510
rect 25115 -528 25137 -510
rect 26790 -510 27035 -507
rect 26790 -528 26814 -510
rect 27013 -528 27035 -510
rect 24788 -832 24812 -595
rect 25322 -832 26658 -646
rect 24788 -837 27155 -832
rect 25176 -839 26847 -837
rect 18163 -905 20530 -900
rect 18551 -907 20222 -905
rect 4960 -925 7327 -920
rect 5348 -927 7019 -925
rect 27939 -1458 28406 -1
rect 32567 -67 32572 49
rect 32910 -67 32918 49
rect 32567 -208 32627 -67
rect 32864 -208 32918 -67
rect 28960 -1038 29321 -1036
rect 28959 -1193 28960 -1038
rect 29320 -1196 29321 -1038
rect 33044 -1455 33576 1506
rect 32225 -1458 33576 -1455
rect 9838 -1720 14271 -1714
rect 16493 -1720 20926 -1706
rect 23115 -1720 27548 -1704
rect 27939 -1720 33576 -1458
rect 1239 -1761 33576 -1720
rect 98 -1798 33576 -1761
rect 98 -1870 28940 -1798
rect 29010 -1870 33576 -1798
rect 98 -1890 33576 -1870
rect 98 -1962 327 -1890
rect 397 -1893 33576 -1890
rect 397 -1922 31106 -1893
rect 397 -1962 5791 -1922
rect 98 -1976 5791 -1962
rect 98 -2002 3309 -1976
rect 1239 -2155 3309 -2002
rect 3508 -2101 5791 -1976
rect 5990 -2101 6938 -1922
rect 7137 -1923 25619 -1922
rect 7137 -1924 18997 -1923
rect 7137 -1978 12342 -1924
rect 7137 -2101 9860 -1978
rect 3508 -2155 9860 -2101
rect 1239 -2157 9860 -2155
rect 10059 -2103 12342 -1978
rect 12541 -2103 13489 -1924
rect 13688 -1977 18997 -1924
rect 13688 -2103 16515 -1977
rect 10059 -2156 16515 -2103
rect 16714 -2102 18997 -1977
rect 19196 -2102 20144 -1923
rect 20343 -1976 25619 -1923
rect 20343 -2102 23137 -1976
rect 16714 -2155 23137 -2102
rect 23336 -2101 25619 -1976
rect 25818 -2101 26766 -1922
rect 26965 -1995 31106 -1922
rect 26965 -2101 28406 -1995
rect 31084 -2072 31106 -1995
rect 31305 -1995 33576 -1893
rect 31305 -2072 31329 -1995
rect 32225 -2000 33576 -1995
rect 31084 -2075 31329 -2072
rect 23336 -2155 28406 -2101
rect 16714 -2156 28406 -2155
rect 10059 -2157 28406 -2156
rect 1239 -2383 28406 -2157
rect 32317 -2268 32703 -2000
rect 32317 -2309 32477 -2268
rect 32319 -2340 32477 -2309
rect 32547 -2309 32703 -2268
rect 32547 -2340 32701 -2309
rect 32319 -2362 32701 -2340
rect 1239 -4518 1917 -2383
rect 92 -4650 1917 -4518
rect 92 -4722 343 -4650
rect 413 -4722 1917 -4650
rect 92 -4759 1917 -4722
rect 1239 -8374 1917 -4759
rect 2768 -3626 3663 -3412
rect 2768 -3805 3323 -3626
rect 3522 -3794 3663 -3626
rect 3522 -3799 4008 -3794
rect 5886 -3799 6233 -3796
rect 7100 -3799 7716 -2383
rect 3522 -3805 7716 -3799
rect 2768 -3969 7716 -3805
rect 2768 -4148 5136 -3969
rect 5335 -4148 7034 -3969
rect 7233 -4148 7716 -3969
rect 2768 -4304 7716 -4148
rect 2768 -5034 2938 -4304
rect 7100 -4309 7716 -4304
rect 9319 -3628 10214 -3414
rect 9319 -3807 9874 -3628
rect 10073 -3796 10214 -3628
rect 10073 -3801 10559 -3796
rect 12437 -3801 12784 -3798
rect 13651 -3801 14267 -2383
rect 10073 -3807 14267 -3801
rect 9319 -3971 14267 -3807
rect 9319 -4150 11687 -3971
rect 11886 -4150 13585 -3971
rect 13784 -4150 14267 -3971
rect 9319 -4306 14267 -4150
rect 2768 -5230 4036 -5034
rect 2768 -5409 3318 -5230
rect 3517 -5409 4036 -5230
rect 2768 -5678 4036 -5409
rect 9319 -5036 9489 -4306
rect 13651 -4311 14267 -4306
rect 15974 -3627 16869 -3413
rect 15974 -3806 16529 -3627
rect 16728 -3795 16869 -3627
rect 16728 -3800 17214 -3795
rect 19092 -3800 19439 -3797
rect 20306 -3800 20922 -2383
rect 16728 -3806 20922 -3800
rect 15974 -3970 20922 -3806
rect 15974 -4149 18342 -3970
rect 18541 -4149 20240 -3970
rect 20439 -4149 20922 -3970
rect 15974 -4305 20922 -4149
rect 15974 -5035 16144 -4305
rect 20306 -4310 20922 -4305
rect 22596 -3626 23491 -3412
rect 22596 -3805 23151 -3626
rect 23350 -3794 23491 -3626
rect 23350 -3799 23836 -3794
rect 25714 -3799 26061 -3796
rect 26928 -3799 27544 -2383
rect 23350 -3805 27544 -3799
rect 22596 -3969 27544 -3805
rect 22596 -4148 24964 -3969
rect 25163 -4148 26862 -3969
rect 27061 -4148 27544 -3969
rect 22596 -4304 27544 -4148
rect 22596 -5034 22766 -4304
rect 26928 -4309 27544 -4304
rect 27939 -4775 28406 -2383
rect 29020 -2959 29383 -2958
rect 29380 -3119 29383 -2959
rect 32571 -3445 32627 -3444
rect 32567 -3446 32627 -3445
rect 32864 -3445 32903 -3444
rect 32864 -3446 32918 -3445
rect 32567 -3562 32572 -3446
rect 32910 -3562 32918 -3446
rect 32567 -3703 32627 -3562
rect 32864 -3703 32918 -3562
rect 30964 -4575 31337 -4505
rect 27939 -4868 29424 -4775
rect 27939 -4940 28937 -4868
rect 29007 -4940 29424 -4868
rect 27939 -5013 29424 -4940
rect 9319 -5232 10587 -5036
rect 9319 -5411 9869 -5232
rect 10068 -5411 10587 -5232
rect 9319 -5680 10587 -5411
rect 15974 -5231 17242 -5035
rect 15974 -5410 16524 -5231
rect 16723 -5410 17242 -5231
rect 15974 -5679 17242 -5410
rect 22596 -5230 23864 -5034
rect 22596 -5409 23146 -5230
rect 23345 -5409 23864 -5230
rect 22596 -5678 23864 -5409
rect 5056 -6378 5301 -6375
rect 5056 -6396 5080 -6378
rect 5279 -6396 5301 -6378
rect 6954 -6378 7199 -6375
rect 6954 -6396 6978 -6378
rect 7177 -6396 7199 -6378
rect 4952 -6700 4976 -6463
rect 5486 -6700 6822 -6514
rect 11607 -6380 11852 -6377
rect 11607 -6398 11631 -6380
rect 11830 -6398 11852 -6380
rect 13505 -6380 13750 -6377
rect 13505 -6398 13529 -6380
rect 13728 -6398 13750 -6380
rect 4952 -6705 7319 -6700
rect 11503 -6702 11527 -6465
rect 12037 -6702 13373 -6516
rect 18262 -6379 18507 -6376
rect 18262 -6397 18286 -6379
rect 18485 -6397 18507 -6379
rect 20160 -6379 20405 -6376
rect 20160 -6397 20184 -6379
rect 20383 -6397 20405 -6379
rect 18158 -6701 18182 -6464
rect 18692 -6701 20028 -6515
rect 24884 -6378 25129 -6375
rect 24884 -6396 24908 -6378
rect 25107 -6396 25129 -6378
rect 26782 -6378 27027 -6375
rect 26782 -6396 26806 -6378
rect 27005 -6396 27027 -6378
rect 24780 -6700 24804 -6463
rect 25314 -6700 26650 -6514
rect 5340 -6707 7011 -6705
rect 11503 -6707 13870 -6702
rect 18158 -6706 20525 -6701
rect 24780 -6705 27147 -6700
rect 11891 -6709 13562 -6707
rect 18546 -6708 20217 -6706
rect 25168 -6707 26839 -6705
rect 27939 -7587 28406 -5013
rect 29015 -6027 29377 -6026
rect 29015 -6201 29016 -6027
rect 29376 -6201 29377 -6027
rect 31373 -6092 32511 -6090
rect 33044 -6092 33576 -2000
rect 31373 -6093 33576 -6092
rect 30899 -6241 33576 -6093
rect 30899 -6339 31106 -6241
rect 31084 -6420 31106 -6339
rect 31305 -6334 33576 -6241
rect 31305 -6339 31756 -6334
rect 32317 -6336 33576 -6334
rect 31305 -6420 31329 -6339
rect 31084 -6423 31329 -6420
rect 32317 -6616 32703 -6336
rect 32317 -6657 32477 -6616
rect 32319 -6688 32477 -6657
rect 32547 -6657 32703 -6616
rect 32547 -6688 32701 -6657
rect 32319 -6710 32701 -6688
rect 27939 -7713 29418 -7587
rect 27939 -7785 28944 -7713
rect 29014 -7785 29418 -7713
rect 27939 -7825 29418 -7785
rect 32571 -7793 32627 -7792
rect 32567 -7794 32627 -7793
rect 32864 -7793 32903 -7792
rect 32864 -7794 32918 -7793
rect 27939 -8374 28406 -7825
rect 32567 -7910 32572 -7794
rect 32910 -7910 32918 -7794
rect 32567 -8051 32627 -7910
rect 32864 -8051 32918 -7910
rect 1234 -8414 28408 -8374
rect 1234 -8419 13607 -8414
rect 1234 -8491 7053 -8419
rect 7123 -8486 13607 -8419
rect 13677 -8426 28408 -8414
rect 13677 -8486 20256 -8426
rect 7123 -8491 20256 -8486
rect 1234 -8498 20256 -8491
rect 20326 -8498 28408 -8426
rect 1234 -8628 28408 -8498
rect 29025 -9038 29026 -8880
rect 29386 -9038 29387 -8880
<< via4 >>
rect 7043 4669 7552 4777
rect 7043 4601 7240 4669
rect 7240 4601 7314 4669
rect 7314 4601 7552 4669
rect 7043 4469 7552 4601
rect 13585 4668 14094 4752
rect 13585 4600 13789 4668
rect 13789 4600 13863 4668
rect 13863 4600 14094 4668
rect 13585 4444 14094 4600
rect 20252 4689 20761 4737
rect 20252 4621 20443 4689
rect 20443 4621 20517 4689
rect 20517 4621 20761 4689
rect 20252 4430 20761 4621
rect 28953 4522 29313 4563
rect 28953 4454 29096 4522
rect 29096 4454 29170 4522
rect 29170 4454 29313 4522
rect 28953 4290 29313 4454
rect 32625 4140 32862 4199
rect 32625 4024 32862 4140
rect 32625 3742 32862 4024
rect 380 2769 888 2839
rect 380 2701 576 2769
rect 576 2701 650 2769
rect 650 2701 888 2769
rect 380 2531 888 2701
rect 3542 2756 4052 2834
rect 3542 2557 3601 2756
rect 3601 2557 3780 2756
rect 3780 2557 4052 2756
rect 3542 2530 4052 2557
rect 5110 2445 5414 2596
rect 355 184 863 257
rect 355 116 568 184
rect 568 116 642 184
rect 642 116 863 184
rect 355 -51 863 116
rect 5110 2266 5144 2445
rect 5144 2266 5343 2445
rect 5343 2266 5414 2445
rect 5110 2086 5414 2266
rect 6244 2443 6548 2606
rect 6244 2264 6286 2443
rect 6286 2264 6485 2443
rect 6485 2264 6548 2443
rect 6244 2096 6548 2264
rect 10091 2844 10601 2922
rect 10091 2645 10150 2844
rect 10150 2645 10329 2844
rect 10329 2645 10601 2844
rect 10091 2618 10601 2645
rect 11659 2533 11963 2684
rect 11659 2354 11693 2533
rect 11693 2354 11892 2533
rect 11892 2354 11963 2533
rect 11659 2174 11963 2354
rect 12793 2531 13097 2694
rect 12793 2352 12835 2531
rect 12835 2352 13034 2531
rect 13034 2352 13097 2531
rect 12793 2184 13097 2352
rect 16745 2776 17255 2854
rect 16745 2577 16804 2776
rect 16804 2577 16983 2776
rect 16983 2577 17255 2776
rect 16745 2550 17255 2577
rect 18313 2465 18617 2616
rect 3536 1106 4046 1174
rect 3536 907 3615 1106
rect 3615 907 3794 1106
rect 3794 907 4046 1106
rect 3536 870 4046 907
rect 18313 2286 18347 2465
rect 18347 2286 18546 2465
rect 18546 2286 18617 2465
rect 18313 2106 18617 2286
rect 19447 2463 19751 2626
rect 19447 2284 19489 2463
rect 19489 2284 19688 2463
rect 19688 2284 19751 2463
rect 19447 2116 19751 2284
rect 23370 2844 23880 2922
rect 23370 2645 23429 2844
rect 23429 2645 23608 2844
rect 23608 2645 23880 2844
rect 23370 2618 23880 2645
rect 24938 2533 25242 2684
rect 10085 1194 10595 1262
rect 10085 995 10164 1194
rect 10164 995 10343 1194
rect 10343 995 10595 1194
rect 10085 958 10595 995
rect 24938 2354 24972 2533
rect 24972 2354 25171 2533
rect 25171 2354 25242 2533
rect 24938 2174 25242 2354
rect 26072 2531 26376 2694
rect 26072 2352 26114 2531
rect 26114 2352 26313 2531
rect 26313 2352 26376 2531
rect 26072 2184 26376 2352
rect 16739 1126 17249 1194
rect 16739 927 16818 1126
rect 16818 927 16997 1126
rect 16997 927 17249 1126
rect 16739 890 17249 927
rect 30962 3348 31335 3350
rect 30962 3153 31025 3348
rect 31025 3153 31291 3348
rect 31291 3153 31335 3348
rect 23364 1194 23874 1262
rect 23364 995 23443 1194
rect 23443 995 23622 1194
rect 23622 995 23874 1194
rect 23364 958 23874 995
rect 30962 3011 31335 3153
rect 28959 1951 29319 2000
rect 28959 1883 29091 1951
rect 29091 1883 29165 1951
rect 29165 1883 29319 1951
rect 28959 1727 29319 1883
rect 32627 49 32864 108
rect 10084 -410 10594 -343
rect 3535 -498 4045 -431
rect 3535 -697 3610 -498
rect 3610 -697 3789 -498
rect 3789 -697 4045 -498
rect 10084 -609 10159 -410
rect 10159 -609 10338 -410
rect 10338 -609 10594 -410
rect 23363 -410 23873 -343
rect 16738 -478 17248 -411
rect 3535 -735 4045 -697
rect 4984 -777 5088 -616
rect 5088 -777 5287 -616
rect 5287 -777 5494 -616
rect 4984 -920 5494 -777
rect 6830 -777 6986 -616
rect 6986 -777 7185 -616
rect 7185 -777 7340 -616
rect 10084 -647 10594 -609
rect 6830 -920 7340 -777
rect 11533 -689 11637 -528
rect 11637 -689 11836 -528
rect 11836 -689 12043 -528
rect 11533 -832 12043 -689
rect 13379 -689 13535 -528
rect 13535 -689 13734 -528
rect 13734 -689 13889 -528
rect 13379 -832 13889 -689
rect 16738 -677 16813 -478
rect 16813 -677 16992 -478
rect 16992 -677 17248 -478
rect 16738 -715 17248 -677
rect 18187 -757 18291 -596
rect 18291 -757 18490 -596
rect 18490 -757 18697 -596
rect 18187 -900 18697 -757
rect 20033 -757 20189 -596
rect 20189 -757 20388 -596
rect 20388 -757 20543 -596
rect 23363 -609 23438 -410
rect 23438 -609 23617 -410
rect 23617 -609 23873 -410
rect 23363 -647 23873 -609
rect 20033 -900 20543 -757
rect 24812 -689 24916 -528
rect 24916 -689 25115 -528
rect 25115 -689 25322 -528
rect 24812 -832 25322 -689
rect 26658 -689 26814 -528
rect 26814 -689 27013 -528
rect 27013 -689 27168 -528
rect 26658 -832 27168 -689
rect 32627 -67 32864 49
rect 32627 -349 32864 -67
rect 30964 -743 31337 -741
rect 30964 -938 31027 -743
rect 31027 -938 31293 -743
rect 31293 -938 31337 -743
rect 28960 -1082 29320 -1038
rect 28960 -1150 29091 -1082
rect 29091 -1150 29165 -1082
rect 29165 -1150 29320 -1082
rect 28960 -1311 29320 -1150
rect 30964 -1080 31337 -938
rect 331 -3094 839 -3048
rect 331 -3162 549 -3094
rect 549 -3162 623 -3094
rect 623 -3162 839 -3094
rect 331 -3356 839 -3162
rect 3534 -3024 4044 -2946
rect 3534 -3223 3593 -3024
rect 3593 -3223 3772 -3024
rect 3772 -3223 4044 -3024
rect 3534 -3250 4044 -3223
rect 5102 -3335 5406 -3184
rect 306 -5854 814 -5812
rect 306 -5922 565 -5854
rect 565 -5922 639 -5854
rect 639 -5922 814 -5854
rect 306 -6120 814 -5922
rect 5102 -3514 5136 -3335
rect 5136 -3514 5335 -3335
rect 5335 -3514 5406 -3335
rect 5102 -3694 5406 -3514
rect 6236 -3337 6540 -3174
rect 6236 -3516 6278 -3337
rect 6278 -3516 6477 -3337
rect 6477 -3516 6540 -3337
rect 6236 -3684 6540 -3516
rect 10085 -3026 10595 -2948
rect 10085 -3225 10144 -3026
rect 10144 -3225 10323 -3026
rect 10323 -3225 10595 -3026
rect 10085 -3252 10595 -3225
rect 11653 -3337 11957 -3186
rect 11653 -3516 11687 -3337
rect 11687 -3516 11886 -3337
rect 11886 -3516 11957 -3337
rect 11653 -3696 11957 -3516
rect 12787 -3339 13091 -3176
rect 12787 -3518 12829 -3339
rect 12829 -3518 13028 -3339
rect 13028 -3518 13091 -3339
rect 12787 -3686 13091 -3518
rect 16740 -3025 17250 -2947
rect 16740 -3224 16799 -3025
rect 16799 -3224 16978 -3025
rect 16978 -3224 17250 -3025
rect 16740 -3251 17250 -3224
rect 18308 -3336 18612 -3185
rect 3528 -4674 4038 -4606
rect 3528 -4873 3607 -4674
rect 3607 -4873 3786 -4674
rect 3786 -4873 4038 -4674
rect 3528 -4910 4038 -4873
rect 18308 -3515 18342 -3336
rect 18342 -3515 18541 -3336
rect 18541 -3515 18612 -3336
rect 18308 -3695 18612 -3515
rect 19442 -3338 19746 -3175
rect 19442 -3517 19484 -3338
rect 19484 -3517 19683 -3338
rect 19683 -3517 19746 -3338
rect 19442 -3685 19746 -3517
rect 23362 -3024 23872 -2946
rect 23362 -3223 23421 -3024
rect 23421 -3223 23600 -3024
rect 23600 -3223 23872 -3024
rect 23362 -3250 23872 -3223
rect 24930 -3335 25234 -3184
rect 10079 -4676 10589 -4608
rect 10079 -4875 10158 -4676
rect 10158 -4875 10337 -4676
rect 10337 -4875 10589 -4676
rect 10079 -4912 10589 -4875
rect 24930 -3514 24964 -3335
rect 24964 -3514 25163 -3335
rect 25163 -3514 25234 -3335
rect 24930 -3694 25234 -3514
rect 26064 -3337 26368 -3174
rect 26064 -3516 26106 -3337
rect 26106 -3516 26305 -3337
rect 26305 -3516 26368 -3337
rect 26064 -3684 26368 -3516
rect 16734 -4675 17244 -4607
rect 16734 -4874 16813 -4675
rect 16813 -4874 16992 -4675
rect 16992 -4874 17244 -4675
rect 16734 -4911 17244 -4874
rect 23356 -4674 23866 -4606
rect 23356 -4873 23435 -4674
rect 23435 -4873 23614 -4674
rect 23614 -4873 23866 -4674
rect 23356 -4910 23866 -4873
rect 29020 -3002 29380 -2959
rect 29020 -3070 29162 -3002
rect 29162 -3070 29236 -3002
rect 29236 -3070 29380 -3002
rect 29020 -3232 29380 -3070
rect 32627 -3446 32864 -3387
rect 32627 -3562 32864 -3446
rect 32627 -3844 32864 -3562
rect 30964 -4238 31337 -4236
rect 30964 -4433 31027 -4238
rect 31027 -4433 31293 -4238
rect 31293 -4433 31337 -4238
rect 30964 -4505 31337 -4433
rect 3527 -6278 4037 -6211
rect 3527 -6477 3602 -6278
rect 3602 -6477 3781 -6278
rect 3781 -6477 4037 -6278
rect 10078 -6280 10588 -6213
rect 3527 -6515 4037 -6477
rect 4976 -6557 5080 -6396
rect 5080 -6557 5279 -6396
rect 5279 -6557 5486 -6396
rect 4976 -6700 5486 -6557
rect 6822 -6557 6978 -6396
rect 6978 -6557 7177 -6396
rect 7177 -6557 7332 -6396
rect 10078 -6479 10153 -6280
rect 10153 -6479 10332 -6280
rect 10332 -6479 10588 -6280
rect 16733 -6279 17243 -6212
rect 10078 -6517 10588 -6479
rect 6822 -6700 7332 -6557
rect 11527 -6559 11631 -6398
rect 11631 -6559 11830 -6398
rect 11830 -6559 12037 -6398
rect 11527 -6702 12037 -6559
rect 13373 -6559 13529 -6398
rect 13529 -6559 13728 -6398
rect 13728 -6559 13883 -6398
rect 16733 -6478 16808 -6279
rect 16808 -6478 16987 -6279
rect 16987 -6478 17243 -6279
rect 23355 -6278 23865 -6211
rect 16733 -6516 17243 -6478
rect 13373 -6702 13883 -6559
rect 18182 -6558 18286 -6397
rect 18286 -6558 18485 -6397
rect 18485 -6558 18692 -6397
rect 18182 -6701 18692 -6558
rect 20028 -6558 20184 -6397
rect 20184 -6558 20383 -6397
rect 20383 -6558 20538 -6397
rect 23355 -6477 23430 -6278
rect 23430 -6477 23609 -6278
rect 23609 -6477 23865 -6278
rect 23355 -6515 23865 -6477
rect 20028 -6701 20538 -6558
rect 24804 -6557 24908 -6396
rect 24908 -6557 25107 -6396
rect 25107 -6557 25314 -6396
rect 24804 -6700 25314 -6557
rect 26650 -6557 26806 -6396
rect 26806 -6557 27005 -6396
rect 27005 -6557 27160 -6396
rect 26650 -6700 27160 -6557
rect 7005 -7219 7513 -7029
rect 7005 -7287 7275 -7219
rect 7275 -7287 7349 -7219
rect 7349 -7287 7513 -7219
rect 7005 -7337 7513 -7287
rect 13544 -7214 14052 -7048
rect 13544 -7282 13829 -7214
rect 13829 -7282 13903 -7214
rect 13903 -7282 14052 -7214
rect 13544 -7356 14052 -7282
rect 20250 -7226 20758 -7073
rect 20250 -7294 20478 -7226
rect 20478 -7294 20552 -7226
rect 20552 -7294 20758 -7226
rect 20250 -7381 20758 -7294
rect 29016 -6072 29376 -6027
rect 29016 -6140 29159 -6072
rect 29159 -6140 29233 -6072
rect 29233 -6140 29376 -6072
rect 29016 -6300 29376 -6140
rect 32627 -7794 32864 -7735
rect 32627 -7910 32864 -7794
rect 32627 -8192 32864 -7910
rect 30964 -8586 31337 -8584
rect 30964 -8781 31027 -8586
rect 31027 -8781 31293 -8586
rect 31293 -8781 31337 -8586
rect 29026 -8917 29386 -8880
rect 29026 -8985 29166 -8917
rect 29166 -8985 29240 -8917
rect 29240 -8985 29386 -8917
rect 29026 -9153 29386 -8985
rect 30964 -8923 31337 -8781
<< metal5 >>
rect -12 4777 33014 5359
rect -12 4469 7043 4777
rect 7552 4752 33014 4777
rect 7552 4469 13585 4752
rect -12 4444 13585 4469
rect 14094 4737 33014 4752
rect 14094 4444 20252 4737
rect -12 4430 20252 4444
rect 20761 4563 33014 4737
rect 20761 4430 28953 4563
rect -12 4290 28953 4430
rect 29313 4290 33014 4563
rect -12 4199 33014 4290
rect -12 3742 32625 4199
rect 32862 3742 33014 4199
rect -12 3350 33014 3742
rect -12 3011 30962 3350
rect 31335 3011 33014 3350
rect -12 2922 33014 3011
rect -12 2839 10091 2922
rect -12 2531 380 2839
rect 888 2834 10091 2839
rect 888 2531 3542 2834
rect -12 2530 3542 2531
rect 4052 2618 10091 2834
rect 10601 2854 23370 2922
rect 10601 2694 16745 2854
rect 10601 2684 12793 2694
rect 10601 2618 11659 2684
rect 4052 2606 11659 2618
rect 4052 2596 6244 2606
rect 4052 2530 5110 2596
rect -12 2086 5110 2530
rect 5414 2096 6244 2596
rect 6548 2174 11659 2606
rect 11963 2184 12793 2684
rect 13097 2550 16745 2694
rect 17255 2626 23370 2854
rect 17255 2616 19447 2626
rect 17255 2550 18313 2616
rect 13097 2184 18313 2550
rect 11963 2174 18313 2184
rect 6548 2106 18313 2174
rect 18617 2116 19447 2616
rect 19751 2618 23370 2626
rect 23880 2694 33014 2922
rect 23880 2684 26072 2694
rect 23880 2618 24938 2684
rect 19751 2174 24938 2618
rect 25242 2184 26072 2684
rect 26376 2184 33014 2694
rect 25242 2174 33014 2184
rect 19751 2116 33014 2174
rect 18617 2106 33014 2116
rect 6548 2096 33014 2106
rect 5414 2086 33014 2096
rect -12 2000 33014 2086
rect -12 1727 28959 2000
rect 29319 1727 33014 2000
rect -12 1262 33014 1727
rect -12 1174 10085 1262
rect -12 870 3536 1174
rect 4046 958 10085 1174
rect 10595 1194 23364 1262
rect 10595 958 16739 1194
rect 4046 890 16739 958
rect 17249 958 23364 1194
rect 23874 958 33014 1262
rect 17249 890 33014 958
rect 4046 870 33014 890
rect -12 257 33014 870
rect -12 -51 355 257
rect 863 108 33014 257
rect 863 -51 32627 108
rect -12 -343 32627 -51
rect -12 -431 10084 -343
rect -12 -735 3535 -431
rect 4045 -616 10084 -431
rect 4045 -735 4984 -616
rect -12 -920 4984 -735
rect 5494 -920 6830 -616
rect 7340 -647 10084 -616
rect 10594 -411 23363 -343
rect 10594 -528 16738 -411
rect 10594 -647 11533 -528
rect 7340 -832 11533 -647
rect 12043 -832 13379 -528
rect 13889 -715 16738 -528
rect 17248 -596 23363 -411
rect 17248 -715 18187 -596
rect 13889 -832 18187 -715
rect 7340 -900 18187 -832
rect 18697 -900 20033 -596
rect 20543 -647 23363 -596
rect 23873 -349 32627 -343
rect 32864 -349 33014 108
rect 23873 -528 33014 -349
rect 23873 -647 24812 -528
rect 20543 -832 24812 -647
rect 25322 -832 26658 -528
rect 27168 -741 33014 -528
rect 27168 -832 30964 -741
rect 20543 -900 30964 -832
rect 7340 -920 30964 -900
rect -12 -1038 30964 -920
rect -12 -1311 28960 -1038
rect 29320 -1080 30964 -1038
rect 31337 -1080 33014 -741
rect 29320 -1311 33014 -1080
rect -12 -2946 33014 -1311
rect -12 -3048 3534 -2946
rect -12 -3356 331 -3048
rect 839 -3250 3534 -3048
rect 4044 -2947 23362 -2946
rect 4044 -2948 16740 -2947
rect 4044 -3174 10085 -2948
rect 4044 -3184 6236 -3174
rect 4044 -3250 5102 -3184
rect 839 -3356 5102 -3250
rect -12 -3694 5102 -3356
rect 5406 -3684 6236 -3184
rect 6540 -3252 10085 -3174
rect 10595 -3176 16740 -2948
rect 10595 -3186 12787 -3176
rect 10595 -3252 11653 -3186
rect 6540 -3684 11653 -3252
rect 5406 -3694 11653 -3684
rect -12 -3696 11653 -3694
rect 11957 -3686 12787 -3186
rect 13091 -3251 16740 -3176
rect 17250 -3175 23362 -2947
rect 17250 -3185 19442 -3175
rect 17250 -3251 18308 -3185
rect 13091 -3686 18308 -3251
rect 11957 -3695 18308 -3686
rect 18612 -3685 19442 -3185
rect 19746 -3250 23362 -3175
rect 23872 -2959 33014 -2946
rect 23872 -3174 29020 -2959
rect 23872 -3184 26064 -3174
rect 23872 -3250 24930 -3184
rect 19746 -3685 24930 -3250
rect 18612 -3694 24930 -3685
rect 25234 -3684 26064 -3184
rect 26368 -3232 29020 -3174
rect 29380 -3232 33014 -2959
rect 26368 -3387 33014 -3232
rect 26368 -3684 32627 -3387
rect 25234 -3694 32627 -3684
rect 18612 -3695 32627 -3694
rect 11957 -3696 32627 -3695
rect -12 -3844 32627 -3696
rect 32864 -3844 33014 -3387
rect -12 -4236 33014 -3844
rect -12 -4505 30964 -4236
rect 31337 -4505 33014 -4236
rect -12 -4606 33014 -4505
rect -12 -4910 3528 -4606
rect 4038 -4607 23356 -4606
rect 4038 -4608 16734 -4607
rect 4038 -4910 10079 -4608
rect -12 -4912 10079 -4910
rect 10589 -4911 16734 -4608
rect 17244 -4910 23356 -4607
rect 23866 -4910 33014 -4606
rect 17244 -4911 33014 -4910
rect 10589 -4912 33014 -4911
rect -12 -5812 33014 -4912
rect -12 -6120 306 -5812
rect 814 -6027 33014 -5812
rect 814 -6120 29016 -6027
rect -12 -6211 29016 -6120
rect -12 -6515 3527 -6211
rect 4037 -6212 23355 -6211
rect 4037 -6213 16733 -6212
rect 4037 -6396 10078 -6213
rect 4037 -6515 4976 -6396
rect -12 -6700 4976 -6515
rect 5486 -6700 6822 -6396
rect 7332 -6517 10078 -6396
rect 10588 -6398 16733 -6213
rect 10588 -6517 11527 -6398
rect 7332 -6700 11527 -6517
rect -12 -6702 11527 -6700
rect 12037 -6702 13373 -6398
rect 13883 -6516 16733 -6398
rect 17243 -6397 23355 -6212
rect 17243 -6516 18182 -6397
rect 13883 -6701 18182 -6516
rect 18692 -6701 20028 -6397
rect 20538 -6515 23355 -6397
rect 23865 -6300 29016 -6211
rect 29376 -6300 33014 -6027
rect 23865 -6396 33014 -6300
rect 23865 -6515 24804 -6396
rect 20538 -6700 24804 -6515
rect 25314 -6700 26650 -6396
rect 27160 -6700 33014 -6396
rect 20538 -6701 33014 -6700
rect 13883 -6702 33014 -6701
rect -12 -7029 33014 -6702
rect -12 -7337 7005 -7029
rect 7513 -7048 33014 -7029
rect 7513 -7337 13544 -7048
rect -12 -7356 13544 -7337
rect 14052 -7073 33014 -7048
rect 14052 -7356 20250 -7073
rect -12 -7381 20250 -7356
rect 20758 -7381 33014 -7073
rect -12 -7735 33014 -7381
rect -12 -8192 32627 -7735
rect 32864 -8192 33014 -7735
rect -12 -8584 33014 -8192
rect -12 -8880 30964 -8584
rect -12 -9153 29026 -8880
rect 29386 -8923 30964 -8880
rect 31337 -8923 33014 -8584
rect 29386 -9153 33014 -8923
rect -12 -9324 33014 -9153
<< labels >>
flabel metal1 27898 -9586 28038 -9452 1 FreeSans 400 0 0 0 Y[5]
port 1 n
flabel metal1 27805 6127 27905 6226 1 FreeSans 400 0 0 0 Y[7]
port 2 n
flabel metal1 27990 6127 28075 6226 1 FreeSans 400 0 0 0 Y[6]
port 3 n
flabel metal1 29723 6128 29802 6221 1 FreeSans 400 0 0 0 Y[0]
port 8 n
flabel metal1 -1114 2912 -1028 3000 1 FreeSans 400 0 0 0 A[1]
port 9 n
flabel metal1 -1114 2723 -1028 2811 1 FreeSans 400 0 0 0 B[1]
port 10 n
flabel metal1 -1113 -5549 -1027 -5465 1 FreeSans 400 0 0 0 B[0]
port 11 n
flabel metal1 -1113 -5677 -1027 -5593 1 FreeSans 400 0 0 0 A[3]
port 12 n
flabel metal1 -1113 102 -1027 186 1 FreeSans 400 0 0 0 A[2]
port 13 n
flabel metal1 -1113 -8770 -1026 -8692 1 FreeSans 400 0 0 0 B[2]
port 14 n
flabel metal1 -1114 -9316 -1026 -9234 1 FreeSans 400 0 0 0 B[3]
port 15 n
flabel metal1 -1114 4277 -1028 4334 1 FreeSans 400 0 0 0 A[0]
port 16 n
flabel metal4 15993 5772 17296 6035 1 FreeSans 2000 0 0 0 VDD
port 17 n
flabel metal5 15993 -7715 17296 -7452 1 FreeSans 2000 0 0 0 VSS
port 18 n
flabel metal1 33660 4285 33769 4384 1 FreeSans 400 0 0 0 Y[2]
port 19 n
flabel metal1 33659 197 33765 291 1 FreeSans 400 0 0 0 Y[1]
port 20 n
flabel metal1 33659 -3294 33769 -3201 1 FreeSans 400 0 0 0 Y[4]
port 21 n
flabel metal1 33660 -7645 33772 -7546 1 FreeSans 400 0 0 0 Y[3]
port 22 n
<< end >>
