magic
tech sky130B
magscale 1 2
timestamp 1736777579
<< nwell >>
rect -471 496 1306 814
rect 2673 496 4450 814
rect 5805 500 7582 818
rect 8949 500 10726 818
rect 12151 496 13928 814
rect 15295 496 17072 814
rect 18427 500 20204 818
rect 21571 500 23348 818
rect -484 95 -420 262
rect 2660 95 2724 262
rect 5792 99 5856 266
rect 8936 99 9000 266
rect -476 62 -420 95
rect 2668 62 2724 95
rect 5800 66 5856 99
rect 8944 66 9000 99
rect 12138 95 12202 262
rect 15282 95 15346 262
rect 18414 99 18478 266
rect 21558 99 21622 266
rect 12146 62 12202 95
rect 15290 62 15346 95
rect 18422 66 18478 99
rect 21566 66 21622 99
<< ndiff >>
rect 115 -1071 167 -871
rect 668 -960 735 -871
rect 667 -987 735 -960
rect 644 -1071 735 -987
rect 3259 -1071 3311 -871
rect 3812 -960 3879 -871
rect 3811 -987 3879 -960
rect 3788 -1071 3879 -987
rect 6391 -1067 6443 -867
rect 6944 -956 7011 -867
rect 6943 -983 7011 -956
rect 6920 -1067 7011 -983
rect 9535 -1067 9587 -867
rect 10088 -956 10155 -867
rect 10087 -983 10155 -956
rect 10064 -1067 10155 -983
rect 12737 -1071 12789 -871
rect 13290 -960 13357 -871
rect 13289 -987 13357 -960
rect 13266 -1071 13357 -987
rect 15881 -1071 15933 -871
rect 16434 -960 16501 -871
rect 16433 -987 16501 -960
rect 16410 -1071 16501 -987
rect 19013 -1067 19065 -867
rect 19566 -956 19633 -867
rect 19565 -983 19633 -956
rect 19542 -1067 19633 -983
rect 22157 -1067 22209 -867
rect 22710 -956 22777 -867
rect 22709 -983 22777 -956
rect 22686 -1067 22777 -983
<< pdiff >>
rect -484 95 -420 262
rect 2660 95 2724 262
rect 5792 99 5856 266
rect 8936 99 9000 266
rect -476 62 -420 95
rect 2668 62 2724 95
rect 5800 66 5856 99
rect 8944 66 9000 99
rect 12138 95 12202 262
rect 15282 95 15346 262
rect 18414 99 18478 266
rect 21558 99 21622 266
rect 12146 62 12202 95
rect 15290 62 15346 95
rect 18422 66 18478 99
rect 21566 66 21622 99
<< psubdiff >>
rect 338 -1526 524 -1502
rect 338 -1572 380 -1526
rect 484 -1572 524 -1526
rect 338 -1608 524 -1572
rect 3482 -1526 3668 -1502
rect 3482 -1572 3524 -1526
rect 3628 -1572 3668 -1526
rect 3482 -1608 3668 -1572
rect 6614 -1522 6800 -1498
rect 6614 -1568 6656 -1522
rect 6760 -1568 6800 -1522
rect 6614 -1604 6800 -1568
rect 9758 -1522 9944 -1498
rect 9758 -1568 9800 -1522
rect 9904 -1568 9944 -1522
rect 9758 -1604 9944 -1568
rect 12960 -1526 13146 -1502
rect 12960 -1572 13002 -1526
rect 13106 -1572 13146 -1526
rect 12960 -1608 13146 -1572
rect 16104 -1526 16290 -1502
rect 16104 -1572 16146 -1526
rect 16250 -1572 16290 -1526
rect 16104 -1608 16290 -1572
rect 19236 -1522 19422 -1498
rect 19236 -1568 19278 -1522
rect 19382 -1568 19422 -1522
rect 19236 -1604 19422 -1568
rect 22380 -1522 22566 -1498
rect 22380 -1568 22422 -1522
rect 22526 -1568 22566 -1522
rect 22380 -1604 22566 -1568
<< nsubdiff >>
rect 268 720 572 776
rect 268 644 322 720
rect 518 644 572 720
rect 268 630 572 644
rect 3412 720 3716 776
rect 3412 644 3466 720
rect 3662 644 3716 720
rect 3412 630 3716 644
rect 6544 724 6848 780
rect 6544 648 6598 724
rect 6794 648 6848 724
rect 6544 634 6848 648
rect 9688 724 9992 780
rect 9688 648 9742 724
rect 9938 648 9992 724
rect 9688 634 9992 648
rect 12890 720 13194 776
rect 12890 644 12944 720
rect 13140 644 13194 720
rect 12890 630 13194 644
rect 16034 720 16338 776
rect 16034 644 16088 720
rect 16284 644 16338 720
rect 16034 630 16338 644
rect 19166 724 19470 780
rect 19166 648 19220 724
rect 19416 648 19470 724
rect 19166 634 19470 648
rect 22310 724 22614 780
rect 22310 648 22364 724
rect 22560 648 22614 724
rect 22310 634 22614 648
<< psubdiffcont >>
rect 380 -1572 484 -1526
rect 3524 -1572 3628 -1526
rect 6656 -1568 6760 -1522
rect 9800 -1568 9904 -1522
rect 13002 -1572 13106 -1526
rect 16146 -1572 16250 -1526
rect 19278 -1568 19382 -1522
rect 22422 -1568 22526 -1522
<< nsubdiffcont >>
rect 322 644 518 720
rect 3466 644 3662 720
rect 6598 648 6794 724
rect 9742 648 9938 724
rect 12944 644 13140 720
rect 16088 644 16284 720
rect 19220 648 19416 724
rect 22364 648 22560 724
<< poly >>
rect -377 477 -81 516
rect 90 477 386 516
rect 444 477 740 516
rect 917 477 1213 516
rect 2767 477 3063 516
rect 3234 477 3530 516
rect 3588 477 3884 516
rect 4061 477 4357 516
rect 5899 481 6195 520
rect 6366 481 6662 520
rect 6720 481 7016 520
rect 7193 481 7489 520
rect 9043 481 9339 520
rect 9510 481 9806 520
rect 9864 481 10160 520
rect 10337 481 10633 520
rect 12245 477 12541 516
rect 12712 477 13008 516
rect 13066 477 13362 516
rect 13539 477 13835 516
rect 15389 477 15685 516
rect 15856 477 16152 516
rect 16210 477 16506 516
rect 16683 477 16979 516
rect 18521 481 18817 520
rect 18988 481 19284 520
rect 19342 481 19638 520
rect 19815 481 20111 520
rect 21665 481 21961 520
rect 22132 481 22428 520
rect 22486 481 22782 520
rect 22959 481 23255 520
rect -818 278 -522 317
rect 1390 278 1686 317
rect 2326 278 2622 317
rect 4534 278 4830 317
rect 5458 282 5754 321
rect 7666 282 7962 321
rect 8602 282 8898 321
rect 10810 282 11106 321
rect 11804 278 12100 317
rect 14012 278 14308 317
rect 14948 278 15244 317
rect 17156 278 17452 317
rect 18080 282 18376 321
rect 20288 282 20584 321
rect 21224 282 21520 321
rect 23432 282 23728 321
rect -818 -224 -758 59
rect -818 -241 -682 -224
rect -818 -296 -759 -241
rect -701 -296 -682 -241
rect -818 -311 -682 -296
rect -818 -623 -758 -311
rect -259 -356 -199 43
rect 209 -124 268 54
rect 209 -125 272 -124
rect 206 -141 272 -125
rect 206 -175 222 -141
rect 256 -175 272 -141
rect 206 -191 272 -175
rect 309 -240 404 -225
rect 309 -295 328 -240
rect 386 -263 404 -240
rect 562 -263 622 43
rect 386 -295 622 -263
rect 309 -312 622 -295
rect -259 -413 268 -356
rect 208 -512 268 -413
rect 197 -525 278 -512
rect 197 -580 210 -525
rect 268 -580 278 -525
rect 197 -591 278 -580
rect -818 -668 76 -623
rect 16 -857 76 -668
rect 208 -857 268 -591
rect 326 -857 386 -312
rect 1035 -354 1095 45
rect 1516 -87 1582 -84
rect 1626 -87 1686 59
rect 1516 -100 1686 -87
rect 1516 -134 1532 -100
rect 1566 -134 1686 -100
rect 1516 -147 1686 -134
rect 1516 -150 1582 -147
rect 557 -371 1095 -354
rect 557 -405 576 -371
rect 610 -405 1095 -371
rect 557 -411 1095 -405
rect 557 -421 626 -411
rect 557 -423 622 -421
rect 441 -761 507 -745
rect 441 -795 457 -761
rect 491 -795 507 -761
rect 441 -811 507 -795
rect 444 -855 504 -811
rect 562 -855 622 -423
rect 1626 -623 1686 -147
rect 758 -668 1686 -623
rect 2326 -224 2386 59
rect 2326 -241 2462 -224
rect 2326 -296 2385 -241
rect 2443 -296 2462 -241
rect 2326 -311 2462 -296
rect 2326 -623 2386 -311
rect 2885 -356 2945 43
rect 3353 -124 3412 54
rect 3353 -125 3416 -124
rect 3350 -141 3416 -125
rect 3350 -175 3366 -141
rect 3400 -175 3416 -141
rect 3350 -191 3416 -175
rect 3453 -240 3548 -225
rect 3453 -295 3472 -240
rect 3530 -263 3548 -240
rect 3706 -263 3766 43
rect 3530 -295 3766 -263
rect 3453 -312 3766 -295
rect 2885 -413 3412 -356
rect 3352 -512 3412 -413
rect 3341 -525 3422 -512
rect 3341 -580 3354 -525
rect 3412 -580 3422 -525
rect 3341 -591 3422 -580
rect 2326 -668 3220 -623
rect 758 -856 818 -668
rect 3160 -857 3220 -668
rect 3352 -857 3412 -591
rect 3470 -857 3530 -312
rect 4179 -354 4239 45
rect 4660 -87 4726 -84
rect 4770 -87 4830 59
rect 4660 -100 4830 -87
rect 4660 -134 4676 -100
rect 4710 -134 4830 -100
rect 4660 -147 4830 -134
rect 4660 -150 4726 -147
rect 3701 -371 4239 -354
rect 3701 -405 3720 -371
rect 3754 -405 4239 -371
rect 3701 -411 4239 -405
rect 3701 -421 3770 -411
rect 3701 -423 3766 -421
rect 3585 -761 3651 -745
rect 3585 -795 3601 -761
rect 3635 -795 3651 -761
rect 3585 -811 3651 -795
rect 3588 -855 3648 -811
rect 3706 -855 3766 -423
rect 4770 -623 4830 -147
rect 3902 -668 4830 -623
rect 5458 -220 5518 63
rect 5458 -237 5594 -220
rect 5458 -292 5517 -237
rect 5575 -292 5594 -237
rect 5458 -307 5594 -292
rect 5458 -619 5518 -307
rect 6017 -352 6077 47
rect 6485 -120 6544 58
rect 6485 -121 6548 -120
rect 6482 -137 6548 -121
rect 6482 -171 6498 -137
rect 6532 -171 6548 -137
rect 6482 -187 6548 -171
rect 6585 -236 6680 -221
rect 6585 -291 6604 -236
rect 6662 -259 6680 -236
rect 6838 -259 6898 47
rect 6662 -291 6898 -259
rect 6585 -308 6898 -291
rect 6017 -409 6544 -352
rect 6484 -508 6544 -409
rect 6473 -521 6554 -508
rect 6473 -576 6486 -521
rect 6544 -576 6554 -521
rect 6473 -587 6554 -576
rect 5458 -664 6352 -619
rect 3902 -856 3962 -668
rect 6292 -853 6352 -664
rect 6484 -853 6544 -587
rect 6602 -853 6662 -308
rect 7311 -350 7371 49
rect 7792 -83 7858 -80
rect 7902 -83 7962 63
rect 7792 -96 7962 -83
rect 7792 -130 7808 -96
rect 7842 -130 7962 -96
rect 7792 -143 7962 -130
rect 7792 -146 7858 -143
rect 6833 -367 7371 -350
rect 6833 -401 6852 -367
rect 6886 -401 7371 -367
rect 6833 -407 7371 -401
rect 6833 -417 6902 -407
rect 6833 -419 6898 -417
rect 6717 -757 6783 -741
rect 6717 -791 6733 -757
rect 6767 -791 6783 -757
rect 6717 -807 6783 -791
rect 6720 -851 6780 -807
rect 6838 -851 6898 -419
rect 7902 -619 7962 -143
rect 7034 -664 7962 -619
rect 8602 -220 8662 63
rect 8602 -237 8738 -220
rect 8602 -292 8661 -237
rect 8719 -292 8738 -237
rect 8602 -307 8738 -292
rect 8602 -619 8662 -307
rect 9161 -352 9221 47
rect 9629 -120 9688 58
rect 9629 -121 9692 -120
rect 9626 -137 9692 -121
rect 9626 -171 9642 -137
rect 9676 -171 9692 -137
rect 9626 -187 9692 -171
rect 9729 -236 9824 -221
rect 9729 -291 9748 -236
rect 9806 -259 9824 -236
rect 9982 -259 10042 47
rect 9806 -291 10042 -259
rect 9729 -308 10042 -291
rect 9161 -409 9688 -352
rect 9628 -508 9688 -409
rect 9617 -521 9698 -508
rect 9617 -576 9630 -521
rect 9688 -576 9698 -521
rect 9617 -587 9698 -576
rect 8602 -664 9496 -619
rect 7034 -852 7094 -664
rect 9436 -853 9496 -664
rect 9628 -853 9688 -587
rect 9746 -853 9806 -308
rect 10455 -350 10515 49
rect 10936 -83 11002 -80
rect 11046 -83 11106 63
rect 10936 -96 11106 -83
rect 10936 -130 10952 -96
rect 10986 -130 11106 -96
rect 10936 -143 11106 -130
rect 10936 -146 11002 -143
rect 9977 -367 10515 -350
rect 9977 -401 9996 -367
rect 10030 -401 10515 -367
rect 9977 -407 10515 -401
rect 9977 -417 10046 -407
rect 9977 -419 10042 -417
rect 9861 -757 9927 -741
rect 9861 -791 9877 -757
rect 9911 -791 9927 -757
rect 9861 -807 9927 -791
rect 9864 -851 9924 -807
rect 9982 -851 10042 -419
rect 11046 -619 11106 -143
rect 10178 -664 11106 -619
rect 11804 -224 11864 59
rect 11804 -241 11940 -224
rect 11804 -296 11863 -241
rect 11921 -296 11940 -241
rect 11804 -311 11940 -296
rect 11804 -623 11864 -311
rect 12363 -356 12423 43
rect 12831 -124 12890 54
rect 12831 -125 12894 -124
rect 12828 -141 12894 -125
rect 12828 -175 12844 -141
rect 12878 -175 12894 -141
rect 12828 -191 12894 -175
rect 12931 -240 13026 -225
rect 12931 -295 12950 -240
rect 13008 -263 13026 -240
rect 13184 -263 13244 43
rect 13008 -295 13244 -263
rect 12931 -312 13244 -295
rect 12363 -413 12890 -356
rect 12830 -512 12890 -413
rect 12819 -525 12900 -512
rect 12819 -580 12832 -525
rect 12890 -580 12900 -525
rect 12819 -591 12900 -580
rect 10178 -852 10238 -664
rect 11804 -668 12698 -623
rect 12638 -857 12698 -668
rect 12830 -857 12890 -591
rect 12948 -857 13008 -312
rect 13657 -354 13717 45
rect 14138 -87 14204 -84
rect 14248 -87 14308 59
rect 14138 -100 14308 -87
rect 14138 -134 14154 -100
rect 14188 -134 14308 -100
rect 14138 -147 14308 -134
rect 14138 -150 14204 -147
rect 13179 -371 13717 -354
rect 13179 -405 13198 -371
rect 13232 -405 13717 -371
rect 13179 -411 13717 -405
rect 13179 -421 13248 -411
rect 13179 -423 13244 -421
rect 13063 -761 13129 -745
rect 13063 -795 13079 -761
rect 13113 -795 13129 -761
rect 13063 -811 13129 -795
rect 13066 -855 13126 -811
rect 13184 -855 13244 -423
rect 14248 -623 14308 -147
rect 13380 -668 14308 -623
rect 14948 -224 15008 59
rect 14948 -241 15084 -224
rect 14948 -296 15007 -241
rect 15065 -296 15084 -241
rect 14948 -311 15084 -296
rect 14948 -623 15008 -311
rect 15507 -356 15567 43
rect 15975 -124 16034 54
rect 15975 -125 16038 -124
rect 15972 -141 16038 -125
rect 15972 -175 15988 -141
rect 16022 -175 16038 -141
rect 15972 -191 16038 -175
rect 16075 -240 16170 -225
rect 16075 -295 16094 -240
rect 16152 -263 16170 -240
rect 16328 -263 16388 43
rect 16152 -295 16388 -263
rect 16075 -312 16388 -295
rect 15507 -413 16034 -356
rect 15974 -512 16034 -413
rect 15963 -525 16044 -512
rect 15963 -580 15976 -525
rect 16034 -580 16044 -525
rect 15963 -591 16044 -580
rect 14948 -668 15842 -623
rect 13380 -856 13440 -668
rect 15782 -857 15842 -668
rect 15974 -857 16034 -591
rect 16092 -857 16152 -312
rect 16801 -354 16861 45
rect 17282 -87 17348 -84
rect 17392 -87 17452 59
rect 17282 -100 17452 -87
rect 17282 -134 17298 -100
rect 17332 -134 17452 -100
rect 17282 -147 17452 -134
rect 17282 -150 17348 -147
rect 16323 -371 16861 -354
rect 16323 -405 16342 -371
rect 16376 -405 16861 -371
rect 16323 -411 16861 -405
rect 16323 -421 16392 -411
rect 16323 -423 16388 -421
rect 16207 -761 16273 -745
rect 16207 -795 16223 -761
rect 16257 -795 16273 -761
rect 16207 -811 16273 -795
rect 16210 -855 16270 -811
rect 16328 -855 16388 -423
rect 17392 -623 17452 -147
rect 16524 -668 17452 -623
rect 18080 -220 18140 63
rect 18080 -237 18216 -220
rect 18080 -292 18139 -237
rect 18197 -292 18216 -237
rect 18080 -307 18216 -292
rect 18080 -619 18140 -307
rect 18639 -352 18699 47
rect 19107 -120 19166 58
rect 19107 -121 19170 -120
rect 19104 -137 19170 -121
rect 19104 -171 19120 -137
rect 19154 -171 19170 -137
rect 19104 -187 19170 -171
rect 19207 -236 19302 -221
rect 19207 -291 19226 -236
rect 19284 -259 19302 -236
rect 19460 -259 19520 47
rect 19284 -291 19520 -259
rect 19207 -308 19520 -291
rect 18639 -409 19166 -352
rect 19106 -508 19166 -409
rect 19095 -521 19176 -508
rect 19095 -576 19108 -521
rect 19166 -576 19176 -521
rect 19095 -587 19176 -576
rect 18080 -664 18974 -619
rect 16524 -856 16584 -668
rect 18914 -853 18974 -664
rect 19106 -853 19166 -587
rect 19224 -853 19284 -308
rect 19933 -350 19993 49
rect 20414 -83 20480 -80
rect 20524 -83 20584 63
rect 20414 -96 20584 -83
rect 20414 -130 20430 -96
rect 20464 -130 20584 -96
rect 20414 -143 20584 -130
rect 20414 -146 20480 -143
rect 19455 -367 19993 -350
rect 19455 -401 19474 -367
rect 19508 -401 19993 -367
rect 19455 -407 19993 -401
rect 19455 -417 19524 -407
rect 19455 -419 19520 -417
rect 19339 -757 19405 -741
rect 19339 -791 19355 -757
rect 19389 -791 19405 -757
rect 19339 -807 19405 -791
rect 19342 -851 19402 -807
rect 19460 -851 19520 -419
rect 20524 -619 20584 -143
rect 19656 -664 20584 -619
rect 21224 -220 21284 63
rect 21224 -237 21360 -220
rect 21224 -292 21283 -237
rect 21341 -292 21360 -237
rect 21224 -307 21360 -292
rect 21224 -619 21284 -307
rect 21783 -352 21843 47
rect 22251 -120 22310 58
rect 22251 -121 22314 -120
rect 22248 -137 22314 -121
rect 22248 -171 22264 -137
rect 22298 -171 22314 -137
rect 22248 -187 22314 -171
rect 22351 -236 22446 -221
rect 22351 -291 22370 -236
rect 22428 -259 22446 -236
rect 22604 -259 22664 47
rect 22428 -291 22664 -259
rect 22351 -308 22664 -291
rect 21783 -409 22310 -352
rect 22250 -508 22310 -409
rect 22239 -521 22320 -508
rect 22239 -576 22252 -521
rect 22310 -576 22320 -521
rect 22239 -587 22320 -576
rect 21224 -664 22118 -619
rect 19656 -852 19716 -664
rect 22058 -853 22118 -664
rect 22250 -853 22310 -587
rect 22368 -853 22428 -308
rect 23077 -350 23137 49
rect 23558 -83 23624 -80
rect 23668 -83 23728 63
rect 23558 -96 23728 -83
rect 23558 -130 23574 -96
rect 23608 -130 23728 -96
rect 23558 -143 23728 -130
rect 23558 -146 23624 -143
rect 22599 -367 23137 -350
rect 22599 -401 22618 -367
rect 22652 -401 23137 -367
rect 22599 -407 23137 -401
rect 22599 -417 22668 -407
rect 22599 -419 22664 -417
rect 22483 -757 22549 -741
rect 22483 -791 22499 -757
rect 22533 -791 22549 -757
rect 22483 -807 22549 -791
rect 22486 -851 22546 -807
rect 22604 -851 22664 -419
rect 23668 -619 23728 -143
rect 22800 -664 23728 -619
rect 22800 -852 22860 -664
rect 383 -1352 449 -1344
rect 758 -1352 818 -1083
rect 383 -1360 818 -1352
rect 383 -1394 399 -1360
rect 433 -1394 818 -1360
rect 383 -1403 818 -1394
rect 3527 -1352 3593 -1344
rect 3902 -1352 3962 -1083
rect 3527 -1360 3962 -1352
rect 3527 -1394 3543 -1360
rect 3577 -1394 3962 -1360
rect 3527 -1403 3962 -1394
rect 6659 -1348 6725 -1340
rect 7034 -1348 7094 -1079
rect 6659 -1356 7094 -1348
rect 6659 -1390 6675 -1356
rect 6709 -1390 7094 -1356
rect 6659 -1399 7094 -1390
rect 9803 -1348 9869 -1340
rect 10178 -1348 10238 -1079
rect 9803 -1356 10238 -1348
rect 9803 -1390 9819 -1356
rect 9853 -1390 10238 -1356
rect 9803 -1399 10238 -1390
rect 13005 -1352 13071 -1344
rect 13380 -1352 13440 -1083
rect 13005 -1360 13440 -1352
rect 13005 -1394 13021 -1360
rect 13055 -1394 13440 -1360
rect 383 -1410 449 -1403
rect 3527 -1410 3593 -1403
rect 6659 -1406 6725 -1399
rect 9803 -1406 9869 -1399
rect 13005 -1403 13440 -1394
rect 16149 -1352 16215 -1344
rect 16524 -1352 16584 -1083
rect 16149 -1360 16584 -1352
rect 16149 -1394 16165 -1360
rect 16199 -1394 16584 -1360
rect 16149 -1403 16584 -1394
rect 19281 -1348 19347 -1340
rect 19656 -1348 19716 -1079
rect 19281 -1356 19716 -1348
rect 19281 -1390 19297 -1356
rect 19331 -1390 19716 -1356
rect 19281 -1399 19716 -1390
rect 22425 -1348 22491 -1340
rect 22800 -1348 22860 -1079
rect 22425 -1356 22860 -1348
rect 22425 -1390 22441 -1356
rect 22475 -1390 22860 -1356
rect 22425 -1399 22860 -1390
rect 13005 -1410 13071 -1403
rect 16149 -1410 16215 -1403
rect 19281 -1406 19347 -1399
rect 22425 -1406 22491 -1399
<< polycont >>
rect -759 -296 -701 -241
rect 222 -175 256 -141
rect 328 -295 386 -240
rect 210 -580 268 -525
rect 1532 -134 1566 -100
rect 576 -405 610 -371
rect 457 -795 491 -761
rect 2385 -296 2443 -241
rect 3366 -175 3400 -141
rect 3472 -295 3530 -240
rect 3354 -580 3412 -525
rect 4676 -134 4710 -100
rect 3720 -405 3754 -371
rect 3601 -795 3635 -761
rect 5517 -292 5575 -237
rect 6498 -171 6532 -137
rect 6604 -291 6662 -236
rect 6486 -576 6544 -521
rect 7808 -130 7842 -96
rect 6852 -401 6886 -367
rect 6733 -791 6767 -757
rect 8661 -292 8719 -237
rect 9642 -171 9676 -137
rect 9748 -291 9806 -236
rect 9630 -576 9688 -521
rect 10952 -130 10986 -96
rect 9996 -401 10030 -367
rect 9877 -791 9911 -757
rect 11863 -296 11921 -241
rect 12844 -175 12878 -141
rect 12950 -295 13008 -240
rect 12832 -580 12890 -525
rect 14154 -134 14188 -100
rect 13198 -405 13232 -371
rect 13079 -795 13113 -761
rect 15007 -296 15065 -241
rect 15988 -175 16022 -141
rect 16094 -295 16152 -240
rect 15976 -580 16034 -525
rect 17298 -134 17332 -100
rect 16342 -405 16376 -371
rect 16223 -795 16257 -761
rect 18139 -292 18197 -237
rect 19120 -171 19154 -137
rect 19226 -291 19284 -236
rect 19108 -576 19166 -521
rect 20430 -130 20464 -96
rect 19474 -401 19508 -367
rect 19355 -791 19389 -757
rect 21283 -292 21341 -237
rect 22264 -171 22298 -137
rect 22370 -291 22428 -236
rect 22252 -576 22310 -521
rect 23574 -130 23608 -96
rect 22618 -401 22652 -367
rect 22499 -791 22533 -757
rect 399 -1394 433 -1360
rect 3543 -1394 3577 -1360
rect 6675 -1390 6709 -1356
rect 9819 -1390 9853 -1356
rect 13021 -1394 13055 -1360
rect 16165 -1394 16199 -1360
rect 19297 -1390 19331 -1356
rect 22441 -1390 22475 -1356
<< locali >>
rect 306 720 534 738
rect 306 644 322 720
rect 518 644 534 720
rect 306 628 534 644
rect 3450 720 3678 738
rect 3450 644 3466 720
rect 3662 644 3678 720
rect 3450 628 3678 644
rect 6582 724 6810 742
rect 6582 648 6598 724
rect 6794 648 6810 724
rect 6582 632 6810 648
rect 9726 724 9954 742
rect 9726 648 9742 724
rect 9938 648 9954 724
rect 9726 632 9954 648
rect 12928 720 13156 738
rect 12928 644 12944 720
rect 13140 644 13156 720
rect 12928 628 13156 644
rect 16072 720 16300 738
rect 16072 644 16088 720
rect 16284 644 16300 720
rect 16072 628 16300 644
rect 19204 724 19432 742
rect 19204 648 19220 724
rect 19416 648 19432 724
rect 19204 632 19432 648
rect 22348 724 22576 742
rect 22348 648 22364 724
rect 22560 648 22576 724
rect 22348 632 22576 648
rect -423 503 -153 542
rect -423 431 -389 503
rect -187 431 -153 503
rect 44 502 314 541
rect 44 430 78 502
rect 280 430 314 502
rect 516 502 786 541
rect 516 430 550 502
rect 752 430 786 502
rect 989 502 1259 541
rect 989 430 1023 502
rect 1225 430 1259 502
rect 2721 503 2991 542
rect 2721 431 2755 503
rect 2957 431 2991 503
rect 3188 502 3458 541
rect 3188 430 3222 502
rect 3424 430 3458 502
rect 3660 502 3930 541
rect 3660 430 3694 502
rect 3896 430 3930 502
rect 4133 502 4403 541
rect 4133 430 4167 502
rect 4369 430 4403 502
rect 5853 507 6123 546
rect 5853 435 5887 507
rect 6089 435 6123 507
rect 6320 506 6590 545
rect 6320 434 6354 506
rect 6556 434 6590 506
rect 6792 506 7062 545
rect 6792 434 6826 506
rect 7028 434 7062 506
rect 7265 506 7535 545
rect 7265 434 7299 506
rect 7501 434 7535 506
rect 8997 507 9267 546
rect 8997 435 9031 507
rect 9233 435 9267 507
rect 9464 506 9734 545
rect 9464 434 9498 506
rect 9700 434 9734 506
rect 9936 506 10206 545
rect 9936 434 9970 506
rect 10172 434 10206 506
rect 10409 506 10679 545
rect 10409 434 10443 506
rect 10645 434 10679 506
rect 12199 503 12469 542
rect 12199 431 12233 503
rect 12435 431 12469 503
rect 12666 502 12936 541
rect 12666 430 12700 502
rect 12902 430 12936 502
rect 13138 502 13408 541
rect 13138 430 13172 502
rect 13374 430 13408 502
rect 13611 502 13881 541
rect 13611 430 13645 502
rect 13847 430 13881 502
rect 15343 503 15613 542
rect 15343 431 15377 503
rect 15579 431 15613 503
rect 15810 502 16080 541
rect 15810 430 15844 502
rect 16046 430 16080 502
rect 16282 502 16552 541
rect 16282 430 16316 502
rect 16518 430 16552 502
rect 16755 502 17025 541
rect 16755 430 16789 502
rect 16991 430 17025 502
rect 18475 507 18745 546
rect 18475 435 18509 507
rect 18711 435 18745 507
rect 18942 506 19212 545
rect 18942 434 18976 506
rect 19178 434 19212 506
rect 19414 506 19684 545
rect 19414 434 19448 506
rect 19650 434 19684 506
rect 19887 506 20157 545
rect 19887 434 19921 506
rect 20123 434 20157 506
rect 21619 507 21889 546
rect 21619 435 21653 507
rect 21855 435 21889 507
rect 22086 506 22356 545
rect 22086 434 22120 506
rect 22322 434 22356 506
rect 22558 506 22828 545
rect 22558 434 22592 506
rect 22794 434 22828 506
rect 23031 506 23301 545
rect 23031 434 23065 506
rect 23267 434 23301 506
rect -864 301 -594 340
rect -864 222 -830 301
rect -628 229 -594 301
rect 1462 300 1732 337
rect 1462 226 1496 300
rect 1698 226 1732 300
rect 2280 301 2550 340
rect 2280 222 2314 301
rect 2516 229 2550 301
rect 4606 300 4876 337
rect 4606 226 4640 300
rect 4842 226 4876 300
rect 5412 305 5682 344
rect 5412 226 5446 305
rect 5648 233 5682 305
rect 7738 304 8008 341
rect 7738 230 7772 304
rect 7974 230 8008 304
rect 8556 305 8826 344
rect 8556 226 8590 305
rect 8792 233 8826 305
rect 10882 304 11152 341
rect 10882 230 10916 304
rect 11118 230 11152 304
rect 11758 301 12028 340
rect 11758 222 11792 301
rect 11994 229 12028 301
rect 14084 300 14354 337
rect 14084 226 14118 300
rect 14320 226 14354 300
rect 14902 301 15172 340
rect 14902 222 14936 301
rect 15138 229 15172 301
rect 17228 300 17498 337
rect 17228 226 17262 300
rect 17464 226 17498 300
rect 18034 305 18304 344
rect 18034 226 18068 305
rect 18270 233 18304 305
rect 20360 304 20630 341
rect 20360 230 20394 304
rect 20596 230 20630 304
rect 21178 305 21448 344
rect 21178 226 21212 305
rect 21414 233 21448 305
rect 23504 304 23774 341
rect 23504 230 23538 304
rect 23740 230 23774 304
rect -746 23 -712 95
rect -510 23 -476 95
rect -746 -16 -476 23
rect -305 23 -271 95
rect -69 23 -35 95
rect 162 23 196 95
rect 398 23 432 95
rect 634 23 668 95
rect 871 23 905 95
rect 1107 23 1141 95
rect -305 -16 1141 23
rect 1344 20 1378 80
rect 1580 20 1614 92
rect 1344 -19 1614 20
rect 2398 23 2432 95
rect 2634 23 2668 95
rect 2398 -16 2668 23
rect 2839 23 2873 95
rect 3075 23 3109 95
rect 3306 23 3340 95
rect 3542 23 3576 95
rect 3778 23 3812 95
rect 4015 23 4049 95
rect 4251 23 4285 95
rect 2839 -16 4285 23
rect 4488 20 4522 80
rect 4724 20 4758 92
rect 4488 -19 4758 20
rect 5530 27 5564 99
rect 5766 27 5800 99
rect 5530 -12 5800 27
rect 5971 27 6005 99
rect 6207 27 6241 99
rect 6438 27 6472 99
rect 6674 27 6708 99
rect 6910 27 6944 99
rect 7147 27 7181 99
rect 7383 27 7417 99
rect 5971 -12 7417 27
rect 7620 24 7654 84
rect 7856 24 7890 96
rect 7620 -15 7890 24
rect 8674 27 8708 99
rect 8910 27 8944 99
rect 8674 -12 8944 27
rect 9115 27 9149 99
rect 9351 27 9385 99
rect 9582 27 9616 99
rect 9818 27 9852 99
rect 10054 27 10088 99
rect 10291 27 10325 99
rect 10527 27 10561 99
rect 9115 -12 10561 27
rect 10764 24 10798 84
rect 11000 24 11034 96
rect 10764 -15 11034 24
rect 11876 23 11910 95
rect 12112 23 12146 95
rect 11876 -16 12146 23
rect 12317 23 12351 95
rect 12553 23 12587 95
rect 12784 23 12818 95
rect 13020 23 13054 95
rect 13256 23 13290 95
rect 13493 23 13527 95
rect 13729 23 13763 95
rect 12317 -16 13763 23
rect 13966 20 14000 80
rect 14202 20 14236 92
rect 13966 -19 14236 20
rect 15020 23 15054 95
rect 15256 23 15290 95
rect 15020 -16 15290 23
rect 15461 23 15495 95
rect 15697 23 15731 95
rect 15928 23 15962 95
rect 16164 23 16198 95
rect 16400 23 16434 95
rect 16637 23 16671 95
rect 16873 23 16907 95
rect 15461 -16 16907 23
rect 17110 20 17144 80
rect 17346 20 17380 92
rect 17110 -19 17380 20
rect 18152 27 18186 99
rect 18388 27 18422 99
rect 18152 -12 18422 27
rect 18593 27 18627 99
rect 18829 27 18863 99
rect 19060 27 19094 99
rect 19296 27 19330 99
rect 19532 27 19566 99
rect 19769 27 19803 99
rect 20005 27 20039 99
rect 18593 -12 20039 27
rect 20242 24 20276 84
rect 20478 24 20512 96
rect 20242 -15 20512 24
rect 21296 27 21330 99
rect 21532 27 21566 99
rect 21296 -12 21566 27
rect 21737 27 21771 99
rect 21973 27 22007 99
rect 22204 27 22238 99
rect 22440 27 22474 99
rect 22676 27 22710 99
rect 22913 27 22947 99
rect 23149 27 23183 99
rect 21737 -12 23183 27
rect 23386 24 23420 84
rect 23622 24 23656 96
rect 23386 -15 23656 24
rect 222 -141 256 -125
rect 1516 -134 1532 -100
rect 1566 -134 1582 -100
rect 222 -191 256 -175
rect 3366 -141 3400 -125
rect 4660 -134 4676 -100
rect 4710 -134 4726 -100
rect 3366 -191 3400 -175
rect 6498 -137 6532 -121
rect 7792 -130 7808 -96
rect 7842 -130 7858 -96
rect 6498 -187 6532 -171
rect 9642 -137 9676 -121
rect 10936 -130 10952 -96
rect 10986 -130 11002 -96
rect 9642 -187 9676 -171
rect 12844 -141 12878 -125
rect 14138 -134 14154 -100
rect 14188 -134 14204 -100
rect 12844 -191 12878 -175
rect 15988 -141 16022 -125
rect 17282 -134 17298 -100
rect 17332 -134 17348 -100
rect 15988 -191 16022 -175
rect 19120 -137 19154 -121
rect 20414 -130 20430 -96
rect 20464 -130 20480 -96
rect 19120 -187 19154 -171
rect 22264 -137 22298 -121
rect 23558 -130 23574 -96
rect 23608 -130 23624 -96
rect 22264 -187 22298 -171
rect -1007 -240 -950 -236
rect -1007 -300 -1003 -240
rect -954 -300 -950 -240
rect -1007 -304 -950 -300
rect -775 -241 -683 -224
rect -775 -296 -759 -241
rect -699 -296 -683 -241
rect -775 -309 -683 -296
rect 310 -240 402 -227
rect 310 -295 326 -240
rect 386 -295 402 -240
rect 310 -312 402 -295
rect 2369 -241 2461 -224
rect 2369 -296 2385 -241
rect 2445 -296 2461 -241
rect 2369 -309 2461 -296
rect 3454 -240 3546 -227
rect 3454 -295 3470 -240
rect 3530 -295 3546 -240
rect 3454 -312 3546 -295
rect 5501 -237 5593 -220
rect 5501 -292 5517 -237
rect 5577 -292 5593 -237
rect 5501 -305 5593 -292
rect 6586 -236 6678 -223
rect 6586 -291 6602 -236
rect 6662 -291 6678 -236
rect 6586 -308 6678 -291
rect 8645 -237 8737 -220
rect 8645 -292 8661 -237
rect 8721 -292 8737 -237
rect 8645 -305 8737 -292
rect 9730 -236 9822 -223
rect 9730 -291 9746 -236
rect 9806 -291 9822 -236
rect 9730 -308 9822 -291
rect 11847 -241 11939 -224
rect 11847 -296 11863 -241
rect 11923 -296 11939 -241
rect 11847 -309 11939 -296
rect 12932 -240 13024 -227
rect 12932 -295 12948 -240
rect 13008 -295 13024 -240
rect 12932 -312 13024 -295
rect 14991 -241 15083 -224
rect 14991 -296 15007 -241
rect 15067 -296 15083 -241
rect 14991 -309 15083 -296
rect 16076 -240 16168 -227
rect 16076 -295 16092 -240
rect 16152 -295 16168 -240
rect 16076 -312 16168 -295
rect 18123 -237 18215 -220
rect 18123 -292 18139 -237
rect 18199 -292 18215 -237
rect 18123 -305 18215 -292
rect 19208 -236 19300 -223
rect 19208 -291 19224 -236
rect 19284 -291 19300 -236
rect 19208 -308 19300 -291
rect 21267 -237 21359 -220
rect 21267 -292 21283 -237
rect 21343 -292 21359 -237
rect 21267 -305 21359 -292
rect 22352 -236 22444 -223
rect 22352 -291 22368 -236
rect 22428 -291 22444 -236
rect 22352 -308 22444 -291
rect 576 -371 610 -355
rect 576 -421 610 -405
rect 2137 -356 2194 -352
rect 2137 -416 2141 -356
rect 2190 -416 2194 -356
rect 2137 -420 2194 -416
rect 3720 -371 3754 -355
rect 3720 -421 3754 -405
rect 6852 -367 6886 -351
rect 6852 -417 6886 -401
rect 8287 -352 8482 -348
rect 8287 -412 8417 -352
rect 8466 -412 8482 -352
rect 8287 -420 8482 -412
rect 9996 -367 10030 -351
rect 14538 -352 14792 -351
rect 17891 -352 17948 -348
rect 9996 -417 10030 -401
rect 13198 -371 13232 -355
rect 8287 -423 8345 -420
rect 13198 -421 13232 -405
rect 14538 -356 14816 -352
rect 14538 -416 14763 -356
rect 14812 -416 14816 -356
rect 14538 -420 14816 -416
rect 16342 -371 16376 -355
rect 8114 -480 8345 -423
rect -1007 -524 -950 -520
rect -1007 -584 -1003 -524
rect -954 -584 -950 -524
rect -1007 -588 -950 -584
rect 192 -525 284 -512
rect 192 -580 208 -525
rect 268 -580 284 -525
rect 192 -597 284 -580
rect 2137 -524 2194 -520
rect 2137 -584 2141 -524
rect 2190 -584 2194 -524
rect 2137 -588 2194 -584
rect 3336 -525 4743 -512
rect 3336 -580 3352 -525
rect 3412 -580 4743 -525
rect 3336 -597 4743 -580
rect 5269 -520 5326 -516
rect 5269 -580 5273 -520
rect 5322 -580 5326 -520
rect 5269 -584 5326 -580
rect 6468 -521 6560 -508
rect 6468 -576 6484 -521
rect 6544 -576 6560 -521
rect 6468 -593 6560 -576
rect 4663 -654 4743 -597
rect 8114 -654 8191 -480
rect 8413 -520 8470 -516
rect 8413 -580 8417 -520
rect 8466 -580 8470 -520
rect 8413 -584 8470 -580
rect 9612 -521 10484 -508
rect 9612 -576 9628 -521
rect 9688 -576 10484 -521
rect 9612 -593 10484 -576
rect 11615 -524 11672 -520
rect 11615 -584 11619 -524
rect 11668 -584 11672 -524
rect 11615 -588 11672 -584
rect 12814 -525 12906 -512
rect 12814 -580 12830 -525
rect 12890 -580 12906 -525
rect 4663 -707 8191 -654
rect 10407 -648 10484 -593
rect 12814 -597 12906 -580
rect 14538 -648 14606 -420
rect 16342 -421 16376 -405
rect 17891 -412 17895 -352
rect 17944 -412 17948 -352
rect 17891 -416 17948 -412
rect 19474 -367 19508 -351
rect 19474 -417 19508 -401
rect 20841 -352 21092 -348
rect 20841 -412 21039 -352
rect 21088 -412 21092 -352
rect 20841 -416 21092 -412
rect 22618 -367 22652 -351
rect 14759 -524 14816 -520
rect 14759 -584 14763 -524
rect 14812 -584 14816 -524
rect 14759 -588 14816 -584
rect 15958 -525 16895 -512
rect 15958 -580 15974 -525
rect 16034 -580 16895 -525
rect 15958 -597 16895 -580
rect 17891 -520 17948 -516
rect 17891 -580 17895 -520
rect 17944 -580 17948 -520
rect 17891 -584 17948 -580
rect 19090 -521 19182 -508
rect 19090 -576 19106 -521
rect 19166 -576 19182 -521
rect 19090 -593 19182 -576
rect 10407 -710 14606 -648
rect 16820 -642 16895 -597
rect 20841 -642 20898 -416
rect 22618 -417 22652 -401
rect 22234 -521 22326 -508
rect 22234 -576 22250 -521
rect 22310 -576 22326 -521
rect 22234 -593 22326 -576
rect 16820 -707 20898 -642
rect 457 -761 491 -745
rect 457 -811 491 -795
rect 3601 -761 3635 -745
rect 3601 -811 3635 -795
rect 6733 -757 6767 -741
rect 6733 -807 6767 -791
rect 9877 -757 9911 -741
rect 9877 -807 9911 -791
rect 13079 -761 13113 -745
rect 13079 -811 13113 -795
rect 16223 -761 16257 -745
rect 16223 -811 16257 -795
rect 19355 -757 19389 -741
rect 19355 -807 19389 -791
rect 22499 -757 22533 -741
rect 22499 -807 22533 -791
rect 115 -1071 167 -871
rect 668 -960 735 -871
rect 667 -987 735 -960
rect 644 -1071 735 -987
rect 3259 -1071 3311 -871
rect 3812 -960 3879 -871
rect 3811 -987 3879 -960
rect 3788 -1071 3879 -987
rect 6391 -1067 6443 -867
rect 6944 -956 7011 -867
rect 6943 -983 7011 -956
rect 6920 -1067 7011 -983
rect 9535 -1067 9587 -867
rect 10088 -956 10155 -867
rect 10087 -983 10155 -956
rect 10064 -1067 10155 -983
rect 12737 -1071 12789 -871
rect 13290 -960 13357 -871
rect 13289 -987 13357 -960
rect 13266 -1071 13357 -987
rect 15881 -1071 15933 -871
rect 16434 -960 16501 -871
rect 16433 -987 16501 -960
rect 16410 -1071 16501 -987
rect 19013 -1067 19065 -867
rect 19566 -956 19633 -867
rect 19565 -983 19633 -956
rect 19542 -1067 19633 -983
rect 22157 -1067 22209 -867
rect 22710 -956 22777 -867
rect 22709 -983 22777 -956
rect 22686 -1067 22777 -983
rect 383 -1394 399 -1360
rect 433 -1394 449 -1360
rect 3527 -1394 3543 -1360
rect 3577 -1394 3593 -1360
rect 6659 -1390 6675 -1356
rect 6709 -1390 6725 -1356
rect 9803 -1390 9819 -1356
rect 9853 -1390 9869 -1356
rect 13005 -1394 13021 -1360
rect 13055 -1394 13071 -1360
rect 16149 -1394 16165 -1360
rect 16199 -1394 16215 -1360
rect 19281 -1390 19297 -1356
rect 19331 -1390 19347 -1356
rect 22425 -1390 22441 -1356
rect 22475 -1390 22491 -1356
rect 6640 -1508 6776 -1504
rect 364 -1512 500 -1508
rect 364 -1526 402 -1512
rect 460 -1526 500 -1512
rect 364 -1572 380 -1526
rect 484 -1572 500 -1526
rect 364 -1594 500 -1572
rect 3508 -1512 3644 -1508
rect 3508 -1526 3546 -1512
rect 3604 -1526 3644 -1512
rect 3508 -1572 3524 -1526
rect 3628 -1572 3644 -1526
rect 3508 -1594 3644 -1572
rect 6640 -1522 6678 -1508
rect 6736 -1522 6776 -1508
rect 6640 -1568 6656 -1522
rect 6760 -1568 6776 -1522
rect 6640 -1590 6776 -1568
rect 9784 -1508 9920 -1504
rect 19262 -1508 19398 -1504
rect 9784 -1522 9822 -1508
rect 9880 -1522 9920 -1508
rect 9784 -1568 9800 -1522
rect 9904 -1568 9920 -1522
rect 9784 -1590 9920 -1568
rect 12986 -1512 13122 -1508
rect 12986 -1526 13024 -1512
rect 13082 -1526 13122 -1512
rect 12986 -1572 13002 -1526
rect 13106 -1572 13122 -1526
rect 12986 -1594 13122 -1572
rect 16130 -1512 16266 -1508
rect 16130 -1526 16168 -1512
rect 16226 -1526 16266 -1512
rect 16130 -1572 16146 -1526
rect 16250 -1572 16266 -1526
rect 16130 -1594 16266 -1572
rect 19262 -1522 19300 -1508
rect 19358 -1522 19398 -1508
rect 19262 -1568 19278 -1522
rect 19382 -1568 19398 -1522
rect 19262 -1590 19398 -1568
rect 22406 -1508 22542 -1504
rect 22406 -1522 22444 -1508
rect 22502 -1522 22542 -1508
rect 22406 -1568 22422 -1522
rect 22526 -1568 22542 -1522
rect 22406 -1590 22542 -1568
<< viali >>
rect 388 646 460 700
rect 3532 646 3604 700
rect 6664 650 6736 704
rect 9808 650 9880 704
rect 13010 646 13082 700
rect 16154 646 16226 700
rect 19286 650 19358 704
rect 22430 650 22502 704
rect 1532 -134 1566 -100
rect 222 -175 256 -141
rect 4676 -134 4710 -100
rect 3366 -175 3400 -141
rect 7808 -130 7842 -96
rect 6498 -171 6532 -137
rect 10952 -130 10986 -96
rect 9642 -171 9676 -137
rect 14154 -134 14188 -100
rect 12844 -175 12878 -141
rect 17298 -134 17332 -100
rect 15988 -175 16022 -141
rect 20430 -130 20464 -96
rect 19120 -171 19154 -137
rect 23574 -130 23608 -96
rect 22264 -171 22298 -137
rect -1003 -300 -954 -240
rect -759 -296 -701 -241
rect -701 -296 -699 -241
rect 326 -295 328 -240
rect 328 -295 386 -240
rect 2385 -296 2443 -241
rect 2443 -296 2445 -241
rect 3470 -295 3472 -240
rect 3472 -295 3530 -240
rect 5517 -292 5575 -237
rect 5575 -292 5577 -237
rect 6602 -291 6604 -236
rect 6604 -291 6662 -236
rect 8661 -292 8719 -237
rect 8719 -292 8721 -237
rect 9746 -291 9748 -236
rect 9748 -291 9806 -236
rect 11863 -296 11921 -241
rect 11921 -296 11923 -241
rect 12948 -295 12950 -240
rect 12950 -295 13008 -240
rect 15007 -296 15065 -241
rect 15065 -296 15067 -241
rect 16092 -295 16094 -240
rect 16094 -295 16152 -240
rect 18139 -292 18197 -237
rect 18197 -292 18199 -237
rect 19224 -291 19226 -236
rect 19226 -291 19284 -236
rect 21283 -292 21341 -237
rect 21341 -292 21343 -237
rect 22368 -291 22370 -236
rect 22370 -291 22428 -236
rect 576 -405 610 -371
rect 2141 -416 2190 -356
rect 3720 -405 3754 -371
rect 6852 -401 6886 -367
rect 8417 -412 8466 -352
rect 9996 -401 10030 -367
rect 13198 -405 13232 -371
rect 14763 -416 14812 -356
rect 16342 -405 16376 -371
rect -1003 -584 -954 -524
rect 208 -580 210 -525
rect 210 -580 268 -525
rect 2141 -584 2190 -524
rect 3352 -580 3354 -525
rect 3354 -580 3412 -525
rect 5273 -580 5322 -520
rect 6484 -576 6486 -521
rect 6486 -576 6544 -521
rect 8417 -580 8466 -520
rect 9628 -576 9630 -521
rect 9630 -576 9688 -521
rect 11619 -584 11668 -524
rect 12830 -580 12832 -525
rect 12832 -580 12890 -525
rect 17895 -412 17944 -352
rect 19474 -401 19508 -367
rect 21039 -412 21088 -352
rect 22618 -401 22652 -367
rect 14763 -584 14812 -524
rect 15974 -580 15976 -525
rect 15976 -580 16034 -525
rect 17895 -580 17944 -520
rect 19106 -576 19108 -521
rect 19108 -576 19166 -521
rect 22250 -576 22252 -521
rect 22252 -576 22310 -521
rect 457 -795 491 -761
rect 3601 -795 3635 -761
rect 6733 -791 6767 -757
rect 9877 -791 9911 -757
rect 13079 -795 13113 -761
rect 16223 -795 16257 -761
rect 19355 -791 19389 -757
rect 22499 -791 22533 -757
rect 399 -1394 433 -1360
rect 3543 -1394 3577 -1360
rect 6675 -1390 6709 -1356
rect 9819 -1390 9853 -1356
rect 13021 -1394 13055 -1360
rect 16165 -1394 16199 -1360
rect 19297 -1390 19331 -1356
rect 22441 -1390 22475 -1356
rect 402 -1526 460 -1512
rect 402 -1558 460 -1526
rect 3546 -1526 3604 -1512
rect 3546 -1558 3604 -1526
rect 6678 -1522 6736 -1508
rect 6678 -1554 6736 -1522
rect 9822 -1522 9880 -1508
rect 9822 -1554 9880 -1522
rect 13024 -1526 13082 -1512
rect 13024 -1558 13082 -1526
rect 16168 -1526 16226 -1512
rect 16168 -1558 16226 -1526
rect 19300 -1522 19358 -1508
rect 19300 -1554 19358 -1522
rect 22444 -1522 22502 -1508
rect 22444 -1554 22502 -1522
<< metal1 >>
rect 374 646 384 706
rect 464 646 474 706
rect 374 606 474 646
rect 3518 646 3528 706
rect 3608 646 3618 706
rect 3518 606 3618 646
rect 6650 650 6660 710
rect 6740 650 6750 710
rect 6650 610 6750 650
rect 9794 650 9804 710
rect 9884 650 9894 710
rect 9794 610 9894 650
rect 12996 646 13006 706
rect 13086 646 13096 706
rect -423 549 1380 606
rect -423 430 -389 549
rect 752 422 786 549
rect -1269 -87 -942 -86
rect -1269 -149 -1006 -87
rect -952 -149 -942 -87
rect -865 -124 -830 110
rect -484 95 -420 262
rect 1343 234 1380 549
rect 2721 549 4524 606
rect 2721 430 2755 549
rect 3896 422 3930 549
rect 1343 189 1364 211
rect -476 62 -420 95
rect 44 -22 78 89
rect 1225 -22 1259 90
rect 44 -64 1259 -22
rect 1225 -84 1259 -64
rect 1225 -100 1582 -84
rect -865 -141 272 -124
rect -865 -175 222 -141
rect 256 -175 272 -141
rect 1225 -134 1532 -100
rect 1566 -134 1582 -100
rect 1225 -150 1582 -134
rect -865 -191 272 -175
rect -1270 -236 -948 -228
rect -1270 -304 -1007 -236
rect -950 -304 -940 -236
rect -1270 -312 -948 -304
rect -1270 -512 -1105 -511
rect -1270 -520 -948 -512
rect -1270 -588 -1007 -520
rect -950 -588 -940 -520
rect -1270 -596 -948 -588
rect -1270 -597 -1105 -596
rect -865 -701 -830 -191
rect -775 -237 -683 -224
rect -775 -300 -763 -237
rect -692 -300 -683 -237
rect -775 -309 -683 -300
rect 310 -237 402 -227
rect 310 -299 322 -237
rect 392 -299 402 -237
rect 310 -312 402 -299
rect 1698 -292 1733 110
rect 2279 -124 2314 110
rect 2660 95 2724 262
rect 4487 234 4524 549
rect 5853 553 7656 610
rect 5853 434 5887 553
rect 7028 426 7062 553
rect 4487 189 4508 211
rect 2668 62 2724 95
rect 3188 -22 3222 89
rect 4369 -22 4403 90
rect 3188 -64 4403 -22
rect 4369 -84 4403 -64
rect 4369 -100 4726 -84
rect 2012 -187 2022 -134
rect 2082 -187 2092 -134
rect 2279 -141 3416 -124
rect 2279 -175 3366 -141
rect 3400 -175 3416 -141
rect 4369 -134 4676 -100
rect 4710 -134 4726 -100
rect 4369 -150 4726 -134
rect 557 -354 622 -351
rect 557 -357 626 -354
rect 557 -417 563 -357
rect 622 -417 632 -357
rect 1698 -410 1879 -292
rect 2020 -344 2083 -187
rect 2279 -191 3416 -175
rect 2020 -352 2196 -344
rect 557 -421 626 -417
rect 557 -423 622 -421
rect 1698 -438 1880 -410
rect 2020 -420 2137 -352
rect 2194 -420 2204 -352
rect 2020 -428 2196 -420
rect 192 -520 284 -512
rect 192 -585 204 -520
rect 272 -585 284 -520
rect 192 -597 284 -585
rect 1698 -700 1733 -438
rect -865 -748 507 -701
rect 829 -747 1733 -700
rect -1270 -762 -943 -761
rect -1270 -824 -1007 -762
rect -953 -824 -943 -762
rect -1270 -897 -943 -896
rect -1270 -959 -1007 -897
rect -953 -959 -943 -897
rect -31 -950 3 -748
rect 441 -761 507 -748
rect 441 -795 457 -761
rect 491 -795 507 -761
rect 441 -811 507 -795
rect -1268 -1009 -941 -1008
rect -1268 -1071 -1005 -1009
rect -951 -1071 -941 -1009
rect 115 -1018 167 -871
rect 668 -960 735 -871
rect 830 -950 864 -747
rect 667 -987 735 -960
rect 88 -1071 167 -1018
rect 644 -1018 735 -987
rect 644 -1071 746 -1018
rect -1268 -1134 -941 -1133
rect -1268 -1196 -1005 -1134
rect -951 -1196 -941 -1134
rect -1263 -1375 -936 -1374
rect -1263 -1437 -1000 -1375
rect -946 -1437 -936 -1375
rect 88 -1438 122 -1071
rect 398 -1344 432 -1242
rect 383 -1360 449 -1344
rect 383 -1394 399 -1360
rect 433 -1394 449 -1360
rect 383 -1410 449 -1394
rect 712 -1438 746 -1071
rect 88 -1490 746 -1438
rect 386 -1512 478 -1490
rect 386 -1564 398 -1512
rect 464 -1564 478 -1512
rect 386 -1568 478 -1564
rect -1266 -1597 -939 -1596
rect -1266 -1659 -1003 -1597
rect -949 -1659 -939 -1597
rect 1819 -1648 1880 -438
rect 2020 -520 2196 -512
rect 2020 -588 2137 -520
rect 2194 -588 2204 -520
rect 2020 -596 2196 -588
rect 2020 -758 2109 -596
rect 2279 -701 2314 -191
rect 2369 -237 2461 -224
rect 2369 -300 2381 -237
rect 2452 -300 2461 -237
rect 2369 -309 2461 -300
rect 3454 -237 3546 -227
rect 3454 -299 3466 -237
rect 3536 -299 3546 -237
rect 3454 -312 3546 -299
rect 4842 -292 4877 110
rect 5411 -120 5446 114
rect 5792 99 5856 266
rect 7619 238 7656 553
rect 8997 553 10800 610
rect 12996 606 13096 646
rect 16140 646 16150 706
rect 16230 646 16240 706
rect 16140 606 16240 646
rect 19272 650 19282 710
rect 19362 650 19372 710
rect 19272 610 19372 650
rect 22416 650 22426 710
rect 22506 650 22516 710
rect 22416 610 22516 650
rect 8997 434 9031 553
rect 10172 426 10206 553
rect 7619 193 7640 215
rect 5800 66 5856 99
rect 6320 -18 6354 93
rect 7501 -18 7535 94
rect 6320 -60 7535 -18
rect 7501 -80 7535 -60
rect 7501 -96 7858 -80
rect 5411 -137 6548 -120
rect 5411 -171 6498 -137
rect 6532 -171 6548 -137
rect 7501 -130 7808 -96
rect 7842 -130 7858 -96
rect 7501 -146 7858 -130
rect 5411 -187 6548 -171
rect 3701 -354 3766 -351
rect 3701 -357 3770 -354
rect 3701 -417 3707 -357
rect 3766 -417 3776 -357
rect 3701 -421 3770 -417
rect 3701 -423 3766 -421
rect 4842 -438 5023 -292
rect 3336 -520 3428 -512
rect 3336 -585 3348 -520
rect 3416 -585 3428 -520
rect 3336 -597 3428 -585
rect 4842 -700 4877 -438
rect 2279 -748 3651 -701
rect 3973 -747 4877 -700
rect 2020 -818 2032 -758
rect 2102 -818 2112 -758
rect 2020 -825 2109 -818
rect 3113 -950 3147 -748
rect 3585 -761 3651 -748
rect 3585 -795 3601 -761
rect 3635 -795 3651 -761
rect 3585 -811 3651 -795
rect 3259 -1018 3311 -871
rect 3812 -960 3879 -871
rect 3974 -950 4008 -747
rect 3811 -987 3879 -960
rect 3232 -1071 3311 -1018
rect 3788 -1018 3879 -987
rect 3788 -1071 3890 -1018
rect 3232 -1438 3266 -1071
rect 3542 -1344 3576 -1242
rect 3527 -1360 3593 -1344
rect 3527 -1394 3543 -1360
rect 3577 -1394 3593 -1360
rect 3527 -1410 3593 -1394
rect 3856 -1438 3890 -1071
rect 4935 -1368 5023 -438
rect 5152 -516 5328 -508
rect 5152 -584 5269 -516
rect 5326 -584 5336 -516
rect 5152 -592 5328 -584
rect 5172 -899 5249 -592
rect 5411 -697 5446 -187
rect 5501 -233 5593 -220
rect 5501 -296 5513 -233
rect 5584 -296 5593 -233
rect 5501 -305 5593 -296
rect 6586 -233 6678 -223
rect 6586 -295 6598 -233
rect 6668 -295 6678 -233
rect 6586 -308 6678 -295
rect 7974 -288 8009 114
rect 8555 -120 8590 114
rect 8936 99 9000 266
rect 10763 238 10800 553
rect 12199 549 14002 606
rect 12199 430 12233 549
rect 13374 422 13408 549
rect 10763 193 10784 215
rect 8944 66 9000 99
rect 9464 -18 9498 93
rect 10645 -18 10679 94
rect 9464 -60 10679 -18
rect 10645 -80 10679 -60
rect 10645 -96 11002 -80
rect 8555 -137 9692 -120
rect 8555 -171 9642 -137
rect 9676 -171 9692 -137
rect 10645 -130 10952 -96
rect 10986 -130 11002 -96
rect 10645 -146 11002 -130
rect 8555 -187 9692 -171
rect 6833 -350 6898 -347
rect 6833 -353 6902 -350
rect 6833 -413 6839 -353
rect 6898 -413 6908 -353
rect 6833 -417 6902 -413
rect 6833 -419 6898 -417
rect 7974 -434 8155 -288
rect 8401 -348 8472 -340
rect 8401 -416 8413 -348
rect 8470 -416 8480 -348
rect 8401 -424 8472 -416
rect 6468 -516 6560 -508
rect 6468 -581 6480 -516
rect 6548 -581 6560 -516
rect 6468 -593 6560 -581
rect 7974 -696 8009 -434
rect 5411 -744 6783 -697
rect 7105 -743 8009 -696
rect 5172 -956 5182 -899
rect 5246 -956 5256 -899
rect 6245 -946 6279 -744
rect 6717 -757 6783 -744
rect 6717 -791 6733 -757
rect 6767 -791 6783 -757
rect 6717 -807 6783 -791
rect 5172 -960 5249 -956
rect 6391 -1014 6443 -867
rect 6944 -956 7011 -867
rect 7106 -946 7140 -743
rect 6943 -983 7011 -956
rect 4904 -1434 4914 -1368
rect 4973 -1434 5023 -1368
rect 6364 -1067 6443 -1014
rect 6920 -1014 7011 -983
rect 6920 -1067 7022 -1014
rect 6364 -1434 6398 -1067
rect 6674 -1340 6708 -1238
rect 6659 -1356 6725 -1340
rect 6659 -1390 6675 -1356
rect 6709 -1390 6725 -1356
rect 6659 -1406 6725 -1390
rect 6988 -1434 7022 -1067
rect 8058 -1251 8155 -434
rect 8296 -516 8472 -508
rect 8296 -584 8413 -516
rect 8470 -584 8480 -516
rect 8296 -592 8472 -584
rect 8301 -1004 8389 -592
rect 8555 -697 8590 -187
rect 8645 -233 8737 -220
rect 8645 -296 8657 -233
rect 8728 -296 8737 -233
rect 8645 -305 8737 -296
rect 9730 -233 9822 -223
rect 9730 -295 9742 -233
rect 9812 -295 9822 -233
rect 9730 -308 9822 -295
rect 11118 -288 11153 114
rect 11757 -124 11792 110
rect 12138 95 12202 262
rect 13965 234 14002 549
rect 15343 549 17146 606
rect 15343 430 15377 549
rect 16518 422 16552 549
rect 13965 189 13986 211
rect 12146 62 12202 95
rect 12666 -22 12700 89
rect 13847 -22 13881 90
rect 12666 -64 13881 -22
rect 13847 -84 13881 -64
rect 13847 -100 14204 -84
rect 11757 -141 12894 -124
rect 11757 -175 12844 -141
rect 12878 -175 12894 -141
rect 13847 -134 14154 -100
rect 14188 -134 14204 -100
rect 13847 -150 14204 -134
rect 11757 -191 12894 -175
rect 9977 -350 10042 -347
rect 9977 -353 10046 -350
rect 9977 -413 9983 -353
rect 10042 -413 10052 -353
rect 9977 -417 10046 -413
rect 9977 -419 10042 -417
rect 11118 -434 11299 -288
rect 9612 -516 9704 -508
rect 9612 -581 9624 -516
rect 9692 -581 9704 -516
rect 9612 -593 9704 -581
rect 11118 -696 11153 -434
rect 8555 -744 9927 -697
rect 10249 -743 11153 -696
rect 9389 -946 9423 -744
rect 9861 -757 9927 -744
rect 9861 -791 9877 -757
rect 9911 -791 9927 -757
rect 9861 -807 9927 -791
rect 8301 -1062 8324 -1004
rect 8378 -1062 8389 -1004
rect 9535 -1014 9587 -867
rect 10088 -956 10155 -867
rect 10250 -946 10284 -743
rect 10087 -983 10155 -956
rect 8301 -1072 8389 -1062
rect 9508 -1067 9587 -1014
rect 10064 -1014 10155 -983
rect 10064 -1067 10166 -1014
rect 8030 -1308 8040 -1251
rect 8099 -1308 8155 -1251
rect 8030 -1309 8155 -1308
rect 3232 -1490 3890 -1438
rect 6364 -1486 7022 -1434
rect 9508 -1434 9542 -1067
rect 9818 -1340 9852 -1238
rect 9803 -1356 9869 -1340
rect 9803 -1390 9819 -1356
rect 9853 -1390 9869 -1356
rect 9803 -1406 9869 -1390
rect 10132 -1434 10166 -1067
rect 11205 -1103 11298 -434
rect 11205 -1171 11215 -1103
rect 11277 -1171 11298 -1103
rect 11205 -1176 11298 -1171
rect 11498 -520 11674 -512
rect 11498 -588 11615 -520
rect 11672 -588 11682 -520
rect 11498 -596 11674 -588
rect 11498 -1228 11564 -596
rect 11757 -701 11792 -191
rect 11847 -237 11939 -224
rect 11847 -300 11859 -237
rect 11930 -300 11939 -237
rect 11847 -309 11939 -300
rect 12932 -237 13024 -227
rect 12932 -299 12944 -237
rect 13014 -299 13024 -237
rect 12932 -312 13024 -299
rect 14320 -292 14355 110
rect 14901 -124 14936 110
rect 15282 95 15346 262
rect 17109 234 17146 549
rect 18475 553 20278 610
rect 18475 434 18509 553
rect 19650 426 19684 553
rect 17109 189 17130 211
rect 15290 62 15346 95
rect 15810 -22 15844 89
rect 16991 -22 17025 90
rect 15810 -64 17025 -22
rect 16991 -84 17025 -64
rect 16991 -100 17348 -84
rect 14901 -141 16038 -124
rect 14901 -175 15988 -141
rect 16022 -175 16038 -141
rect 16991 -134 17298 -100
rect 17332 -134 17348 -100
rect 16991 -150 17348 -134
rect 14901 -191 16038 -175
rect 13179 -354 13244 -351
rect 13179 -357 13248 -354
rect 13179 -417 13185 -357
rect 13244 -417 13254 -357
rect 13179 -421 13248 -417
rect 13179 -423 13244 -421
rect 14320 -438 14501 -292
rect 14747 -352 14818 -347
rect 14747 -420 14759 -352
rect 14816 -420 14826 -352
rect 14747 -426 14818 -420
rect 12814 -520 12906 -512
rect 12814 -585 12826 -520
rect 12894 -585 12906 -520
rect 12814 -597 12906 -585
rect 14320 -700 14355 -438
rect 11757 -748 13129 -701
rect 13451 -747 14355 -700
rect 12591 -950 12625 -748
rect 13063 -761 13129 -748
rect 13063 -795 13079 -761
rect 13113 -795 13129 -761
rect 13063 -811 13129 -795
rect 12737 -1018 12789 -871
rect 13290 -960 13357 -871
rect 13452 -950 13486 -747
rect 14431 -952 14501 -438
rect 14642 -520 14818 -512
rect 14642 -588 14759 -520
rect 14816 -588 14826 -520
rect 14642 -596 14818 -588
rect 13289 -987 13357 -960
rect 12710 -1071 12789 -1018
rect 13266 -1018 13357 -987
rect 13266 -1071 13368 -1018
rect 14430 -1021 14440 -952
rect 14496 -1021 14506 -952
rect 14431 -1027 14501 -1021
rect 11484 -1289 11494 -1228
rect 11563 -1289 11573 -1228
rect 11484 -1297 11573 -1289
rect 9508 -1486 10166 -1434
rect 12710 -1438 12744 -1071
rect 13020 -1344 13054 -1242
rect 13005 -1360 13071 -1344
rect 13005 -1394 13021 -1360
rect 13055 -1394 13071 -1360
rect 13005 -1410 13071 -1394
rect 13334 -1438 13368 -1071
rect 14642 -1363 14725 -596
rect 14901 -701 14936 -191
rect 14991 -237 15083 -224
rect 14991 -300 15003 -237
rect 15074 -300 15083 -237
rect 14991 -309 15083 -300
rect 16076 -237 16168 -227
rect 16076 -299 16088 -237
rect 16158 -299 16168 -237
rect 16076 -312 16168 -299
rect 17464 -292 17499 110
rect 18033 -120 18068 114
rect 18414 99 18478 266
rect 20241 238 20278 553
rect 21619 553 23422 610
rect 21619 434 21653 553
rect 22794 426 22828 553
rect 20241 193 20262 215
rect 18422 66 18478 99
rect 18942 -18 18976 93
rect 20123 -18 20157 94
rect 18942 -60 20157 -18
rect 20123 -80 20157 -60
rect 20123 -96 20480 -80
rect 18033 -137 19170 -120
rect 18033 -171 19120 -137
rect 19154 -171 19170 -137
rect 20123 -130 20430 -96
rect 20464 -130 20480 -96
rect 20123 -146 20480 -130
rect 18033 -187 19170 -171
rect 16323 -354 16388 -351
rect 16323 -357 16392 -354
rect 16323 -417 16329 -357
rect 16388 -417 16398 -357
rect 16323 -421 16392 -417
rect 16323 -423 16388 -421
rect 17464 -438 17645 -292
rect 17880 -348 17950 -343
rect 17880 -416 17891 -348
rect 17948 -416 17958 -348
rect 17880 -422 17950 -416
rect 15958 -520 16050 -512
rect 15958 -585 15970 -520
rect 16038 -585 16050 -520
rect 15958 -597 16050 -585
rect 17464 -700 17499 -438
rect 14901 -748 16273 -701
rect 16595 -747 17499 -700
rect 15735 -950 15769 -748
rect 16207 -761 16273 -748
rect 16207 -795 16223 -761
rect 16257 -795 16273 -761
rect 16207 -811 16273 -795
rect 15881 -1018 15933 -871
rect 16434 -960 16501 -871
rect 16596 -950 16630 -747
rect 17573 -799 17645 -438
rect 17774 -516 17950 -508
rect 17774 -584 17891 -516
rect 17948 -584 17958 -516
rect 17774 -592 17950 -584
rect 17566 -858 17576 -799
rect 17640 -858 17650 -799
rect 16433 -987 16501 -960
rect 14635 -1430 14645 -1363
rect 14702 -1427 14725 -1363
rect 15854 -1071 15933 -1018
rect 16410 -1018 16501 -987
rect 16410 -1071 16512 -1018
rect 14702 -1430 14712 -1427
rect 3530 -1512 3622 -1490
rect 3530 -1564 3542 -1512
rect 3608 -1564 3622 -1512
rect 6662 -1508 6754 -1486
rect 6662 -1560 6674 -1508
rect 6740 -1560 6754 -1508
rect 6662 -1564 6754 -1560
rect 9806 -1508 9898 -1486
rect 12710 -1490 13368 -1438
rect 15854 -1438 15888 -1071
rect 16164 -1344 16198 -1242
rect 16149 -1360 16215 -1344
rect 16149 -1394 16165 -1360
rect 16199 -1394 16215 -1360
rect 16149 -1410 16215 -1394
rect 16478 -1438 16512 -1071
rect 15854 -1490 16512 -1438
rect 9806 -1560 9818 -1508
rect 9884 -1560 9898 -1508
rect 9806 -1564 9898 -1560
rect 13008 -1512 13100 -1490
rect 13008 -1564 13020 -1512
rect 13086 -1564 13100 -1512
rect 3530 -1568 3622 -1564
rect 13008 -1568 13100 -1564
rect 16152 -1512 16244 -1490
rect 16152 -1564 16164 -1512
rect 16230 -1564 16244 -1512
rect 16152 -1568 16244 -1564
rect 17774 -1579 17847 -592
rect 18033 -697 18068 -187
rect 18123 -233 18215 -220
rect 18123 -296 18135 -233
rect 18206 -296 18215 -233
rect 18123 -305 18215 -296
rect 19208 -233 19300 -223
rect 19208 -295 19220 -233
rect 19290 -295 19300 -233
rect 19208 -308 19300 -295
rect 20596 -288 20631 114
rect 21177 -120 21212 114
rect 21558 99 21622 266
rect 23385 238 23422 553
rect 23385 193 23406 215
rect 21566 66 21622 99
rect 22086 -18 22120 93
rect 23267 -18 23301 94
rect 22086 -60 23301 -18
rect 23267 -80 23301 -60
rect 23267 -96 23624 -80
rect 21177 -137 22314 -120
rect 21177 -171 22264 -137
rect 22298 -171 22314 -137
rect 23267 -130 23574 -96
rect 23608 -130 23624 -96
rect 23267 -146 23624 -130
rect 21177 -187 22314 -171
rect 19455 -350 19520 -347
rect 19455 -353 19524 -350
rect 19455 -413 19461 -353
rect 19520 -413 19530 -353
rect 20596 -383 20777 -288
rect 21024 -348 21094 -343
rect 19455 -417 19524 -413
rect 19455 -419 19520 -417
rect 20596 -434 20778 -383
rect 21024 -416 21035 -348
rect 21092 -416 21102 -348
rect 21024 -422 21094 -416
rect 19090 -516 19182 -508
rect 19090 -581 19102 -516
rect 19170 -581 19182 -516
rect 19090 -593 19182 -581
rect 20596 -696 20631 -434
rect 18033 -744 19405 -697
rect 19727 -743 20631 -696
rect 20683 -672 20778 -434
rect 20683 -729 20721 -672
rect 20774 -729 20784 -672
rect 21177 -697 21212 -187
rect 21267 -233 21359 -220
rect 21267 -296 21279 -233
rect 21350 -296 21359 -233
rect 21267 -305 21359 -296
rect 22352 -233 22444 -223
rect 22352 -295 22364 -233
rect 22434 -295 22444 -233
rect 22352 -308 22444 -295
rect 23740 -288 23775 114
rect 22599 -350 22664 -347
rect 22599 -353 22668 -350
rect 22599 -413 22605 -353
rect 22664 -413 22674 -353
rect 23740 -376 24354 -288
rect 22599 -417 22668 -413
rect 22599 -419 22664 -417
rect 22234 -516 22326 -508
rect 22234 -581 22246 -516
rect 22314 -581 22326 -516
rect 22234 -593 22326 -581
rect 23740 -696 23775 -376
rect 20683 -737 20778 -729
rect 18867 -946 18901 -744
rect 19339 -757 19405 -744
rect 19339 -791 19355 -757
rect 19389 -791 19405 -757
rect 19339 -807 19405 -791
rect 19013 -1014 19065 -867
rect 19566 -956 19633 -867
rect 19728 -946 19762 -743
rect 21177 -744 22549 -697
rect 22871 -743 23775 -696
rect 24206 -664 24355 -652
rect 24206 -735 24219 -664
rect 24290 -735 24355 -664
rect 22011 -946 22045 -744
rect 22483 -757 22549 -744
rect 22483 -791 22499 -757
rect 22533 -791 22549 -757
rect 22483 -807 22549 -791
rect 19565 -983 19633 -956
rect 18986 -1067 19065 -1014
rect 19542 -1014 19633 -983
rect 22157 -1014 22209 -867
rect 22710 -956 22777 -867
rect 22872 -946 22906 -743
rect 24206 -746 24355 -735
rect 24197 -800 24356 -789
rect 24197 -860 24207 -800
rect 24273 -860 24356 -800
rect 24197 -871 24356 -860
rect 22709 -983 22777 -956
rect 19542 -1067 19644 -1014
rect 18986 -1434 19020 -1067
rect 19296 -1340 19330 -1238
rect 19281 -1356 19347 -1340
rect 19281 -1390 19297 -1356
rect 19331 -1390 19347 -1356
rect 19281 -1406 19347 -1390
rect 19610 -1434 19644 -1067
rect 18986 -1486 19644 -1434
rect 22130 -1067 22209 -1014
rect 22686 -1014 22777 -983
rect 24186 -958 24356 -947
rect 22686 -1067 22788 -1014
rect 24186 -1027 24197 -958
rect 24261 -1027 24356 -958
rect 24186 -1038 24356 -1027
rect 22130 -1434 22164 -1067
rect 22440 -1340 22474 -1238
rect 22425 -1356 22491 -1340
rect 22425 -1390 22441 -1356
rect 22475 -1390 22491 -1356
rect 22425 -1406 22491 -1390
rect 22754 -1434 22788 -1067
rect 24186 -1104 24356 -1093
rect 24186 -1173 24197 -1104
rect 24261 -1173 24356 -1104
rect 24186 -1184 24356 -1173
rect 24186 -1244 24356 -1233
rect 24186 -1313 24197 -1244
rect 24261 -1313 24356 -1244
rect 24186 -1324 24356 -1313
rect 22130 -1486 22788 -1434
rect 24185 -1383 24355 -1372
rect 24185 -1452 24196 -1383
rect 24260 -1452 24355 -1383
rect 24185 -1463 24355 -1452
rect 19284 -1508 19376 -1486
rect 19284 -1560 19296 -1508
rect 19362 -1560 19376 -1508
rect 19284 -1564 19376 -1560
rect 22428 -1508 22520 -1486
rect 22428 -1560 22440 -1508
rect 22506 -1560 22520 -1508
rect 22428 -1564 22520 -1560
rect 1771 -1729 1781 -1648
rect 1854 -1729 1880 -1648
rect 17764 -1655 17774 -1579
rect 17844 -1655 17854 -1579
rect 24185 -1651 24355 -1640
rect 1819 -1730 1880 -1729
rect 24185 -1720 24196 -1651
rect 24260 -1720 24355 -1651
rect 24185 -1731 24355 -1720
<< via1 >>
rect 384 700 464 706
rect 384 646 388 700
rect 388 646 460 700
rect 460 646 464 700
rect 3528 700 3608 706
rect 3528 646 3532 700
rect 3532 646 3604 700
rect 3604 646 3608 700
rect 6660 704 6740 710
rect 6660 650 6664 704
rect 6664 650 6736 704
rect 6736 650 6740 704
rect 9804 704 9884 710
rect 9804 650 9808 704
rect 9808 650 9880 704
rect 9880 650 9884 704
rect 13006 700 13086 706
rect 13006 646 13010 700
rect 13010 646 13082 700
rect 13082 646 13086 700
rect -1006 -149 -952 -87
rect -1007 -240 -950 -236
rect -1007 -300 -1003 -240
rect -1003 -300 -954 -240
rect -954 -300 -950 -240
rect -1007 -304 -950 -300
rect -1007 -524 -950 -520
rect -1007 -584 -1003 -524
rect -1003 -584 -954 -524
rect -954 -584 -950 -524
rect -1007 -588 -950 -584
rect -763 -241 -692 -237
rect -763 -296 -759 -241
rect -759 -296 -699 -241
rect -699 -296 -692 -241
rect -763 -300 -692 -296
rect 322 -240 392 -237
rect 322 -295 326 -240
rect 326 -295 386 -240
rect 386 -295 392 -240
rect 322 -299 392 -295
rect 2022 -187 2082 -134
rect 563 -371 622 -357
rect 563 -405 576 -371
rect 576 -405 610 -371
rect 610 -405 622 -371
rect 563 -417 622 -405
rect 2137 -356 2194 -352
rect 2137 -416 2141 -356
rect 2141 -416 2190 -356
rect 2190 -416 2194 -356
rect 2137 -420 2194 -416
rect 204 -525 272 -520
rect 204 -580 208 -525
rect 208 -580 268 -525
rect 268 -580 272 -525
rect 204 -585 272 -580
rect -1007 -824 -953 -762
rect -1007 -959 -953 -897
rect -1005 -1071 -951 -1009
rect -1005 -1196 -951 -1134
rect -1000 -1437 -946 -1375
rect 398 -1558 402 -1512
rect 402 -1558 460 -1512
rect 460 -1558 464 -1512
rect 398 -1564 464 -1558
rect -1003 -1659 -949 -1597
rect 2137 -524 2194 -520
rect 2137 -584 2141 -524
rect 2141 -584 2190 -524
rect 2190 -584 2194 -524
rect 2137 -588 2194 -584
rect 2381 -241 2452 -237
rect 2381 -296 2385 -241
rect 2385 -296 2445 -241
rect 2445 -296 2452 -241
rect 2381 -300 2452 -296
rect 3466 -240 3536 -237
rect 3466 -295 3470 -240
rect 3470 -295 3530 -240
rect 3530 -295 3536 -240
rect 3466 -299 3536 -295
rect 16150 700 16230 706
rect 16150 646 16154 700
rect 16154 646 16226 700
rect 16226 646 16230 700
rect 19282 704 19362 710
rect 19282 650 19286 704
rect 19286 650 19358 704
rect 19358 650 19362 704
rect 22426 704 22506 710
rect 22426 650 22430 704
rect 22430 650 22502 704
rect 22502 650 22506 704
rect 3707 -371 3766 -357
rect 3707 -405 3720 -371
rect 3720 -405 3754 -371
rect 3754 -405 3766 -371
rect 3707 -417 3766 -405
rect 3348 -525 3416 -520
rect 3348 -580 3352 -525
rect 3352 -580 3412 -525
rect 3412 -580 3416 -525
rect 3348 -585 3416 -580
rect 2032 -818 2102 -758
rect 5269 -520 5326 -516
rect 5269 -580 5273 -520
rect 5273 -580 5322 -520
rect 5322 -580 5326 -520
rect 5269 -584 5326 -580
rect 5513 -237 5584 -233
rect 5513 -292 5517 -237
rect 5517 -292 5577 -237
rect 5577 -292 5584 -237
rect 5513 -296 5584 -292
rect 6598 -236 6668 -233
rect 6598 -291 6602 -236
rect 6602 -291 6662 -236
rect 6662 -291 6668 -236
rect 6598 -295 6668 -291
rect 6839 -367 6898 -353
rect 6839 -401 6852 -367
rect 6852 -401 6886 -367
rect 6886 -401 6898 -367
rect 6839 -413 6898 -401
rect 8413 -352 8470 -348
rect 8413 -412 8417 -352
rect 8417 -412 8466 -352
rect 8466 -412 8470 -352
rect 8413 -416 8470 -412
rect 6480 -521 6548 -516
rect 6480 -576 6484 -521
rect 6484 -576 6544 -521
rect 6544 -576 6548 -521
rect 6480 -581 6548 -576
rect 5182 -956 5246 -899
rect 4914 -1434 4973 -1368
rect 8413 -520 8470 -516
rect 8413 -580 8417 -520
rect 8417 -580 8466 -520
rect 8466 -580 8470 -520
rect 8413 -584 8470 -580
rect 8657 -237 8728 -233
rect 8657 -292 8661 -237
rect 8661 -292 8721 -237
rect 8721 -292 8728 -237
rect 8657 -296 8728 -292
rect 9742 -236 9812 -233
rect 9742 -291 9746 -236
rect 9746 -291 9806 -236
rect 9806 -291 9812 -236
rect 9742 -295 9812 -291
rect 9983 -367 10042 -353
rect 9983 -401 9996 -367
rect 9996 -401 10030 -367
rect 10030 -401 10042 -367
rect 9983 -413 10042 -401
rect 9624 -521 9692 -516
rect 9624 -576 9628 -521
rect 9628 -576 9688 -521
rect 9688 -576 9692 -521
rect 9624 -581 9692 -576
rect 8324 -1062 8378 -1004
rect 8040 -1308 8099 -1251
rect 11215 -1171 11277 -1103
rect 11615 -524 11672 -520
rect 11615 -584 11619 -524
rect 11619 -584 11668 -524
rect 11668 -584 11672 -524
rect 11615 -588 11672 -584
rect 11859 -241 11930 -237
rect 11859 -296 11863 -241
rect 11863 -296 11923 -241
rect 11923 -296 11930 -241
rect 11859 -300 11930 -296
rect 12944 -240 13014 -237
rect 12944 -295 12948 -240
rect 12948 -295 13008 -240
rect 13008 -295 13014 -240
rect 12944 -299 13014 -295
rect 13185 -371 13244 -357
rect 13185 -405 13198 -371
rect 13198 -405 13232 -371
rect 13232 -405 13244 -371
rect 13185 -417 13244 -405
rect 14759 -356 14816 -352
rect 14759 -416 14763 -356
rect 14763 -416 14812 -356
rect 14812 -416 14816 -356
rect 14759 -420 14816 -416
rect 12826 -525 12894 -520
rect 12826 -580 12830 -525
rect 12830 -580 12890 -525
rect 12890 -580 12894 -525
rect 12826 -585 12894 -580
rect 14759 -524 14816 -520
rect 14759 -584 14763 -524
rect 14763 -584 14812 -524
rect 14812 -584 14816 -524
rect 14759 -588 14816 -584
rect 14440 -1021 14496 -952
rect 11494 -1289 11563 -1228
rect 15003 -241 15074 -237
rect 15003 -296 15007 -241
rect 15007 -296 15067 -241
rect 15067 -296 15074 -241
rect 15003 -300 15074 -296
rect 16088 -240 16158 -237
rect 16088 -295 16092 -240
rect 16092 -295 16152 -240
rect 16152 -295 16158 -240
rect 16088 -299 16158 -295
rect 16329 -371 16388 -357
rect 16329 -405 16342 -371
rect 16342 -405 16376 -371
rect 16376 -405 16388 -371
rect 16329 -417 16388 -405
rect 17891 -352 17948 -348
rect 17891 -412 17895 -352
rect 17895 -412 17944 -352
rect 17944 -412 17948 -352
rect 17891 -416 17948 -412
rect 15970 -525 16038 -520
rect 15970 -580 15974 -525
rect 15974 -580 16034 -525
rect 16034 -580 16038 -525
rect 15970 -585 16038 -580
rect 17891 -520 17948 -516
rect 17891 -580 17895 -520
rect 17895 -580 17944 -520
rect 17944 -580 17948 -520
rect 17891 -584 17948 -580
rect 17576 -858 17640 -799
rect 14645 -1430 14702 -1363
rect 3542 -1558 3546 -1512
rect 3546 -1558 3604 -1512
rect 3604 -1558 3608 -1512
rect 3542 -1564 3608 -1558
rect 6674 -1554 6678 -1508
rect 6678 -1554 6736 -1508
rect 6736 -1554 6740 -1508
rect 6674 -1560 6740 -1554
rect 9818 -1554 9822 -1508
rect 9822 -1554 9880 -1508
rect 9880 -1554 9884 -1508
rect 9818 -1560 9884 -1554
rect 13020 -1558 13024 -1512
rect 13024 -1558 13082 -1512
rect 13082 -1558 13086 -1512
rect 13020 -1564 13086 -1558
rect 16164 -1558 16168 -1512
rect 16168 -1558 16226 -1512
rect 16226 -1558 16230 -1512
rect 16164 -1564 16230 -1558
rect 18135 -237 18206 -233
rect 18135 -292 18139 -237
rect 18139 -292 18199 -237
rect 18199 -292 18206 -237
rect 18135 -296 18206 -292
rect 19220 -236 19290 -233
rect 19220 -291 19224 -236
rect 19224 -291 19284 -236
rect 19284 -291 19290 -236
rect 19220 -295 19290 -291
rect 19461 -367 19520 -353
rect 19461 -401 19474 -367
rect 19474 -401 19508 -367
rect 19508 -401 19520 -367
rect 19461 -413 19520 -401
rect 21035 -352 21092 -348
rect 21035 -412 21039 -352
rect 21039 -412 21088 -352
rect 21088 -412 21092 -352
rect 21035 -416 21092 -412
rect 19102 -521 19170 -516
rect 19102 -576 19106 -521
rect 19106 -576 19166 -521
rect 19166 -576 19170 -521
rect 19102 -581 19170 -576
rect 20721 -729 20774 -672
rect 21279 -237 21350 -233
rect 21279 -292 21283 -237
rect 21283 -292 21343 -237
rect 21343 -292 21350 -237
rect 21279 -296 21350 -292
rect 22364 -236 22434 -233
rect 22364 -291 22368 -236
rect 22368 -291 22428 -236
rect 22428 -291 22434 -236
rect 22364 -295 22434 -291
rect 22605 -367 22664 -353
rect 22605 -401 22618 -367
rect 22618 -401 22652 -367
rect 22652 -401 22664 -367
rect 22605 -413 22664 -401
rect 22246 -521 22314 -516
rect 22246 -576 22250 -521
rect 22250 -576 22310 -521
rect 22310 -576 22314 -521
rect 22246 -581 22314 -576
rect 24219 -735 24290 -664
rect 24207 -860 24273 -800
rect 24197 -1027 24261 -958
rect 24197 -1173 24261 -1104
rect 24197 -1313 24261 -1244
rect 24196 -1452 24260 -1383
rect 19296 -1554 19300 -1508
rect 19300 -1554 19358 -1508
rect 19358 -1554 19362 -1508
rect 19296 -1560 19362 -1554
rect 22440 -1554 22444 -1508
rect 22444 -1554 22502 -1508
rect 22502 -1554 22506 -1508
rect 22440 -1560 22506 -1554
rect 1781 -1729 1854 -1648
rect 17774 -1655 17844 -1579
rect 24196 -1720 24260 -1651
<< metal2 >>
rect 372 734 472 744
rect 372 632 472 642
rect 3516 734 3616 744
rect 3516 632 3616 642
rect 6648 738 6748 748
rect 6648 636 6748 646
rect 9792 738 9892 748
rect 9792 636 9892 646
rect 12994 734 13094 744
rect 12994 632 13094 642
rect 16138 734 16238 744
rect 16138 632 16238 642
rect 19270 738 19370 748
rect 19270 636 19370 646
rect 22414 738 22514 748
rect 22414 636 22514 646
rect -1006 -85 -952 -77
rect -1017 -87 2082 -85
rect -1017 -149 -1006 -87
rect -952 -134 2082 -87
rect -952 -149 2022 -134
rect -1017 -150 -938 -149
rect -1006 -159 -952 -150
rect 2022 -197 2082 -187
rect 5502 -223 5595 -221
rect 8646 -223 8739 -221
rect 18124 -223 18217 -221
rect 21268 -223 21361 -221
rect -1007 -227 -950 -226
rect -774 -227 -681 -225
rect 2370 -227 2463 -225
rect 3413 -227 9821 -223
rect 11848 -227 11941 -225
rect 14992 -227 15085 -225
rect 16076 -227 22443 -223
rect -1015 -228 401 -227
rect 2196 -228 22443 -227
rect -1018 -233 22443 -228
rect -1018 -236 5513 -233
rect -1018 -304 -1007 -236
rect -950 -237 5513 -236
rect -950 -300 -763 -237
rect -692 -299 322 -237
rect 392 -299 2381 -237
rect -692 -300 2381 -299
rect 2452 -299 3466 -237
rect 3536 -296 5513 -237
rect 5584 -295 6598 -233
rect 6668 -295 8657 -233
rect 5584 -296 8657 -295
rect 8728 -295 9742 -233
rect 9812 -237 18135 -233
rect 9812 -295 11859 -237
rect 8728 -296 11859 -295
rect 3536 -299 11859 -296
rect 2452 -300 11859 -299
rect 11930 -299 12944 -237
rect 13014 -299 15003 -237
rect 11930 -300 15003 -299
rect 15074 -299 16088 -237
rect 16158 -296 18135 -237
rect 18206 -295 19220 -233
rect 19290 -295 21279 -233
rect 18206 -296 21279 -295
rect 21350 -295 22364 -233
rect 22434 -295 22443 -233
rect 21350 -296 22443 -295
rect 16158 -299 22443 -296
rect 15074 -300 22443 -299
rect -950 -304 22443 -300
rect -1018 -307 22443 -304
rect -1018 -308 5336 -307
rect -1018 -311 5226 -308
rect 11604 -311 17955 -307
rect -1018 -312 -940 -311
rect 358 -312 2204 -311
rect 12932 -312 14826 -311
rect -1007 -314 -950 -312
rect 8413 -340 8470 -338
rect 2137 -344 2194 -342
rect 8402 -343 8498 -340
rect 2126 -347 2222 -344
rect -1018 -357 622 -347
rect -1018 -361 563 -357
rect -1018 -417 -1008 -361
rect -952 -417 563 -361
rect -1018 -426 622 -417
rect -1008 -427 -952 -426
rect 563 -427 622 -426
rect 2126 -352 3766 -347
rect 2126 -420 2137 -352
rect 2194 -357 3766 -352
rect 2194 -417 3707 -357
rect 2194 -420 3766 -417
rect 2126 -426 3766 -420
rect 2126 -429 2222 -426
rect 3707 -427 3766 -426
rect 5080 -353 6898 -343
rect 5080 -413 6839 -353
rect 5080 -422 6898 -413
rect 2137 -430 2194 -429
rect 5080 -466 5137 -422
rect 6839 -423 6898 -422
rect 8402 -348 10042 -343
rect 8402 -416 8413 -348
rect 8470 -353 10042 -348
rect 8470 -413 9983 -353
rect 8470 -416 10042 -413
rect 8402 -422 10042 -416
rect 8402 -425 8498 -422
rect 9983 -423 10042 -422
rect 11337 -357 13244 -347
rect 11337 -417 13185 -357
rect 8413 -426 8470 -425
rect 11337 -426 13244 -417
rect 14748 -352 16388 -347
rect 14748 -420 14759 -352
rect 14816 -357 16388 -352
rect 14816 -417 16329 -357
rect 14816 -420 16388 -417
rect 14748 -426 16388 -420
rect -1007 -511 -950 -510
rect 2137 -511 2194 -510
rect 4922 -511 5137 -466
rect 5269 -507 5326 -506
rect 8413 -507 8470 -506
rect 5258 -508 5354 -507
rect 8402 -508 8498 -507
rect -1018 -512 -922 -511
rect 2126 -512 2222 -511
rect -1018 -520 1815 -512
rect -1018 -588 -1007 -520
rect -950 -585 204 -520
rect 272 -585 1815 -520
rect -950 -588 1815 -585
rect -1018 -596 1815 -588
rect 2126 -520 3427 -512
rect 2126 -588 2137 -520
rect 2194 -585 3348 -520
rect 3416 -585 3427 -520
rect 2194 -588 3427 -585
rect 2126 -596 3427 -588
rect -1007 -598 -950 -596
rect 1740 -637 1815 -596
rect 2137 -598 2194 -596
rect 4922 -637 4994 -511
rect 5258 -516 8036 -508
rect 5258 -584 5269 -516
rect 5326 -581 6480 -516
rect 6548 -581 8036 -516
rect 5326 -584 8036 -581
rect 5258 -592 8036 -584
rect 8402 -516 9703 -508
rect 8402 -584 8413 -516
rect 8470 -581 9624 -516
rect 9692 -581 9703 -516
rect 8470 -584 9703 -581
rect 8402 -592 9703 -584
rect 5269 -594 5326 -592
rect 1740 -702 4994 -637
rect 7957 -675 8036 -592
rect 8413 -594 8470 -592
rect 11337 -675 11427 -426
rect 13185 -427 13244 -426
rect 16329 -427 16388 -426
rect 17658 -348 19520 -343
rect 17658 -416 17891 -348
rect 17948 -353 19520 -348
rect 17948 -413 19461 -353
rect 17948 -416 19520 -413
rect 17658 -422 19520 -416
rect 21024 -348 22664 -343
rect 21024 -416 21035 -348
rect 21092 -353 22664 -348
rect 21092 -413 22605 -353
rect 21092 -416 22664 -413
rect 21024 -422 22664 -416
rect 11615 -511 11672 -510
rect 14759 -511 14816 -510
rect 11604 -512 11700 -511
rect 14748 -512 14844 -511
rect 11604 -520 12906 -512
rect 11604 -588 11615 -520
rect 11672 -585 12826 -520
rect 12894 -585 12906 -520
rect 11672 -588 12906 -585
rect 11604 -596 12906 -588
rect 14748 -520 16049 -512
rect 14748 -588 14759 -520
rect 14816 -585 15970 -520
rect 16038 -585 16049 -520
rect 14816 -588 16049 -585
rect 14748 -596 16049 -588
rect 11615 -598 11672 -596
rect 7957 -743 11427 -675
rect 12825 -653 12906 -596
rect 14759 -598 14816 -596
rect 17658 -653 17739 -422
rect 19461 -423 19520 -422
rect 22605 -423 22664 -422
rect 21024 -506 21103 -496
rect 17891 -507 17948 -506
rect 17880 -508 17976 -507
rect 17880 -516 19181 -508
rect 17880 -584 17891 -516
rect 17948 -581 19102 -516
rect 19170 -581 19181 -516
rect 17948 -584 19181 -581
rect 17880 -592 19181 -584
rect 17891 -594 17948 -592
rect 21103 -508 21120 -507
rect 21103 -516 22325 -508
rect 21103 -581 22246 -516
rect 22314 -581 22325 -516
rect 21103 -592 22325 -581
rect 21024 -605 21103 -595
rect 12825 -732 17739 -653
rect 20721 -654 24255 -653
rect 20721 -664 24290 -654
rect 20721 -672 24219 -664
rect 20774 -729 24219 -672
rect 20721 -735 24219 -729
rect 20721 -743 24290 -735
rect 24219 -745 24290 -743
rect -1007 -761 -953 -752
rect 2032 -758 2102 -748
rect -1018 -762 2032 -761
rect -1018 -824 -1007 -762
rect -953 -818 2032 -762
rect 2102 -818 2109 -761
rect -953 -824 2109 -818
rect -1018 -825 2109 -824
rect 17576 -799 17640 -789
rect -1007 -834 -953 -825
rect 2032 -828 2102 -825
rect 17576 -868 17640 -858
rect 24207 -800 24273 -790
rect 24207 -870 24273 -860
rect -1007 -896 -953 -887
rect 5182 -896 5246 -889
rect -1018 -897 5246 -896
rect -1018 -959 -1007 -897
rect -953 -899 5246 -897
rect -953 -956 5182 -899
rect -953 -959 5246 -956
rect -1018 -960 5246 -959
rect -1007 -969 -953 -960
rect 5182 -966 5246 -960
rect 14440 -952 14496 -942
rect -1005 -1008 -951 -999
rect 8324 -1004 8378 -994
rect -1016 -1009 8324 -1008
rect -1016 -1071 -1005 -1009
rect -951 -1062 8324 -1009
rect 14440 -1031 14496 -1021
rect 24197 -958 24261 -948
rect 24197 -1037 24261 -1027
rect -951 -1071 8378 -1062
rect -1016 -1072 8378 -1071
rect -1005 -1081 -951 -1072
rect 11215 -1103 11277 -1093
rect -1005 -1133 -951 -1124
rect -1016 -1134 -789 -1133
rect -1016 -1196 -1005 -1134
rect -951 -1196 11091 -1134
rect 11215 -1181 11277 -1171
rect 24197 -1104 24261 -1094
rect 24197 -1183 24261 -1173
rect -1016 -1197 11091 -1196
rect -1005 -1206 -951 -1197
rect 11023 -1232 11091 -1197
rect 11494 -1228 11563 -1218
rect 8040 -1251 8099 -1241
rect 4688 -1327 5135 -1263
rect 11023 -1289 11494 -1232
rect 11023 -1296 11563 -1289
rect 11494 -1299 11563 -1296
rect 24197 -1244 24261 -1234
rect 8040 -1318 8099 -1308
rect 24197 -1323 24261 -1313
rect -1000 -1367 -946 -1365
rect 4688 -1367 4752 -1327
rect -1017 -1375 4752 -1367
rect -1017 -1432 -1000 -1375
rect -1011 -1437 -1000 -1432
rect -946 -1432 4752 -1375
rect 4914 -1368 4973 -1358
rect -946 -1437 -935 -1432
rect -1011 -1438 -935 -1437
rect 5071 -1368 5135 -1327
rect 14645 -1363 14702 -1353
rect 5071 -1430 14645 -1368
rect 5071 -1432 14702 -1430
rect -1000 -1447 -946 -1438
rect 4914 -1444 4973 -1434
rect 14645 -1440 14702 -1432
rect 24196 -1383 24260 -1373
rect 24196 -1462 24260 -1452
rect 392 -1510 468 -1500
rect 392 -1578 468 -1568
rect 3536 -1510 3612 -1500
rect 3536 -1578 3612 -1568
rect 6668 -1506 6744 -1496
rect 6668 -1574 6744 -1564
rect 9812 -1506 9888 -1496
rect 9812 -1574 9888 -1564
rect 13014 -1510 13090 -1500
rect 13014 -1578 13090 -1568
rect 16158 -1510 16234 -1500
rect 16158 -1578 16234 -1568
rect 19290 -1506 19366 -1496
rect 17774 -1579 17844 -1569
rect 19290 -1574 19366 -1564
rect 22434 -1506 22510 -1496
rect 22434 -1574 22510 -1564
rect -1003 -1596 -949 -1589
rect -1014 -1597 -896 -1596
rect -1014 -1659 -1003 -1597
rect -949 -1607 -896 -1597
rect -949 -1659 1642 -1607
rect -1014 -1660 1642 -1659
rect -1003 -1669 -949 -1660
rect 1578 -1768 1642 -1660
rect 1781 -1648 1854 -1638
rect 1913 -1655 17774 -1606
rect 1913 -1660 17844 -1655
rect 1913 -1665 1976 -1660
rect 17774 -1665 17844 -1660
rect 24196 -1651 24260 -1641
rect 1781 -1739 1854 -1729
rect 1912 -1768 1976 -1665
rect 24196 -1730 24260 -1720
rect 1578 -1796 1976 -1768
<< via2 >>
rect 372 706 472 734
rect 372 646 384 706
rect 384 646 464 706
rect 464 646 472 706
rect 372 642 472 646
rect 3516 706 3616 734
rect 3516 646 3528 706
rect 3528 646 3608 706
rect 3608 646 3616 706
rect 3516 642 3616 646
rect 6648 710 6748 738
rect 6648 650 6660 710
rect 6660 650 6740 710
rect 6740 650 6748 710
rect 6648 646 6748 650
rect 9792 710 9892 738
rect 9792 650 9804 710
rect 9804 650 9884 710
rect 9884 650 9892 710
rect 9792 646 9892 650
rect 12994 706 13094 734
rect 12994 646 13006 706
rect 13006 646 13086 706
rect 13086 646 13094 706
rect 12994 642 13094 646
rect 16138 706 16238 734
rect 16138 646 16150 706
rect 16150 646 16230 706
rect 16230 646 16238 706
rect 16138 642 16238 646
rect 19270 710 19370 738
rect 19270 650 19282 710
rect 19282 650 19362 710
rect 19362 650 19370 710
rect 19270 646 19370 650
rect 22414 710 22514 738
rect 22414 650 22426 710
rect 22426 650 22506 710
rect 22506 650 22514 710
rect 22414 646 22514 650
rect -1008 -417 -952 -361
rect 21024 -595 21103 -506
rect 17576 -858 17640 -799
rect 24207 -860 24273 -800
rect 14440 -1021 14496 -952
rect 24197 -1027 24261 -958
rect 11215 -1171 11277 -1103
rect 24197 -1173 24261 -1104
rect 8040 -1308 8099 -1251
rect 24197 -1313 24261 -1244
rect 4914 -1434 4973 -1368
rect 24196 -1452 24260 -1383
rect 392 -1512 468 -1510
rect 392 -1564 398 -1512
rect 398 -1564 464 -1512
rect 464 -1564 468 -1512
rect 392 -1568 468 -1564
rect 3536 -1512 3612 -1510
rect 3536 -1564 3542 -1512
rect 3542 -1564 3608 -1512
rect 3608 -1564 3612 -1512
rect 3536 -1568 3612 -1564
rect 6668 -1508 6744 -1506
rect 6668 -1560 6674 -1508
rect 6674 -1560 6740 -1508
rect 6740 -1560 6744 -1508
rect 6668 -1564 6744 -1560
rect 9812 -1508 9888 -1506
rect 9812 -1560 9818 -1508
rect 9818 -1560 9884 -1508
rect 9884 -1560 9888 -1508
rect 9812 -1564 9888 -1560
rect 13014 -1512 13090 -1510
rect 13014 -1564 13020 -1512
rect 13020 -1564 13086 -1512
rect 13086 -1564 13090 -1512
rect 13014 -1568 13090 -1564
rect 16158 -1512 16234 -1510
rect 16158 -1564 16164 -1512
rect 16164 -1564 16230 -1512
rect 16230 -1564 16234 -1512
rect 16158 -1568 16234 -1564
rect 19290 -1508 19366 -1506
rect 19290 -1560 19296 -1508
rect 19296 -1560 19362 -1508
rect 19362 -1560 19366 -1508
rect 19290 -1564 19366 -1560
rect 22434 -1508 22510 -1506
rect 22434 -1560 22440 -1508
rect 22440 -1560 22506 -1508
rect 22506 -1560 22510 -1508
rect 22434 -1564 22510 -1560
rect 1781 -1729 1854 -1648
rect 24196 -1720 24260 -1651
<< metal3 >>
rect 362 734 482 739
rect 362 640 372 734
rect 472 640 482 734
rect 362 637 482 640
rect 3506 734 3626 739
rect 3506 640 3516 734
rect 3616 640 3626 734
rect 6638 738 6758 743
rect 6638 644 6648 738
rect 6748 644 6758 738
rect 6638 641 6758 644
rect 9782 738 9902 743
rect 9782 644 9792 738
rect 9892 644 9902 738
rect 9782 641 9902 644
rect 12984 734 13104 739
rect 3506 637 3626 640
rect 12984 640 12994 734
rect 13094 640 13104 734
rect 12984 637 13104 640
rect 16128 734 16248 739
rect 16128 640 16138 734
rect 16238 640 16248 734
rect 19260 738 19380 743
rect 19260 644 19270 738
rect 19370 644 19380 738
rect 19260 641 19380 644
rect 22404 738 22524 743
rect 22404 644 22414 738
rect 22514 644 22524 738
rect 22404 641 22524 644
rect 16128 637 16248 640
rect -1028 -347 -931 -346
rect -1028 -430 -1018 -347
rect -941 -430 -931 -347
rect -1028 -449 -931 -430
rect 21003 -605 21013 -496
rect 21113 -605 21123 -496
rect 17566 -795 24279 -794
rect 17566 -799 24283 -795
rect 17566 -858 17576 -799
rect 17640 -800 24283 -799
rect 17640 -858 24207 -800
rect 17566 -860 24207 -858
rect 24273 -860 24283 -800
rect 17566 -863 24283 -860
rect 24197 -865 24283 -863
rect 14430 -952 14506 -947
rect 14430 -1021 14440 -952
rect 14496 -958 14506 -952
rect 24187 -958 24271 -953
rect 14496 -1021 24197 -958
rect 14430 -1026 24197 -1021
rect 24187 -1027 24197 -1026
rect 24261 -1027 24271 -958
rect 24187 -1032 24271 -1027
rect 11205 -1103 11287 -1098
rect 11205 -1171 11215 -1103
rect 11277 -1104 11287 -1103
rect 24187 -1104 24271 -1099
rect 11277 -1171 24197 -1104
rect 11205 -1172 24197 -1171
rect 11205 -1176 11287 -1172
rect 24187 -1173 24197 -1172
rect 24261 -1173 24271 -1104
rect 24187 -1178 24271 -1173
rect 24187 -1244 24271 -1239
rect 8085 -1246 24197 -1244
rect 8030 -1251 24197 -1246
rect 8030 -1308 8040 -1251
rect 8099 -1308 24197 -1251
rect 8030 -1312 24197 -1308
rect 8030 -1313 8109 -1312
rect 24187 -1313 24197 -1312
rect 24261 -1313 24271 -1244
rect 24187 -1318 24271 -1313
rect 4904 -1368 4983 -1363
rect 4904 -1434 4914 -1368
rect 4973 -1377 4983 -1368
rect 22650 -1377 24059 -1372
rect 4973 -1382 24059 -1377
rect 24126 -1382 24270 -1378
rect 4973 -1383 24270 -1382
rect 4973 -1434 24196 -1383
rect 4904 -1438 24196 -1434
rect 4904 -1439 4983 -1438
rect 22650 -1446 24196 -1438
rect 24094 -1451 24196 -1446
rect 24186 -1452 24196 -1451
rect 24260 -1452 24270 -1383
rect 24186 -1457 24270 -1452
rect 352 -1510 518 -1502
rect 352 -1578 386 -1510
rect 470 -1578 518 -1510
rect 352 -1582 518 -1578
rect 3496 -1510 3662 -1502
rect 3496 -1578 3530 -1510
rect 3614 -1578 3662 -1510
rect 6628 -1506 6794 -1498
rect 6628 -1574 6662 -1506
rect 6746 -1574 6794 -1506
rect 6628 -1578 6794 -1574
rect 9772 -1506 9938 -1498
rect 9772 -1574 9806 -1506
rect 9890 -1574 9938 -1506
rect 9772 -1578 9938 -1574
rect 12974 -1510 13140 -1502
rect 12974 -1578 13008 -1510
rect 13092 -1578 13140 -1510
rect 3496 -1582 3662 -1578
rect 12974 -1582 13140 -1578
rect 16118 -1510 16284 -1502
rect 16118 -1578 16152 -1510
rect 16236 -1578 16284 -1510
rect 19250 -1506 19416 -1498
rect 19250 -1574 19284 -1506
rect 19368 -1574 19416 -1506
rect 19250 -1578 19416 -1574
rect 22394 -1506 22560 -1498
rect 22394 -1574 22428 -1506
rect 22512 -1574 22560 -1506
rect 22394 -1578 22560 -1574
rect 16118 -1582 16284 -1578
rect 1771 -1648 1864 -1643
rect 24103 -1648 24270 -1646
rect 1771 -1729 1781 -1648
rect 1854 -1651 24270 -1648
rect 1854 -1720 24196 -1651
rect 24260 -1720 24270 -1651
rect 1854 -1725 24270 -1720
rect 1854 -1728 24210 -1725
rect 1854 -1729 1864 -1728
rect 1771 -1734 1864 -1729
<< via3 >>
rect 372 642 472 732
rect 372 640 472 642
rect 3516 642 3616 732
rect 3516 640 3616 642
rect 6648 646 6748 736
rect 6648 644 6748 646
rect 9792 646 9892 736
rect 9792 644 9892 646
rect 12994 642 13094 732
rect 12994 640 13094 642
rect 16138 642 16238 732
rect 16138 640 16238 642
rect 19270 646 19370 736
rect 19270 644 19370 646
rect 22414 646 22514 736
rect 22414 644 22514 646
rect -1018 -361 -941 -347
rect -1018 -417 -1008 -361
rect -1008 -417 -952 -361
rect -952 -417 -941 -361
rect -1018 -430 -941 -417
rect 21013 -506 21113 -496
rect 21013 -595 21024 -506
rect 21024 -595 21103 -506
rect 21103 -595 21113 -506
rect 21013 -605 21113 -595
rect 386 -1568 392 -1510
rect 392 -1568 468 -1510
rect 468 -1568 470 -1510
rect 386 -1578 470 -1568
rect 3530 -1568 3536 -1510
rect 3536 -1568 3612 -1510
rect 3612 -1568 3614 -1510
rect 3530 -1578 3614 -1568
rect 6662 -1564 6668 -1506
rect 6668 -1564 6744 -1506
rect 6744 -1564 6746 -1506
rect 6662 -1574 6746 -1564
rect 9806 -1564 9812 -1506
rect 9812 -1564 9888 -1506
rect 9888 -1564 9890 -1506
rect 9806 -1574 9890 -1564
rect 13008 -1568 13014 -1510
rect 13014 -1568 13090 -1510
rect 13090 -1568 13092 -1510
rect 13008 -1578 13092 -1568
rect 16152 -1568 16158 -1510
rect 16158 -1568 16234 -1510
rect 16234 -1568 16236 -1510
rect 16152 -1578 16236 -1568
rect 19284 -1564 19290 -1506
rect 19290 -1564 19366 -1506
rect 19366 -1564 19368 -1506
rect 19284 -1574 19368 -1564
rect 22428 -1564 22434 -1506
rect 22434 -1564 22510 -1506
rect 22510 -1564 22512 -1506
rect 22428 -1574 22512 -1564
<< metal4 >>
rect -484 736 23446 842
rect -484 732 6648 736
rect -484 640 372 732
rect 472 640 3516 732
rect 3616 644 6648 732
rect 6748 644 9792 736
rect 9892 732 19270 736
rect 9892 644 12994 732
rect 3616 640 12994 644
rect 13094 640 16138 732
rect 16238 644 19270 732
rect 19370 644 22414 736
rect 22514 644 23446 736
rect 16238 640 23446 644
rect -484 608 23446 640
rect -1028 -347 -940 -346
rect -1028 -430 -1018 -347
rect -941 -430 -940 -347
rect -1028 -1499 -940 -430
rect 21003 -496 21124 -495
rect 21003 -605 21013 -496
rect 21113 -605 21124 -496
rect 21003 -1498 21124 -605
rect -504 -1499 22870 -1498
rect -1028 -1506 22870 -1499
rect -1028 -1510 6662 -1506
rect -1028 -1578 386 -1510
rect 470 -1578 3530 -1510
rect 3614 -1574 6662 -1510
rect 6746 -1574 9806 -1506
rect 9890 -1510 19284 -1506
rect 9890 -1574 13008 -1510
rect 3614 -1578 13008 -1574
rect 13092 -1578 16152 -1510
rect 16236 -1574 19284 -1510
rect 19368 -1574 22428 -1506
rect 22512 -1574 22870 -1506
rect 16236 -1578 22870 -1574
rect -1028 -1678 22870 -1578
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_0
timestamp 1736594632
transform 1 0 3190 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_1
timestamp 1736594632
transform 1 0 3932 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_2
timestamp 1736594632
transform 1 0 788 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_3
timestamp 1736594632
transform 1 0 46 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_4
timestamp 1736594632
transform 1 0 7064 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_5
timestamp 1736594632
transform 1 0 6322 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_6
timestamp 1736594632
transform 1 0 9466 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_7
timestamp 1736594632
transform 1 0 10208 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_8
timestamp 1736594632
transform 1 0 12668 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_9
timestamp 1736594632
transform 1 0 13410 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_10
timestamp 1736594632
transform 1 0 15812 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_11
timestamp 1736594632
transform 1 0 16554 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_12
timestamp 1736594632
transform 1 0 19686 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_13
timestamp 1736594632
transform 1 0 18944 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_14
timestamp 1736594632
transform 1 0 22830 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_15
timestamp 1736594632
transform 1 0 22088 0 1 -967
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_0
timestamp 1736594632
transform 1 0 3559 0 1 -1071
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_1
timestamp 1736594632
transform 1 0 415 0 1 -1071
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_2
timestamp 1736594632
transform 1 0 6691 0 1 -1067
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_3
timestamp 1736594632
transform 1 0 9835 0 1 -1067
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_4
timestamp 1736594632
transform 1 0 13037 0 1 -1071
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_5
timestamp 1736594632
transform 1 0 16181 0 1 -1071
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_6
timestamp 1736594632
transform 1 0 19313 0 1 -1067
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_7
timestamp 1736594632
transform 1 0 22457 0 1 -1067
box -265 -226 265 226
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_0
timestamp 1736594632
transform 1 0 3559 0 1 262
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_1
timestamp 1736594632
transform 1 0 415 0 1 262
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_2
timestamp 1736594632
transform 1 0 6691 0 1 266
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_3
timestamp 1736594632
transform 1 0 9835 0 1 266
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_4
timestamp 1736594632
transform 1 0 13037 0 1 262
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_5
timestamp 1736594632
transform 1 0 16181 0 1 262
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_6
timestamp 1736594632
transform 1 0 19313 0 1 266
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_7
timestamp 1736594632
transform 1 0 22457 0 1 266
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_0
timestamp 1736594632
transform 1 0 4209 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_1
timestamp 1736594632
transform 1 0 2915 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_2
timestamp 1736594632
transform 1 0 -229 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_3
timestamp 1736594632
transform 1 0 1065 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_4
timestamp 1736594632
transform 1 0 6047 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_5
timestamp 1736594632
transform 1 0 7341 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_6
timestamp 1736594632
transform 1 0 9191 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_7
timestamp 1736594632
transform 1 0 10485 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_8
timestamp 1736594632
transform 1 0 12393 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_9
timestamp 1736594632
transform 1 0 13687 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_10
timestamp 1736594632
transform 1 0 15537 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_11
timestamp 1736594632
transform 1 0 16831 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_12
timestamp 1736594632
transform 1 0 19963 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_13
timestamp 1736594632
transform 1 0 18669 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_14
timestamp 1736594632
transform 1 0 21813 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_15
timestamp 1736594632
transform 1 0 23107 0 1 266
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_0
timestamp 1736594632
transform 1 0 4682 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_1
timestamp 1736594632
transform 1 0 -670 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_2
timestamp 1736594632
transform 1 0 2474 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_3
timestamp 1736594632
transform 1 0 1538 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_4
timestamp 1736594632
transform 1 0 5606 0 1 166
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_5
timestamp 1736594632
transform 1 0 7814 0 1 166
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_6
timestamp 1736594632
transform 1 0 8750 0 1 166
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_7
timestamp 1736594632
transform 1 0 10958 0 1 166
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_8
timestamp 1736594632
transform 1 0 11952 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_9
timestamp 1736594632
transform 1 0 14160 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_10
timestamp 1736594632
transform 1 0 15096 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_11
timestamp 1736594632
transform 1 0 18228 0 1 166
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_12
timestamp 1736594632
transform 1 0 17304 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_13
timestamp 1736594632
transform 1 0 21372 0 1 166
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_14
timestamp 1736594632
transform 1 0 20436 0 1 166
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_15
timestamp 1736594632
transform 1 0 23580 0 1 166
box -242 -162 242 162
<< labels >>
flabel metal4 11190 624 11552 788 1 FreeSerif 960 0 0 0 VDD
port 1 n
flabel metal4 11162 -1670 11548 -1542 1 FreeSerif 960 0 0 0 VSS
port 2 n
flabel metal1 24275 -373 24351 -293 1 FreeSerif 720 0 0 0 Y[7]
port 20 n
flabel metal1 24303 -734 24345 -666 1 FreeSerif 720 0 0 0 Y[6]
port 21 n
flabel metal1 24301 -863 24346 -803 1 FreeSerif 720 0 0 0 Y[5]
port 22 n
flabel metal1 24294 -1028 24347 -959 1 FreeSerif 720 0 0 0 Y[4]
port 23 n
flabel metal1 24287 -1181 24348 -1105 1 FreeSerif 720 0 0 0 Y[3]
port 15 n
flabel metal1 24279 -1323 24354 -1240 1 FreeSerif 720 0 0 0 Y[2]
port 24 n
flabel metal1 24276 -1455 24349 -1378 1 FreeSerif 720 0 0 0 Y[1]
port 17 n
flabel metal1 24287 -1724 24343 -1657 1 FreeSerif 720 0 0 0 Y[0]
port 25 n
flabel metal1 -1266 -309 -1200 -233 1 FreeSerif 720 0 0 0 dir
port 26 n
flabel metal1 -1263 -591 -1194 -521 1 FreeSerif 720 0 0 0 A[1]
port 27 n
flabel metal1 -1261 -819 -1197 -769 1 FreeSerif 720 0 0 0 A[2]
port 5 n
flabel metal1 -1262 -955 -1200 -903 1 FreeSerif 720 0 0 0 A[3]
port 6 n
flabel metal1 -1262 -1065 -1212 -1015 1 FreeSerif 720 0 0 0 A[4]
port 7 n
flabel metal1 -1255 -1431 -1209 -1383 1 FreeSerif 720 0 0 0 A[6]
port 9 n
flabel metal1 -1265 -1194 -1209 -1138 1 FreeSerif 720 0 0 0 A[5]
port 8 n
flabel metal1 -1253 -1647 -1180 -1612 1 FreeSerif 720 0 0 0 A[7]
port 28 n
flabel metal1 -1266 -148 -1184 -94 1 FreeSerif 720 0 0 0 A[0]
port 29 n
<< end >>
