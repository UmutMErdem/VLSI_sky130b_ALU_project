magic
tech sky130B
magscale 1 2
timestamp 1736520155
<< nwell >>
rect -1146 1370 -649 1827
rect -1792 1124 1192 1370
rect -1792 803 1193 1124
rect -1365 110 -527 803
rect 1 800 1193 803
<< nmos >>
rect 332 225 392 625
rect 450 225 510 625
rect 685 425 745 625
rect -1573 -360 -1513 -160
rect -1153 -560 -1093 -160
rect -1035 -560 -975 -160
rect -917 -560 -857 -160
rect -799 -560 -739 -160
rect -275 -360 -215 -160
<< pmos >>
rect -1698 865 -1638 1065
rect -1580 865 -1520 1065
rect -1462 865 -1402 1065
rect -1214 865 -1154 1265
rect -1096 865 -1036 1265
rect -978 865 -918 1265
rect -860 865 -800 1265
rect -742 865 -682 1265
rect -624 865 -564 1265
rect -377 865 -317 1065
rect -259 865 -199 1065
rect -141 865 -81 1065
rect 95 862 155 1062
rect 213 862 273 1062
rect 331 862 391 1062
rect 449 862 509 1062
rect 567 862 627 1062
rect 685 862 745 1062
rect 803 862 863 1062
rect 921 862 981 1062
rect 1039 862 1099 1062
rect -1271 172 -1211 572
rect -1153 172 -1093 572
rect -1035 172 -975 572
rect -917 172 -857 572
rect -799 172 -739 572
rect -681 172 -621 572
<< ndiff >>
rect 274 613 332 625
rect 274 237 286 613
rect 320 237 332 613
rect 274 225 332 237
rect 392 613 450 625
rect 392 237 404 613
rect 438 237 450 613
rect 392 225 450 237
rect 510 613 568 625
rect 510 237 522 613
rect 556 237 568 613
rect 627 613 685 625
rect 627 437 639 613
rect 673 437 685 613
rect 627 425 685 437
rect 745 613 803 625
rect 745 437 757 613
rect 791 437 803 613
rect 745 425 803 437
rect 510 225 568 237
rect -1631 -172 -1573 -160
rect -1631 -348 -1619 -172
rect -1585 -348 -1573 -172
rect -1631 -360 -1573 -348
rect -1513 -172 -1455 -160
rect -1513 -348 -1501 -172
rect -1467 -348 -1455 -172
rect -1513 -360 -1455 -348
rect -1211 -172 -1153 -160
rect -1211 -548 -1199 -172
rect -1165 -548 -1153 -172
rect -1211 -560 -1153 -548
rect -1093 -172 -1035 -160
rect -1093 -548 -1081 -172
rect -1047 -548 -1035 -172
rect -1093 -560 -1035 -548
rect -975 -172 -917 -160
rect -975 -548 -963 -172
rect -929 -548 -917 -172
rect -975 -560 -917 -548
rect -857 -172 -799 -160
rect -857 -548 -845 -172
rect -811 -548 -799 -172
rect -857 -560 -799 -548
rect -739 -172 -681 -160
rect -739 -548 -727 -172
rect -693 -548 -681 -172
rect -333 -172 -275 -160
rect -333 -348 -321 -172
rect -287 -348 -275 -172
rect -333 -360 -275 -348
rect -215 -172 -157 -160
rect -215 -348 -203 -172
rect -169 -348 -157 -172
rect -215 -360 -157 -348
rect -739 -560 -681 -548
<< pdiff >>
rect -1272 1253 -1214 1265
rect -1756 1053 -1698 1065
rect -1756 877 -1744 1053
rect -1710 877 -1698 1053
rect -1756 865 -1698 877
rect -1638 1053 -1580 1065
rect -1638 877 -1626 1053
rect -1592 877 -1580 1053
rect -1638 865 -1580 877
rect -1520 1053 -1462 1065
rect -1520 877 -1508 1053
rect -1474 877 -1462 1053
rect -1520 865 -1462 877
rect -1402 1053 -1344 1065
rect -1402 877 -1390 1053
rect -1356 877 -1344 1053
rect -1402 865 -1344 877
rect -1272 877 -1260 1253
rect -1226 877 -1214 1253
rect -1272 865 -1214 877
rect -1154 1253 -1096 1265
rect -1154 877 -1142 1253
rect -1108 877 -1096 1253
rect -1154 865 -1096 877
rect -1036 1253 -978 1265
rect -1036 877 -1024 1253
rect -990 877 -978 1253
rect -1036 865 -978 877
rect -918 1253 -860 1265
rect -918 877 -906 1253
rect -872 877 -860 1253
rect -918 865 -860 877
rect -800 1253 -742 1265
rect -800 877 -788 1253
rect -754 877 -742 1253
rect -800 865 -742 877
rect -682 1253 -624 1265
rect -682 877 -670 1253
rect -636 877 -624 1253
rect -682 865 -624 877
rect -564 1253 -506 1265
rect -564 877 -552 1253
rect -518 877 -506 1253
rect -564 865 -506 877
rect -435 1053 -377 1065
rect -435 877 -423 1053
rect -389 877 -377 1053
rect -435 865 -377 877
rect -317 1053 -259 1065
rect -317 877 -305 1053
rect -271 877 -259 1053
rect -317 865 -259 877
rect -199 1053 -141 1065
rect -199 877 -187 1053
rect -153 877 -141 1053
rect -199 865 -141 877
rect -81 1053 -23 1065
rect -81 877 -69 1053
rect -35 877 -23 1053
rect -81 865 -23 877
rect 37 1050 95 1062
rect 37 874 49 1050
rect 83 874 95 1050
rect 37 862 95 874
rect 155 1050 213 1062
rect 155 874 167 1050
rect 201 874 213 1050
rect 155 862 213 874
rect 273 1050 331 1062
rect 273 874 285 1050
rect 319 874 331 1050
rect 273 862 331 874
rect 391 1050 449 1062
rect 391 874 403 1050
rect 437 874 449 1050
rect 391 862 449 874
rect 509 1050 567 1062
rect 509 874 521 1050
rect 555 874 567 1050
rect 509 862 567 874
rect 627 1050 685 1062
rect 627 874 639 1050
rect 673 874 685 1050
rect 627 862 685 874
rect 745 1050 803 1062
rect 745 874 757 1050
rect 791 874 803 1050
rect 745 862 803 874
rect 863 1050 921 1062
rect 863 874 875 1050
rect 909 874 921 1050
rect 863 862 921 874
rect 981 1050 1039 1062
rect 981 874 993 1050
rect 1027 874 1039 1050
rect 981 862 1039 874
rect 1099 1050 1157 1062
rect 1099 874 1111 1050
rect 1145 874 1157 1050
rect 1099 862 1157 874
rect -1329 560 -1271 572
rect -1329 184 -1317 560
rect -1283 184 -1271 560
rect -1329 172 -1271 184
rect -1211 560 -1153 572
rect -1211 184 -1199 560
rect -1165 184 -1153 560
rect -1211 172 -1153 184
rect -1093 560 -1035 572
rect -1093 184 -1081 560
rect -1047 184 -1035 560
rect -1093 172 -1035 184
rect -975 560 -917 572
rect -975 184 -963 560
rect -929 184 -917 560
rect -975 172 -917 184
rect -857 560 -799 572
rect -857 184 -845 560
rect -811 184 -799 560
rect -857 172 -799 184
rect -739 560 -681 572
rect -739 184 -727 560
rect -693 184 -681 560
rect -739 172 -681 184
rect -621 560 -563 572
rect -621 184 -609 560
rect -575 184 -563 560
rect -621 172 -563 184
<< ndiffc >>
rect 286 237 320 613
rect 404 237 438 613
rect 522 237 556 613
rect 639 437 673 613
rect 757 437 791 613
rect -1619 -348 -1585 -172
rect -1501 -348 -1467 -172
rect -1199 -548 -1165 -172
rect -1081 -548 -1047 -172
rect -963 -548 -929 -172
rect -845 -548 -811 -172
rect -727 -548 -693 -172
rect -321 -348 -287 -172
rect -203 -348 -169 -172
<< pdiffc >>
rect -1744 877 -1710 1053
rect -1626 877 -1592 1053
rect -1508 877 -1474 1053
rect -1390 877 -1356 1053
rect -1260 877 -1226 1253
rect -1142 877 -1108 1253
rect -1024 877 -990 1253
rect -906 877 -872 1253
rect -788 877 -754 1253
rect -670 877 -636 1253
rect -552 877 -518 1253
rect -423 877 -389 1053
rect -305 877 -271 1053
rect -187 877 -153 1053
rect -69 877 -35 1053
rect 49 874 83 1050
rect 167 874 201 1050
rect 285 874 319 1050
rect 403 874 437 1050
rect 521 874 555 1050
rect 639 874 673 1050
rect 757 874 791 1050
rect 875 874 909 1050
rect 993 874 1027 1050
rect 1111 874 1145 1050
rect -1317 184 -1283 560
rect -1199 184 -1165 560
rect -1081 184 -1047 560
rect -963 184 -929 560
rect -845 184 -811 560
rect -727 184 -693 560
rect -609 184 -575 560
<< psubdiff >>
rect 538 82 750 112
rect 538 26 578 82
rect 712 26 750 82
rect 538 4 750 26
rect -1052 -719 -810 -707
rect -1052 -821 -1005 -719
rect -870 -821 -810 -719
rect -1052 -838 -810 -821
<< nsubdiff >>
rect -1110 1757 -689 1791
rect -1110 1612 -1047 1757
rect -738 1612 -689 1757
rect -1110 1591 -689 1612
rect 298 1290 542 1328
rect 298 1220 354 1290
rect 490 1220 542 1290
rect 298 1198 542 1220
<< psubdiffcont >>
rect 578 26 712 82
rect -1005 -821 -870 -719
<< nsubdiffcont >>
rect -1047 1612 -738 1757
rect 354 1220 490 1290
<< poly >>
rect -1214 1280 -918 1331
rect -1214 1265 -1154 1280
rect -1096 1265 -1036 1280
rect -978 1265 -918 1280
rect -860 1265 -800 1291
rect -742 1265 -682 1291
rect -624 1265 -564 1291
rect -1698 1065 -1638 1091
rect -1580 1065 -1520 1091
rect -1462 1065 -1402 1091
rect -377 1082 -81 1133
rect -377 1065 -317 1082
rect -259 1065 -199 1082
rect -141 1065 -81 1082
rect 95 1083 391 1119
rect 95 1062 155 1083
rect 213 1062 273 1083
rect 331 1062 391 1083
rect 449 1082 745 1118
rect 449 1062 509 1082
rect 567 1062 627 1082
rect 685 1062 745 1082
rect 803 1082 1099 1118
rect 803 1062 863 1082
rect 921 1062 981 1082
rect 1039 1062 1099 1082
rect -1698 848 -1638 865
rect -1580 848 -1520 865
rect -1462 848 -1402 865
rect -1214 848 -1154 865
rect -1698 797 -1154 848
rect -1096 839 -1036 865
rect -978 839 -918 865
rect -860 846 -800 865
rect -742 846 -682 865
rect -624 846 -564 865
rect -377 846 -317 865
rect -259 846 -199 865
rect -1573 593 -1513 797
rect -860 795 -317 846
rect -275 839 -199 846
rect -141 839 -81 865
rect -275 795 -200 839
rect 95 836 155 862
rect 213 836 273 862
rect 331 836 391 862
rect 449 842 509 862
rect 449 836 510 842
rect 567 836 627 862
rect 685 836 745 862
rect -275 713 -215 795
rect -275 695 -41 713
rect -275 661 -92 695
rect -58 661 -41 695
rect -1271 595 -975 655
rect -1573 576 -1442 593
rect -1573 542 -1492 576
rect -1458 542 -1442 576
rect -1271 572 -1211 595
rect -1153 572 -1093 595
rect -1035 572 -975 595
rect -917 596 -621 656
rect -917 572 -857 596
rect -799 572 -739 596
rect -681 572 -621 596
rect -275 645 -41 661
rect 332 651 390 836
rect -1573 525 -1442 542
rect -1573 -55 -1513 525
rect -1271 146 -1211 172
rect -1303 5 -1236 12
rect -1153 5 -1093 172
rect -1035 146 -975 172
rect -917 146 -857 172
rect -1303 -4 -1093 5
rect -1303 -38 -1287 -4
rect -1253 -38 -1093 -4
rect -1303 -54 -1093 -38
rect -1573 -71 -1422 -55
rect -1573 -105 -1472 -71
rect -1438 -105 -1422 -71
rect -1573 -121 -1422 -105
rect -1573 -160 -1513 -121
rect -1153 -160 -1093 -54
rect -799 5 -739 172
rect -681 146 -621 172
rect -656 5 -589 12
rect -799 -4 -589 5
rect -799 -38 -639 -4
rect -605 -38 -589 -4
rect -799 -54 -589 -38
rect -1037 -88 -971 -72
rect -1037 -122 -1021 -88
rect -987 -122 -971 -88
rect -1037 -138 -971 -122
rect -919 -87 -853 -72
rect -919 -121 -903 -87
rect -869 -121 -853 -87
rect -919 -137 -853 -121
rect -1035 -160 -975 -138
rect -917 -160 -857 -137
rect -799 -160 -739 -54
rect -275 -56 -215 645
rect 332 625 392 651
rect 450 625 510 836
rect 803 830 863 862
rect 921 836 981 862
rect 1039 836 1099 862
rect 800 814 866 830
rect 800 780 816 814
rect 850 780 866 814
rect 800 764 866 780
rect 682 697 748 713
rect 682 663 698 697
rect 732 663 748 697
rect 682 647 748 663
rect 685 625 745 647
rect 685 399 745 425
rect 332 203 392 225
rect 450 203 510 225
rect 329 187 395 203
rect 329 153 345 187
rect 379 153 395 187
rect 329 137 395 153
rect 447 187 513 203
rect 447 153 463 187
rect 497 153 513 187
rect 447 137 513 153
rect -365 -72 -215 -56
rect -365 -106 -349 -72
rect -315 -106 -215 -72
rect -365 -122 -215 -106
rect -275 -160 -215 -122
rect -1573 -386 -1513 -360
rect -275 -386 -215 -360
rect -1153 -586 -1093 -560
rect -1035 -586 -975 -560
rect -917 -586 -857 -560
rect -799 -586 -739 -560
<< polycont >>
rect -92 661 -58 695
rect -1492 542 -1458 576
rect -1287 -38 -1253 -4
rect -1472 -105 -1438 -71
rect -639 -38 -605 -4
rect -1021 -122 -987 -88
rect -903 -121 -869 -87
rect 816 780 850 814
rect 698 663 732 697
rect 345 153 379 187
rect 463 153 497 187
rect -349 -106 -315 -72
<< locali >>
rect -1121 1791 -677 1797
rect -1121 1591 -1110 1791
rect -689 1591 -677 1791
rect -1121 1585 -677 1591
rect -906 1306 -636 1341
rect -1260 1253 -1226 1269
rect -1744 1107 -1474 1142
rect -1744 1053 -1710 1107
rect -1744 861 -1710 877
rect -1626 1053 -1592 1069
rect -1626 861 -1592 877
rect -1508 1053 -1474 1107
rect -1508 861 -1474 877
rect -1390 1053 -1356 1069
rect -1390 861 -1356 877
rect -1260 861 -1226 877
rect -1142 1253 -1108 1269
rect -1142 861 -1108 877
rect -1024 1253 -990 1269
rect -1024 861 -990 877
rect -906 1253 -872 1306
rect -906 861 -872 877
rect -788 1253 -754 1269
rect -788 861 -754 877
rect -670 1253 -636 1306
rect 338 1290 506 1306
rect -670 861 -636 877
rect -552 1253 -518 1269
rect 338 1220 354 1290
rect 490 1220 506 1290
rect 338 1204 506 1220
rect 875 1100 1145 1134
rect -552 861 -518 877
rect -423 1053 -389 1069
rect -423 861 -389 877
rect -305 1053 -271 1069
rect -305 861 -271 877
rect -187 1053 -153 1069
rect -187 861 -153 877
rect -69 1053 -35 1069
rect -69 861 -35 877
rect 49 1050 83 1066
rect 49 858 83 874
rect 167 1050 201 1066
rect 167 858 201 874
rect 285 1050 319 1066
rect 285 858 319 874
rect 403 1050 437 1066
rect 403 858 437 874
rect 521 1050 555 1066
rect 521 858 555 874
rect 639 1050 673 1066
rect 639 858 673 874
rect 757 1050 791 1066
rect 757 858 791 874
rect 875 1050 909 1100
rect 875 858 909 874
rect 993 1050 1027 1066
rect 993 858 1027 874
rect 1111 1050 1145 1100
rect 1111 858 1145 874
rect 800 780 816 814
rect 850 780 866 814
rect -92 695 -58 711
rect 682 663 698 697
rect 732 663 748 697
rect -92 645 -58 661
rect 286 613 320 629
rect -1498 576 -1442 593
rect -1498 542 -1492 576
rect -1458 542 -1442 576
rect -1498 525 -1442 542
rect -1317 560 -1283 576
rect -1199 560 -1165 576
rect -1317 168 -1283 184
rect -1200 184 -1199 231
rect -1081 560 -1047 576
rect -1165 184 -1164 231
rect -1200 126 -1164 184
rect -963 560 -929 576
rect -1081 168 -1047 184
rect -965 184 -963 231
rect -965 126 -929 184
rect -845 560 -811 576
rect -845 168 -811 184
rect -727 560 -693 576
rect -609 560 -575 576
rect -693 184 -691 230
rect -727 126 -691 184
rect -447 355 -377 359
rect -447 264 -443 355
rect -381 264 -377 355
rect -447 259 -377 264
rect -609 168 -575 184
rect -432 126 -391 259
rect 286 221 320 237
rect 404 613 438 629
rect 404 221 438 237
rect 522 613 556 629
rect 639 613 673 629
rect 639 421 673 437
rect 757 613 791 629
rect 757 421 791 437
rect 522 221 556 237
rect 329 153 345 187
rect 379 153 395 187
rect 447 153 463 187
rect 497 153 513 187
rect -1200 86 -391 126
rect -1181 85 -391 86
rect -1303 -4 -1236 12
rect -1303 -38 -1287 -4
rect -1253 -38 -1236 -4
rect -1303 -54 -1236 -38
rect -1472 -71 -1438 -55
rect -1472 -121 -1438 -105
rect -1126 -156 -1092 85
rect 562 82 730 100
rect 562 26 578 82
rect 712 26 730 82
rect -656 -4 -589 12
rect 562 10 730 26
rect -656 -38 -639 -4
rect -605 -38 -589 -4
rect -656 -54 -589 -38
rect -349 -72 -315 -56
rect -1037 -122 -1021 -88
rect -987 -122 -971 -88
rect -919 -121 -903 -87
rect -869 -121 -853 -87
rect -349 -122 -315 -106
rect -1619 -172 -1585 -156
rect -1619 -364 -1585 -348
rect -1501 -172 -1467 -156
rect -1501 -364 -1467 -348
rect -1199 -172 -1165 -156
rect -1126 -172 -1047 -156
rect -1126 -202 -1081 -172
rect -1199 -615 -1164 -548
rect -1081 -564 -1047 -548
rect -963 -172 -929 -156
rect -963 -564 -929 -548
rect -845 -172 -811 -156
rect -727 -172 -693 -156
rect -321 -172 -287 -156
rect -321 -364 -287 -348
rect -203 -172 -169 -156
rect -203 -364 -169 -348
rect -845 -564 -811 -548
rect -728 -615 -693 -548
rect -1199 -650 -693 -615
rect -1052 -719 -810 -707
rect -1052 -821 -1005 -719
rect -870 -821 -810 -719
rect -1052 -838 -810 -821
<< viali >>
rect -1110 1757 -689 1791
rect -1110 1612 -1047 1757
rect -1047 1612 -738 1757
rect -738 1612 -689 1757
rect -1110 1591 -689 1612
rect -1744 877 -1710 1053
rect -1626 877 -1592 1053
rect -1508 877 -1474 1053
rect -1390 877 -1356 1053
rect -1260 877 -1226 1253
rect -1142 877 -1108 1253
rect -1024 877 -990 1253
rect -906 877 -872 1253
rect -788 877 -754 1253
rect -670 877 -636 1253
rect -552 877 -518 1253
rect 390 1226 450 1288
rect -423 877 -389 1053
rect -305 877 -271 1053
rect -187 877 -153 1053
rect -69 877 -35 1053
rect 49 874 83 1050
rect 167 874 201 1050
rect 285 874 319 1050
rect 403 874 437 1050
rect 521 874 555 1050
rect 639 874 673 1050
rect 757 874 791 1050
rect 875 874 909 1050
rect 993 874 1027 1050
rect 1111 874 1145 1050
rect 816 780 850 814
rect -92 661 -58 695
rect 698 663 732 697
rect -1492 542 -1458 576
rect -1317 184 -1283 560
rect -1199 184 -1165 560
rect -1081 184 -1047 560
rect -963 184 -929 560
rect -845 184 -811 560
rect -727 184 -693 560
rect -609 184 -575 560
rect -443 264 -381 355
rect 286 237 320 613
rect 404 237 438 613
rect 522 237 556 613
rect 639 437 673 613
rect 757 437 791 613
rect 345 153 379 187
rect 463 153 497 187
rect -1287 -38 -1253 -4
rect -1472 -105 -1438 -71
rect 618 30 670 76
rect -639 -38 -605 -4
rect -1021 -122 -987 -88
rect -903 -121 -869 -87
rect -349 -106 -315 -72
rect -1619 -348 -1585 -172
rect -1501 -348 -1467 -172
rect -1199 -548 -1165 -172
rect -1081 -548 -1047 -172
rect -963 -548 -929 -172
rect -845 -548 -811 -172
rect -727 -548 -693 -172
rect -321 -348 -287 -172
rect -203 -348 -169 -172
rect -1005 -821 -870 -719
<< metal1 >>
rect -1122 1791 -677 1797
rect -1122 1591 -1110 1791
rect -689 1591 -677 1791
rect -1122 1585 -954 1591
rect -964 1517 -954 1585
rect -822 1585 -677 1591
rect -822 1517 -812 1585
rect -954 1477 -822 1517
rect -955 1411 -822 1477
rect -1626 1368 -153 1411
rect -1626 1065 -1592 1368
rect -1260 1265 -1226 1368
rect -1024 1265 -990 1368
rect -788 1265 -754 1368
rect -552 1265 -518 1368
rect -1266 1253 -1220 1265
rect -1750 1053 -1704 1065
rect -1750 877 -1744 1053
rect -1710 877 -1704 1053
rect -1750 865 -1704 877
rect -1632 1053 -1586 1065
rect -1632 877 -1626 1053
rect -1592 877 -1586 1053
rect -1632 865 -1586 877
rect -1514 1053 -1468 1065
rect -1514 877 -1508 1053
rect -1474 877 -1468 1053
rect -1514 865 -1468 877
rect -1396 1053 -1350 1065
rect -1266 1053 -1260 1253
rect -1396 877 -1390 1053
rect -1356 877 -1260 1053
rect -1226 877 -1220 1253
rect -1396 865 -1350 877
rect -1266 865 -1220 877
rect -1148 1253 -1102 1265
rect -1148 877 -1142 1253
rect -1108 877 -1102 1253
rect -1148 865 -1102 877
rect -1030 1253 -984 1265
rect -1030 877 -1024 1253
rect -990 877 -984 1253
rect -1030 865 -984 877
rect -912 1253 -866 1265
rect -912 877 -906 1253
rect -872 877 -866 1253
rect -912 865 -866 877
rect -794 1253 -748 1265
rect -794 877 -788 1253
rect -754 877 -748 1253
rect -794 865 -748 877
rect -676 1253 -630 1265
rect -676 877 -670 1253
rect -636 877 -630 1253
rect -676 865 -630 877
rect -558 1253 -512 1265
rect -558 877 -552 1253
rect -518 1053 -512 1253
rect -187 1065 -153 1368
rect 354 1288 490 1308
rect 354 1226 390 1288
rect 450 1226 490 1288
rect 354 1198 490 1226
rect 50 1168 1027 1198
rect -429 1053 -383 1065
rect -518 877 -423 1053
rect -389 877 -383 1053
rect -558 865 -512 877
rect -429 865 -383 877
rect -311 1053 -265 1065
rect -311 877 -305 1053
rect -271 877 -265 1053
rect -311 865 -265 877
rect -193 1053 -147 1065
rect -193 877 -187 1053
rect -153 877 -147 1053
rect -193 865 -147 877
rect -75 1053 -29 1065
rect 50 1062 82 1168
rect 286 1062 318 1168
rect 522 1062 554 1168
rect 758 1062 790 1168
rect 993 1062 1027 1168
rect -75 877 -69 1053
rect -35 877 -29 1053
rect -75 865 -29 877
rect 43 1050 89 1062
rect 43 874 49 1050
rect 83 874 89 1050
rect -1744 831 -1710 865
rect -1142 831 -1108 865
rect -906 831 -872 865
rect -1744 796 -1585 831
rect -1142 796 -872 831
rect -305 831 -271 865
rect -69 831 -35 865
rect 43 862 89 874
rect 161 1050 207 1062
rect 161 874 167 1050
rect 201 874 207 1050
rect 161 862 207 874
rect 279 1050 325 1062
rect 279 874 285 1050
rect 319 874 325 1050
rect 279 862 325 874
rect 397 1050 443 1062
rect 397 874 403 1050
rect 437 874 443 1050
rect 397 862 443 874
rect 515 1050 561 1062
rect 515 874 521 1050
rect 555 874 561 1050
rect 515 862 561 874
rect 633 1050 679 1062
rect 633 874 639 1050
rect 673 874 679 1050
rect 633 862 679 874
rect 751 1050 797 1062
rect 751 874 757 1050
rect 791 874 797 1050
rect 751 862 797 874
rect 869 1050 915 1062
rect 869 874 875 1050
rect 909 874 915 1050
rect 869 862 915 874
rect 987 1050 1033 1062
rect 987 874 993 1050
rect 1027 874 1033 1050
rect 987 862 1033 874
rect 1105 1050 1151 1062
rect 1105 874 1111 1050
rect 1145 874 1151 1050
rect 1105 862 1151 874
rect -305 796 -35 831
rect -1792 648 -1757 711
rect -1690 648 -1680 711
rect -1792 522 -1757 585
rect -1690 522 -1680 585
rect -1619 12 -1585 796
rect -906 734 -872 796
rect -1317 696 -575 734
rect -1507 525 -1497 593
rect -1442 525 -1432 593
rect -1317 572 -1283 696
rect -1081 572 -1047 696
rect -845 572 -811 696
rect -609 572 -575 696
rect -1323 560 -1277 572
rect -1323 184 -1317 560
rect -1283 184 -1277 560
rect -1323 172 -1277 184
rect -1205 560 -1159 572
rect -1205 184 -1199 560
rect -1165 184 -1159 560
rect -1205 172 -1159 184
rect -1087 560 -1041 572
rect -1087 184 -1081 560
rect -1047 184 -1041 560
rect -1087 172 -1041 184
rect -969 560 -923 572
rect -969 184 -963 560
rect -929 184 -923 560
rect -969 172 -923 184
rect -851 560 -805 572
rect -851 184 -845 560
rect -811 184 -805 560
rect -851 172 -805 184
rect -733 560 -687 572
rect -733 184 -727 560
rect -693 184 -687 560
rect -733 172 -687 184
rect -615 560 -569 572
rect -615 184 -609 560
rect -575 184 -569 560
rect -449 355 -375 367
rect -453 264 -443 355
rect -381 264 -371 355
rect -449 252 -375 264
rect -615 172 -569 184
rect -203 13 -169 796
rect 166 768 202 862
rect 402 768 438 862
rect 638 769 674 862
rect 800 814 866 821
rect 800 780 816 814
rect 850 780 866 814
rect 800 769 866 780
rect 638 768 866 769
rect 166 739 866 768
rect 166 738 748 739
rect -108 706 -32 711
rect -111 650 -101 706
rect -48 705 -32 706
rect -48 650 218 705
rect -108 645 218 650
rect 13 603 104 608
rect 13 514 23 603
rect 96 514 104 603
rect 13 502 104 514
rect 50 108 104 502
rect 164 193 218 645
rect 286 625 320 738
rect 682 697 748 738
rect 682 663 698 697
rect 732 663 748 697
rect 682 656 748 663
rect 1110 629 1145 862
rect 756 625 1145 629
rect 280 613 326 625
rect 280 237 286 613
rect 320 237 326 613
rect 280 225 326 237
rect 398 613 444 625
rect 398 237 404 613
rect 438 237 444 613
rect 398 225 444 237
rect 516 613 562 625
rect 516 237 522 613
rect 556 264 562 613
rect 633 613 679 625
rect 633 437 639 613
rect 673 437 679 613
rect 633 430 679 437
rect 751 613 1145 625
rect 751 437 757 613
rect 791 600 1145 613
rect 791 437 797 600
rect 970 511 1145 600
rect 633 425 682 430
rect 751 425 797 437
rect 639 264 682 425
rect 556 237 682 264
rect 905 262 915 353
rect 1048 262 1146 353
rect 516 225 682 237
rect 522 221 682 225
rect 164 187 395 193
rect 164 153 345 187
rect 379 153 395 187
rect 164 137 395 153
rect 447 187 513 193
rect 447 153 463 187
rect 497 153 513 187
rect 447 108 513 153
rect 50 100 513 108
rect 50 68 514 100
rect 606 84 682 221
rect 602 24 612 84
rect 674 24 684 84
rect -476 12 -169 13
rect -1619 7 -1303 12
rect -589 7 -169 12
rect -1619 -4 -1236 7
rect -1619 -31 -1287 -4
rect -1619 -160 -1585 -31
rect -1303 -38 -1287 -31
rect -1253 -38 -1236 -4
rect -1303 -44 -1236 -38
rect -656 -4 -169 7
rect 610 -2 680 24
rect -656 -38 -639 -4
rect -605 -31 -169 -4
rect -605 -38 -589 -31
rect -476 -32 -169 -31
rect -656 -44 -589 -38
rect -1478 -71 -1422 -59
rect -1478 -105 -1472 -71
rect -1438 -72 -1422 -71
rect -365 -72 -309 -60
rect -1438 -88 -971 -72
rect -1438 -105 -1021 -88
rect -1478 -121 -1021 -105
rect -1037 -122 -1021 -121
rect -987 -122 -971 -88
rect -1037 -129 -971 -122
rect -919 -87 -349 -72
rect -919 -121 -903 -87
rect -869 -106 -349 -87
rect -315 -106 -309 -72
rect -869 -121 -309 -106
rect -919 -131 -852 -121
rect -365 -122 -309 -121
rect -203 -160 -169 -32
rect -1625 -172 -1579 -160
rect -1625 -348 -1619 -172
rect -1585 -348 -1579 -172
rect -1625 -360 -1579 -348
rect -1507 -172 -1461 -160
rect -1507 -348 -1501 -172
rect -1467 -348 -1461 -172
rect -1507 -360 -1461 -348
rect -1205 -172 -1159 -160
rect -1502 -654 -1468 -360
rect -1205 -548 -1199 -172
rect -1165 -548 -1159 -172
rect -1205 -560 -1159 -548
rect -1087 -172 -1041 -160
rect -1087 -548 -1081 -172
rect -1047 -548 -1041 -172
rect -1087 -560 -1041 -548
rect -969 -172 -923 -160
rect -969 -548 -963 -172
rect -929 -548 -923 -172
rect -969 -560 -923 -548
rect -851 -172 -805 -160
rect -851 -548 -845 -172
rect -811 -548 -805 -172
rect -851 -560 -805 -548
rect -733 -172 -687 -160
rect -733 -548 -727 -172
rect -693 -548 -687 -172
rect -327 -172 -281 -160
rect -327 -348 -321 -172
rect -287 -348 -281 -172
rect -327 -360 -281 -348
rect -209 -172 -163 -160
rect -209 -348 -203 -172
rect -169 -348 -163 -172
rect -209 -360 -163 -348
rect -733 -560 -687 -548
rect -845 -654 -811 -560
rect -321 -654 -288 -360
rect -1502 -686 -288 -654
rect -1136 -710 -730 -686
rect -1136 -833 -1024 -710
rect -850 -833 -730 -710
rect -1136 -877 -730 -833
<< via1 >>
rect -954 1591 -822 1625
rect -954 1517 -822 1591
rect 390 1226 450 1288
rect -1757 648 -1690 711
rect -1757 522 -1690 585
rect -1497 576 -1442 593
rect -1497 542 -1492 576
rect -1492 542 -1458 576
rect -1458 542 -1442 576
rect -1497 525 -1442 542
rect -443 264 -381 355
rect -101 695 -48 706
rect -101 661 -92 695
rect -92 661 -58 695
rect -58 661 -48 695
rect -101 650 -48 661
rect 23 514 96 603
rect 915 262 1048 353
rect 612 76 674 84
rect 612 30 618 76
rect 618 30 670 76
rect 670 30 674 76
rect 612 24 674 30
rect -1024 -719 -850 -710
rect -1024 -821 -1005 -719
rect -1005 -821 -870 -719
rect -870 -821 -850 -719
rect -1024 -833 -850 -821
<< metal2 >>
rect -965 1636 -812 1646
rect -965 1497 -812 1507
rect 390 1288 450 1298
rect 390 1216 450 1226
rect -1757 716 -1690 721
rect -1764 711 -48 716
rect -1764 648 -1757 711
rect -1690 706 -48 711
rect -1690 650 -101 706
rect -1690 648 -48 650
rect -1764 640 -48 648
rect -1757 638 -1690 640
rect 23 603 96 613
rect -1757 594 -1690 595
rect -1497 594 23 603
rect -1765 593 23 594
rect -1765 585 -1497 593
rect -1765 522 -1757 585
rect -1690 525 -1497 585
rect -1442 525 23 593
rect -1690 522 23 525
rect -1765 515 23 522
rect -1764 514 -1675 515
rect -1757 512 -1690 514
rect 23 504 96 514
rect -443 355 1048 365
rect -381 353 1048 355
rect -381 264 915 353
rect -443 262 915 264
rect -443 254 1048 262
rect 915 252 1048 254
rect 612 92 674 94
rect 612 84 676 92
rect 674 82 676 84
rect 612 10 676 20
rect -1043 -694 -832 -684
rect -1043 -861 -832 -851
<< via2 >>
rect -965 1625 -812 1636
rect -965 1517 -954 1625
rect -954 1517 -822 1625
rect -822 1517 -812 1625
rect -965 1507 -812 1517
rect 390 1226 450 1288
rect 612 24 674 82
rect 674 24 676 82
rect 612 20 676 24
rect -1043 -710 -832 -694
rect -1043 -833 -1024 -710
rect -1024 -833 -850 -710
rect -850 -833 -832 -710
rect -1043 -851 -832 -833
<< metal3 >>
rect -997 1488 -987 1667
rect -788 1488 -778 1667
rect 374 1292 472 1310
rect 374 1220 384 1292
rect 454 1220 472 1292
rect 374 1212 472 1220
rect 469 -2 479 114
rect 817 -2 827 114
rect -1076 -873 -1066 -678
rect -800 -873 -790 -678
<< via3 >>
rect -987 1636 -788 1667
rect -987 1507 -965 1636
rect -965 1507 -812 1636
rect -812 1507 -788 1636
rect -987 1488 -788 1507
rect 384 1288 454 1292
rect 384 1226 390 1288
rect 390 1226 450 1288
rect 450 1226 454 1288
rect 384 1220 454 1226
rect 479 82 817 114
rect 479 20 612 82
rect 612 20 676 82
rect 676 20 817 82
rect 479 -2 817 20
rect -1066 -694 -800 -678
rect -1066 -851 -1043 -694
rect -1043 -851 -832 -694
rect -832 -851 -800 -694
rect -1066 -873 -800 -851
<< metal4 >>
rect -720 1816 418 1818
rect -720 1815 610 1816
rect -1129 1667 610 1815
rect -1129 1573 -987 1667
rect -1009 1488 -987 1573
rect -788 1574 610 1667
rect -788 1573 -660 1574
rect -788 1488 -764 1573
rect -1009 1485 -764 1488
rect 224 1292 610 1574
rect 224 1251 384 1292
rect 226 1220 384 1251
rect 454 1251 610 1292
rect 454 1220 608 1251
rect 226 1198 608 1220
rect 478 115 534 116
rect 474 114 534 115
rect 771 115 810 116
rect 771 114 825 115
rect 474 -2 479 114
rect 817 -2 825 114
rect 474 -143 534 -2
rect 771 -143 825 -2
<< via4 >>
rect 534 114 771 173
rect 534 -2 771 114
rect 534 -284 771 -2
rect -1129 -678 -756 -676
rect -1129 -873 -1066 -678
rect -1066 -873 -800 -678
rect -800 -873 -756 -678
rect -1129 -1015 -756 -873
<< metal5 >>
rect 472 173 829 200
rect 472 -284 534 173
rect 771 -284 829 173
rect -1201 -676 -553 -652
rect -1201 -773 -1129 -676
rect -1202 -1015 -1129 -773
rect -756 -773 -553 -676
rect 472 -773 829 -284
rect -756 -1008 829 -773
rect -756 -1015 826 -1008
rect -1202 -1094 826 -1015
<< labels >>
flabel metal1 -1785 655 -1685 704 1 FreeSans 400 0 0 0 A
port 3 n
flabel metal1 -1785 529 -1685 578 1 FreeSans 400 0 0 0 B
port 4 n
flabel metal5 -399 -936 220 -810 1 FreeSans 1040 0 0 0 VSS
port 7 n
flabel metal1 993 268 1097 346 1 FreeSans 400 0 0 0 Y
port 6 n
flabel metal1 980 519 1135 615 1 FreeSans 400 0 0 0 carry_out
port 5 n
flabel metal4 -381 1609 222 1769 1 FreeSans 1040 0 0 0 VDD
port 1 n
<< end >>
