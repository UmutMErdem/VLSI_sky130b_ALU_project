magic
tech sky130B
timestamp 1736004884
<< nwell >>
rect 0 121 242 274
rect 369 120 611 273
rect 738 120 980 273
rect 1109 120 1351 273
rect 1479 120 1721 273
rect 1848 120 2090 273
rect 2217 120 2459 273
rect 2586 120 2828 273
<< psubdiff >>
rect 22 -214 152 -191
rect 22 -249 53 -214
rect 125 -249 152 -214
rect 22 -266 152 -249
rect 391 -215 521 -192
rect 391 -250 422 -215
rect 494 -250 521 -215
rect 391 -267 521 -250
rect 760 -215 890 -192
rect 760 -250 791 -215
rect 863 -250 890 -215
rect 760 -267 890 -250
rect 1131 -215 1261 -192
rect 1131 -250 1162 -215
rect 1234 -250 1261 -215
rect 1131 -267 1261 -250
rect 1501 -215 1631 -192
rect 1501 -250 1532 -215
rect 1604 -250 1631 -215
rect 1501 -267 1631 -250
rect 1870 -215 2000 -192
rect 1870 -250 1901 -215
rect 1973 -250 2000 -215
rect 1870 -267 2000 -250
rect 2239 -215 2369 -192
rect 2239 -250 2270 -215
rect 2342 -250 2369 -215
rect 2239 -267 2369 -250
rect 2608 -215 2738 -192
rect 2608 -250 2639 -215
rect 2711 -250 2738 -215
rect 2608 -267 2738 -250
<< nsubdiff >>
rect 47 226 195 233
rect 47 195 86 226
rect 156 195 195 226
rect 47 167 195 195
rect 416 225 564 232
rect 416 194 455 225
rect 525 194 564 225
rect 416 166 564 194
rect 785 225 933 232
rect 785 194 824 225
rect 894 194 933 225
rect 785 166 933 194
rect 1156 225 1304 232
rect 1156 194 1195 225
rect 1265 194 1304 225
rect 1156 166 1304 194
rect 1526 225 1674 232
rect 1526 194 1565 225
rect 1635 194 1674 225
rect 1526 166 1674 194
rect 1895 225 2043 232
rect 1895 194 1934 225
rect 2004 194 2043 225
rect 1895 166 2043 194
rect 2264 225 2412 232
rect 2264 194 2303 225
rect 2373 194 2412 225
rect 2264 166 2412 194
rect 2633 225 2781 232
rect 2633 194 2672 225
rect 2742 194 2781 225
rect 2633 166 2781 194
<< psubdiffcont >>
rect 53 -249 125 -214
rect 422 -250 494 -215
rect 791 -250 863 -215
rect 1162 -250 1234 -215
rect 1532 -250 1604 -215
rect 1901 -250 1973 -215
rect 2270 -250 2342 -215
rect 2639 -250 2711 -215
<< nsubdiffcont >>
rect 86 195 156 226
rect 455 194 525 225
rect 824 194 894 225
rect 1195 194 1265 225
rect 1565 194 1635 225
rect 1934 194 2004 225
rect 2303 194 2373 225
rect 2672 194 2742 225
<< poly >>
rect 47 3 195 21
rect 106 -18 136 3
rect 416 2 564 20
rect 785 2 933 20
rect 1156 2 1304 20
rect 1526 2 1674 20
rect 1895 2 2043 20
rect 2264 2 2412 20
rect 2633 2 2781 20
rect 106 -35 112 -18
rect 129 -35 136 -18
rect 106 -56 136 -35
rect 475 -19 505 2
rect 475 -36 481 -19
rect 498 -36 505 -19
rect 475 -57 505 -36
rect 844 -19 874 2
rect 844 -36 850 -19
rect 867 -36 874 -19
rect 844 -57 874 -36
rect 1215 -19 1245 2
rect 1215 -36 1221 -19
rect 1238 -36 1245 -19
rect 1215 -57 1245 -36
rect 1585 -19 1615 2
rect 1585 -36 1591 -19
rect 1608 -36 1615 -19
rect 1585 -57 1615 -36
rect 1954 -19 1984 2
rect 1954 -36 1960 -19
rect 1977 -36 1984 -19
rect 1954 -57 1984 -36
rect 2323 -19 2353 2
rect 2323 -36 2329 -19
rect 2346 -36 2353 -19
rect 2323 -57 2353 -36
rect 2692 -19 2722 2
rect 2692 -36 2698 -19
rect 2715 -36 2722 -19
rect 2692 -57 2722 -36
<< polycont >>
rect 112 -35 129 -18
rect 481 -36 498 -19
rect 850 -36 867 -19
rect 1221 -36 1238 -19
rect 1591 -36 1608 -19
rect 1960 -36 1977 -19
rect 2329 -36 2346 -19
rect 2698 -36 2715 -19
<< locali >>
rect 69 226 176 228
rect 69 195 86 226
rect 156 195 176 226
rect 69 186 176 195
rect 438 225 545 227
rect 438 194 455 225
rect 525 194 545 225
rect 438 185 545 194
rect 807 225 914 227
rect 807 194 824 225
rect 894 194 914 225
rect 807 185 914 194
rect 1178 225 1285 227
rect 1178 194 1195 225
rect 1265 194 1285 225
rect 1178 185 1285 194
rect 1548 225 1655 227
rect 1548 194 1565 225
rect 1635 194 1655 225
rect 1548 185 1655 194
rect 1917 225 2024 227
rect 1917 194 1934 225
rect 2004 194 2024 225
rect 1917 185 2024 194
rect 2286 225 2393 227
rect 2286 194 2303 225
rect 2373 194 2393 225
rect 2286 185 2393 194
rect 2655 225 2762 227
rect 2655 194 2672 225
rect 2742 194 2762 225
rect 2655 185 2762 194
rect 83 151 218 168
rect 83 129 100 151
rect 201 129 218 151
rect 452 150 587 167
rect 452 128 469 150
rect 570 128 587 150
rect 821 150 956 167
rect 821 128 838 150
rect 939 128 956 150
rect 1192 150 1327 167
rect 1192 128 1209 150
rect 1310 128 1327 150
rect 1562 150 1697 167
rect 1562 128 1579 150
rect 1680 128 1697 150
rect 1931 150 2066 167
rect 1931 128 1948 150
rect 2049 128 2066 150
rect 2300 150 2435 167
rect 2300 128 2317 150
rect 2418 128 2435 150
rect 2669 150 2804 167
rect 2669 128 2686 150
rect 2787 128 2804 150
rect 104 -35 112 -18
rect 129 -35 137 -18
rect 473 -36 481 -19
rect 498 -36 506 -19
rect 842 -36 850 -19
rect 867 -36 875 -19
rect 1213 -36 1221 -19
rect 1238 -36 1246 -19
rect 1583 -36 1591 -19
rect 1608 -36 1616 -19
rect 1952 -36 1960 -19
rect 1977 -36 1985 -19
rect 2321 -36 2329 -19
rect 2346 -36 2354 -19
rect 2690 -36 2698 -19
rect 2715 -36 2723 -19
rect 43 -214 135 -204
rect 43 -249 53 -214
rect 125 -249 135 -214
rect 43 -252 135 -249
rect 412 -215 504 -205
rect 412 -250 422 -215
rect 494 -250 504 -215
rect 412 -253 504 -250
rect 781 -215 873 -205
rect 781 -250 791 -215
rect 863 -250 873 -215
rect 781 -253 873 -250
rect 1152 -215 1244 -205
rect 1152 -250 1162 -215
rect 1234 -250 1244 -215
rect 1152 -253 1244 -250
rect 1522 -215 1614 -205
rect 1522 -250 1532 -215
rect 1604 -250 1614 -215
rect 1522 -253 1614 -250
rect 1891 -215 1983 -205
rect 1891 -250 1901 -215
rect 1973 -250 1983 -215
rect 1891 -253 1983 -250
rect 2260 -215 2352 -205
rect 2260 -250 2270 -215
rect 2342 -250 2352 -215
rect 2260 -253 2352 -250
rect 2629 -215 2721 -205
rect 2629 -250 2639 -215
rect 2711 -250 2721 -215
rect 2629 -253 2721 -250
<< viali >>
rect 96 198 144 216
rect 465 197 513 215
rect 834 197 882 215
rect 1205 197 1253 215
rect 1575 197 1623 215
rect 1944 197 1992 215
rect 2313 197 2361 215
rect 2682 197 2730 215
rect 112 -35 129 -18
rect 481 -36 498 -19
rect 850 -36 867 -19
rect 1221 -36 1238 -19
rect 1591 -36 1608 -19
rect 1960 -36 1977 -19
rect 2329 -36 2346 -19
rect 2698 -36 2715 -19
rect 71 -245 110 -218
rect 440 -246 479 -219
rect 809 -246 848 -219
rect 1180 -246 1219 -219
rect 1550 -246 1589 -219
rect 1919 -246 1958 -219
rect 2288 -246 2327 -219
rect 2657 -246 2696 -219
<< metal1 >>
rect 98 219 103 226
rect 83 216 103 219
rect 141 219 146 226
rect 141 216 162 219
rect 467 218 472 225
rect 83 198 96 216
rect 144 198 162 216
rect 83 189 103 198
rect 141 189 162 198
rect 83 169 162 189
rect 21 146 162 169
rect 452 215 472 218
rect 510 218 515 225
rect 836 218 841 225
rect 510 215 531 218
rect 452 197 465 215
rect 513 197 531 215
rect 452 188 472 197
rect 510 188 531 197
rect 452 168 531 188
rect 821 215 841 218
rect 879 218 884 225
rect 1207 218 1212 225
rect 879 215 900 218
rect 821 197 834 215
rect 882 197 900 215
rect 821 188 841 197
rect 879 188 900 197
rect 821 168 900 188
rect 1192 215 1212 218
rect 1250 218 1255 225
rect 1577 218 1582 225
rect 1250 215 1271 218
rect 1192 197 1205 215
rect 1253 197 1271 215
rect 1192 188 1212 197
rect 1250 188 1271 197
rect 1192 168 1271 188
rect 1562 215 1582 218
rect 1620 218 1625 225
rect 1946 218 1951 225
rect 1620 215 1641 218
rect 1562 197 1575 215
rect 1623 197 1641 215
rect 1562 188 1582 197
rect 1620 188 1641 197
rect 1562 168 1641 188
rect 1931 215 1951 218
rect 1989 218 1994 225
rect 2315 218 2320 225
rect 1989 215 2010 218
rect 1931 197 1944 215
rect 1992 197 2010 215
rect 1931 188 1951 197
rect 1989 188 2010 197
rect 1931 168 2010 188
rect 2300 215 2320 218
rect 2358 218 2363 225
rect 2684 218 2689 225
rect 2358 215 2379 218
rect 2300 197 2313 215
rect 2361 197 2379 215
rect 2300 188 2320 197
rect 2358 188 2379 197
rect 2300 168 2379 188
rect 2669 215 2689 218
rect 2727 218 2732 225
rect 2727 215 2748 218
rect 2669 197 2682 215
rect 2730 197 2748 215
rect 2669 188 2689 197
rect 2727 188 2748 197
rect 2669 168 2748 188
rect 21 128 44 146
rect 139 128 162 146
rect 390 145 531 168
rect 390 127 413 145
rect 508 127 531 145
rect 759 145 900 168
rect 759 127 782 145
rect 877 127 900 145
rect 1130 145 1271 168
rect 1130 127 1153 145
rect 1248 127 1271 145
rect 1500 145 1641 168
rect 1500 127 1523 145
rect 1618 127 1641 145
rect 1869 145 2010 168
rect 1869 127 1892 145
rect 1987 127 2010 145
rect 2238 145 2379 168
rect 2238 127 2261 145
rect 2356 127 2379 145
rect 2607 145 2748 168
rect 2607 127 2630 145
rect 2725 127 2748 145
rect 20 -15 39 -12
rect 198 -13 222 34
rect 20 -18 135 -15
rect 20 -35 112 -18
rect 129 -35 135 -18
rect 196 -32 224 -13
rect 389 -16 408 -13
rect 567 -14 591 33
rect 389 -19 504 -16
rect 20 -38 135 -35
rect 20 -40 39 -38
rect 198 -62 222 -32
rect 389 -36 481 -19
rect 498 -36 504 -19
rect 565 -33 593 -14
rect 758 -16 777 -13
rect 936 -14 960 33
rect 758 -19 873 -16
rect 389 -39 504 -36
rect 389 -41 408 -39
rect 139 -77 222 -62
rect 567 -63 591 -33
rect 758 -36 850 -19
rect 867 -36 873 -19
rect 934 -33 962 -14
rect 1129 -16 1148 -13
rect 1307 -14 1331 33
rect 1129 -19 1244 -16
rect 758 -39 873 -36
rect 758 -41 777 -39
rect 936 -63 960 -33
rect 1129 -36 1221 -19
rect 1238 -36 1244 -19
rect 1305 -33 1333 -14
rect 1499 -16 1518 -13
rect 1677 -14 1701 33
rect 1499 -19 1614 -16
rect 1129 -39 1244 -36
rect 1129 -41 1148 -39
rect 1307 -63 1331 -33
rect 1499 -36 1591 -19
rect 1608 -36 1614 -19
rect 1675 -33 1703 -14
rect 1868 -16 1887 -13
rect 2046 -14 2070 33
rect 1868 -19 1983 -16
rect 1499 -39 1614 -36
rect 1499 -41 1518 -39
rect 1677 -63 1701 -33
rect 1868 -36 1960 -19
rect 1977 -36 1983 -19
rect 2044 -33 2072 -14
rect 2237 -16 2256 -13
rect 2415 -14 2439 33
rect 2237 -19 2352 -16
rect 1868 -39 1983 -36
rect 1868 -41 1887 -39
rect 2046 -63 2070 -33
rect 2237 -36 2329 -19
rect 2346 -36 2352 -19
rect 2413 -33 2441 -14
rect 2606 -16 2625 -13
rect 2784 -14 2808 33
rect 2606 -19 2721 -16
rect 2237 -39 2352 -36
rect 2237 -41 2256 -39
rect 2415 -63 2439 -33
rect 2606 -36 2698 -19
rect 2715 -36 2721 -19
rect 2782 -33 2810 -14
rect 2606 -39 2721 -36
rect 2606 -41 2625 -39
rect 2784 -63 2808 -33
rect 508 -78 591 -63
rect 877 -78 960 -63
rect 1248 -78 1331 -63
rect 1618 -78 1701 -63
rect 1987 -78 2070 -63
rect 2356 -78 2439 -63
rect 2725 -78 2808 -63
rect 80 -215 103 -160
rect 60 -248 65 -215
rect 116 -248 121 -215
rect 449 -216 472 -161
rect 818 -216 841 -161
rect 1189 -216 1212 -161
rect 1559 -216 1582 -161
rect 1928 -216 1951 -161
rect 2297 -216 2320 -161
rect 2666 -216 2689 -161
rect 429 -249 434 -216
rect 485 -249 490 -216
rect 798 -249 803 -216
rect 854 -249 859 -216
rect 1169 -249 1174 -216
rect 1225 -249 1230 -216
rect 1539 -249 1544 -216
rect 1595 -249 1600 -216
rect 1908 -249 1913 -216
rect 1964 -249 1969 -216
rect 2277 -249 2282 -216
rect 2333 -249 2338 -216
rect 2646 -249 2651 -216
rect 2702 -249 2707 -216
<< via1 >>
rect 103 216 141 226
rect 103 198 141 216
rect 103 189 141 198
rect 472 215 510 225
rect 472 197 510 215
rect 472 188 510 197
rect 841 215 879 225
rect 841 197 879 215
rect 841 188 879 197
rect 1212 215 1250 225
rect 1212 197 1250 215
rect 1212 188 1250 197
rect 1582 215 1620 225
rect 1582 197 1620 215
rect 1582 188 1620 197
rect 1951 215 1989 225
rect 1951 197 1989 215
rect 1951 188 1989 197
rect 2320 215 2358 225
rect 2320 197 2358 215
rect 2320 188 2358 197
rect 2689 215 2727 225
rect 2689 197 2727 215
rect 2689 188 2727 197
rect 65 -218 116 -215
rect 65 -245 71 -218
rect 71 -245 110 -218
rect 110 -245 116 -218
rect 65 -248 116 -245
rect 434 -219 485 -216
rect 434 -246 440 -219
rect 440 -246 479 -219
rect 479 -246 485 -219
rect 434 -249 485 -246
rect 803 -219 854 -216
rect 803 -246 809 -219
rect 809 -246 848 -219
rect 848 -246 854 -219
rect 803 -249 854 -246
rect 1174 -219 1225 -216
rect 1174 -246 1180 -219
rect 1180 -246 1219 -219
rect 1219 -246 1225 -219
rect 1174 -249 1225 -246
rect 1544 -219 1595 -216
rect 1544 -246 1550 -219
rect 1550 -246 1589 -219
rect 1589 -246 1595 -219
rect 1544 -249 1595 -246
rect 1913 -219 1964 -216
rect 1913 -246 1919 -219
rect 1919 -246 1958 -219
rect 1958 -246 1964 -219
rect 1913 -249 1964 -246
rect 2282 -219 2333 -216
rect 2282 -246 2288 -219
rect 2288 -246 2327 -219
rect 2327 -246 2333 -219
rect 2282 -249 2333 -246
rect 2651 -219 2702 -216
rect 2651 -246 2657 -219
rect 2657 -246 2696 -219
rect 2696 -246 2702 -219
rect 2651 -249 2702 -246
<< metal2 >>
rect 99 231 146 236
rect 99 184 146 189
rect 468 230 515 235
rect 468 183 515 188
rect 837 230 884 235
rect 837 183 884 188
rect 1208 230 1255 235
rect 1208 183 1255 188
rect 1578 230 1625 235
rect 1578 183 1625 188
rect 1947 230 1994 235
rect 1947 183 1994 188
rect 2316 230 2363 235
rect 2316 183 2363 188
rect 2685 230 2732 235
rect 2685 183 2732 188
rect 65 -213 116 -210
rect 65 -215 117 -213
rect 116 -248 117 -215
rect 65 -252 117 -248
rect 434 -214 485 -211
rect 803 -214 854 -211
rect 1174 -214 1225 -211
rect 1544 -214 1595 -211
rect 1913 -214 1964 -211
rect 2282 -214 2333 -211
rect 2651 -214 2702 -211
rect 434 -216 486 -214
rect 485 -249 486 -216
rect 65 -253 116 -252
rect 434 -253 486 -249
rect 803 -216 855 -214
rect 854 -249 855 -216
rect 803 -253 855 -249
rect 1174 -216 1226 -214
rect 1225 -249 1226 -216
rect 1174 -253 1226 -249
rect 1544 -216 1596 -214
rect 1595 -249 1596 -216
rect 1544 -253 1596 -249
rect 1913 -216 1965 -214
rect 1964 -249 1965 -216
rect 1913 -253 1965 -249
rect 2282 -216 2334 -214
rect 2333 -249 2334 -216
rect 2282 -253 2334 -249
rect 2651 -216 2703 -214
rect 2702 -249 2703 -216
rect 2651 -253 2703 -249
rect 434 -254 485 -253
rect 803 -254 854 -253
rect 1174 -254 1225 -253
rect 1544 -254 1595 -253
rect 1913 -254 1964 -253
rect 2282 -254 2333 -253
rect 2651 -254 2702 -253
<< via2 >>
rect 99 226 146 231
rect 99 189 103 226
rect 103 189 141 226
rect 141 189 146 226
rect 468 225 515 230
rect 468 188 472 225
rect 472 188 510 225
rect 510 188 515 225
rect 837 225 884 230
rect 837 188 841 225
rect 841 188 879 225
rect 879 188 884 225
rect 1208 225 1255 230
rect 1208 188 1212 225
rect 1212 188 1250 225
rect 1250 188 1255 225
rect 1578 225 1625 230
rect 1578 188 1582 225
rect 1582 188 1620 225
rect 1620 188 1625 225
rect 1947 225 1994 230
rect 1947 188 1951 225
rect 1951 188 1989 225
rect 1989 188 1994 225
rect 2316 225 2363 230
rect 2316 188 2320 225
rect 2320 188 2358 225
rect 2358 188 2363 225
rect 2685 225 2732 230
rect 2685 188 2689 225
rect 2689 188 2727 225
rect 2727 188 2732 225
rect 73 -247 106 -218
rect 442 -248 475 -219
rect 811 -248 844 -219
rect 1182 -248 1215 -219
rect 1552 -248 1585 -219
rect 1921 -248 1954 -219
rect 2290 -248 2323 -219
rect 2659 -248 2692 -219
<< metal3 >>
rect 21 238 218 241
rect 21 184 95 238
rect 150 184 218 238
rect 21 166 218 184
rect 390 237 587 240
rect 390 183 464 237
rect 519 183 587 237
rect 390 165 587 183
rect 759 237 956 240
rect 759 183 833 237
rect 888 183 956 237
rect 759 165 956 183
rect 1130 237 1327 240
rect 1130 183 1204 237
rect 1259 183 1327 237
rect 1130 165 1327 183
rect 1500 237 1697 240
rect 1500 183 1574 237
rect 1629 183 1697 237
rect 1500 165 1697 183
rect 1869 237 2066 240
rect 1869 183 1943 237
rect 1998 183 2066 237
rect 1869 165 2066 183
rect 2238 237 2435 240
rect 2238 183 2312 237
rect 2367 183 2435 237
rect 2238 165 2435 183
rect 2607 237 2804 240
rect 2607 183 2681 237
rect 2736 183 2804 237
rect 2607 165 2804 183
rect 50 -208 130 -207
rect 50 -213 65 -208
rect 49 -254 65 -213
rect 50 -258 65 -254
rect 116 -258 130 -208
rect 419 -209 499 -208
rect 419 -214 434 -209
rect 418 -255 434 -214
rect 50 -261 130 -258
rect 419 -259 434 -255
rect 485 -259 499 -209
rect 788 -209 868 -208
rect 788 -214 803 -209
rect 787 -255 803 -214
rect 419 -262 499 -259
rect 788 -259 803 -255
rect 854 -259 868 -209
rect 1159 -209 1239 -208
rect 1159 -214 1174 -209
rect 1158 -255 1174 -214
rect 788 -262 868 -259
rect 1159 -259 1174 -255
rect 1225 -259 1239 -209
rect 1529 -209 1609 -208
rect 1529 -214 1544 -209
rect 1528 -255 1544 -214
rect 1159 -262 1239 -259
rect 1529 -259 1544 -255
rect 1595 -259 1609 -209
rect 1898 -209 1978 -208
rect 1898 -214 1913 -209
rect 1897 -255 1913 -214
rect 1529 -262 1609 -259
rect 1898 -259 1913 -255
rect 1964 -259 1978 -209
rect 2267 -209 2347 -208
rect 2267 -214 2282 -209
rect 2266 -255 2282 -214
rect 1898 -262 1978 -259
rect 2267 -259 2282 -255
rect 2333 -259 2347 -209
rect 2636 -209 2716 -208
rect 2636 -214 2651 -209
rect 2635 -255 2651 -214
rect 2267 -262 2347 -259
rect 2636 -259 2651 -255
rect 2702 -259 2716 -209
rect 2636 -262 2716 -259
<< via3 >>
rect 95 231 150 238
rect 95 189 99 231
rect 99 189 146 231
rect 146 189 150 231
rect 95 184 150 189
rect 464 230 519 237
rect 464 188 468 230
rect 468 188 515 230
rect 515 188 519 230
rect 464 183 519 188
rect 833 230 888 237
rect 833 188 837 230
rect 837 188 884 230
rect 884 188 888 230
rect 833 183 888 188
rect 1204 230 1259 237
rect 1204 188 1208 230
rect 1208 188 1255 230
rect 1255 188 1259 230
rect 1204 183 1259 188
rect 1574 230 1629 237
rect 1574 188 1578 230
rect 1578 188 1625 230
rect 1625 188 1629 230
rect 1574 183 1629 188
rect 1943 230 1998 237
rect 1943 188 1947 230
rect 1947 188 1994 230
rect 1994 188 1998 230
rect 1943 183 1998 188
rect 2312 230 2367 237
rect 2312 188 2316 230
rect 2316 188 2363 230
rect 2363 188 2367 230
rect 2312 183 2367 188
rect 2681 230 2736 237
rect 2681 188 2685 230
rect 2685 188 2732 230
rect 2732 188 2736 230
rect 2681 183 2736 188
rect 65 -218 116 -208
rect 65 -247 73 -218
rect 73 -247 106 -218
rect 106 -247 116 -218
rect 65 -258 116 -247
rect 434 -219 485 -209
rect 434 -248 442 -219
rect 442 -248 475 -219
rect 475 -248 485 -219
rect 434 -259 485 -248
rect 803 -219 854 -209
rect 803 -248 811 -219
rect 811 -248 844 -219
rect 844 -248 854 -219
rect 803 -259 854 -248
rect 1174 -219 1225 -209
rect 1174 -248 1182 -219
rect 1182 -248 1215 -219
rect 1215 -248 1225 -219
rect 1174 -259 1225 -248
rect 1544 -219 1595 -209
rect 1544 -248 1552 -219
rect 1552 -248 1585 -219
rect 1585 -248 1595 -219
rect 1544 -259 1595 -248
rect 1913 -219 1964 -209
rect 1913 -248 1921 -219
rect 1921 -248 1954 -219
rect 1954 -248 1964 -219
rect 1913 -259 1964 -248
rect 2282 -219 2333 -209
rect 2282 -248 2290 -219
rect 2290 -248 2323 -219
rect 2323 -248 2333 -219
rect 2282 -259 2333 -248
rect 2651 -219 2702 -209
rect 2651 -248 2659 -219
rect 2659 -248 2692 -219
rect 2692 -248 2702 -219
rect 2651 -259 2702 -248
<< metal4 >>
rect 0 238 2830 275
rect 0 184 95 238
rect 150 237 2830 238
rect 150 184 464 237
rect 0 183 464 184
rect 519 183 833 237
rect 888 183 1204 237
rect 1259 183 1574 237
rect 1629 183 1943 237
rect 1998 183 2312 237
rect 2367 183 2681 237
rect 2736 183 2830 237
rect 0 180 2830 183
rect -1 -208 2829 -180
rect -1 -258 65 -208
rect 116 -209 2829 -208
rect 116 -258 434 -209
rect -1 -259 434 -258
rect 485 -259 803 -209
rect 854 -259 1174 -209
rect 1225 -259 1544 -209
rect 1595 -259 1913 -209
rect 1964 -259 2282 -209
rect 2333 -259 2651 -209
rect 2702 -259 2829 -209
rect -1 -275 2829 -259
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_0
timestamp 1735996060
transform 1 0 490 0 1 -113
box -44 -63 44 63
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_1
timestamp 1735996060
transform 1 0 859 0 1 -115
box -44 -63 44 63
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_2
timestamp 1735996060
transform 1 0 1230 0 1 -115
box -44 -63 44 63
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_3
timestamp 1735996060
transform 1 0 1600 0 1 -115
box -44 -63 44 63
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_4
timestamp 1735996060
transform 1 0 2707 0 1 -113
box -44 -63 44 63
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_5
timestamp 1735996060
transform 1 0 1969 0 1 -115
box -44 -63 44 63
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_6
timestamp 1735996060
transform 1 0 2338 0 1 -113
box -44 -63 44 63
use sky130_fd_pr__nfet_01v8_CH4TXP  sky130_fd_pr__nfet_01v8_CH4TXP_7
timestamp 1735996060
transform 1 0 121 0 1 -114
box -44 -63 44 63
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_0
timestamp 1735996060
transform 1 0 490 0 1 81
box -121 -81 121 81
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_1
timestamp 1735996060
transform 1 0 859 0 1 79
box -121 -81 121 81
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_2
timestamp 1735996060
transform 1 0 1230 0 1 78
box -121 -81 121 81
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_3
timestamp 1735996060
transform 1 0 1600 0 1 78
box -121 -81 121 81
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_4
timestamp 1735996060
transform 1 0 2707 0 1 78
box -121 -81 121 81
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_5
timestamp 1735996060
transform 1 0 1969 0 1 78
box -121 -81 121 81
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_6
timestamp 1735996060
transform 1 0 2338 0 1 78
box -121 -81 121 81
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_7
timestamp 1735996060
transform 1 0 121 0 1 79
box -121 -81 121 81
<< labels >>
flabel metal1 20 -40 39 -12 1 FreeSerif 160 0 0 0 A[0]
port 3 n
flabel metal1 389 -41 408 -13 1 FreeSerif 160 0 0 0 A[1]
port 4 n
flabel metal1 758 -41 777 -13 1 FreeSerif 160 0 0 0 A[2]
port 5 n
flabel metal1 1129 -41 1148 -13 1 FreeSerif 160 0 0 0 A[3]
port 6 n
flabel metal1 1499 -41 1518 -13 1 FreeSerif 160 0 0 0 A[4]
port 7 n
flabel metal1 1868 -41 1887 -13 1 FreeSerif 160 0 0 0 A[5]
port 8 n
flabel metal1 2237 -41 2256 -13 1 FreeSerif 160 0 0 0 A[6]
port 9 n
flabel metal1 2606 -41 2625 -13 1 FreeSerif 160 0 0 0 A[7]
port 10 n
flabel metal1 2782 -33 2810 -14 1 FreeSerif 160 0 0 0 Y[7]
port 11 n
flabel metal1 2413 -33 2441 -14 1 FreeSerif 160 0 0 0 Y[6]
port 12 n
flabel metal1 2044 -33 2072 -14 1 FreeSerif 160 0 0 0 Y[5]
port 13 n
flabel metal1 1675 -33 1703 -14 1 FreeSerif 160 0 0 0 Y[4]
port 14 n
flabel metal1 1305 -33 1333 -14 1 FreeSerif 160 0 0 0 Y[3]
port 15 n
flabel metal1 934 -33 962 -14 1 FreeSerif 160 0 0 0 Y[2]
port 16 n
flabel metal1 565 -33 593 -14 1 FreeSerif 160 0 0 0 Y[1]
port 17 n
flabel metal1 196 -32 224 -13 1 FreeSerif 160 0 0 0 Y[0]
port 18 n
flabel metal4 1306 181 1497 275 1 FreeSerif 400 0 0 0 VDD
port 19 n
flabel metal4 1305 -275 1507 -193 1 FreeSerif 400 0 0 0 VSS
port 20 n
<< end >>
