magic
tech sky130B
magscale 1 2
timestamp 1736531572
<< nwell >>
rect 546 772 1022 964
rect 356 476 1200 772
rect -31 181 265 198
rect -77 153 265 181
rect 807 173 1096 196
rect 302 -60 1140 173
<< psubdiff >>
rect 600 -1386 852 -1366
rect 600 -1442 658 -1386
rect 790 -1442 852 -1386
rect 600 -1464 852 -1442
<< nsubdiff >>
rect 584 874 984 926
rect 584 830 708 874
rect 830 830 984 874
rect 584 782 984 830
<< psubdiffcont >>
rect 658 -1442 790 -1386
<< nsubdiffcont >>
rect 708 830 830 874
<< poly >>
rect 453 630 749 681
rect 1290 432 1586 483
rect -31 147 513 198
rect 1408 196 1467 214
rect 94 -132 154 147
rect 807 145 1350 196
rect 1392 145 1467 196
rect 1392 58 1452 145
rect 1324 48 1452 58
rect 1324 14 1340 48
rect 1374 14 1452 48
rect 396 -55 692 5
rect 750 -54 1046 6
rect 1324 4 1452 14
rect 750 -55 810 -54
rect 868 -55 928 -54
rect 986 -55 1046 -54
rect -70 -146 154 -132
rect -70 -180 -54 -146
rect -20 -180 154 -146
rect -70 -192 154 -180
rect 94 -705 154 -192
rect 364 -645 431 -638
rect 514 -645 574 -497
rect 364 -654 574 -645
rect 364 -688 380 -654
rect 414 -688 574 -654
rect 364 -704 574 -688
rect 94 -721 245 -705
rect 94 -755 195 -721
rect 229 -755 245 -721
rect 94 -771 245 -755
rect 94 -800 154 -771
rect 514 -801 574 -704
rect 868 -645 928 -497
rect 1011 -645 1078 -638
rect 868 -654 1078 -645
rect 868 -688 1028 -654
rect 1062 -688 1078 -654
rect 868 -704 1078 -688
rect 630 -738 696 -722
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 630 -788 696 -772
rect 748 -737 814 -722
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 748 -787 814 -771
rect 632 -800 692 -788
rect 750 -799 810 -787
rect 868 -801 928 -704
rect 1392 -706 1452 4
rect 1302 -722 1452 -706
rect 1302 -756 1318 -722
rect 1352 -756 1452 -722
rect 1302 -772 1452 -756
rect 1392 -800 1452 -772
<< polycont >>
rect 1340 14 1374 48
rect -54 -180 -20 -146
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1028 -688 1062 -654
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 1318 -756 1352 -722
<< locali >>
rect 674 874 876 894
rect 674 830 708 874
rect 830 830 876 874
rect 674 820 760 830
rect 798 820 876 830
rect 674 802 876 820
rect 761 656 1031 691
rect 761 613 795 656
rect 997 613 1031 656
rect -77 457 193 492
rect -77 415 -43 457
rect 159 415 193 457
rect 1324 14 1330 48
rect 1384 14 1390 48
rect 467 -524 503 -419
rect 702 -524 738 -419
rect 940 -524 976 -420
rect 467 -564 1562 -524
rect 486 -565 1562 -564
rect 364 -654 431 -638
rect 364 -688 380 -654
rect 414 -688 431 -654
rect 364 -704 431 -688
rect 195 -721 229 -705
rect 195 -771 229 -755
rect 541 -806 575 -565
rect 1011 -654 1078 -638
rect 1011 -688 1028 -654
rect 1062 -688 1078 -654
rect 1011 -704 1078 -688
rect 1318 -722 1352 -706
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 1318 -772 1352 -756
rect 541 -809 613 -806
rect 541 -852 620 -809
rect 468 -1265 503 -1198
rect 939 -1265 974 -1198
rect 468 -1300 974 -1265
rect 642 -1386 698 -1370
rect 748 -1386 806 -1370
rect 642 -1442 658 -1386
rect 790 -1442 806 -1386
rect 642 -1458 806 -1442
<< viali >>
rect 760 830 798 858
rect 760 820 798 830
rect 1330 48 1384 58
rect 1330 14 1340 48
rect 1340 14 1374 48
rect 1374 14 1384 48
rect 1330 4 1384 14
rect -70 -146 -4 -132
rect -70 -180 -54 -146
rect -54 -180 -20 -146
rect -20 -180 -4 -146
rect -70 -192 -4 -180
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1562 -596 1664 -494
rect 1028 -688 1062 -654
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 1318 -756 1352 -722
rect 698 -1386 748 -1364
rect 698 -1406 748 -1386
<< metal1 >>
rect 740 844 750 866
rect 712 812 750 844
rect 804 844 814 866
rect 804 812 846 844
rect 712 761 846 812
rect 41 718 1514 761
rect 41 415 75 718
rect 407 613 441 718
rect 643 613 677 718
rect 879 613 913 718
rect 1115 613 1149 718
rect 1480 415 1514 718
rect 186 378 193 403
rect 311 378 410 403
rect -77 181 -43 235
rect 304 227 410 378
rect 761 247 795 337
rect 525 235 565 247
rect 637 235 683 247
rect 755 235 795 247
rect 525 181 559 235
rect 761 181 795 235
rect 1143 227 1247 403
rect -77 146 82 181
rect 525 146 795 181
rect 1362 181 1396 249
rect 1598 181 1632 249
rect 1362 146 1632 181
rect -132 -2 -58 64
rect 8 -2 18 64
rect -132 -132 8 -126
rect -132 -192 -70 -132
rect -4 -192 8 -132
rect -132 -198 8 -192
rect 48 -638 82 146
rect 761 84 795 146
rect 350 46 1092 84
rect 350 -92 384 46
rect 586 -96 620 46
rect 822 -98 856 46
rect 1058 -98 1092 46
rect 1318 58 1396 64
rect 1318 4 1330 58
rect 1384 4 1396 58
rect 1318 -2 1396 4
rect 350 -393 385 -359
rect 585 -393 620 -359
rect 822 -393 857 -359
rect 1058 -381 1092 -359
rect 1464 -637 1498 146
rect 1550 -494 1676 -488
rect 1550 -596 1562 -494
rect 1664 -596 1676 -494
rect 1550 -602 1676 -596
rect 1191 -638 1498 -637
rect 48 -643 364 -638
rect 1078 -643 1498 -638
rect 48 -654 431 -643
rect 48 -681 380 -654
rect 48 -828 82 -681
rect 364 -688 380 -681
rect 414 -688 431 -654
rect 364 -694 431 -688
rect 1011 -654 1498 -643
rect 1011 -688 1028 -654
rect 1062 -681 1498 -654
rect 1062 -688 1078 -681
rect 1191 -682 1498 -681
rect 1011 -694 1078 -688
rect 189 -721 245 -709
rect 189 -755 195 -721
rect 229 -722 245 -721
rect 1302 -722 1358 -710
rect 229 -738 696 -722
rect 229 -755 646 -738
rect 189 -771 646 -755
rect 630 -772 646 -771
rect 680 -772 696 -738
rect 630 -779 696 -772
rect 748 -737 1318 -722
rect 748 -771 764 -737
rect 798 -756 1318 -737
rect 1352 -756 1358 -722
rect 798 -771 1358 -756
rect 748 -781 815 -771
rect 1302 -772 1358 -771
rect 1464 -828 1498 -682
rect 165 -1304 199 -995
rect 822 -1304 856 -1198
rect 1346 -1304 1379 -982
rect 165 -1336 1379 -1304
rect 658 -1358 790 -1336
rect 658 -1416 692 -1358
rect 754 -1416 790 -1358
rect 658 -1421 790 -1416
<< via1 >>
rect 750 858 804 866
rect 750 820 760 858
rect 760 820 798 858
rect 798 820 804 858
rect 750 812 804 820
rect -58 -2 8 64
rect 1330 4 1384 58
rect 692 -1364 754 -1358
rect 692 -1406 698 -1364
rect 698 -1406 748 -1364
rect 748 -1406 754 -1364
rect 692 -1416 754 -1406
<< metal2 >>
rect 738 874 816 884
rect 738 794 816 804
rect -64 -2 -58 64
rect 8 58 1384 64
rect 8 4 1330 58
rect 8 -2 1384 4
rect 686 -1356 758 -1346
rect 686 -1436 758 -1426
<< via2 >>
rect 738 866 816 874
rect 738 812 750 866
rect 750 812 804 866
rect 804 812 816 866
rect 738 804 816 812
rect 686 -1358 758 -1356
rect 686 -1416 692 -1358
rect 692 -1416 754 -1358
rect 754 -1416 758 -1358
rect 686 -1426 758 -1416
<< metal3 >>
rect 668 876 882 880
rect 668 804 738 876
rect 814 874 882 876
rect 816 804 882 874
rect 668 802 882 804
rect 728 799 826 802
rect 648 -1342 800 -1340
rect 646 -1346 800 -1342
rect 646 -1434 676 -1346
rect 770 -1434 800 -1346
rect 646 -1440 800 -1434
rect 648 -1450 800 -1440
<< via3 >>
rect 738 874 814 876
rect 738 810 814 874
rect 676 -1356 770 -1346
rect 676 -1426 686 -1356
rect 686 -1426 758 -1356
rect 758 -1426 770 -1356
rect 676 -1434 770 -1426
<< metal4 >>
rect -106 876 1652 932
rect -106 810 738 876
rect 814 810 1652 876
rect -106 768 1652 810
rect 50 -1346 1414 -1340
rect 50 -1434 676 -1346
rect 770 -1434 1414 -1346
rect 50 -1464 1414 -1434
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_0
timestamp 1736499154
transform 1 0 721 0 1 -1010
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_0
timestamp 1736499154
transform 1 0 1422 0 1 -910
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_1
timestamp 1736499154
transform 1 0 124 0 1 -910
box -88 -126 88 126
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_0
timestamp 1736499154
transform 1 0 721 0 1 -278
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_1
timestamp 1736499154
transform 1 0 778 0 1 415
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_0
timestamp 1736499154
transform 1 0 1438 0 1 315
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_1
timestamp 1736499154
transform 1 0 117 0 1 315
box -242 -162 242 162
<< labels >>
flabel metal4 672 -1440 772 -1366 1 FreeSerif 640 0 0 0 VSS
port 11 n
flabel metal4 700 798 860 916 1 FreeSerif 640 0 0 0 VDD
port 14 n
flabel metal1 1554 -600 1674 -492 1 FreeSerif 400 0 0 0 Y
port 15 n
flabel metal1 -132 -198 -72 -132 1 FreeSerif 480 0 0 0 A
port 16 n
flabel metal1 -132 -2 -72 56 1 FreeSerif 480 0 0 0 B
port 17 n
<< end >>
