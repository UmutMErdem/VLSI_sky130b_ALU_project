magic
tech sky130B
magscale 1 2
timestamp 1736520267
<< nwell >>
rect 0 330 1192 576
rect 1448 330 2640 576
rect 2946 332 4138 578
rect 4394 332 5586 578
rect 0 318 1193 330
rect 1448 318 2641 330
rect 2946 320 4139 332
rect 4394 320 5587 332
rect 1 6 1193 318
rect 1449 6 2641 318
rect 2947 8 4139 320
rect 4395 8 5587 320
rect 5914 330 7106 576
rect 7362 330 8554 576
rect 8860 332 10052 578
rect 10308 332 11500 578
rect 5914 318 7107 330
rect 7362 318 8555 330
rect 8860 320 10053 332
rect 10308 320 11501 332
rect 5915 6 7107 318
rect 7363 6 8555 318
rect 8861 8 10053 320
rect 10309 8 11501 320
<< nmos >>
rect 332 -569 392 -169
rect 450 -569 510 -169
rect 685 -369 745 -169
rect 1780 -569 1840 -169
rect 1898 -569 1958 -169
rect 2133 -369 2193 -169
rect 3278 -567 3338 -167
rect 3396 -567 3456 -167
rect 3631 -367 3691 -167
rect 4726 -567 4786 -167
rect 4844 -567 4904 -167
rect 5079 -367 5139 -167
rect 6246 -569 6306 -169
rect 6364 -569 6424 -169
rect 6599 -369 6659 -169
rect 7694 -569 7754 -169
rect 7812 -569 7872 -169
rect 8047 -369 8107 -169
rect 9192 -567 9252 -167
rect 9310 -567 9370 -167
rect 9545 -367 9605 -167
rect 10640 -567 10700 -167
rect 10758 -567 10818 -167
rect 10993 -367 11053 -167
<< pmos >>
rect 95 68 155 268
rect 213 68 273 268
rect 331 68 391 268
rect 449 68 509 268
rect 567 68 627 268
rect 685 68 745 268
rect 803 68 863 268
rect 921 68 981 268
rect 1039 68 1099 268
rect 1543 68 1603 268
rect 1661 68 1721 268
rect 1779 68 1839 268
rect 1897 68 1957 268
rect 2015 68 2075 268
rect 2133 68 2193 268
rect 2251 68 2311 268
rect 2369 68 2429 268
rect 2487 68 2547 268
rect 3041 70 3101 270
rect 3159 70 3219 270
rect 3277 70 3337 270
rect 3395 70 3455 270
rect 3513 70 3573 270
rect 3631 70 3691 270
rect 3749 70 3809 270
rect 3867 70 3927 270
rect 3985 70 4045 270
rect 4489 70 4549 270
rect 4607 70 4667 270
rect 4725 70 4785 270
rect 4843 70 4903 270
rect 4961 70 5021 270
rect 5079 70 5139 270
rect 5197 70 5257 270
rect 5315 70 5375 270
rect 5433 70 5493 270
rect 6009 68 6069 268
rect 6127 68 6187 268
rect 6245 68 6305 268
rect 6363 68 6423 268
rect 6481 68 6541 268
rect 6599 68 6659 268
rect 6717 68 6777 268
rect 6835 68 6895 268
rect 6953 68 7013 268
rect 7457 68 7517 268
rect 7575 68 7635 268
rect 7693 68 7753 268
rect 7811 68 7871 268
rect 7929 68 7989 268
rect 8047 68 8107 268
rect 8165 68 8225 268
rect 8283 68 8343 268
rect 8401 68 8461 268
rect 8955 70 9015 270
rect 9073 70 9133 270
rect 9191 70 9251 270
rect 9309 70 9369 270
rect 9427 70 9487 270
rect 9545 70 9605 270
rect 9663 70 9723 270
rect 9781 70 9841 270
rect 9899 70 9959 270
rect 10403 70 10463 270
rect 10521 70 10581 270
rect 10639 70 10699 270
rect 10757 70 10817 270
rect 10875 70 10935 270
rect 10993 70 11053 270
rect 11111 70 11171 270
rect 11229 70 11289 270
rect 11347 70 11407 270
<< ndiff >>
rect 274 -181 332 -169
rect 274 -557 286 -181
rect 320 -557 332 -181
rect 274 -569 332 -557
rect 392 -181 450 -169
rect 392 -557 404 -181
rect 438 -557 450 -181
rect 392 -569 450 -557
rect 510 -181 568 -169
rect 510 -557 522 -181
rect 556 -557 568 -181
rect 627 -181 685 -169
rect 627 -357 639 -181
rect 673 -357 685 -181
rect 627 -369 685 -357
rect 745 -181 803 -169
rect 745 -357 757 -181
rect 791 -357 803 -181
rect 745 -369 803 -357
rect 1722 -181 1780 -169
rect 510 -569 568 -557
rect 1722 -557 1734 -181
rect 1768 -557 1780 -181
rect 1722 -569 1780 -557
rect 1840 -181 1898 -169
rect 1840 -557 1852 -181
rect 1886 -557 1898 -181
rect 1840 -569 1898 -557
rect 1958 -181 2016 -169
rect 1958 -557 1970 -181
rect 2004 -557 2016 -181
rect 2075 -181 2133 -169
rect 2075 -357 2087 -181
rect 2121 -357 2133 -181
rect 2075 -369 2133 -357
rect 2193 -181 2251 -169
rect 2193 -357 2205 -181
rect 2239 -357 2251 -181
rect 2193 -369 2251 -357
rect 3220 -179 3278 -167
rect 1958 -569 2016 -557
rect 3220 -555 3232 -179
rect 3266 -555 3278 -179
rect 3220 -567 3278 -555
rect 3338 -179 3396 -167
rect 3338 -555 3350 -179
rect 3384 -555 3396 -179
rect 3338 -567 3396 -555
rect 3456 -179 3514 -167
rect 3456 -555 3468 -179
rect 3502 -555 3514 -179
rect 3573 -179 3631 -167
rect 3573 -355 3585 -179
rect 3619 -355 3631 -179
rect 3573 -367 3631 -355
rect 3691 -179 3749 -167
rect 3691 -355 3703 -179
rect 3737 -355 3749 -179
rect 3691 -367 3749 -355
rect 4668 -179 4726 -167
rect 3456 -567 3514 -555
rect 4668 -555 4680 -179
rect 4714 -555 4726 -179
rect 4668 -567 4726 -555
rect 4786 -179 4844 -167
rect 4786 -555 4798 -179
rect 4832 -555 4844 -179
rect 4786 -567 4844 -555
rect 4904 -179 4962 -167
rect 4904 -555 4916 -179
rect 4950 -555 4962 -179
rect 5021 -179 5079 -167
rect 5021 -355 5033 -179
rect 5067 -355 5079 -179
rect 5021 -367 5079 -355
rect 5139 -179 5197 -167
rect 5139 -355 5151 -179
rect 5185 -355 5197 -179
rect 5139 -367 5197 -355
rect 6188 -181 6246 -169
rect 4904 -567 4962 -555
rect 6188 -557 6200 -181
rect 6234 -557 6246 -181
rect 6188 -569 6246 -557
rect 6306 -181 6364 -169
rect 6306 -557 6318 -181
rect 6352 -557 6364 -181
rect 6306 -569 6364 -557
rect 6424 -181 6482 -169
rect 6424 -557 6436 -181
rect 6470 -557 6482 -181
rect 6541 -181 6599 -169
rect 6541 -357 6553 -181
rect 6587 -357 6599 -181
rect 6541 -369 6599 -357
rect 6659 -181 6717 -169
rect 6659 -357 6671 -181
rect 6705 -357 6717 -181
rect 6659 -369 6717 -357
rect 7636 -181 7694 -169
rect 6424 -569 6482 -557
rect 7636 -557 7648 -181
rect 7682 -557 7694 -181
rect 7636 -569 7694 -557
rect 7754 -181 7812 -169
rect 7754 -557 7766 -181
rect 7800 -557 7812 -181
rect 7754 -569 7812 -557
rect 7872 -181 7930 -169
rect 7872 -557 7884 -181
rect 7918 -557 7930 -181
rect 7989 -181 8047 -169
rect 7989 -357 8001 -181
rect 8035 -357 8047 -181
rect 7989 -369 8047 -357
rect 8107 -181 8165 -169
rect 8107 -357 8119 -181
rect 8153 -357 8165 -181
rect 8107 -369 8165 -357
rect 9134 -179 9192 -167
rect 7872 -569 7930 -557
rect 9134 -555 9146 -179
rect 9180 -555 9192 -179
rect 9134 -567 9192 -555
rect 9252 -179 9310 -167
rect 9252 -555 9264 -179
rect 9298 -555 9310 -179
rect 9252 -567 9310 -555
rect 9370 -179 9428 -167
rect 9370 -555 9382 -179
rect 9416 -555 9428 -179
rect 9487 -179 9545 -167
rect 9487 -355 9499 -179
rect 9533 -355 9545 -179
rect 9487 -367 9545 -355
rect 9605 -179 9663 -167
rect 9605 -355 9617 -179
rect 9651 -355 9663 -179
rect 9605 -367 9663 -355
rect 10582 -179 10640 -167
rect 9370 -567 9428 -555
rect 10582 -555 10594 -179
rect 10628 -555 10640 -179
rect 10582 -567 10640 -555
rect 10700 -179 10758 -167
rect 10700 -555 10712 -179
rect 10746 -555 10758 -179
rect 10700 -567 10758 -555
rect 10818 -179 10876 -167
rect 10818 -555 10830 -179
rect 10864 -555 10876 -179
rect 10935 -179 10993 -167
rect 10935 -355 10947 -179
rect 10981 -355 10993 -179
rect 10935 -367 10993 -355
rect 11053 -179 11111 -167
rect 11053 -355 11065 -179
rect 11099 -355 11111 -179
rect 11053 -367 11111 -355
rect 10818 -567 10876 -555
<< pdiff >>
rect 37 256 95 268
rect 37 80 49 256
rect 83 80 95 256
rect 37 68 95 80
rect 155 256 213 268
rect 155 80 167 256
rect 201 80 213 256
rect 155 68 213 80
rect 273 256 331 268
rect 273 80 285 256
rect 319 80 331 256
rect 273 68 331 80
rect 391 256 449 268
rect 391 80 403 256
rect 437 80 449 256
rect 391 68 449 80
rect 509 256 567 268
rect 509 80 521 256
rect 555 80 567 256
rect 509 68 567 80
rect 627 256 685 268
rect 627 80 639 256
rect 673 80 685 256
rect 627 68 685 80
rect 745 256 803 268
rect 745 80 757 256
rect 791 80 803 256
rect 745 68 803 80
rect 863 256 921 268
rect 863 80 875 256
rect 909 80 921 256
rect 863 68 921 80
rect 981 256 1039 268
rect 981 80 993 256
rect 1027 80 1039 256
rect 981 68 1039 80
rect 1099 256 1157 268
rect 1099 80 1111 256
rect 1145 80 1157 256
rect 1099 68 1157 80
rect 1485 256 1543 268
rect 1485 80 1497 256
rect 1531 80 1543 256
rect 1485 68 1543 80
rect 1603 256 1661 268
rect 1603 80 1615 256
rect 1649 80 1661 256
rect 1603 68 1661 80
rect 1721 256 1779 268
rect 1721 80 1733 256
rect 1767 80 1779 256
rect 1721 68 1779 80
rect 1839 256 1897 268
rect 1839 80 1851 256
rect 1885 80 1897 256
rect 1839 68 1897 80
rect 1957 256 2015 268
rect 1957 80 1969 256
rect 2003 80 2015 256
rect 1957 68 2015 80
rect 2075 256 2133 268
rect 2075 80 2087 256
rect 2121 80 2133 256
rect 2075 68 2133 80
rect 2193 256 2251 268
rect 2193 80 2205 256
rect 2239 80 2251 256
rect 2193 68 2251 80
rect 2311 256 2369 268
rect 2311 80 2323 256
rect 2357 80 2369 256
rect 2311 68 2369 80
rect 2429 256 2487 268
rect 2429 80 2441 256
rect 2475 80 2487 256
rect 2429 68 2487 80
rect 2547 256 2605 268
rect 2547 80 2559 256
rect 2593 80 2605 256
rect 2547 68 2605 80
rect 2983 258 3041 270
rect 2983 82 2995 258
rect 3029 82 3041 258
rect 2983 70 3041 82
rect 3101 258 3159 270
rect 3101 82 3113 258
rect 3147 82 3159 258
rect 3101 70 3159 82
rect 3219 258 3277 270
rect 3219 82 3231 258
rect 3265 82 3277 258
rect 3219 70 3277 82
rect 3337 258 3395 270
rect 3337 82 3349 258
rect 3383 82 3395 258
rect 3337 70 3395 82
rect 3455 258 3513 270
rect 3455 82 3467 258
rect 3501 82 3513 258
rect 3455 70 3513 82
rect 3573 258 3631 270
rect 3573 82 3585 258
rect 3619 82 3631 258
rect 3573 70 3631 82
rect 3691 258 3749 270
rect 3691 82 3703 258
rect 3737 82 3749 258
rect 3691 70 3749 82
rect 3809 258 3867 270
rect 3809 82 3821 258
rect 3855 82 3867 258
rect 3809 70 3867 82
rect 3927 258 3985 270
rect 3927 82 3939 258
rect 3973 82 3985 258
rect 3927 70 3985 82
rect 4045 258 4103 270
rect 4045 82 4057 258
rect 4091 82 4103 258
rect 4045 70 4103 82
rect 4431 258 4489 270
rect 4431 82 4443 258
rect 4477 82 4489 258
rect 4431 70 4489 82
rect 4549 258 4607 270
rect 4549 82 4561 258
rect 4595 82 4607 258
rect 4549 70 4607 82
rect 4667 258 4725 270
rect 4667 82 4679 258
rect 4713 82 4725 258
rect 4667 70 4725 82
rect 4785 258 4843 270
rect 4785 82 4797 258
rect 4831 82 4843 258
rect 4785 70 4843 82
rect 4903 258 4961 270
rect 4903 82 4915 258
rect 4949 82 4961 258
rect 4903 70 4961 82
rect 5021 258 5079 270
rect 5021 82 5033 258
rect 5067 82 5079 258
rect 5021 70 5079 82
rect 5139 258 5197 270
rect 5139 82 5151 258
rect 5185 82 5197 258
rect 5139 70 5197 82
rect 5257 258 5315 270
rect 5257 82 5269 258
rect 5303 82 5315 258
rect 5257 70 5315 82
rect 5375 258 5433 270
rect 5375 82 5387 258
rect 5421 82 5433 258
rect 5375 70 5433 82
rect 5493 258 5551 270
rect 5493 82 5505 258
rect 5539 82 5551 258
rect 5493 70 5551 82
rect 5951 256 6009 268
rect 5951 80 5963 256
rect 5997 80 6009 256
rect 5951 68 6009 80
rect 6069 256 6127 268
rect 6069 80 6081 256
rect 6115 80 6127 256
rect 6069 68 6127 80
rect 6187 256 6245 268
rect 6187 80 6199 256
rect 6233 80 6245 256
rect 6187 68 6245 80
rect 6305 256 6363 268
rect 6305 80 6317 256
rect 6351 80 6363 256
rect 6305 68 6363 80
rect 6423 256 6481 268
rect 6423 80 6435 256
rect 6469 80 6481 256
rect 6423 68 6481 80
rect 6541 256 6599 268
rect 6541 80 6553 256
rect 6587 80 6599 256
rect 6541 68 6599 80
rect 6659 256 6717 268
rect 6659 80 6671 256
rect 6705 80 6717 256
rect 6659 68 6717 80
rect 6777 256 6835 268
rect 6777 80 6789 256
rect 6823 80 6835 256
rect 6777 68 6835 80
rect 6895 256 6953 268
rect 6895 80 6907 256
rect 6941 80 6953 256
rect 6895 68 6953 80
rect 7013 256 7071 268
rect 7013 80 7025 256
rect 7059 80 7071 256
rect 7013 68 7071 80
rect 7399 256 7457 268
rect 7399 80 7411 256
rect 7445 80 7457 256
rect 7399 68 7457 80
rect 7517 256 7575 268
rect 7517 80 7529 256
rect 7563 80 7575 256
rect 7517 68 7575 80
rect 7635 256 7693 268
rect 7635 80 7647 256
rect 7681 80 7693 256
rect 7635 68 7693 80
rect 7753 256 7811 268
rect 7753 80 7765 256
rect 7799 80 7811 256
rect 7753 68 7811 80
rect 7871 256 7929 268
rect 7871 80 7883 256
rect 7917 80 7929 256
rect 7871 68 7929 80
rect 7989 256 8047 268
rect 7989 80 8001 256
rect 8035 80 8047 256
rect 7989 68 8047 80
rect 8107 256 8165 268
rect 8107 80 8119 256
rect 8153 80 8165 256
rect 8107 68 8165 80
rect 8225 256 8283 268
rect 8225 80 8237 256
rect 8271 80 8283 256
rect 8225 68 8283 80
rect 8343 256 8401 268
rect 8343 80 8355 256
rect 8389 80 8401 256
rect 8343 68 8401 80
rect 8461 256 8519 268
rect 8461 80 8473 256
rect 8507 80 8519 256
rect 8461 68 8519 80
rect 8897 258 8955 270
rect 8897 82 8909 258
rect 8943 82 8955 258
rect 8897 70 8955 82
rect 9015 258 9073 270
rect 9015 82 9027 258
rect 9061 82 9073 258
rect 9015 70 9073 82
rect 9133 258 9191 270
rect 9133 82 9145 258
rect 9179 82 9191 258
rect 9133 70 9191 82
rect 9251 258 9309 270
rect 9251 82 9263 258
rect 9297 82 9309 258
rect 9251 70 9309 82
rect 9369 258 9427 270
rect 9369 82 9381 258
rect 9415 82 9427 258
rect 9369 70 9427 82
rect 9487 258 9545 270
rect 9487 82 9499 258
rect 9533 82 9545 258
rect 9487 70 9545 82
rect 9605 258 9663 270
rect 9605 82 9617 258
rect 9651 82 9663 258
rect 9605 70 9663 82
rect 9723 258 9781 270
rect 9723 82 9735 258
rect 9769 82 9781 258
rect 9723 70 9781 82
rect 9841 258 9899 270
rect 9841 82 9853 258
rect 9887 82 9899 258
rect 9841 70 9899 82
rect 9959 258 10017 270
rect 9959 82 9971 258
rect 10005 82 10017 258
rect 9959 70 10017 82
rect 10345 258 10403 270
rect 10345 82 10357 258
rect 10391 82 10403 258
rect 10345 70 10403 82
rect 10463 258 10521 270
rect 10463 82 10475 258
rect 10509 82 10521 258
rect 10463 70 10521 82
rect 10581 258 10639 270
rect 10581 82 10593 258
rect 10627 82 10639 258
rect 10581 70 10639 82
rect 10699 258 10757 270
rect 10699 82 10711 258
rect 10745 82 10757 258
rect 10699 70 10757 82
rect 10817 258 10875 270
rect 10817 82 10829 258
rect 10863 82 10875 258
rect 10817 70 10875 82
rect 10935 258 10993 270
rect 10935 82 10947 258
rect 10981 82 10993 258
rect 10935 70 10993 82
rect 11053 258 11111 270
rect 11053 82 11065 258
rect 11099 82 11111 258
rect 11053 70 11111 82
rect 11171 258 11229 270
rect 11171 82 11183 258
rect 11217 82 11229 258
rect 11171 70 11229 82
rect 11289 258 11347 270
rect 11289 82 11301 258
rect 11335 82 11347 258
rect 11289 70 11347 82
rect 11407 258 11465 270
rect 11407 82 11419 258
rect 11453 82 11465 258
rect 11407 70 11465 82
<< ndiffc >>
rect 286 -557 320 -181
rect 404 -557 438 -181
rect 522 -557 556 -181
rect 639 -357 673 -181
rect 757 -357 791 -181
rect 1734 -557 1768 -181
rect 1852 -557 1886 -181
rect 1970 -557 2004 -181
rect 2087 -357 2121 -181
rect 2205 -357 2239 -181
rect 3232 -555 3266 -179
rect 3350 -555 3384 -179
rect 3468 -555 3502 -179
rect 3585 -355 3619 -179
rect 3703 -355 3737 -179
rect 4680 -555 4714 -179
rect 4798 -555 4832 -179
rect 4916 -555 4950 -179
rect 5033 -355 5067 -179
rect 5151 -355 5185 -179
rect 6200 -557 6234 -181
rect 6318 -557 6352 -181
rect 6436 -557 6470 -181
rect 6553 -357 6587 -181
rect 6671 -357 6705 -181
rect 7648 -557 7682 -181
rect 7766 -557 7800 -181
rect 7884 -557 7918 -181
rect 8001 -357 8035 -181
rect 8119 -357 8153 -181
rect 9146 -555 9180 -179
rect 9264 -555 9298 -179
rect 9382 -555 9416 -179
rect 9499 -355 9533 -179
rect 9617 -355 9651 -179
rect 10594 -555 10628 -179
rect 10712 -555 10746 -179
rect 10830 -555 10864 -179
rect 10947 -355 10981 -179
rect 11065 -355 11099 -179
<< pdiffc >>
rect 49 80 83 256
rect 167 80 201 256
rect 285 80 319 256
rect 403 80 437 256
rect 521 80 555 256
rect 639 80 673 256
rect 757 80 791 256
rect 875 80 909 256
rect 993 80 1027 256
rect 1111 80 1145 256
rect 1497 80 1531 256
rect 1615 80 1649 256
rect 1733 80 1767 256
rect 1851 80 1885 256
rect 1969 80 2003 256
rect 2087 80 2121 256
rect 2205 80 2239 256
rect 2323 80 2357 256
rect 2441 80 2475 256
rect 2559 80 2593 256
rect 2995 82 3029 258
rect 3113 82 3147 258
rect 3231 82 3265 258
rect 3349 82 3383 258
rect 3467 82 3501 258
rect 3585 82 3619 258
rect 3703 82 3737 258
rect 3821 82 3855 258
rect 3939 82 3973 258
rect 4057 82 4091 258
rect 4443 82 4477 258
rect 4561 82 4595 258
rect 4679 82 4713 258
rect 4797 82 4831 258
rect 4915 82 4949 258
rect 5033 82 5067 258
rect 5151 82 5185 258
rect 5269 82 5303 258
rect 5387 82 5421 258
rect 5505 82 5539 258
rect 5963 80 5997 256
rect 6081 80 6115 256
rect 6199 80 6233 256
rect 6317 80 6351 256
rect 6435 80 6469 256
rect 6553 80 6587 256
rect 6671 80 6705 256
rect 6789 80 6823 256
rect 6907 80 6941 256
rect 7025 80 7059 256
rect 7411 80 7445 256
rect 7529 80 7563 256
rect 7647 80 7681 256
rect 7765 80 7799 256
rect 7883 80 7917 256
rect 8001 80 8035 256
rect 8119 80 8153 256
rect 8237 80 8271 256
rect 8355 80 8389 256
rect 8473 80 8507 256
rect 8909 82 8943 258
rect 9027 82 9061 258
rect 9145 82 9179 258
rect 9263 82 9297 258
rect 9381 82 9415 258
rect 9499 82 9533 258
rect 9617 82 9651 258
rect 9735 82 9769 258
rect 9853 82 9887 258
rect 9971 82 10005 258
rect 10357 82 10391 258
rect 10475 82 10509 258
rect 10593 82 10627 258
rect 10711 82 10745 258
rect 10829 82 10863 258
rect 10947 82 10981 258
rect 11065 82 11099 258
rect 11183 82 11217 258
rect 11301 82 11335 258
rect 11419 82 11453 258
<< psubdiff >>
rect 538 -712 750 -682
rect 538 -768 578 -712
rect 712 -768 750 -712
rect 538 -790 750 -768
rect 1986 -712 2198 -682
rect 1986 -768 2026 -712
rect 2160 -768 2198 -712
rect 1986 -790 2198 -768
rect 3484 -710 3696 -680
rect 3484 -766 3524 -710
rect 3658 -766 3696 -710
rect 3484 -788 3696 -766
rect 4932 -710 5144 -680
rect 4932 -766 4972 -710
rect 5106 -766 5144 -710
rect 4932 -788 5144 -766
rect 6452 -712 6664 -682
rect 6452 -768 6492 -712
rect 6626 -768 6664 -712
rect 6452 -790 6664 -768
rect 7900 -712 8112 -682
rect 7900 -768 7940 -712
rect 8074 -768 8112 -712
rect 7900 -790 8112 -768
rect 9398 -710 9610 -680
rect 9398 -766 9438 -710
rect 9572 -766 9610 -710
rect 9398 -788 9610 -766
rect 10846 -710 11058 -680
rect 10846 -766 10886 -710
rect 11020 -766 11058 -710
rect 10846 -788 11058 -766
<< nsubdiff >>
rect 298 496 542 534
rect 298 426 354 496
rect 490 426 542 496
rect 298 404 542 426
rect 1746 496 1990 534
rect 1746 426 1802 496
rect 1938 426 1990 496
rect 1746 404 1990 426
rect 3244 498 3488 536
rect 3244 428 3300 498
rect 3436 428 3488 498
rect 3244 406 3488 428
rect 4692 498 4936 536
rect 4692 428 4748 498
rect 4884 428 4936 498
rect 4692 406 4936 428
rect 6212 496 6456 534
rect 6212 426 6268 496
rect 6404 426 6456 496
rect 6212 404 6456 426
rect 7660 496 7904 534
rect 7660 426 7716 496
rect 7852 426 7904 496
rect 7660 404 7904 426
rect 9158 498 9402 536
rect 9158 428 9214 498
rect 9350 428 9402 498
rect 9158 406 9402 428
rect 10606 498 10850 536
rect 10606 428 10662 498
rect 10798 428 10850 498
rect 10606 406 10850 428
<< psubdiffcont >>
rect 578 -768 712 -712
rect 2026 -768 2160 -712
rect 3524 -766 3658 -710
rect 4972 -766 5106 -710
rect 6492 -768 6626 -712
rect 7940 -768 8074 -712
rect 9438 -766 9572 -710
rect 10886 -766 11020 -710
<< nsubdiffcont >>
rect 354 426 490 496
rect 1802 426 1938 496
rect 3300 428 3436 498
rect 4748 428 4884 498
rect 6268 426 6404 496
rect 7716 426 7852 496
rect 9214 428 9350 498
rect 10662 428 10798 498
<< poly >>
rect 95 289 391 325
rect 95 268 155 289
rect 213 268 273 289
rect 331 268 391 289
rect 449 288 745 324
rect 449 268 509 288
rect 567 268 627 288
rect 685 268 745 288
rect 803 288 1099 324
rect 803 268 863 288
rect 921 268 981 288
rect 1039 268 1099 288
rect 1543 289 1839 325
rect 1543 268 1603 289
rect 1661 268 1721 289
rect 1779 268 1839 289
rect 1897 288 2193 324
rect 1897 268 1957 288
rect 2015 268 2075 288
rect 2133 268 2193 288
rect 2251 288 2547 324
rect 2251 268 2311 288
rect 2369 268 2429 288
rect 2487 268 2547 288
rect 3041 291 3337 327
rect 3041 270 3101 291
rect 3159 270 3219 291
rect 3277 270 3337 291
rect 3395 290 3691 326
rect 3395 270 3455 290
rect 3513 270 3573 290
rect 3631 270 3691 290
rect 3749 290 4045 326
rect 3749 270 3809 290
rect 3867 270 3927 290
rect 3985 270 4045 290
rect 4489 291 4785 327
rect 4489 270 4549 291
rect 4607 270 4667 291
rect 4725 270 4785 291
rect 4843 290 5139 326
rect 4843 270 4903 290
rect 4961 270 5021 290
rect 5079 270 5139 290
rect 5197 290 5493 326
rect 5197 270 5257 290
rect 5315 270 5375 290
rect 5433 270 5493 290
rect 6009 289 6305 325
rect 6009 268 6069 289
rect 6127 268 6187 289
rect 6245 268 6305 289
rect 6363 288 6659 324
rect 6363 268 6423 288
rect 6481 268 6541 288
rect 6599 268 6659 288
rect 6717 288 7013 324
rect 6717 268 6777 288
rect 6835 268 6895 288
rect 6953 268 7013 288
rect 7457 289 7753 325
rect 7457 268 7517 289
rect 7575 268 7635 289
rect 7693 268 7753 289
rect 7811 288 8107 324
rect 7811 268 7871 288
rect 7929 268 7989 288
rect 8047 268 8107 288
rect 8165 288 8461 324
rect 8165 268 8225 288
rect 8283 268 8343 288
rect 8401 268 8461 288
rect 8955 291 9251 327
rect 8955 270 9015 291
rect 9073 270 9133 291
rect 9191 270 9251 291
rect 9309 290 9605 326
rect 9309 270 9369 290
rect 9427 270 9487 290
rect 9545 270 9605 290
rect 9663 290 9959 326
rect 9663 270 9723 290
rect 9781 270 9841 290
rect 9899 270 9959 290
rect 10403 291 10699 327
rect 10403 270 10463 291
rect 10521 270 10581 291
rect 10639 270 10699 291
rect 10757 290 11053 326
rect 10757 270 10817 290
rect 10875 270 10935 290
rect 10993 270 11053 290
rect 11111 290 11407 326
rect 11111 270 11171 290
rect 11229 270 11289 290
rect 11347 270 11407 290
rect 95 42 155 68
rect 213 42 273 68
rect 331 42 391 68
rect 449 48 509 68
rect 449 42 510 48
rect 567 42 627 68
rect 685 42 745 68
rect 332 -143 390 42
rect 332 -169 392 -143
rect 450 -169 510 42
rect 803 36 863 68
rect 921 42 981 68
rect 1039 42 1099 68
rect 1543 42 1603 68
rect 1661 42 1721 68
rect 1779 42 1839 68
rect 1897 48 1957 68
rect 1897 42 1958 48
rect 2015 42 2075 68
rect 2133 42 2193 68
rect 800 20 866 36
rect 800 -14 816 20
rect 850 -14 866 20
rect 800 -30 866 -14
rect 682 -97 748 -81
rect 682 -131 698 -97
rect 732 -131 748 -97
rect 682 -147 748 -131
rect 1780 -143 1838 42
rect 685 -169 745 -147
rect 1780 -169 1840 -143
rect 1898 -169 1958 42
rect 2251 36 2311 68
rect 2369 42 2429 68
rect 2487 42 2547 68
rect 3041 44 3101 70
rect 3159 44 3219 70
rect 3277 44 3337 70
rect 3395 50 3455 70
rect 3395 44 3456 50
rect 3513 44 3573 70
rect 3631 44 3691 70
rect 2248 20 2314 36
rect 2248 -14 2264 20
rect 2298 -14 2314 20
rect 2248 -30 2314 -14
rect 2130 -97 2196 -81
rect 2130 -131 2146 -97
rect 2180 -131 2196 -97
rect 2130 -147 2196 -131
rect 3278 -141 3336 44
rect 2133 -169 2193 -147
rect 3278 -167 3338 -141
rect 3396 -167 3456 44
rect 3749 38 3809 70
rect 3867 44 3927 70
rect 3985 44 4045 70
rect 4489 44 4549 70
rect 4607 44 4667 70
rect 4725 44 4785 70
rect 4843 50 4903 70
rect 4843 44 4904 50
rect 4961 44 5021 70
rect 5079 44 5139 70
rect 3746 22 3812 38
rect 3746 -12 3762 22
rect 3796 -12 3812 22
rect 3746 -28 3812 -12
rect 3628 -95 3694 -79
rect 3628 -129 3644 -95
rect 3678 -129 3694 -95
rect 3628 -145 3694 -129
rect 4726 -141 4784 44
rect 3631 -167 3691 -145
rect 4726 -167 4786 -141
rect 4844 -167 4904 44
rect 5197 38 5257 70
rect 5315 44 5375 70
rect 5433 44 5493 70
rect 6009 42 6069 68
rect 6127 42 6187 68
rect 6245 42 6305 68
rect 6363 48 6423 68
rect 6363 42 6424 48
rect 6481 42 6541 68
rect 6599 42 6659 68
rect 5194 22 5260 38
rect 5194 -12 5210 22
rect 5244 -12 5260 22
rect 5194 -28 5260 -12
rect 5076 -95 5142 -79
rect 5076 -129 5092 -95
rect 5126 -129 5142 -95
rect 5076 -145 5142 -129
rect 6246 -143 6304 42
rect 5079 -167 5139 -145
rect 685 -395 745 -369
rect 2133 -395 2193 -369
rect 3631 -393 3691 -367
rect 6246 -169 6306 -143
rect 6364 -169 6424 42
rect 6717 36 6777 68
rect 6835 42 6895 68
rect 6953 42 7013 68
rect 7457 42 7517 68
rect 7575 42 7635 68
rect 7693 42 7753 68
rect 7811 48 7871 68
rect 7811 42 7872 48
rect 7929 42 7989 68
rect 8047 42 8107 68
rect 6714 20 6780 36
rect 6714 -14 6730 20
rect 6764 -14 6780 20
rect 6714 -30 6780 -14
rect 6596 -97 6662 -81
rect 6596 -131 6612 -97
rect 6646 -131 6662 -97
rect 6596 -147 6662 -131
rect 7694 -143 7752 42
rect 6599 -169 6659 -147
rect 7694 -169 7754 -143
rect 7812 -169 7872 42
rect 8165 36 8225 68
rect 8283 42 8343 68
rect 8401 42 8461 68
rect 8955 44 9015 70
rect 9073 44 9133 70
rect 9191 44 9251 70
rect 9309 50 9369 70
rect 9309 44 9370 50
rect 9427 44 9487 70
rect 9545 44 9605 70
rect 8162 20 8228 36
rect 8162 -14 8178 20
rect 8212 -14 8228 20
rect 8162 -30 8228 -14
rect 8044 -97 8110 -81
rect 8044 -131 8060 -97
rect 8094 -131 8110 -97
rect 8044 -147 8110 -131
rect 9192 -141 9250 44
rect 8047 -169 8107 -147
rect 9192 -167 9252 -141
rect 9310 -167 9370 44
rect 9663 38 9723 70
rect 9781 44 9841 70
rect 9899 44 9959 70
rect 10403 44 10463 70
rect 10521 44 10581 70
rect 10639 44 10699 70
rect 10757 50 10817 70
rect 10757 44 10818 50
rect 10875 44 10935 70
rect 10993 44 11053 70
rect 9660 22 9726 38
rect 9660 -12 9676 22
rect 9710 -12 9726 22
rect 9660 -28 9726 -12
rect 9542 -95 9608 -79
rect 9542 -129 9558 -95
rect 9592 -129 9608 -95
rect 9542 -145 9608 -129
rect 10640 -141 10698 44
rect 9545 -167 9605 -145
rect 10640 -167 10700 -141
rect 10758 -167 10818 44
rect 11111 38 11171 70
rect 11229 44 11289 70
rect 11347 44 11407 70
rect 11108 22 11174 38
rect 11108 -12 11124 22
rect 11158 -12 11174 22
rect 11108 -28 11174 -12
rect 10990 -95 11056 -79
rect 10990 -129 11006 -95
rect 11040 -129 11056 -95
rect 10990 -145 11056 -129
rect 10993 -167 11053 -145
rect 5079 -393 5139 -367
rect 332 -591 392 -569
rect 450 -591 510 -569
rect 1780 -591 1840 -569
rect 1898 -591 1958 -569
rect 3278 -589 3338 -567
rect 3396 -589 3456 -567
rect 4726 -589 4786 -567
rect 4844 -589 4904 -567
rect 6599 -395 6659 -369
rect 8047 -395 8107 -369
rect 9545 -393 9605 -367
rect 10993 -393 11053 -367
rect 329 -607 395 -591
rect 329 -641 345 -607
rect 379 -641 395 -607
rect 329 -657 395 -641
rect 447 -607 513 -591
rect 447 -641 463 -607
rect 497 -641 513 -607
rect 447 -657 513 -641
rect 1777 -607 1843 -591
rect 1777 -641 1793 -607
rect 1827 -641 1843 -607
rect 1777 -657 1843 -641
rect 1895 -607 1961 -591
rect 1895 -641 1911 -607
rect 1945 -641 1961 -607
rect 1895 -657 1961 -641
rect 3275 -605 3341 -589
rect 3275 -639 3291 -605
rect 3325 -639 3341 -605
rect 3275 -655 3341 -639
rect 3393 -605 3459 -589
rect 3393 -639 3409 -605
rect 3443 -639 3459 -605
rect 3393 -655 3459 -639
rect 4723 -605 4789 -589
rect 4723 -639 4739 -605
rect 4773 -639 4789 -605
rect 4723 -655 4789 -639
rect 4841 -605 4907 -589
rect 6246 -591 6306 -569
rect 6364 -591 6424 -569
rect 7694 -591 7754 -569
rect 7812 -591 7872 -569
rect 9192 -589 9252 -567
rect 9310 -589 9370 -567
rect 10640 -589 10700 -567
rect 10758 -589 10818 -567
rect 4841 -639 4857 -605
rect 4891 -639 4907 -605
rect 4841 -655 4907 -639
rect 6243 -607 6309 -591
rect 6243 -641 6259 -607
rect 6293 -641 6309 -607
rect 6243 -657 6309 -641
rect 6361 -607 6427 -591
rect 6361 -641 6377 -607
rect 6411 -641 6427 -607
rect 6361 -657 6427 -641
rect 7691 -607 7757 -591
rect 7691 -641 7707 -607
rect 7741 -641 7757 -607
rect 7691 -657 7757 -641
rect 7809 -607 7875 -591
rect 7809 -641 7825 -607
rect 7859 -641 7875 -607
rect 7809 -657 7875 -641
rect 9189 -605 9255 -589
rect 9189 -639 9205 -605
rect 9239 -639 9255 -605
rect 9189 -655 9255 -639
rect 9307 -605 9373 -589
rect 9307 -639 9323 -605
rect 9357 -639 9373 -605
rect 9307 -655 9373 -639
rect 10637 -605 10703 -589
rect 10637 -639 10653 -605
rect 10687 -639 10703 -605
rect 10637 -655 10703 -639
rect 10755 -605 10821 -589
rect 10755 -639 10771 -605
rect 10805 -639 10821 -605
rect 10755 -655 10821 -639
<< polycont >>
rect 816 -14 850 20
rect 698 -131 732 -97
rect 2264 -14 2298 20
rect 2146 -131 2180 -97
rect 3762 -12 3796 22
rect 3644 -129 3678 -95
rect 5210 -12 5244 22
rect 5092 -129 5126 -95
rect 6730 -14 6764 20
rect 6612 -131 6646 -97
rect 8178 -14 8212 20
rect 8060 -131 8094 -97
rect 9676 -12 9710 22
rect 9558 -129 9592 -95
rect 11124 -12 11158 22
rect 11006 -129 11040 -95
rect 345 -641 379 -607
rect 463 -641 497 -607
rect 1793 -641 1827 -607
rect 1911 -641 1945 -607
rect 3291 -639 3325 -605
rect 3409 -639 3443 -605
rect 4739 -639 4773 -605
rect 4857 -639 4891 -605
rect 6259 -641 6293 -607
rect 6377 -641 6411 -607
rect 7707 -641 7741 -607
rect 7825 -641 7859 -607
rect 9205 -639 9239 -605
rect 9323 -639 9357 -605
rect 10653 -639 10687 -605
rect 10771 -639 10805 -605
<< locali >>
rect 338 496 506 512
rect 338 426 354 496
rect 490 426 506 496
rect 338 410 506 426
rect 1786 496 1954 512
rect 1786 426 1802 496
rect 1938 426 1954 496
rect 1786 410 1954 426
rect 3284 498 3452 514
rect 3284 428 3300 498
rect 3436 428 3452 498
rect 3284 412 3452 428
rect 4732 498 4900 514
rect 4732 428 4748 498
rect 4884 428 4900 498
rect 4732 412 4900 428
rect 6252 496 6420 512
rect 6252 426 6268 496
rect 6404 426 6420 496
rect 6252 410 6420 426
rect 7700 496 7868 512
rect 7700 426 7716 496
rect 7852 426 7868 496
rect 7700 410 7868 426
rect 9198 498 9366 514
rect 9198 428 9214 498
rect 9350 428 9366 498
rect 9198 412 9366 428
rect 10646 498 10814 514
rect 10646 428 10662 498
rect 10798 428 10814 498
rect 10646 412 10814 428
rect 875 306 1145 340
rect 49 256 83 272
rect 49 64 83 80
rect 167 256 201 272
rect 167 64 201 80
rect 285 256 319 272
rect 285 64 319 80
rect 403 256 437 272
rect 403 64 437 80
rect 521 256 555 272
rect 521 64 555 80
rect 639 256 673 272
rect 639 64 673 80
rect 757 256 791 272
rect 757 64 791 80
rect 875 256 909 306
rect 875 64 909 80
rect 993 256 1027 272
rect 993 64 1027 80
rect 1111 256 1145 306
rect 2323 306 2593 340
rect 1111 64 1145 80
rect 1497 256 1531 272
rect 1497 64 1531 80
rect 1615 256 1649 272
rect 1615 64 1649 80
rect 1733 256 1767 272
rect 1733 64 1767 80
rect 1851 256 1885 272
rect 1851 64 1885 80
rect 1969 256 2003 272
rect 1969 64 2003 80
rect 2087 256 2121 272
rect 2087 64 2121 80
rect 2205 256 2239 272
rect 2205 64 2239 80
rect 2323 256 2357 306
rect 2323 64 2357 80
rect 2441 256 2475 272
rect 2441 64 2475 80
rect 2559 256 2593 306
rect 3821 308 4091 342
rect 2559 64 2593 80
rect 2995 258 3029 274
rect 2995 66 3029 82
rect 3113 258 3147 274
rect 3113 66 3147 82
rect 3231 258 3265 274
rect 3231 66 3265 82
rect 3349 258 3383 274
rect 3349 66 3383 82
rect 3467 258 3501 274
rect 3467 66 3501 82
rect 3585 258 3619 274
rect 3585 66 3619 82
rect 3703 258 3737 274
rect 3703 66 3737 82
rect 3821 258 3855 308
rect 3821 66 3855 82
rect 3939 258 3973 274
rect 3939 66 3973 82
rect 4057 258 4091 308
rect 5269 308 5539 342
rect 4057 66 4091 82
rect 4443 258 4477 274
rect 4443 66 4477 82
rect 4561 258 4595 274
rect 4561 66 4595 82
rect 4679 258 4713 274
rect 4679 66 4713 82
rect 4797 258 4831 274
rect 4797 66 4831 82
rect 4915 258 4949 274
rect 4915 66 4949 82
rect 5033 258 5067 274
rect 5033 66 5067 82
rect 5151 258 5185 274
rect 5151 66 5185 82
rect 5269 258 5303 308
rect 5269 66 5303 82
rect 5387 258 5421 274
rect 5387 66 5421 82
rect 5505 258 5539 308
rect 6789 306 7059 340
rect 5505 66 5539 82
rect 5963 256 5997 272
rect 5963 64 5997 80
rect 6081 256 6115 272
rect 6081 64 6115 80
rect 6199 256 6233 272
rect 6199 64 6233 80
rect 6317 256 6351 272
rect 6317 64 6351 80
rect 6435 256 6469 272
rect 6435 64 6469 80
rect 6553 256 6587 272
rect 6553 64 6587 80
rect 6671 256 6705 272
rect 6671 64 6705 80
rect 6789 256 6823 306
rect 6789 64 6823 80
rect 6907 256 6941 272
rect 6907 64 6941 80
rect 7025 256 7059 306
rect 8237 306 8507 340
rect 7025 64 7059 80
rect 7411 256 7445 272
rect 7411 64 7445 80
rect 7529 256 7563 272
rect 7529 64 7563 80
rect 7647 256 7681 272
rect 7647 64 7681 80
rect 7765 256 7799 272
rect 7765 64 7799 80
rect 7883 256 7917 272
rect 7883 64 7917 80
rect 8001 256 8035 272
rect 8001 64 8035 80
rect 8119 256 8153 272
rect 8119 64 8153 80
rect 8237 256 8271 306
rect 8237 64 8271 80
rect 8355 256 8389 272
rect 8355 64 8389 80
rect 8473 256 8507 306
rect 9735 308 10005 342
rect 8473 64 8507 80
rect 8909 258 8943 274
rect 8909 66 8943 82
rect 9027 258 9061 274
rect 9027 66 9061 82
rect 9145 258 9179 274
rect 9145 66 9179 82
rect 9263 258 9297 274
rect 9263 66 9297 82
rect 9381 258 9415 274
rect 9381 66 9415 82
rect 9499 258 9533 274
rect 9499 66 9533 82
rect 9617 258 9651 274
rect 9617 66 9651 82
rect 9735 258 9769 308
rect 9735 66 9769 82
rect 9853 258 9887 274
rect 9853 66 9887 82
rect 9971 258 10005 308
rect 11183 308 11453 342
rect 9971 66 10005 82
rect 10357 258 10391 274
rect 10357 66 10391 82
rect 10475 258 10509 274
rect 10475 66 10509 82
rect 10593 258 10627 274
rect 10593 66 10627 82
rect 10711 258 10745 274
rect 10711 66 10745 82
rect 10829 258 10863 274
rect 10829 66 10863 82
rect 10947 258 10981 274
rect 10947 66 10981 82
rect 11065 258 11099 274
rect 11065 66 11099 82
rect 11183 258 11217 308
rect 11183 66 11217 82
rect 11301 258 11335 274
rect 11301 66 11335 82
rect 11419 258 11453 308
rect 11419 66 11453 82
rect 800 -14 816 20
rect 850 -14 866 20
rect 2248 -14 2264 20
rect 2298 -14 2314 20
rect 3746 -12 3762 22
rect 3796 -12 3812 22
rect 5194 -12 5210 22
rect 5244 -12 5260 22
rect 6714 -14 6730 20
rect 6764 -14 6780 20
rect 8162 -14 8178 20
rect 8212 -14 8228 20
rect 9660 -12 9676 22
rect 9710 -12 9726 22
rect 11108 -12 11124 22
rect 11158 -12 11174 22
rect 682 -131 698 -97
rect 732 -131 748 -97
rect 2130 -131 2146 -97
rect 2180 -131 2196 -97
rect 3628 -129 3644 -95
rect 3678 -129 3694 -95
rect 5076 -129 5092 -95
rect 5126 -129 5142 -95
rect 6596 -131 6612 -97
rect 6646 -131 6662 -97
rect 8044 -131 8060 -97
rect 8094 -131 8110 -97
rect 9542 -129 9558 -95
rect 9592 -129 9608 -95
rect 10990 -129 11006 -95
rect 11040 -129 11056 -95
rect 286 -181 320 -165
rect 286 -573 320 -557
rect 404 -181 438 -165
rect 404 -573 438 -557
rect 522 -181 556 -165
rect 639 -181 673 -165
rect 639 -373 673 -357
rect 757 -181 791 -165
rect 757 -373 791 -357
rect 1734 -181 1768 -165
rect 522 -573 556 -557
rect 1734 -573 1768 -557
rect 1852 -181 1886 -165
rect 1852 -573 1886 -557
rect 1970 -181 2004 -165
rect 2087 -181 2121 -165
rect 2087 -373 2121 -357
rect 2205 -181 2239 -165
rect 2205 -373 2239 -357
rect 3232 -179 3266 -163
rect 1970 -573 2004 -557
rect 3232 -571 3266 -555
rect 3350 -179 3384 -163
rect 3350 -571 3384 -555
rect 3468 -179 3502 -163
rect 3585 -179 3619 -163
rect 3585 -371 3619 -355
rect 3703 -179 3737 -163
rect 3703 -371 3737 -355
rect 4680 -179 4714 -163
rect 3468 -571 3502 -555
rect 4680 -571 4714 -555
rect 4798 -179 4832 -163
rect 4798 -571 4832 -555
rect 4916 -179 4950 -163
rect 5033 -179 5067 -163
rect 5033 -371 5067 -355
rect 5151 -179 5185 -163
rect 5151 -371 5185 -355
rect 6200 -181 6234 -165
rect 4916 -571 4950 -555
rect 6200 -573 6234 -557
rect 6318 -181 6352 -165
rect 6318 -573 6352 -557
rect 6436 -181 6470 -165
rect 6553 -181 6587 -165
rect 6553 -373 6587 -357
rect 6671 -181 6705 -165
rect 6671 -373 6705 -357
rect 7648 -181 7682 -165
rect 6436 -573 6470 -557
rect 7648 -573 7682 -557
rect 7766 -181 7800 -165
rect 7766 -573 7800 -557
rect 7884 -181 7918 -165
rect 8001 -181 8035 -165
rect 8001 -373 8035 -357
rect 8119 -181 8153 -165
rect 8119 -373 8153 -357
rect 9146 -179 9180 -163
rect 7884 -573 7918 -557
rect 9146 -571 9180 -555
rect 9264 -179 9298 -163
rect 9264 -571 9298 -555
rect 9382 -179 9416 -163
rect 9499 -179 9533 -163
rect 9499 -371 9533 -355
rect 9617 -179 9651 -163
rect 9617 -371 9651 -355
rect 10594 -179 10628 -163
rect 9382 -571 9416 -555
rect 10594 -571 10628 -555
rect 10712 -179 10746 -163
rect 10712 -571 10746 -555
rect 10830 -179 10864 -163
rect 10947 -179 10981 -163
rect 10947 -371 10981 -355
rect 11065 -179 11099 -163
rect 11065 -371 11099 -355
rect 10830 -571 10864 -555
rect 329 -641 345 -607
rect 379 -641 395 -607
rect 447 -641 463 -607
rect 497 -641 513 -607
rect 1777 -641 1793 -607
rect 1827 -641 1843 -607
rect 1895 -641 1911 -607
rect 1945 -641 1961 -607
rect 3275 -639 3291 -605
rect 3325 -639 3341 -605
rect 3393 -639 3409 -605
rect 3443 -639 3459 -605
rect 4723 -639 4739 -605
rect 4773 -639 4789 -605
rect 4841 -639 4857 -605
rect 4891 -639 4907 -605
rect 6243 -641 6259 -607
rect 6293 -641 6309 -607
rect 6361 -641 6377 -607
rect 6411 -641 6427 -607
rect 7691 -641 7707 -607
rect 7741 -641 7757 -607
rect 7809 -641 7825 -607
rect 7859 -641 7875 -607
rect 9189 -639 9205 -605
rect 9239 -639 9255 -605
rect 9307 -639 9323 -605
rect 9357 -639 9373 -605
rect 10637 -639 10653 -605
rect 10687 -639 10703 -605
rect 10755 -639 10771 -605
rect 10805 -639 10821 -605
rect 562 -712 730 -694
rect 562 -768 578 -712
rect 712 -768 730 -712
rect 562 -784 730 -768
rect 2010 -712 2178 -694
rect 2010 -768 2026 -712
rect 2160 -768 2178 -712
rect 2010 -784 2178 -768
rect 3508 -710 3676 -692
rect 3508 -766 3524 -710
rect 3658 -766 3676 -710
rect 3508 -782 3676 -766
rect 4956 -710 5124 -692
rect 4956 -766 4972 -710
rect 5106 -766 5124 -710
rect 4956 -782 5124 -766
rect 6476 -712 6644 -694
rect 6476 -768 6492 -712
rect 6626 -768 6644 -712
rect 6476 -784 6644 -768
rect 7924 -712 8092 -694
rect 7924 -768 7940 -712
rect 8074 -768 8092 -712
rect 7924 -784 8092 -768
rect 9422 -710 9590 -692
rect 9422 -766 9438 -710
rect 9572 -766 9590 -710
rect 9422 -782 9590 -766
rect 10870 -710 11038 -692
rect 10870 -766 10886 -710
rect 11020 -766 11038 -710
rect 10870 -782 11038 -766
<< viali >>
rect 390 432 450 494
rect 1838 432 1898 494
rect 3336 434 3396 496
rect 4784 434 4844 496
rect 6304 432 6364 494
rect 7752 432 7812 494
rect 9250 434 9310 496
rect 10698 434 10758 496
rect 49 80 83 256
rect 167 80 201 256
rect 285 80 319 256
rect 403 80 437 256
rect 521 80 555 256
rect 639 80 673 256
rect 757 80 791 256
rect 875 80 909 256
rect 993 80 1027 256
rect 1111 80 1145 256
rect 1497 80 1531 256
rect 1615 80 1649 256
rect 1733 80 1767 256
rect 1851 80 1885 256
rect 1969 80 2003 256
rect 2087 80 2121 256
rect 2205 80 2239 256
rect 2323 80 2357 256
rect 2441 80 2475 256
rect 2559 80 2593 256
rect 2995 82 3029 258
rect 3113 82 3147 258
rect 3231 82 3265 258
rect 3349 82 3383 258
rect 3467 82 3501 258
rect 3585 82 3619 258
rect 3703 82 3737 258
rect 3821 82 3855 258
rect 3939 82 3973 258
rect 4057 82 4091 258
rect 4443 82 4477 258
rect 4561 82 4595 258
rect 4679 82 4713 258
rect 4797 82 4831 258
rect 4915 82 4949 258
rect 5033 82 5067 258
rect 5151 82 5185 258
rect 5269 82 5303 258
rect 5387 82 5421 258
rect 5505 82 5539 258
rect 5963 80 5997 256
rect 6081 80 6115 256
rect 6199 80 6233 256
rect 6317 80 6351 256
rect 6435 80 6469 256
rect 6553 80 6587 256
rect 6671 80 6705 256
rect 6789 80 6823 256
rect 6907 80 6941 256
rect 7025 80 7059 256
rect 7411 80 7445 256
rect 7529 80 7563 256
rect 7647 80 7681 256
rect 7765 80 7799 256
rect 7883 80 7917 256
rect 8001 80 8035 256
rect 8119 80 8153 256
rect 8237 80 8271 256
rect 8355 80 8389 256
rect 8473 80 8507 256
rect 8909 82 8943 258
rect 9027 82 9061 258
rect 9145 82 9179 258
rect 9263 82 9297 258
rect 9381 82 9415 258
rect 9499 82 9533 258
rect 9617 82 9651 258
rect 9735 82 9769 258
rect 9853 82 9887 258
rect 9971 82 10005 258
rect 10357 82 10391 258
rect 10475 82 10509 258
rect 10593 82 10627 258
rect 10711 82 10745 258
rect 10829 82 10863 258
rect 10947 82 10981 258
rect 11065 82 11099 258
rect 11183 82 11217 258
rect 11301 82 11335 258
rect 11419 82 11453 258
rect 816 -14 850 20
rect 2264 -14 2298 20
rect 3762 -12 3796 22
rect 5210 -12 5244 22
rect 6730 -14 6764 20
rect 8178 -14 8212 20
rect 9676 -12 9710 22
rect 11124 -12 11158 22
rect 698 -131 732 -97
rect 2146 -131 2180 -97
rect 3644 -129 3678 -95
rect 5092 -129 5126 -95
rect 6612 -131 6646 -97
rect 8060 -131 8094 -97
rect 9558 -129 9592 -95
rect 11006 -129 11040 -95
rect 286 -557 320 -181
rect 404 -557 438 -181
rect 522 -557 556 -181
rect 639 -357 673 -181
rect 757 -357 791 -181
rect 1734 -557 1768 -181
rect 1852 -557 1886 -181
rect 1970 -557 2004 -181
rect 2087 -357 2121 -181
rect 2205 -357 2239 -181
rect 3232 -555 3266 -179
rect 3350 -555 3384 -179
rect 3468 -555 3502 -179
rect 3585 -355 3619 -179
rect 3703 -355 3737 -179
rect 4680 -555 4714 -179
rect 4798 -555 4832 -179
rect 4916 -555 4950 -179
rect 5033 -355 5067 -179
rect 5151 -355 5185 -179
rect 6200 -557 6234 -181
rect 6318 -557 6352 -181
rect 6436 -557 6470 -181
rect 6553 -357 6587 -181
rect 6671 -357 6705 -181
rect 7648 -557 7682 -181
rect 7766 -557 7800 -181
rect 7884 -557 7918 -181
rect 8001 -357 8035 -181
rect 8119 -357 8153 -181
rect 9146 -555 9180 -179
rect 9264 -555 9298 -179
rect 9382 -555 9416 -179
rect 9499 -355 9533 -179
rect 9617 -355 9651 -179
rect 10594 -555 10628 -179
rect 10712 -555 10746 -179
rect 10830 -555 10864 -179
rect 10947 -355 10981 -179
rect 11065 -355 11099 -179
rect 345 -641 379 -607
rect 463 -641 497 -607
rect 1793 -641 1827 -607
rect 1911 -641 1945 -607
rect 3291 -639 3325 -605
rect 3409 -639 3443 -605
rect 4739 -639 4773 -605
rect 4857 -639 4891 -605
rect 6259 -641 6293 -607
rect 6377 -641 6411 -607
rect 7707 -641 7741 -607
rect 7825 -641 7859 -607
rect 9205 -639 9239 -605
rect 9323 -639 9357 -605
rect 10653 -639 10687 -605
rect 10771 -639 10805 -605
rect 618 -764 670 -718
rect 2066 -764 2118 -718
rect 3564 -762 3616 -716
rect 5012 -762 5064 -716
rect 6532 -764 6584 -718
rect 7980 -764 8032 -718
rect 9478 -762 9530 -716
rect 10926 -762 10978 -716
<< metal1 >>
rect 354 494 490 514
rect 354 432 390 494
rect 450 432 490 494
rect 354 404 490 432
rect 1802 494 1938 514
rect 1802 432 1838 494
rect 1898 432 1938 494
rect 1802 404 1938 432
rect 3300 496 3436 516
rect 3300 434 3336 496
rect 3396 434 3436 496
rect 3300 406 3436 434
rect 4748 496 4884 516
rect 4748 434 4784 496
rect 4844 434 4884 496
rect 4748 406 4884 434
rect 6268 494 6404 514
rect 6268 432 6304 494
rect 6364 432 6404 494
rect 50 374 1027 404
rect 50 268 82 374
rect 286 268 318 374
rect 522 268 554 374
rect 758 268 790 374
rect 993 268 1027 374
rect 1498 374 2475 404
rect 1498 268 1530 374
rect 1734 268 1766 374
rect 1970 268 2002 374
rect 2206 268 2238 374
rect 2441 268 2475 374
rect 2996 376 3973 406
rect 2996 270 3028 376
rect 3232 270 3264 376
rect 3468 270 3500 376
rect 3704 270 3736 376
rect 3939 270 3973 376
rect 4444 376 5421 406
rect 6268 404 6404 432
rect 7716 494 7852 514
rect 7716 432 7752 494
rect 7812 432 7852 494
rect 7716 404 7852 432
rect 9214 496 9350 516
rect 9214 434 9250 496
rect 9310 434 9350 496
rect 9214 406 9350 434
rect 10662 496 10798 516
rect 10662 434 10698 496
rect 10758 434 10798 496
rect 10662 406 10798 434
rect 4444 270 4476 376
rect 4680 270 4712 376
rect 4916 270 4948 376
rect 5152 270 5184 376
rect 5387 270 5421 376
rect 5964 374 6941 404
rect 43 256 89 268
rect 43 80 49 256
rect 83 80 89 256
rect 43 68 89 80
rect 161 256 207 268
rect 161 80 167 256
rect 201 80 207 256
rect 161 68 207 80
rect 279 256 325 268
rect 279 80 285 256
rect 319 80 325 256
rect 279 68 325 80
rect 397 256 443 268
rect 397 80 403 256
rect 437 80 443 256
rect 397 68 443 80
rect 515 256 561 268
rect 515 80 521 256
rect 555 80 561 256
rect 515 68 561 80
rect 633 256 679 268
rect 633 80 639 256
rect 673 80 679 256
rect 633 68 679 80
rect 751 256 797 268
rect 751 80 757 256
rect 791 80 797 256
rect 751 68 797 80
rect 869 256 915 268
rect 869 80 875 256
rect 909 80 915 256
rect 869 68 915 80
rect 987 256 1033 268
rect 987 80 993 256
rect 1027 80 1033 256
rect 987 68 1033 80
rect 1105 256 1151 268
rect 1105 80 1111 256
rect 1145 80 1151 256
rect 1105 68 1151 80
rect 1491 256 1537 268
rect 1491 80 1497 256
rect 1531 80 1537 256
rect 1491 68 1537 80
rect 1609 256 1655 268
rect 1609 80 1615 256
rect 1649 80 1655 256
rect 1609 68 1655 80
rect 1727 256 1773 268
rect 1727 80 1733 256
rect 1767 80 1773 256
rect 1727 68 1773 80
rect 1845 256 1891 268
rect 1845 80 1851 256
rect 1885 80 1891 256
rect 1845 68 1891 80
rect 1963 256 2009 268
rect 1963 80 1969 256
rect 2003 80 2009 256
rect 1963 68 2009 80
rect 2081 256 2127 268
rect 2081 80 2087 256
rect 2121 80 2127 256
rect 2081 68 2127 80
rect 2199 256 2245 268
rect 2199 80 2205 256
rect 2239 80 2245 256
rect 2199 68 2245 80
rect 2317 256 2363 268
rect 2317 80 2323 256
rect 2357 80 2363 256
rect 2317 68 2363 80
rect 2435 256 2481 268
rect 2435 80 2441 256
rect 2475 80 2481 256
rect 2435 68 2481 80
rect 2553 256 2599 268
rect 2553 80 2559 256
rect 2593 80 2599 256
rect 2553 68 2599 80
rect 2989 258 3035 270
rect 2989 82 2995 258
rect 3029 82 3035 258
rect 2989 70 3035 82
rect 3107 258 3153 270
rect 3107 82 3113 258
rect 3147 82 3153 258
rect 3107 70 3153 82
rect 3225 258 3271 270
rect 3225 82 3231 258
rect 3265 82 3271 258
rect 3225 70 3271 82
rect 3343 258 3389 270
rect 3343 82 3349 258
rect 3383 82 3389 258
rect 3343 70 3389 82
rect 3461 258 3507 270
rect 3461 82 3467 258
rect 3501 82 3507 258
rect 3461 70 3507 82
rect 3579 258 3625 270
rect 3579 82 3585 258
rect 3619 82 3625 258
rect 3579 70 3625 82
rect 3697 258 3743 270
rect 3697 82 3703 258
rect 3737 82 3743 258
rect 3697 70 3743 82
rect 3815 258 3861 270
rect 3815 82 3821 258
rect 3855 82 3861 258
rect 3815 70 3861 82
rect 3933 258 3979 270
rect 3933 82 3939 258
rect 3973 82 3979 258
rect 3933 70 3979 82
rect 4051 258 4097 270
rect 4051 82 4057 258
rect 4091 82 4097 258
rect 4051 70 4097 82
rect 4437 258 4483 270
rect 4437 82 4443 258
rect 4477 82 4483 258
rect 4437 70 4483 82
rect 4555 258 4601 270
rect 4555 82 4561 258
rect 4595 82 4601 258
rect 4555 70 4601 82
rect 4673 258 4719 270
rect 4673 82 4679 258
rect 4713 82 4719 258
rect 4673 70 4719 82
rect 4791 258 4837 270
rect 4791 82 4797 258
rect 4831 82 4837 258
rect 4791 70 4837 82
rect 4909 258 4955 270
rect 4909 82 4915 258
rect 4949 82 4955 258
rect 4909 70 4955 82
rect 5027 258 5073 270
rect 5027 82 5033 258
rect 5067 82 5073 258
rect 5027 70 5073 82
rect 5145 258 5191 270
rect 5145 82 5151 258
rect 5185 82 5191 258
rect 5145 70 5191 82
rect 5263 258 5309 270
rect 5263 82 5269 258
rect 5303 82 5309 258
rect 5263 70 5309 82
rect 5381 258 5427 270
rect 5381 82 5387 258
rect 5421 82 5427 258
rect 5381 70 5427 82
rect 5499 258 5545 270
rect 5964 268 5996 374
rect 6200 268 6232 374
rect 6436 268 6468 374
rect 6672 268 6704 374
rect 6907 268 6941 374
rect 7412 374 8389 404
rect 7412 268 7444 374
rect 7648 268 7680 374
rect 7884 268 7916 374
rect 8120 268 8152 374
rect 8355 268 8389 374
rect 8910 376 9887 406
rect 8910 270 8942 376
rect 9146 270 9178 376
rect 9382 270 9414 376
rect 9618 270 9650 376
rect 9853 270 9887 376
rect 10358 376 11335 406
rect 10358 270 10390 376
rect 10594 270 10626 376
rect 10830 270 10862 376
rect 11066 270 11098 376
rect 11301 270 11335 376
rect 5499 82 5505 258
rect 5539 82 5545 258
rect 5499 70 5545 82
rect 5957 256 6003 268
rect 5957 80 5963 256
rect 5997 80 6003 256
rect 166 -26 202 68
rect 402 -26 438 68
rect 638 -25 674 68
rect 800 20 866 27
rect 800 -14 816 20
rect 850 -14 866 20
rect 800 -25 866 -14
rect 638 -26 866 -25
rect 166 -55 866 -26
rect 166 -56 748 -55
rect 286 -169 320 -56
rect 682 -97 748 -56
rect 682 -131 698 -97
rect 732 -131 748 -97
rect 682 -138 748 -131
rect 1110 -165 1145 68
rect 1614 -26 1650 68
rect 1850 -26 1886 68
rect 2086 -25 2122 68
rect 2248 20 2314 27
rect 2248 -14 2264 20
rect 2298 -14 2314 20
rect 2248 -25 2314 -14
rect 2086 -26 2314 -25
rect 1614 -55 2314 -26
rect 1614 -56 2196 -55
rect 756 -169 1145 -165
rect 1734 -169 1768 -56
rect 2130 -97 2196 -56
rect 2130 -131 2146 -97
rect 2180 -131 2196 -97
rect 2130 -138 2196 -131
rect 2558 -165 2593 68
rect 3112 -24 3148 70
rect 3348 -24 3384 70
rect 3584 -23 3620 70
rect 3746 22 3812 29
rect 3746 -12 3762 22
rect 3796 -12 3812 22
rect 3746 -23 3812 -12
rect 3584 -24 3812 -23
rect 3112 -53 3812 -24
rect 3112 -54 3694 -53
rect 2204 -169 2593 -165
rect 3232 -167 3266 -54
rect 3628 -95 3694 -54
rect 3628 -129 3644 -95
rect 3678 -129 3694 -95
rect 3628 -136 3694 -129
rect 4056 -163 4091 70
rect 4560 -24 4596 70
rect 4796 -24 4832 70
rect 5032 -23 5068 70
rect 5194 22 5260 29
rect 5194 -12 5210 22
rect 5244 -12 5260 22
rect 5194 -23 5260 -12
rect 5032 -24 5260 -23
rect 4560 -53 5260 -24
rect 4560 -54 5142 -53
rect 3702 -167 4091 -163
rect 4680 -167 4714 -54
rect 5076 -95 5142 -54
rect 5076 -129 5092 -95
rect 5126 -129 5142 -95
rect 5076 -136 5142 -129
rect 5504 -163 5539 70
rect 5957 68 6003 80
rect 6075 256 6121 268
rect 6075 80 6081 256
rect 6115 80 6121 256
rect 6075 68 6121 80
rect 6193 256 6239 268
rect 6193 80 6199 256
rect 6233 80 6239 256
rect 6193 68 6239 80
rect 6311 256 6357 268
rect 6311 80 6317 256
rect 6351 80 6357 256
rect 6311 68 6357 80
rect 6429 256 6475 268
rect 6429 80 6435 256
rect 6469 80 6475 256
rect 6429 68 6475 80
rect 6547 256 6593 268
rect 6547 80 6553 256
rect 6587 80 6593 256
rect 6547 68 6593 80
rect 6665 256 6711 268
rect 6665 80 6671 256
rect 6705 80 6711 256
rect 6665 68 6711 80
rect 6783 256 6829 268
rect 6783 80 6789 256
rect 6823 80 6829 256
rect 6783 68 6829 80
rect 6901 256 6947 268
rect 6901 80 6907 256
rect 6941 80 6947 256
rect 6901 68 6947 80
rect 7019 256 7065 268
rect 7019 80 7025 256
rect 7059 80 7065 256
rect 7019 68 7065 80
rect 7405 256 7451 268
rect 7405 80 7411 256
rect 7445 80 7451 256
rect 7405 68 7451 80
rect 7523 256 7569 268
rect 7523 80 7529 256
rect 7563 80 7569 256
rect 7523 68 7569 80
rect 7641 256 7687 268
rect 7641 80 7647 256
rect 7681 80 7687 256
rect 7641 68 7687 80
rect 7759 256 7805 268
rect 7759 80 7765 256
rect 7799 80 7805 256
rect 7759 68 7805 80
rect 7877 256 7923 268
rect 7877 80 7883 256
rect 7917 80 7923 256
rect 7877 68 7923 80
rect 7995 256 8041 268
rect 7995 80 8001 256
rect 8035 80 8041 256
rect 7995 68 8041 80
rect 8113 256 8159 268
rect 8113 80 8119 256
rect 8153 80 8159 256
rect 8113 68 8159 80
rect 8231 256 8277 268
rect 8231 80 8237 256
rect 8271 80 8277 256
rect 8231 68 8277 80
rect 8349 256 8395 268
rect 8349 80 8355 256
rect 8389 80 8395 256
rect 8349 68 8395 80
rect 8467 256 8513 268
rect 8467 80 8473 256
rect 8507 80 8513 256
rect 8467 68 8513 80
rect 8903 258 8949 270
rect 8903 82 8909 258
rect 8943 82 8949 258
rect 8903 70 8949 82
rect 9021 258 9067 270
rect 9021 82 9027 258
rect 9061 82 9067 258
rect 9021 70 9067 82
rect 9139 258 9185 270
rect 9139 82 9145 258
rect 9179 82 9185 258
rect 9139 70 9185 82
rect 9257 258 9303 270
rect 9257 82 9263 258
rect 9297 82 9303 258
rect 9257 70 9303 82
rect 9375 258 9421 270
rect 9375 82 9381 258
rect 9415 82 9421 258
rect 9375 70 9421 82
rect 9493 258 9539 270
rect 9493 82 9499 258
rect 9533 82 9539 258
rect 9493 70 9539 82
rect 9611 258 9657 270
rect 9611 82 9617 258
rect 9651 82 9657 258
rect 9611 70 9657 82
rect 9729 258 9775 270
rect 9729 82 9735 258
rect 9769 82 9775 258
rect 9729 70 9775 82
rect 9847 258 9893 270
rect 9847 82 9853 258
rect 9887 82 9893 258
rect 9847 70 9893 82
rect 9965 258 10011 270
rect 9965 82 9971 258
rect 10005 82 10011 258
rect 9965 70 10011 82
rect 10351 258 10397 270
rect 10351 82 10357 258
rect 10391 82 10397 258
rect 10351 70 10397 82
rect 10469 258 10515 270
rect 10469 82 10475 258
rect 10509 82 10515 258
rect 10469 70 10515 82
rect 10587 258 10633 270
rect 10587 82 10593 258
rect 10627 82 10633 258
rect 10587 70 10633 82
rect 10705 258 10751 270
rect 10705 82 10711 258
rect 10745 82 10751 258
rect 10705 70 10751 82
rect 10823 258 10869 270
rect 10823 82 10829 258
rect 10863 82 10869 258
rect 10823 70 10869 82
rect 10941 258 10987 270
rect 10941 82 10947 258
rect 10981 82 10987 258
rect 10941 70 10987 82
rect 11059 258 11105 270
rect 11059 82 11065 258
rect 11099 82 11105 258
rect 11059 70 11105 82
rect 11177 258 11223 270
rect 11177 82 11183 258
rect 11217 82 11223 258
rect 11177 70 11223 82
rect 11295 258 11341 270
rect 11295 82 11301 258
rect 11335 82 11341 258
rect 11295 70 11341 82
rect 11413 258 11459 270
rect 11413 82 11419 258
rect 11453 82 11459 258
rect 11413 70 11459 82
rect 6080 -26 6116 68
rect 6316 -26 6352 68
rect 6552 -25 6588 68
rect 6714 20 6780 27
rect 6714 -14 6730 20
rect 6764 -14 6780 20
rect 6714 -25 6780 -14
rect 6552 -26 6780 -25
rect 6080 -55 6780 -26
rect 6080 -56 6662 -55
rect 5150 -167 5539 -163
rect 280 -181 326 -169
rect 140 -409 240 -309
rect 28 -537 128 -437
rect 50 -686 104 -537
rect 164 -601 218 -409
rect 280 -557 286 -181
rect 320 -557 326 -181
rect 280 -569 326 -557
rect 398 -181 444 -169
rect 398 -557 404 -181
rect 438 -557 444 -181
rect 398 -569 444 -557
rect 516 -181 562 -169
rect 516 -557 522 -181
rect 556 -530 562 -181
rect 633 -181 679 -169
rect 633 -357 639 -181
rect 673 -357 679 -181
rect 633 -364 679 -357
rect 751 -181 1145 -169
rect 751 -357 757 -181
rect 791 -194 1145 -181
rect 791 -357 797 -194
rect 1041 -274 1145 -194
rect 1728 -181 1774 -169
rect 633 -369 682 -364
rect 751 -369 797 -357
rect 639 -530 682 -369
rect 1588 -409 1688 -309
rect 556 -557 682 -530
rect 1476 -537 1576 -437
rect 516 -569 682 -557
rect 522 -573 682 -569
rect 164 -607 395 -601
rect 164 -641 345 -607
rect 379 -641 395 -607
rect 164 -657 395 -641
rect 447 -607 513 -601
rect 447 -641 463 -607
rect 497 -641 513 -607
rect 447 -686 513 -641
rect 50 -694 513 -686
rect 50 -726 514 -694
rect 606 -710 682 -573
rect 1498 -686 1552 -537
rect 1612 -601 1666 -409
rect 1728 -557 1734 -181
rect 1768 -557 1774 -181
rect 1728 -569 1774 -557
rect 1846 -181 1892 -169
rect 1846 -557 1852 -181
rect 1886 -557 1892 -181
rect 1846 -569 1892 -557
rect 1964 -181 2010 -169
rect 1964 -557 1970 -181
rect 2004 -530 2010 -181
rect 2081 -181 2127 -169
rect 2081 -357 2087 -181
rect 2121 -357 2127 -181
rect 2081 -364 2127 -357
rect 2199 -181 2593 -169
rect 2199 -357 2205 -181
rect 2239 -194 2593 -181
rect 2239 -357 2245 -194
rect 2489 -274 2593 -194
rect 3226 -179 3272 -167
rect 2081 -369 2130 -364
rect 2199 -369 2245 -357
rect 2087 -530 2130 -369
rect 3086 -407 3186 -307
rect 2004 -557 2130 -530
rect 2974 -535 3074 -435
rect 1964 -569 2130 -557
rect 1970 -573 2130 -569
rect 1612 -607 1843 -601
rect 1612 -641 1793 -607
rect 1827 -641 1843 -607
rect 1612 -657 1843 -641
rect 1895 -607 1961 -601
rect 1895 -641 1911 -607
rect 1945 -641 1961 -607
rect 1895 -686 1961 -641
rect 1498 -694 1961 -686
rect 602 -770 612 -710
rect 674 -770 684 -710
rect 1498 -726 1962 -694
rect 2054 -710 2130 -573
rect 2996 -684 3050 -535
rect 3110 -599 3164 -407
rect 3226 -555 3232 -179
rect 3266 -555 3272 -179
rect 3226 -567 3272 -555
rect 3344 -179 3390 -167
rect 3344 -555 3350 -179
rect 3384 -555 3390 -179
rect 3344 -567 3390 -555
rect 3462 -179 3508 -167
rect 3462 -555 3468 -179
rect 3502 -528 3508 -179
rect 3579 -179 3625 -167
rect 3579 -355 3585 -179
rect 3619 -355 3625 -179
rect 3579 -362 3625 -355
rect 3697 -179 4091 -167
rect 3697 -355 3703 -179
rect 3737 -192 4091 -179
rect 3737 -355 3743 -192
rect 3987 -272 4091 -192
rect 4674 -179 4720 -167
rect 3579 -367 3628 -362
rect 3697 -367 3743 -355
rect 3585 -528 3628 -367
rect 4534 -407 4634 -307
rect 3502 -555 3628 -528
rect 4422 -535 4522 -435
rect 3462 -567 3628 -555
rect 3468 -571 3628 -567
rect 3110 -605 3341 -599
rect 3110 -639 3291 -605
rect 3325 -639 3341 -605
rect 3110 -655 3341 -639
rect 3393 -605 3459 -599
rect 3393 -639 3409 -605
rect 3443 -639 3459 -605
rect 3393 -684 3459 -639
rect 2996 -692 3459 -684
rect 2050 -770 2060 -710
rect 2122 -770 2132 -710
rect 2996 -724 3460 -692
rect 3552 -708 3628 -571
rect 4444 -684 4498 -535
rect 4558 -599 4612 -407
rect 4674 -555 4680 -179
rect 4714 -555 4720 -179
rect 4674 -567 4720 -555
rect 4792 -179 4838 -167
rect 4792 -555 4798 -179
rect 4832 -555 4838 -179
rect 4792 -567 4838 -555
rect 4910 -179 4956 -167
rect 4910 -555 4916 -179
rect 4950 -528 4956 -179
rect 5027 -179 5073 -167
rect 5027 -355 5033 -179
rect 5067 -355 5073 -179
rect 5027 -362 5073 -355
rect 5145 -179 5539 -167
rect 6200 -169 6234 -56
rect 6596 -97 6662 -56
rect 6596 -131 6612 -97
rect 6646 -131 6662 -97
rect 6596 -138 6662 -131
rect 7024 -165 7059 68
rect 7528 -26 7564 68
rect 7764 -26 7800 68
rect 8000 -25 8036 68
rect 8162 20 8228 27
rect 8162 -14 8178 20
rect 8212 -14 8228 20
rect 8162 -25 8228 -14
rect 8000 -26 8228 -25
rect 7528 -55 8228 -26
rect 7528 -56 8110 -55
rect 6670 -169 7059 -165
rect 7648 -169 7682 -56
rect 8044 -97 8110 -56
rect 8044 -131 8060 -97
rect 8094 -131 8110 -97
rect 8044 -138 8110 -131
rect 8472 -165 8507 68
rect 9026 -24 9062 70
rect 9262 -24 9298 70
rect 9498 -23 9534 70
rect 9660 22 9726 29
rect 9660 -12 9676 22
rect 9710 -12 9726 22
rect 9660 -23 9726 -12
rect 9498 -24 9726 -23
rect 9026 -53 9726 -24
rect 9026 -54 9608 -53
rect 8118 -169 8507 -165
rect 9146 -167 9180 -54
rect 9542 -95 9608 -54
rect 9542 -129 9558 -95
rect 9592 -129 9608 -95
rect 9542 -136 9608 -129
rect 9970 -163 10005 70
rect 10474 -24 10510 70
rect 10710 -24 10746 70
rect 10946 -23 10982 70
rect 11108 22 11174 29
rect 11108 -12 11124 22
rect 11158 -12 11174 22
rect 11108 -23 11174 -12
rect 10946 -24 11174 -23
rect 10474 -53 11174 -24
rect 10474 -54 11056 -53
rect 9616 -167 10005 -163
rect 10594 -167 10628 -54
rect 10990 -95 11056 -54
rect 10990 -129 11006 -95
rect 11040 -129 11056 -95
rect 10990 -136 11056 -129
rect 11418 -163 11453 70
rect 11064 -167 11453 -163
rect 5145 -355 5151 -179
rect 5185 -192 5539 -179
rect 5185 -355 5191 -192
rect 5435 -272 5539 -192
rect 6194 -181 6240 -169
rect 5027 -367 5076 -362
rect 5145 -367 5191 -355
rect 5033 -528 5076 -367
rect 6054 -409 6154 -309
rect 4950 -555 5076 -528
rect 5942 -537 6042 -437
rect 4910 -567 5076 -555
rect 4916 -571 5076 -567
rect 4558 -605 4789 -599
rect 4558 -639 4739 -605
rect 4773 -639 4789 -605
rect 4558 -655 4789 -639
rect 4841 -605 4907 -599
rect 4841 -639 4857 -605
rect 4891 -639 4907 -605
rect 4841 -684 4907 -639
rect 4444 -692 4907 -684
rect 3548 -768 3558 -708
rect 3620 -768 3630 -708
rect 4444 -724 4908 -692
rect 5000 -708 5076 -571
rect 5964 -686 6018 -537
rect 6078 -601 6132 -409
rect 6194 -557 6200 -181
rect 6234 -557 6240 -181
rect 6194 -569 6240 -557
rect 6312 -181 6358 -169
rect 6312 -557 6318 -181
rect 6352 -557 6358 -181
rect 6312 -569 6358 -557
rect 6430 -181 6476 -169
rect 6430 -557 6436 -181
rect 6470 -530 6476 -181
rect 6547 -181 6593 -169
rect 6547 -357 6553 -181
rect 6587 -357 6593 -181
rect 6547 -364 6593 -357
rect 6665 -181 7059 -169
rect 6665 -357 6671 -181
rect 6705 -194 7059 -181
rect 6705 -357 6711 -194
rect 6955 -274 7059 -194
rect 7642 -181 7688 -169
rect 6547 -369 6596 -364
rect 6665 -369 6711 -357
rect 6553 -530 6596 -369
rect 7502 -409 7602 -309
rect 6470 -557 6596 -530
rect 7390 -537 7490 -437
rect 6430 -569 6596 -557
rect 6436 -573 6596 -569
rect 6078 -607 6309 -601
rect 6078 -641 6259 -607
rect 6293 -641 6309 -607
rect 6078 -657 6309 -641
rect 6361 -607 6427 -601
rect 6361 -641 6377 -607
rect 6411 -641 6427 -607
rect 6361 -686 6427 -641
rect 5964 -694 6427 -686
rect 4996 -768 5006 -708
rect 5068 -768 5078 -708
rect 5964 -726 6428 -694
rect 6520 -710 6596 -573
rect 7412 -686 7466 -537
rect 7526 -601 7580 -409
rect 7642 -557 7648 -181
rect 7682 -557 7688 -181
rect 7642 -569 7688 -557
rect 7760 -181 7806 -169
rect 7760 -557 7766 -181
rect 7800 -557 7806 -181
rect 7760 -569 7806 -557
rect 7878 -181 7924 -169
rect 7878 -557 7884 -181
rect 7918 -530 7924 -181
rect 7995 -181 8041 -169
rect 7995 -357 8001 -181
rect 8035 -357 8041 -181
rect 7995 -364 8041 -357
rect 8113 -181 8507 -169
rect 8113 -357 8119 -181
rect 8153 -194 8507 -181
rect 8153 -357 8159 -194
rect 8403 -274 8507 -194
rect 9140 -179 9186 -167
rect 7995 -369 8044 -364
rect 8113 -369 8159 -357
rect 8001 -530 8044 -369
rect 9000 -407 9100 -307
rect 7918 -557 8044 -530
rect 8888 -535 8988 -435
rect 7878 -569 8044 -557
rect 7884 -573 8044 -569
rect 7526 -607 7757 -601
rect 7526 -641 7707 -607
rect 7741 -641 7757 -607
rect 7526 -657 7757 -641
rect 7809 -607 7875 -601
rect 7809 -641 7825 -607
rect 7859 -641 7875 -607
rect 7809 -686 7875 -641
rect 7412 -694 7875 -686
rect 6516 -770 6526 -710
rect 6588 -770 6598 -710
rect 7412 -726 7876 -694
rect 7968 -710 8044 -573
rect 8910 -684 8964 -535
rect 9024 -599 9078 -407
rect 9140 -555 9146 -179
rect 9180 -555 9186 -179
rect 9140 -567 9186 -555
rect 9258 -179 9304 -167
rect 9258 -555 9264 -179
rect 9298 -555 9304 -179
rect 9258 -567 9304 -555
rect 9376 -179 9422 -167
rect 9376 -555 9382 -179
rect 9416 -528 9422 -179
rect 9493 -179 9539 -167
rect 9493 -355 9499 -179
rect 9533 -355 9539 -179
rect 9493 -362 9539 -355
rect 9611 -179 10005 -167
rect 9611 -355 9617 -179
rect 9651 -192 10005 -179
rect 9651 -355 9657 -192
rect 9901 -272 10005 -192
rect 10588 -179 10634 -167
rect 9493 -367 9542 -362
rect 9611 -367 9657 -355
rect 9499 -528 9542 -367
rect 10448 -407 10548 -307
rect 9416 -555 9542 -528
rect 10336 -535 10436 -435
rect 9376 -567 9542 -555
rect 9382 -571 9542 -567
rect 9024 -605 9255 -599
rect 9024 -639 9205 -605
rect 9239 -639 9255 -605
rect 9024 -655 9255 -639
rect 9307 -605 9373 -599
rect 9307 -639 9323 -605
rect 9357 -639 9373 -605
rect 9307 -684 9373 -639
rect 8910 -692 9373 -684
rect 7964 -770 7974 -710
rect 8036 -770 8046 -710
rect 8910 -724 9374 -692
rect 9466 -708 9542 -571
rect 10358 -684 10412 -535
rect 10472 -599 10526 -407
rect 10588 -555 10594 -179
rect 10628 -555 10634 -179
rect 10588 -567 10634 -555
rect 10706 -179 10752 -167
rect 10706 -555 10712 -179
rect 10746 -555 10752 -179
rect 10706 -567 10752 -555
rect 10824 -179 10870 -167
rect 10824 -555 10830 -179
rect 10864 -528 10870 -179
rect 10941 -179 10987 -167
rect 10941 -355 10947 -179
rect 10981 -355 10987 -179
rect 10941 -362 10987 -355
rect 11059 -179 11453 -167
rect 11059 -355 11065 -179
rect 11099 -192 11453 -179
rect 11099 -355 11105 -192
rect 11349 -272 11453 -192
rect 10941 -367 10990 -362
rect 11059 -367 11105 -355
rect 10947 -528 10990 -367
rect 10864 -555 10990 -528
rect 10824 -567 10990 -555
rect 10830 -571 10990 -567
rect 10472 -605 10703 -599
rect 10472 -639 10653 -605
rect 10687 -639 10703 -605
rect 10472 -655 10703 -639
rect 10755 -605 10821 -599
rect 10755 -639 10771 -605
rect 10805 -639 10821 -605
rect 10755 -684 10821 -639
rect 10358 -692 10821 -684
rect 9462 -768 9472 -708
rect 9534 -768 9544 -708
rect 10358 -724 10822 -692
rect 10914 -708 10990 -571
rect 10910 -768 10920 -708
rect 10982 -768 10992 -708
<< via1 >>
rect 390 432 450 494
rect 1838 432 1898 494
rect 3336 434 3396 496
rect 4784 434 4844 496
rect 6304 432 6364 494
rect 7752 432 7812 494
rect 9250 434 9310 496
rect 10698 434 10758 496
rect 612 -718 674 -710
rect 612 -764 618 -718
rect 618 -764 670 -718
rect 670 -764 674 -718
rect 612 -770 674 -764
rect 2060 -718 2122 -710
rect 2060 -764 2066 -718
rect 2066 -764 2118 -718
rect 2118 -764 2122 -718
rect 2060 -770 2122 -764
rect 3558 -716 3620 -708
rect 3558 -762 3564 -716
rect 3564 -762 3616 -716
rect 3616 -762 3620 -716
rect 3558 -768 3620 -762
rect 5006 -716 5068 -708
rect 5006 -762 5012 -716
rect 5012 -762 5064 -716
rect 5064 -762 5068 -716
rect 5006 -768 5068 -762
rect 6526 -718 6588 -710
rect 6526 -764 6532 -718
rect 6532 -764 6584 -718
rect 6584 -764 6588 -718
rect 6526 -770 6588 -764
rect 7974 -718 8036 -710
rect 7974 -764 7980 -718
rect 7980 -764 8032 -718
rect 8032 -764 8036 -718
rect 7974 -770 8036 -764
rect 9472 -716 9534 -708
rect 9472 -762 9478 -716
rect 9478 -762 9530 -716
rect 9530 -762 9534 -716
rect 9472 -768 9534 -762
rect 10920 -716 10982 -708
rect 10920 -762 10926 -716
rect 10926 -762 10978 -716
rect 10978 -762 10982 -716
rect 10920 -768 10982 -762
<< metal2 >>
rect 390 494 450 504
rect 390 422 450 432
rect 1838 494 1898 504
rect 1838 422 1898 432
rect 3336 496 3396 506
rect 3336 424 3396 434
rect 4784 496 4844 506
rect 4784 424 4844 434
rect 6304 494 6364 504
rect 6304 422 6364 432
rect 7752 494 7812 504
rect 7752 422 7812 432
rect 9250 496 9310 506
rect 9250 424 9310 434
rect 10698 496 10758 506
rect 10698 424 10758 434
rect 3558 -700 3620 -698
rect 5006 -700 5068 -698
rect 9472 -700 9534 -698
rect 10920 -700 10982 -698
rect 612 -702 674 -700
rect 2060 -702 2122 -700
rect 612 -710 676 -702
rect 674 -712 676 -710
rect 612 -784 676 -774
rect 2060 -710 2124 -702
rect 2122 -712 2124 -710
rect 2060 -784 2124 -774
rect 3558 -708 3622 -700
rect 3620 -710 3622 -708
rect 3558 -782 3622 -772
rect 5006 -708 5070 -700
rect 5068 -710 5070 -708
rect 5006 -782 5070 -772
rect 6526 -702 6588 -700
rect 7974 -702 8036 -700
rect 6526 -710 6590 -702
rect 6588 -712 6590 -710
rect 6526 -784 6590 -774
rect 7974 -710 8038 -702
rect 8036 -712 8038 -710
rect 7974 -784 8038 -774
rect 9472 -708 9536 -700
rect 9534 -710 9536 -708
rect 9472 -782 9536 -772
rect 10920 -708 10984 -700
rect 10982 -710 10984 -708
rect 10920 -782 10984 -772
<< via2 >>
rect 390 432 450 494
rect 1838 432 1898 494
rect 3336 434 3396 496
rect 4784 434 4844 496
rect 6304 432 6364 494
rect 7752 432 7812 494
rect 9250 434 9310 496
rect 10698 434 10758 496
rect 612 -770 674 -712
rect 674 -770 676 -712
rect 612 -774 676 -770
rect 2060 -770 2122 -712
rect 2122 -770 2124 -712
rect 2060 -774 2124 -770
rect 3558 -768 3620 -710
rect 3620 -768 3622 -710
rect 3558 -772 3622 -768
rect 5006 -768 5068 -710
rect 5068 -768 5070 -710
rect 5006 -772 5070 -768
rect 6526 -770 6588 -712
rect 6588 -770 6590 -712
rect 6526 -774 6590 -770
rect 7974 -770 8036 -712
rect 8036 -770 8038 -712
rect 7974 -774 8038 -770
rect 9472 -768 9534 -710
rect 9534 -768 9536 -710
rect 9472 -772 9536 -768
rect 10920 -768 10982 -710
rect 10982 -768 10984 -710
rect 10920 -772 10984 -768
<< metal3 >>
rect 374 498 472 516
rect 374 426 384 498
rect 454 426 472 498
rect 374 418 472 426
rect 1822 498 1920 516
rect 1822 426 1832 498
rect 1902 426 1920 498
rect 1822 418 1920 426
rect 3320 500 3418 518
rect 3320 428 3330 500
rect 3400 428 3418 500
rect 3320 420 3418 428
rect 4768 500 4866 518
rect 4768 428 4778 500
rect 4848 428 4866 500
rect 4768 420 4866 428
rect 6288 498 6386 516
rect 6288 426 6298 498
rect 6368 426 6386 498
rect 6288 418 6386 426
rect 7736 498 7834 516
rect 7736 426 7746 498
rect 7816 426 7834 498
rect 7736 418 7834 426
rect 9234 500 9332 518
rect 9234 428 9244 500
rect 9314 428 9332 500
rect 9234 420 9332 428
rect 10682 500 10780 518
rect 10682 428 10692 500
rect 10762 428 10780 500
rect 10682 420 10780 428
rect 592 -706 694 -690
rect 592 -774 606 -706
rect 680 -774 694 -706
rect 592 -788 694 -774
rect 2040 -706 2142 -690
rect 2040 -774 2054 -706
rect 2128 -774 2142 -706
rect 2040 -788 2142 -774
rect 3538 -704 3640 -688
rect 3538 -772 3552 -704
rect 3626 -772 3640 -704
rect 3538 -786 3640 -772
rect 4986 -704 5088 -688
rect 4986 -772 5000 -704
rect 5074 -772 5088 -704
rect 4986 -786 5088 -772
rect 6506 -706 6608 -690
rect 6506 -774 6520 -706
rect 6594 -774 6608 -706
rect 6506 -788 6608 -774
rect 7954 -706 8056 -690
rect 7954 -774 7968 -706
rect 8042 -774 8056 -706
rect 7954 -788 8056 -774
rect 9452 -704 9554 -688
rect 9452 -772 9466 -704
rect 9540 -772 9554 -704
rect 9452 -786 9554 -772
rect 10900 -704 11002 -688
rect 10900 -772 10914 -704
rect 10988 -772 11002 -704
rect 10900 -786 11002 -772
<< via3 >>
rect 384 494 454 498
rect 384 432 390 494
rect 390 432 450 494
rect 450 432 454 494
rect 384 426 454 432
rect 1832 494 1902 498
rect 1832 432 1838 494
rect 1838 432 1898 494
rect 1898 432 1902 494
rect 1832 426 1902 432
rect 3330 496 3400 500
rect 3330 434 3336 496
rect 3336 434 3396 496
rect 3396 434 3400 496
rect 3330 428 3400 434
rect 4778 496 4848 500
rect 4778 434 4784 496
rect 4784 434 4844 496
rect 4844 434 4848 496
rect 4778 428 4848 434
rect 6298 494 6368 498
rect 6298 432 6304 494
rect 6304 432 6364 494
rect 6364 432 6368 494
rect 6298 426 6368 432
rect 7746 494 7816 498
rect 7746 432 7752 494
rect 7752 432 7812 494
rect 7812 432 7816 494
rect 7746 426 7816 432
rect 9244 496 9314 500
rect 9244 434 9250 496
rect 9250 434 9310 496
rect 9310 434 9314 496
rect 9244 428 9314 434
rect 10692 496 10762 500
rect 10692 434 10698 496
rect 10698 434 10758 496
rect 10758 434 10762 496
rect 10692 428 10762 434
rect 606 -712 680 -706
rect 606 -774 612 -712
rect 612 -774 676 -712
rect 676 -774 680 -712
rect 2054 -712 2128 -706
rect 2054 -774 2060 -712
rect 2060 -774 2124 -712
rect 2124 -774 2128 -712
rect 3552 -710 3626 -704
rect 3552 -772 3558 -710
rect 3558 -772 3622 -710
rect 3622 -772 3626 -710
rect 5000 -710 5074 -704
rect 5000 -772 5006 -710
rect 5006 -772 5070 -710
rect 5070 -772 5074 -710
rect 6520 -712 6594 -706
rect 6520 -774 6526 -712
rect 6526 -774 6590 -712
rect 6590 -774 6594 -712
rect 7968 -712 8042 -706
rect 7968 -774 7974 -712
rect 7974 -774 8038 -712
rect 8038 -774 8042 -712
rect 9466 -710 9540 -704
rect 9466 -772 9472 -710
rect 9472 -772 9536 -710
rect 9536 -772 9540 -710
rect 10914 -710 10988 -704
rect 10914 -772 10920 -710
rect 10920 -772 10984 -710
rect 10984 -772 10988 -710
<< metal4 >>
rect 28 500 11162 556
rect 28 498 3330 500
rect 28 426 384 498
rect 454 426 1832 498
rect 1902 428 3330 498
rect 3400 428 4778 500
rect 4848 498 9244 500
rect 4848 428 6298 498
rect 1902 426 6298 428
rect 6368 426 7746 498
rect 7816 428 9244 498
rect 9314 428 10692 500
rect 10762 428 11162 500
rect 7816 426 11162 428
rect 28 398 11162 426
rect 3424 -678 3756 -676
rect 4872 -678 5204 -676
rect 9338 -678 9670 -676
rect 10786 -678 11118 -676
rect 32 -704 11156 -678
rect 32 -706 3552 -704
rect 32 -774 606 -706
rect 680 -774 2054 -706
rect 2128 -772 3552 -706
rect 3626 -772 5000 -704
rect 5074 -706 9466 -704
rect 5074 -772 6520 -706
rect 2128 -774 6520 -772
rect 6594 -774 7968 -706
rect 8042 -772 9466 -706
rect 9540 -772 10914 -704
rect 10988 -772 11156 -704
rect 8042 -774 11156 -772
rect 32 -812 11156 -774
<< labels >>
flabel metal4 5504 -790 5734 -706 1 FreeSerif 640 0 0 0 VSS
port 1 n
flabel metal4 5566 432 5778 540 1 FreeSerif 640 0 0 0 VDD
port 2 n
flabel metal1 152 -390 228 -320 1 FreeSerif 400 0 0 0 A[0]
port 3 n
flabel metal1 1600 -396 1676 -326 1 FreeSerif 400 0 0 0 A[1]
port 4 n
flabel metal1 3102 -390 3178 -320 1 FreeSerif 400 0 0 0 A[2]
port 5 n
flabel metal1 4548 -392 4624 -322 1 FreeSerif 400 0 0 0 A[3]
port 6 n
flabel metal1 6070 -390 6146 -320 1 FreeSerif 400 0 0 0 A[4]
port 7 n
flabel metal1 7520 -386 7596 -316 1 FreeSerif 400 0 0 0 A[5]
port 8 n
flabel metal1 9014 -392 9090 -322 1 FreeSerif 400 0 0 0 A[6]
port 9 n
flabel metal1 10460 -392 10536 -322 1 FreeSerif 400 0 0 0 A[7]
port 10 n
flabel metal1 10348 -516 10424 -446 1 FreeSerif 400 0 0 0 B[7]
port 11 n
flabel metal1 8900 -516 8976 -446 1 FreeSerif 400 0 0 0 B[6]
port 12 n
flabel metal1 7400 -520 7476 -450 1 FreeSerif 400 0 0 0 B[5]
port 13 n
flabel metal1 4434 -518 4510 -448 1 FreeSerif 400 0 0 0 B[3]
port 14 n
flabel metal1 5952 -518 6028 -448 1 FreeSerif 400 0 0 0 B[4]
port 15 n
flabel metal1 2988 -520 3064 -450 1 FreeSerif 400 0 0 0 B[2]
port 16 n
flabel metal1 1492 -518 1568 -448 1 FreeSerif 400 0 0 0 B[1]
port 17 n
flabel metal1 44 -518 120 -448 1 FreeSerif 400 0 0 0 B[0]
port 18 n
flabel metal1 1058 -258 1134 -188 1 FreeSerif 400 0 0 0 Y[0]
port 19 n
flabel metal1 2500 -254 2576 -184 1 FreeSerif 400 0 0 0 Y[1]
port 20 n
flabel metal1 4004 -252 4080 -182 1 FreeSerif 400 0 0 0 Y[2]
port 21 n
flabel metal1 5454 -254 5530 -184 1 FreeSerif 400 0 0 0 Y[3]
port 22 n
flabel metal1 6970 -252 7046 -182 1 FreeSerif 400 0 0 0 Y[4]
port 23 n
flabel metal1 8422 -254 8498 -184 1 FreeSerif 400 0 0 0 Y[5]
port 24 n
flabel metal1 9912 -262 9988 -192 1 FreeSerif 400 0 0 0 Y[6]
port 25 n
flabel metal1 11362 -256 11438 -186 1 FreeSerif 400 0 0 0 Y[7]
port 26 n
<< end >>
