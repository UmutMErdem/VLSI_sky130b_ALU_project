magic
tech sky130B
magscale 1 2
timestamp 1736542143
<< nwell >>
rect 546 772 1022 964
rect 2614 774 3090 964
rect 356 477 1200 772
rect 2424 479 3268 774
rect 4683 772 5159 964
rect 6751 774 7227 964
rect 8820 774 9296 966
rect 10888 776 11364 966
rect -125 153 1680 477
rect 1943 155 3748 479
rect 4493 477 5337 772
rect 6561 479 7405 774
rect 8630 479 9474 774
rect 10698 481 11542 776
rect 12957 774 13433 966
rect 15025 776 15501 966
rect 302 -540 1140 153
rect 2370 -538 3208 155
rect 4012 153 5817 477
rect 6080 155 7885 479
rect 8149 155 9954 479
rect 10217 157 12022 481
rect 12767 479 13611 774
rect 14835 481 15679 776
rect 4439 -540 5277 153
rect 6507 -538 7345 155
rect 8576 -538 9414 155
rect 10644 -536 11482 157
rect 12286 155 14091 479
rect 14354 157 16159 481
rect 12713 -538 13551 155
rect 14781 -536 15619 157
<< nmos >>
rect 94 -1010 154 -810
rect 514 -1210 574 -810
rect 632 -1210 692 -810
rect 750 -1210 810 -810
rect 868 -1210 928 -810
rect 1392 -1010 1452 -810
rect 2162 -1008 2222 -808
rect 2582 -1208 2642 -808
rect 2700 -1208 2760 -808
rect 2818 -1208 2878 -808
rect 2936 -1208 2996 -808
rect 3460 -1008 3520 -808
rect 4231 -1010 4291 -810
rect 4651 -1210 4711 -810
rect 4769 -1210 4829 -810
rect 4887 -1210 4947 -810
rect 5005 -1210 5065 -810
rect 5529 -1010 5589 -810
rect 6299 -1008 6359 -808
rect 6719 -1208 6779 -808
rect 6837 -1208 6897 -808
rect 6955 -1208 7015 -808
rect 7073 -1208 7133 -808
rect 7597 -1008 7657 -808
rect 8368 -1008 8428 -808
rect 8788 -1208 8848 -808
rect 8906 -1208 8966 -808
rect 9024 -1208 9084 -808
rect 9142 -1208 9202 -808
rect 9666 -1008 9726 -808
rect 10436 -1006 10496 -806
rect 10856 -1206 10916 -806
rect 10974 -1206 11034 -806
rect 11092 -1206 11152 -806
rect 11210 -1206 11270 -806
rect 11734 -1006 11794 -806
rect 12505 -1008 12565 -808
rect 12925 -1208 12985 -808
rect 13043 -1208 13103 -808
rect 13161 -1208 13221 -808
rect 13279 -1208 13339 -808
rect 13803 -1008 13863 -808
rect 14573 -1006 14633 -806
rect 14993 -1206 15053 -806
rect 15111 -1206 15171 -806
rect 15229 -1206 15289 -806
rect 15347 -1206 15407 -806
rect 15871 -1006 15931 -806
<< pmos >>
rect -31 215 29 415
rect 87 215 147 415
rect 205 215 265 415
rect 453 215 513 615
rect 571 215 631 615
rect 689 215 749 615
rect 807 215 867 615
rect 925 215 985 615
rect 1043 215 1103 615
rect 1290 215 1350 415
rect 1408 215 1468 415
rect 1526 215 1586 415
rect 2037 217 2097 417
rect 2155 217 2215 417
rect 2273 217 2333 417
rect 2521 217 2581 617
rect 2639 217 2699 617
rect 2757 217 2817 617
rect 2875 217 2935 617
rect 2993 217 3053 617
rect 3111 217 3171 617
rect 3358 217 3418 417
rect 3476 217 3536 417
rect 3594 217 3654 417
rect 396 -478 456 -78
rect 514 -478 574 -78
rect 632 -478 692 -78
rect 750 -478 810 -78
rect 868 -478 928 -78
rect 986 -478 1046 -78
rect 4106 215 4166 415
rect 4224 215 4284 415
rect 4342 215 4402 415
rect 4590 215 4650 615
rect 4708 215 4768 615
rect 4826 215 4886 615
rect 4944 215 5004 615
rect 5062 215 5122 615
rect 5180 215 5240 615
rect 5427 215 5487 415
rect 5545 215 5605 415
rect 5663 215 5723 415
rect 6174 217 6234 417
rect 6292 217 6352 417
rect 6410 217 6470 417
rect 6658 217 6718 617
rect 6776 217 6836 617
rect 6894 217 6954 617
rect 7012 217 7072 617
rect 7130 217 7190 617
rect 7248 217 7308 617
rect 7495 217 7555 417
rect 7613 217 7673 417
rect 7731 217 7791 417
rect 8243 217 8303 417
rect 8361 217 8421 417
rect 8479 217 8539 417
rect 8727 217 8787 617
rect 8845 217 8905 617
rect 8963 217 9023 617
rect 9081 217 9141 617
rect 9199 217 9259 617
rect 9317 217 9377 617
rect 9564 217 9624 417
rect 9682 217 9742 417
rect 9800 217 9860 417
rect 10311 219 10371 419
rect 10429 219 10489 419
rect 10547 219 10607 419
rect 10795 219 10855 619
rect 10913 219 10973 619
rect 11031 219 11091 619
rect 11149 219 11209 619
rect 11267 219 11327 619
rect 11385 219 11445 619
rect 11632 219 11692 419
rect 11750 219 11810 419
rect 11868 219 11928 419
rect 2464 -476 2524 -76
rect 2582 -476 2642 -76
rect 2700 -476 2760 -76
rect 2818 -476 2878 -76
rect 2936 -476 2996 -76
rect 3054 -476 3114 -76
rect 4533 -478 4593 -78
rect 4651 -478 4711 -78
rect 4769 -478 4829 -78
rect 4887 -478 4947 -78
rect 5005 -478 5065 -78
rect 5123 -478 5183 -78
rect 6601 -476 6661 -76
rect 6719 -476 6779 -76
rect 6837 -476 6897 -76
rect 6955 -476 7015 -76
rect 7073 -476 7133 -76
rect 7191 -476 7251 -76
rect 8670 -476 8730 -76
rect 8788 -476 8848 -76
rect 8906 -476 8966 -76
rect 9024 -476 9084 -76
rect 9142 -476 9202 -76
rect 9260 -476 9320 -76
rect 12380 217 12440 417
rect 12498 217 12558 417
rect 12616 217 12676 417
rect 12864 217 12924 617
rect 12982 217 13042 617
rect 13100 217 13160 617
rect 13218 217 13278 617
rect 13336 217 13396 617
rect 13454 217 13514 617
rect 13701 217 13761 417
rect 13819 217 13879 417
rect 13937 217 13997 417
rect 14448 219 14508 419
rect 14566 219 14626 419
rect 14684 219 14744 419
rect 14932 219 14992 619
rect 15050 219 15110 619
rect 15168 219 15228 619
rect 15286 219 15346 619
rect 15404 219 15464 619
rect 15522 219 15582 619
rect 15769 219 15829 419
rect 15887 219 15947 419
rect 16005 219 16065 419
rect 10738 -474 10798 -74
rect 10856 -474 10916 -74
rect 10974 -474 11034 -74
rect 11092 -474 11152 -74
rect 11210 -474 11270 -74
rect 11328 -474 11388 -74
rect 12807 -476 12867 -76
rect 12925 -476 12985 -76
rect 13043 -476 13103 -76
rect 13161 -476 13221 -76
rect 13279 -476 13339 -76
rect 13397 -476 13457 -76
rect 14875 -474 14935 -74
rect 14993 -474 15053 -74
rect 15111 -474 15171 -74
rect 15229 -474 15289 -74
rect 15347 -474 15407 -74
rect 15465 -474 15525 -74
<< ndiff >>
rect 36 -822 94 -810
rect 36 -998 48 -822
rect 82 -998 94 -822
rect 36 -1010 94 -998
rect 154 -822 212 -810
rect 154 -998 166 -822
rect 200 -998 212 -822
rect 154 -1010 212 -998
rect 456 -822 514 -810
rect 456 -1198 468 -822
rect 502 -1198 514 -822
rect 456 -1210 514 -1198
rect 574 -822 632 -810
rect 574 -1198 586 -822
rect 620 -1198 632 -822
rect 574 -1210 632 -1198
rect 692 -822 750 -810
rect 692 -1198 704 -822
rect 738 -1198 750 -822
rect 692 -1210 750 -1198
rect 810 -822 868 -810
rect 810 -1198 822 -822
rect 856 -1198 868 -822
rect 810 -1210 868 -1198
rect 928 -822 986 -810
rect 928 -1198 940 -822
rect 974 -1198 986 -822
rect 1334 -822 1392 -810
rect 1334 -998 1346 -822
rect 1380 -998 1392 -822
rect 1334 -1010 1392 -998
rect 1452 -822 1510 -810
rect 1452 -998 1464 -822
rect 1498 -998 1510 -822
rect 1452 -1010 1510 -998
rect 2104 -820 2162 -808
rect 2104 -996 2116 -820
rect 2150 -996 2162 -820
rect 2104 -1008 2162 -996
rect 2222 -820 2280 -808
rect 2222 -996 2234 -820
rect 2268 -996 2280 -820
rect 2222 -1008 2280 -996
rect 2524 -820 2582 -808
rect 928 -1210 986 -1198
rect 2524 -1196 2536 -820
rect 2570 -1196 2582 -820
rect 2524 -1208 2582 -1196
rect 2642 -820 2700 -808
rect 2642 -1196 2654 -820
rect 2688 -1196 2700 -820
rect 2642 -1208 2700 -1196
rect 2760 -820 2818 -808
rect 2760 -1196 2772 -820
rect 2806 -1196 2818 -820
rect 2760 -1208 2818 -1196
rect 2878 -820 2936 -808
rect 2878 -1196 2890 -820
rect 2924 -1196 2936 -820
rect 2878 -1208 2936 -1196
rect 2996 -820 3054 -808
rect 2996 -1196 3008 -820
rect 3042 -1196 3054 -820
rect 3402 -820 3460 -808
rect 3402 -996 3414 -820
rect 3448 -996 3460 -820
rect 3402 -1008 3460 -996
rect 3520 -820 3578 -808
rect 3520 -996 3532 -820
rect 3566 -996 3578 -820
rect 3520 -1008 3578 -996
rect 4173 -822 4231 -810
rect 4173 -998 4185 -822
rect 4219 -998 4231 -822
rect 4173 -1010 4231 -998
rect 4291 -822 4349 -810
rect 4291 -998 4303 -822
rect 4337 -998 4349 -822
rect 4291 -1010 4349 -998
rect 4593 -822 4651 -810
rect 2996 -1208 3054 -1196
rect 4593 -1198 4605 -822
rect 4639 -1198 4651 -822
rect 4593 -1210 4651 -1198
rect 4711 -822 4769 -810
rect 4711 -1198 4723 -822
rect 4757 -1198 4769 -822
rect 4711 -1210 4769 -1198
rect 4829 -822 4887 -810
rect 4829 -1198 4841 -822
rect 4875 -1198 4887 -822
rect 4829 -1210 4887 -1198
rect 4947 -822 5005 -810
rect 4947 -1198 4959 -822
rect 4993 -1198 5005 -822
rect 4947 -1210 5005 -1198
rect 5065 -822 5123 -810
rect 5065 -1198 5077 -822
rect 5111 -1198 5123 -822
rect 5471 -822 5529 -810
rect 5471 -998 5483 -822
rect 5517 -998 5529 -822
rect 5471 -1010 5529 -998
rect 5589 -822 5647 -810
rect 5589 -998 5601 -822
rect 5635 -998 5647 -822
rect 5589 -1010 5647 -998
rect 6241 -820 6299 -808
rect 6241 -996 6253 -820
rect 6287 -996 6299 -820
rect 6241 -1008 6299 -996
rect 6359 -820 6417 -808
rect 6359 -996 6371 -820
rect 6405 -996 6417 -820
rect 6359 -1008 6417 -996
rect 6661 -820 6719 -808
rect 5065 -1210 5123 -1198
rect 6661 -1196 6673 -820
rect 6707 -1196 6719 -820
rect 6661 -1208 6719 -1196
rect 6779 -820 6837 -808
rect 6779 -1196 6791 -820
rect 6825 -1196 6837 -820
rect 6779 -1208 6837 -1196
rect 6897 -820 6955 -808
rect 6897 -1196 6909 -820
rect 6943 -1196 6955 -820
rect 6897 -1208 6955 -1196
rect 7015 -820 7073 -808
rect 7015 -1196 7027 -820
rect 7061 -1196 7073 -820
rect 7015 -1208 7073 -1196
rect 7133 -820 7191 -808
rect 7133 -1196 7145 -820
rect 7179 -1196 7191 -820
rect 7539 -820 7597 -808
rect 7539 -996 7551 -820
rect 7585 -996 7597 -820
rect 7539 -1008 7597 -996
rect 7657 -820 7715 -808
rect 7657 -996 7669 -820
rect 7703 -996 7715 -820
rect 7657 -1008 7715 -996
rect 8310 -820 8368 -808
rect 8310 -996 8322 -820
rect 8356 -996 8368 -820
rect 8310 -1008 8368 -996
rect 8428 -820 8486 -808
rect 8428 -996 8440 -820
rect 8474 -996 8486 -820
rect 8428 -1008 8486 -996
rect 8730 -820 8788 -808
rect 7133 -1208 7191 -1196
rect 8730 -1196 8742 -820
rect 8776 -1196 8788 -820
rect 8730 -1208 8788 -1196
rect 8848 -820 8906 -808
rect 8848 -1196 8860 -820
rect 8894 -1196 8906 -820
rect 8848 -1208 8906 -1196
rect 8966 -820 9024 -808
rect 8966 -1196 8978 -820
rect 9012 -1196 9024 -820
rect 8966 -1208 9024 -1196
rect 9084 -820 9142 -808
rect 9084 -1196 9096 -820
rect 9130 -1196 9142 -820
rect 9084 -1208 9142 -1196
rect 9202 -820 9260 -808
rect 9202 -1196 9214 -820
rect 9248 -1196 9260 -820
rect 9608 -820 9666 -808
rect 9608 -996 9620 -820
rect 9654 -996 9666 -820
rect 9608 -1008 9666 -996
rect 9726 -820 9784 -808
rect 9726 -996 9738 -820
rect 9772 -996 9784 -820
rect 9726 -1008 9784 -996
rect 10378 -818 10436 -806
rect 10378 -994 10390 -818
rect 10424 -994 10436 -818
rect 10378 -1006 10436 -994
rect 10496 -818 10554 -806
rect 10496 -994 10508 -818
rect 10542 -994 10554 -818
rect 10496 -1006 10554 -994
rect 10798 -818 10856 -806
rect 9202 -1208 9260 -1196
rect 10798 -1194 10810 -818
rect 10844 -1194 10856 -818
rect 10798 -1206 10856 -1194
rect 10916 -818 10974 -806
rect 10916 -1194 10928 -818
rect 10962 -1194 10974 -818
rect 10916 -1206 10974 -1194
rect 11034 -818 11092 -806
rect 11034 -1194 11046 -818
rect 11080 -1194 11092 -818
rect 11034 -1206 11092 -1194
rect 11152 -818 11210 -806
rect 11152 -1194 11164 -818
rect 11198 -1194 11210 -818
rect 11152 -1206 11210 -1194
rect 11270 -818 11328 -806
rect 11270 -1194 11282 -818
rect 11316 -1194 11328 -818
rect 11676 -818 11734 -806
rect 11676 -994 11688 -818
rect 11722 -994 11734 -818
rect 11676 -1006 11734 -994
rect 11794 -818 11852 -806
rect 11794 -994 11806 -818
rect 11840 -994 11852 -818
rect 11794 -1006 11852 -994
rect 12447 -820 12505 -808
rect 12447 -996 12459 -820
rect 12493 -996 12505 -820
rect 12447 -1008 12505 -996
rect 12565 -820 12623 -808
rect 12565 -996 12577 -820
rect 12611 -996 12623 -820
rect 12565 -1008 12623 -996
rect 12867 -820 12925 -808
rect 11270 -1206 11328 -1194
rect 12867 -1196 12879 -820
rect 12913 -1196 12925 -820
rect 12867 -1208 12925 -1196
rect 12985 -820 13043 -808
rect 12985 -1196 12997 -820
rect 13031 -1196 13043 -820
rect 12985 -1208 13043 -1196
rect 13103 -820 13161 -808
rect 13103 -1196 13115 -820
rect 13149 -1196 13161 -820
rect 13103 -1208 13161 -1196
rect 13221 -820 13279 -808
rect 13221 -1196 13233 -820
rect 13267 -1196 13279 -820
rect 13221 -1208 13279 -1196
rect 13339 -820 13397 -808
rect 13339 -1196 13351 -820
rect 13385 -1196 13397 -820
rect 13745 -820 13803 -808
rect 13745 -996 13757 -820
rect 13791 -996 13803 -820
rect 13745 -1008 13803 -996
rect 13863 -820 13921 -808
rect 13863 -996 13875 -820
rect 13909 -996 13921 -820
rect 13863 -1008 13921 -996
rect 14515 -818 14573 -806
rect 14515 -994 14527 -818
rect 14561 -994 14573 -818
rect 14515 -1006 14573 -994
rect 14633 -818 14691 -806
rect 14633 -994 14645 -818
rect 14679 -994 14691 -818
rect 14633 -1006 14691 -994
rect 14935 -818 14993 -806
rect 13339 -1208 13397 -1196
rect 14935 -1194 14947 -818
rect 14981 -1194 14993 -818
rect 14935 -1206 14993 -1194
rect 15053 -818 15111 -806
rect 15053 -1194 15065 -818
rect 15099 -1194 15111 -818
rect 15053 -1206 15111 -1194
rect 15171 -818 15229 -806
rect 15171 -1194 15183 -818
rect 15217 -1194 15229 -818
rect 15171 -1206 15229 -1194
rect 15289 -818 15347 -806
rect 15289 -1194 15301 -818
rect 15335 -1194 15347 -818
rect 15289 -1206 15347 -1194
rect 15407 -818 15465 -806
rect 15407 -1194 15419 -818
rect 15453 -1194 15465 -818
rect 15813 -818 15871 -806
rect 15813 -994 15825 -818
rect 15859 -994 15871 -818
rect 15813 -1006 15871 -994
rect 15931 -818 15989 -806
rect 15931 -994 15943 -818
rect 15977 -994 15989 -818
rect 15931 -1006 15989 -994
rect 15407 -1206 15465 -1194
<< pdiff >>
rect 395 603 453 615
rect -89 403 -31 415
rect -89 227 -77 403
rect -43 227 -31 403
rect -89 215 -31 227
rect 29 403 87 415
rect 29 227 41 403
rect 75 227 87 403
rect 29 215 87 227
rect 147 403 205 415
rect 147 227 159 403
rect 193 227 205 403
rect 147 215 205 227
rect 265 403 323 415
rect 265 227 277 403
rect 311 227 323 403
rect 265 215 323 227
rect 395 227 407 603
rect 441 227 453 603
rect 395 215 453 227
rect 513 603 571 615
rect 513 227 525 603
rect 559 227 571 603
rect 513 215 571 227
rect 631 603 689 615
rect 631 227 643 603
rect 677 227 689 603
rect 631 215 689 227
rect 749 603 807 615
rect 749 227 761 603
rect 795 227 807 603
rect 749 215 807 227
rect 867 603 925 615
rect 867 227 879 603
rect 913 227 925 603
rect 867 215 925 227
rect 985 603 1043 615
rect 985 227 997 603
rect 1031 227 1043 603
rect 985 215 1043 227
rect 1103 603 1161 615
rect 1103 227 1115 603
rect 1149 227 1161 603
rect 2463 605 2521 617
rect 1103 215 1161 227
rect 1232 403 1290 415
rect 1232 227 1244 403
rect 1278 227 1290 403
rect 1232 215 1290 227
rect 1350 403 1408 415
rect 1350 227 1362 403
rect 1396 227 1408 403
rect 1350 215 1408 227
rect 1468 403 1526 415
rect 1468 227 1480 403
rect 1514 227 1526 403
rect 1468 215 1526 227
rect 1586 403 1644 415
rect 1586 227 1598 403
rect 1632 227 1644 403
rect 1586 215 1644 227
rect 1979 405 2037 417
rect 1979 229 1991 405
rect 2025 229 2037 405
rect 1979 217 2037 229
rect 2097 405 2155 417
rect 2097 229 2109 405
rect 2143 229 2155 405
rect 2097 217 2155 229
rect 2215 405 2273 417
rect 2215 229 2227 405
rect 2261 229 2273 405
rect 2215 217 2273 229
rect 2333 405 2391 417
rect 2333 229 2345 405
rect 2379 229 2391 405
rect 2333 217 2391 229
rect 2463 229 2475 605
rect 2509 229 2521 605
rect 2463 217 2521 229
rect 2581 605 2639 617
rect 2581 229 2593 605
rect 2627 229 2639 605
rect 2581 217 2639 229
rect 2699 605 2757 617
rect 2699 229 2711 605
rect 2745 229 2757 605
rect 2699 217 2757 229
rect 2817 605 2875 617
rect 2817 229 2829 605
rect 2863 229 2875 605
rect 2817 217 2875 229
rect 2935 605 2993 617
rect 2935 229 2947 605
rect 2981 229 2993 605
rect 2935 217 2993 229
rect 3053 605 3111 617
rect 3053 229 3065 605
rect 3099 229 3111 605
rect 3053 217 3111 229
rect 3171 605 3229 617
rect 3171 229 3183 605
rect 3217 229 3229 605
rect 4532 603 4590 615
rect 3171 217 3229 229
rect 3300 405 3358 417
rect 3300 229 3312 405
rect 3346 229 3358 405
rect 3300 217 3358 229
rect 3418 405 3476 417
rect 3418 229 3430 405
rect 3464 229 3476 405
rect 3418 217 3476 229
rect 3536 405 3594 417
rect 3536 229 3548 405
rect 3582 229 3594 405
rect 3536 217 3594 229
rect 3654 405 3712 417
rect 3654 229 3666 405
rect 3700 229 3712 405
rect 3654 217 3712 229
rect 4048 403 4106 415
rect 4048 227 4060 403
rect 4094 227 4106 403
rect 338 -90 396 -78
rect 338 -466 350 -90
rect 384 -466 396 -90
rect 338 -478 396 -466
rect 456 -90 514 -78
rect 456 -466 468 -90
rect 502 -466 514 -90
rect 456 -478 514 -466
rect 574 -90 632 -78
rect 574 -466 586 -90
rect 620 -466 632 -90
rect 574 -478 632 -466
rect 692 -90 750 -78
rect 692 -466 704 -90
rect 738 -466 750 -90
rect 692 -478 750 -466
rect 810 -90 868 -78
rect 810 -466 822 -90
rect 856 -466 868 -90
rect 810 -478 868 -466
rect 928 -90 986 -78
rect 928 -466 940 -90
rect 974 -466 986 -90
rect 928 -478 986 -466
rect 1046 -90 1104 -78
rect 1046 -466 1058 -90
rect 1092 -466 1104 -90
rect 1046 -478 1104 -466
rect 4048 215 4106 227
rect 4166 403 4224 415
rect 4166 227 4178 403
rect 4212 227 4224 403
rect 4166 215 4224 227
rect 4284 403 4342 415
rect 4284 227 4296 403
rect 4330 227 4342 403
rect 4284 215 4342 227
rect 4402 403 4460 415
rect 4402 227 4414 403
rect 4448 227 4460 403
rect 4402 215 4460 227
rect 4532 227 4544 603
rect 4578 227 4590 603
rect 4532 215 4590 227
rect 4650 603 4708 615
rect 4650 227 4662 603
rect 4696 227 4708 603
rect 4650 215 4708 227
rect 4768 603 4826 615
rect 4768 227 4780 603
rect 4814 227 4826 603
rect 4768 215 4826 227
rect 4886 603 4944 615
rect 4886 227 4898 603
rect 4932 227 4944 603
rect 4886 215 4944 227
rect 5004 603 5062 615
rect 5004 227 5016 603
rect 5050 227 5062 603
rect 5004 215 5062 227
rect 5122 603 5180 615
rect 5122 227 5134 603
rect 5168 227 5180 603
rect 5122 215 5180 227
rect 5240 603 5298 615
rect 5240 227 5252 603
rect 5286 227 5298 603
rect 6600 605 6658 617
rect 5240 215 5298 227
rect 5369 403 5427 415
rect 5369 227 5381 403
rect 5415 227 5427 403
rect 5369 215 5427 227
rect 5487 403 5545 415
rect 5487 227 5499 403
rect 5533 227 5545 403
rect 5487 215 5545 227
rect 5605 403 5663 415
rect 5605 227 5617 403
rect 5651 227 5663 403
rect 5605 215 5663 227
rect 5723 403 5781 415
rect 5723 227 5735 403
rect 5769 227 5781 403
rect 5723 215 5781 227
rect 6116 405 6174 417
rect 6116 229 6128 405
rect 6162 229 6174 405
rect 6116 217 6174 229
rect 6234 405 6292 417
rect 6234 229 6246 405
rect 6280 229 6292 405
rect 6234 217 6292 229
rect 6352 405 6410 417
rect 6352 229 6364 405
rect 6398 229 6410 405
rect 6352 217 6410 229
rect 6470 405 6528 417
rect 6470 229 6482 405
rect 6516 229 6528 405
rect 6470 217 6528 229
rect 6600 229 6612 605
rect 6646 229 6658 605
rect 6600 217 6658 229
rect 6718 605 6776 617
rect 6718 229 6730 605
rect 6764 229 6776 605
rect 6718 217 6776 229
rect 6836 605 6894 617
rect 6836 229 6848 605
rect 6882 229 6894 605
rect 6836 217 6894 229
rect 6954 605 7012 617
rect 6954 229 6966 605
rect 7000 229 7012 605
rect 6954 217 7012 229
rect 7072 605 7130 617
rect 7072 229 7084 605
rect 7118 229 7130 605
rect 7072 217 7130 229
rect 7190 605 7248 617
rect 7190 229 7202 605
rect 7236 229 7248 605
rect 7190 217 7248 229
rect 7308 605 7366 617
rect 7308 229 7320 605
rect 7354 229 7366 605
rect 8669 605 8727 617
rect 7308 217 7366 229
rect 7437 405 7495 417
rect 7437 229 7449 405
rect 7483 229 7495 405
rect 7437 217 7495 229
rect 7555 405 7613 417
rect 7555 229 7567 405
rect 7601 229 7613 405
rect 7555 217 7613 229
rect 7673 405 7731 417
rect 7673 229 7685 405
rect 7719 229 7731 405
rect 7673 217 7731 229
rect 7791 405 7849 417
rect 7791 229 7803 405
rect 7837 229 7849 405
rect 7791 217 7849 229
rect 8185 405 8243 417
rect 8185 229 8197 405
rect 8231 229 8243 405
rect 8185 217 8243 229
rect 8303 405 8361 417
rect 8303 229 8315 405
rect 8349 229 8361 405
rect 8303 217 8361 229
rect 8421 405 8479 417
rect 8421 229 8433 405
rect 8467 229 8479 405
rect 8421 217 8479 229
rect 8539 405 8597 417
rect 8539 229 8551 405
rect 8585 229 8597 405
rect 8539 217 8597 229
rect 8669 229 8681 605
rect 8715 229 8727 605
rect 8669 217 8727 229
rect 8787 605 8845 617
rect 8787 229 8799 605
rect 8833 229 8845 605
rect 8787 217 8845 229
rect 8905 605 8963 617
rect 8905 229 8917 605
rect 8951 229 8963 605
rect 8905 217 8963 229
rect 9023 605 9081 617
rect 9023 229 9035 605
rect 9069 229 9081 605
rect 9023 217 9081 229
rect 9141 605 9199 617
rect 9141 229 9153 605
rect 9187 229 9199 605
rect 9141 217 9199 229
rect 9259 605 9317 617
rect 9259 229 9271 605
rect 9305 229 9317 605
rect 9259 217 9317 229
rect 9377 605 9435 617
rect 9377 229 9389 605
rect 9423 229 9435 605
rect 10737 607 10795 619
rect 9377 217 9435 229
rect 9506 405 9564 417
rect 9506 229 9518 405
rect 9552 229 9564 405
rect 9506 217 9564 229
rect 9624 405 9682 417
rect 9624 229 9636 405
rect 9670 229 9682 405
rect 9624 217 9682 229
rect 9742 405 9800 417
rect 9742 229 9754 405
rect 9788 229 9800 405
rect 9742 217 9800 229
rect 9860 405 9918 417
rect 9860 229 9872 405
rect 9906 229 9918 405
rect 9860 217 9918 229
rect 10253 407 10311 419
rect 10253 231 10265 407
rect 10299 231 10311 407
rect 10253 219 10311 231
rect 10371 407 10429 419
rect 10371 231 10383 407
rect 10417 231 10429 407
rect 10371 219 10429 231
rect 10489 407 10547 419
rect 10489 231 10501 407
rect 10535 231 10547 407
rect 10489 219 10547 231
rect 10607 407 10665 419
rect 10607 231 10619 407
rect 10653 231 10665 407
rect 10607 219 10665 231
rect 10737 231 10749 607
rect 10783 231 10795 607
rect 10737 219 10795 231
rect 10855 607 10913 619
rect 10855 231 10867 607
rect 10901 231 10913 607
rect 10855 219 10913 231
rect 10973 607 11031 619
rect 10973 231 10985 607
rect 11019 231 11031 607
rect 10973 219 11031 231
rect 11091 607 11149 619
rect 11091 231 11103 607
rect 11137 231 11149 607
rect 11091 219 11149 231
rect 11209 607 11267 619
rect 11209 231 11221 607
rect 11255 231 11267 607
rect 11209 219 11267 231
rect 11327 607 11385 619
rect 11327 231 11339 607
rect 11373 231 11385 607
rect 11327 219 11385 231
rect 11445 607 11503 619
rect 11445 231 11457 607
rect 11491 231 11503 607
rect 12806 605 12864 617
rect 11445 219 11503 231
rect 11574 407 11632 419
rect 11574 231 11586 407
rect 11620 231 11632 407
rect 11574 219 11632 231
rect 11692 407 11750 419
rect 11692 231 11704 407
rect 11738 231 11750 407
rect 11692 219 11750 231
rect 11810 407 11868 419
rect 11810 231 11822 407
rect 11856 231 11868 407
rect 11810 219 11868 231
rect 11928 407 11986 419
rect 11928 231 11940 407
rect 11974 231 11986 407
rect 11928 219 11986 231
rect 12322 405 12380 417
rect 12322 229 12334 405
rect 12368 229 12380 405
rect 2406 -88 2464 -76
rect 2406 -464 2418 -88
rect 2452 -464 2464 -88
rect 2406 -476 2464 -464
rect 2524 -88 2582 -76
rect 2524 -464 2536 -88
rect 2570 -464 2582 -88
rect 2524 -476 2582 -464
rect 2642 -88 2700 -76
rect 2642 -464 2654 -88
rect 2688 -464 2700 -88
rect 2642 -476 2700 -464
rect 2760 -88 2818 -76
rect 2760 -464 2772 -88
rect 2806 -464 2818 -88
rect 2760 -476 2818 -464
rect 2878 -88 2936 -76
rect 2878 -464 2890 -88
rect 2924 -464 2936 -88
rect 2878 -476 2936 -464
rect 2996 -88 3054 -76
rect 2996 -464 3008 -88
rect 3042 -464 3054 -88
rect 2996 -476 3054 -464
rect 3114 -88 3172 -76
rect 3114 -464 3126 -88
rect 3160 -464 3172 -88
rect 3114 -476 3172 -464
rect 4475 -90 4533 -78
rect 4475 -466 4487 -90
rect 4521 -466 4533 -90
rect 4475 -478 4533 -466
rect 4593 -90 4651 -78
rect 4593 -466 4605 -90
rect 4639 -466 4651 -90
rect 4593 -478 4651 -466
rect 4711 -90 4769 -78
rect 4711 -466 4723 -90
rect 4757 -466 4769 -90
rect 4711 -478 4769 -466
rect 4829 -90 4887 -78
rect 4829 -466 4841 -90
rect 4875 -466 4887 -90
rect 4829 -478 4887 -466
rect 4947 -90 5005 -78
rect 4947 -466 4959 -90
rect 4993 -466 5005 -90
rect 4947 -478 5005 -466
rect 5065 -90 5123 -78
rect 5065 -466 5077 -90
rect 5111 -466 5123 -90
rect 5065 -478 5123 -466
rect 5183 -90 5241 -78
rect 5183 -466 5195 -90
rect 5229 -466 5241 -90
rect 5183 -478 5241 -466
rect 6543 -88 6601 -76
rect 6543 -464 6555 -88
rect 6589 -464 6601 -88
rect 6543 -476 6601 -464
rect 6661 -88 6719 -76
rect 6661 -464 6673 -88
rect 6707 -464 6719 -88
rect 6661 -476 6719 -464
rect 6779 -88 6837 -76
rect 6779 -464 6791 -88
rect 6825 -464 6837 -88
rect 6779 -476 6837 -464
rect 6897 -88 6955 -76
rect 6897 -464 6909 -88
rect 6943 -464 6955 -88
rect 6897 -476 6955 -464
rect 7015 -88 7073 -76
rect 7015 -464 7027 -88
rect 7061 -464 7073 -88
rect 7015 -476 7073 -464
rect 7133 -88 7191 -76
rect 7133 -464 7145 -88
rect 7179 -464 7191 -88
rect 7133 -476 7191 -464
rect 7251 -88 7309 -76
rect 7251 -464 7263 -88
rect 7297 -464 7309 -88
rect 7251 -476 7309 -464
rect 8612 -88 8670 -76
rect 8612 -464 8624 -88
rect 8658 -464 8670 -88
rect 8612 -476 8670 -464
rect 8730 -88 8788 -76
rect 8730 -464 8742 -88
rect 8776 -464 8788 -88
rect 8730 -476 8788 -464
rect 8848 -88 8906 -76
rect 8848 -464 8860 -88
rect 8894 -464 8906 -88
rect 8848 -476 8906 -464
rect 8966 -88 9024 -76
rect 8966 -464 8978 -88
rect 9012 -464 9024 -88
rect 8966 -476 9024 -464
rect 9084 -88 9142 -76
rect 9084 -464 9096 -88
rect 9130 -464 9142 -88
rect 9084 -476 9142 -464
rect 9202 -88 9260 -76
rect 9202 -464 9214 -88
rect 9248 -464 9260 -88
rect 9202 -476 9260 -464
rect 9320 -88 9378 -76
rect 9320 -464 9332 -88
rect 9366 -464 9378 -88
rect 9320 -476 9378 -464
rect 12322 217 12380 229
rect 12440 405 12498 417
rect 12440 229 12452 405
rect 12486 229 12498 405
rect 12440 217 12498 229
rect 12558 405 12616 417
rect 12558 229 12570 405
rect 12604 229 12616 405
rect 12558 217 12616 229
rect 12676 405 12734 417
rect 12676 229 12688 405
rect 12722 229 12734 405
rect 12676 217 12734 229
rect 12806 229 12818 605
rect 12852 229 12864 605
rect 12806 217 12864 229
rect 12924 605 12982 617
rect 12924 229 12936 605
rect 12970 229 12982 605
rect 12924 217 12982 229
rect 13042 605 13100 617
rect 13042 229 13054 605
rect 13088 229 13100 605
rect 13042 217 13100 229
rect 13160 605 13218 617
rect 13160 229 13172 605
rect 13206 229 13218 605
rect 13160 217 13218 229
rect 13278 605 13336 617
rect 13278 229 13290 605
rect 13324 229 13336 605
rect 13278 217 13336 229
rect 13396 605 13454 617
rect 13396 229 13408 605
rect 13442 229 13454 605
rect 13396 217 13454 229
rect 13514 605 13572 617
rect 13514 229 13526 605
rect 13560 229 13572 605
rect 14874 607 14932 619
rect 13514 217 13572 229
rect 13643 405 13701 417
rect 13643 229 13655 405
rect 13689 229 13701 405
rect 13643 217 13701 229
rect 13761 405 13819 417
rect 13761 229 13773 405
rect 13807 229 13819 405
rect 13761 217 13819 229
rect 13879 405 13937 417
rect 13879 229 13891 405
rect 13925 229 13937 405
rect 13879 217 13937 229
rect 13997 405 14055 417
rect 13997 229 14009 405
rect 14043 229 14055 405
rect 13997 217 14055 229
rect 14390 407 14448 419
rect 14390 231 14402 407
rect 14436 231 14448 407
rect 14390 219 14448 231
rect 14508 407 14566 419
rect 14508 231 14520 407
rect 14554 231 14566 407
rect 14508 219 14566 231
rect 14626 407 14684 419
rect 14626 231 14638 407
rect 14672 231 14684 407
rect 14626 219 14684 231
rect 14744 407 14802 419
rect 14744 231 14756 407
rect 14790 231 14802 407
rect 14744 219 14802 231
rect 14874 231 14886 607
rect 14920 231 14932 607
rect 14874 219 14932 231
rect 14992 607 15050 619
rect 14992 231 15004 607
rect 15038 231 15050 607
rect 14992 219 15050 231
rect 15110 607 15168 619
rect 15110 231 15122 607
rect 15156 231 15168 607
rect 15110 219 15168 231
rect 15228 607 15286 619
rect 15228 231 15240 607
rect 15274 231 15286 607
rect 15228 219 15286 231
rect 15346 607 15404 619
rect 15346 231 15358 607
rect 15392 231 15404 607
rect 15346 219 15404 231
rect 15464 607 15522 619
rect 15464 231 15476 607
rect 15510 231 15522 607
rect 15464 219 15522 231
rect 15582 607 15640 619
rect 15582 231 15594 607
rect 15628 231 15640 607
rect 15582 219 15640 231
rect 15711 407 15769 419
rect 15711 231 15723 407
rect 15757 231 15769 407
rect 15711 219 15769 231
rect 15829 407 15887 419
rect 15829 231 15841 407
rect 15875 231 15887 407
rect 15829 219 15887 231
rect 15947 407 16005 419
rect 15947 231 15959 407
rect 15993 231 16005 407
rect 15947 219 16005 231
rect 16065 407 16123 419
rect 16065 231 16077 407
rect 16111 231 16123 407
rect 16065 219 16123 231
rect 10680 -86 10738 -74
rect 10680 -462 10692 -86
rect 10726 -462 10738 -86
rect 10680 -474 10738 -462
rect 10798 -86 10856 -74
rect 10798 -462 10810 -86
rect 10844 -462 10856 -86
rect 10798 -474 10856 -462
rect 10916 -86 10974 -74
rect 10916 -462 10928 -86
rect 10962 -462 10974 -86
rect 10916 -474 10974 -462
rect 11034 -86 11092 -74
rect 11034 -462 11046 -86
rect 11080 -462 11092 -86
rect 11034 -474 11092 -462
rect 11152 -86 11210 -74
rect 11152 -462 11164 -86
rect 11198 -462 11210 -86
rect 11152 -474 11210 -462
rect 11270 -86 11328 -74
rect 11270 -462 11282 -86
rect 11316 -462 11328 -86
rect 11270 -474 11328 -462
rect 11388 -86 11446 -74
rect 11388 -462 11400 -86
rect 11434 -462 11446 -86
rect 11388 -474 11446 -462
rect 12749 -88 12807 -76
rect 12749 -464 12761 -88
rect 12795 -464 12807 -88
rect 12749 -476 12807 -464
rect 12867 -88 12925 -76
rect 12867 -464 12879 -88
rect 12913 -464 12925 -88
rect 12867 -476 12925 -464
rect 12985 -88 13043 -76
rect 12985 -464 12997 -88
rect 13031 -464 13043 -88
rect 12985 -476 13043 -464
rect 13103 -88 13161 -76
rect 13103 -464 13115 -88
rect 13149 -464 13161 -88
rect 13103 -476 13161 -464
rect 13221 -88 13279 -76
rect 13221 -464 13233 -88
rect 13267 -464 13279 -88
rect 13221 -476 13279 -464
rect 13339 -88 13397 -76
rect 13339 -464 13351 -88
rect 13385 -464 13397 -88
rect 13339 -476 13397 -464
rect 13457 -88 13515 -76
rect 13457 -464 13469 -88
rect 13503 -464 13515 -88
rect 13457 -476 13515 -464
rect 14817 -86 14875 -74
rect 14817 -462 14829 -86
rect 14863 -462 14875 -86
rect 14817 -474 14875 -462
rect 14935 -86 14993 -74
rect 14935 -462 14947 -86
rect 14981 -462 14993 -86
rect 14935 -474 14993 -462
rect 15053 -86 15111 -74
rect 15053 -462 15065 -86
rect 15099 -462 15111 -86
rect 15053 -474 15111 -462
rect 15171 -86 15229 -74
rect 15171 -462 15183 -86
rect 15217 -462 15229 -86
rect 15171 -474 15229 -462
rect 15289 -86 15347 -74
rect 15289 -462 15301 -86
rect 15335 -462 15347 -86
rect 15289 -474 15347 -462
rect 15407 -86 15465 -74
rect 15407 -462 15419 -86
rect 15453 -462 15465 -86
rect 15407 -474 15465 -462
rect 15525 -86 15583 -74
rect 15525 -462 15537 -86
rect 15571 -462 15583 -86
rect 15525 -474 15583 -462
<< ndiffc >>
rect 48 -998 82 -822
rect 166 -998 200 -822
rect 468 -1198 502 -822
rect 586 -1198 620 -822
rect 704 -1198 738 -822
rect 822 -1198 856 -822
rect 940 -1198 974 -822
rect 1346 -998 1380 -822
rect 1464 -998 1498 -822
rect 2116 -996 2150 -820
rect 2234 -996 2268 -820
rect 2536 -1196 2570 -820
rect 2654 -1196 2688 -820
rect 2772 -1196 2806 -820
rect 2890 -1196 2924 -820
rect 3008 -1196 3042 -820
rect 3414 -996 3448 -820
rect 3532 -996 3566 -820
rect 4185 -998 4219 -822
rect 4303 -998 4337 -822
rect 4605 -1198 4639 -822
rect 4723 -1198 4757 -822
rect 4841 -1198 4875 -822
rect 4959 -1198 4993 -822
rect 5077 -1198 5111 -822
rect 5483 -998 5517 -822
rect 5601 -998 5635 -822
rect 6253 -996 6287 -820
rect 6371 -996 6405 -820
rect 6673 -1196 6707 -820
rect 6791 -1196 6825 -820
rect 6909 -1196 6943 -820
rect 7027 -1196 7061 -820
rect 7145 -1196 7179 -820
rect 7551 -996 7585 -820
rect 7669 -996 7703 -820
rect 8322 -996 8356 -820
rect 8440 -996 8474 -820
rect 8742 -1196 8776 -820
rect 8860 -1196 8894 -820
rect 8978 -1196 9012 -820
rect 9096 -1196 9130 -820
rect 9214 -1196 9248 -820
rect 9620 -996 9654 -820
rect 9738 -996 9772 -820
rect 10390 -994 10424 -818
rect 10508 -994 10542 -818
rect 10810 -1194 10844 -818
rect 10928 -1194 10962 -818
rect 11046 -1194 11080 -818
rect 11164 -1194 11198 -818
rect 11282 -1194 11316 -818
rect 11688 -994 11722 -818
rect 11806 -994 11840 -818
rect 12459 -996 12493 -820
rect 12577 -996 12611 -820
rect 12879 -1196 12913 -820
rect 12997 -1196 13031 -820
rect 13115 -1196 13149 -820
rect 13233 -1196 13267 -820
rect 13351 -1196 13385 -820
rect 13757 -996 13791 -820
rect 13875 -996 13909 -820
rect 14527 -994 14561 -818
rect 14645 -994 14679 -818
rect 14947 -1194 14981 -818
rect 15065 -1194 15099 -818
rect 15183 -1194 15217 -818
rect 15301 -1194 15335 -818
rect 15419 -1194 15453 -818
rect 15825 -994 15859 -818
rect 15943 -994 15977 -818
<< pdiffc >>
rect -77 227 -43 403
rect 41 227 75 403
rect 159 227 193 403
rect 277 227 311 403
rect 407 227 441 603
rect 525 227 559 603
rect 643 227 677 603
rect 761 227 795 603
rect 879 227 913 603
rect 997 227 1031 603
rect 1115 227 1149 603
rect 1244 227 1278 403
rect 1362 227 1396 403
rect 1480 227 1514 403
rect 1598 227 1632 403
rect 1991 229 2025 405
rect 2109 229 2143 405
rect 2227 229 2261 405
rect 2345 229 2379 405
rect 2475 229 2509 605
rect 2593 229 2627 605
rect 2711 229 2745 605
rect 2829 229 2863 605
rect 2947 229 2981 605
rect 3065 229 3099 605
rect 3183 229 3217 605
rect 3312 229 3346 405
rect 3430 229 3464 405
rect 3548 229 3582 405
rect 3666 229 3700 405
rect 4060 227 4094 403
rect 350 -466 384 -90
rect 468 -466 502 -90
rect 586 -466 620 -90
rect 704 -466 738 -90
rect 822 -466 856 -90
rect 940 -466 974 -90
rect 1058 -466 1092 -90
rect 4178 227 4212 403
rect 4296 227 4330 403
rect 4414 227 4448 403
rect 4544 227 4578 603
rect 4662 227 4696 603
rect 4780 227 4814 603
rect 4898 227 4932 603
rect 5016 227 5050 603
rect 5134 227 5168 603
rect 5252 227 5286 603
rect 5381 227 5415 403
rect 5499 227 5533 403
rect 5617 227 5651 403
rect 5735 227 5769 403
rect 6128 229 6162 405
rect 6246 229 6280 405
rect 6364 229 6398 405
rect 6482 229 6516 405
rect 6612 229 6646 605
rect 6730 229 6764 605
rect 6848 229 6882 605
rect 6966 229 7000 605
rect 7084 229 7118 605
rect 7202 229 7236 605
rect 7320 229 7354 605
rect 7449 229 7483 405
rect 7567 229 7601 405
rect 7685 229 7719 405
rect 7803 229 7837 405
rect 8197 229 8231 405
rect 8315 229 8349 405
rect 8433 229 8467 405
rect 8551 229 8585 405
rect 8681 229 8715 605
rect 8799 229 8833 605
rect 8917 229 8951 605
rect 9035 229 9069 605
rect 9153 229 9187 605
rect 9271 229 9305 605
rect 9389 229 9423 605
rect 9518 229 9552 405
rect 9636 229 9670 405
rect 9754 229 9788 405
rect 9872 229 9906 405
rect 10265 231 10299 407
rect 10383 231 10417 407
rect 10501 231 10535 407
rect 10619 231 10653 407
rect 10749 231 10783 607
rect 10867 231 10901 607
rect 10985 231 11019 607
rect 11103 231 11137 607
rect 11221 231 11255 607
rect 11339 231 11373 607
rect 11457 231 11491 607
rect 11586 231 11620 407
rect 11704 231 11738 407
rect 11822 231 11856 407
rect 11940 231 11974 407
rect 12334 229 12368 405
rect 2418 -464 2452 -88
rect 2536 -464 2570 -88
rect 2654 -464 2688 -88
rect 2772 -464 2806 -88
rect 2890 -464 2924 -88
rect 3008 -464 3042 -88
rect 3126 -464 3160 -88
rect 4487 -466 4521 -90
rect 4605 -466 4639 -90
rect 4723 -466 4757 -90
rect 4841 -466 4875 -90
rect 4959 -466 4993 -90
rect 5077 -466 5111 -90
rect 5195 -466 5229 -90
rect 6555 -464 6589 -88
rect 6673 -464 6707 -88
rect 6791 -464 6825 -88
rect 6909 -464 6943 -88
rect 7027 -464 7061 -88
rect 7145 -464 7179 -88
rect 7263 -464 7297 -88
rect 8624 -464 8658 -88
rect 8742 -464 8776 -88
rect 8860 -464 8894 -88
rect 8978 -464 9012 -88
rect 9096 -464 9130 -88
rect 9214 -464 9248 -88
rect 9332 -464 9366 -88
rect 12452 229 12486 405
rect 12570 229 12604 405
rect 12688 229 12722 405
rect 12818 229 12852 605
rect 12936 229 12970 605
rect 13054 229 13088 605
rect 13172 229 13206 605
rect 13290 229 13324 605
rect 13408 229 13442 605
rect 13526 229 13560 605
rect 13655 229 13689 405
rect 13773 229 13807 405
rect 13891 229 13925 405
rect 14009 229 14043 405
rect 14402 231 14436 407
rect 14520 231 14554 407
rect 14638 231 14672 407
rect 14756 231 14790 407
rect 14886 231 14920 607
rect 15004 231 15038 607
rect 15122 231 15156 607
rect 15240 231 15274 607
rect 15358 231 15392 607
rect 15476 231 15510 607
rect 15594 231 15628 607
rect 15723 231 15757 407
rect 15841 231 15875 407
rect 15959 231 15993 407
rect 16077 231 16111 407
rect 10692 -462 10726 -86
rect 10810 -462 10844 -86
rect 10928 -462 10962 -86
rect 11046 -462 11080 -86
rect 11164 -462 11198 -86
rect 11282 -462 11316 -86
rect 11400 -462 11434 -86
rect 12761 -464 12795 -88
rect 12879 -464 12913 -88
rect 12997 -464 13031 -88
rect 13115 -464 13149 -88
rect 13233 -464 13267 -88
rect 13351 -464 13385 -88
rect 13469 -464 13503 -88
rect 14829 -462 14863 -86
rect 14947 -462 14981 -86
rect 15065 -462 15099 -86
rect 15183 -462 15217 -86
rect 15301 -462 15335 -86
rect 15419 -462 15453 -86
rect 15537 -462 15571 -86
<< psubdiff >>
rect 600 -1386 852 -1366
rect 600 -1442 658 -1386
rect 790 -1442 852 -1386
rect 600 -1464 852 -1442
rect 2668 -1384 2920 -1364
rect 2668 -1440 2726 -1384
rect 2858 -1440 2920 -1384
rect 2668 -1462 2920 -1440
rect 4737 -1386 4989 -1366
rect 4737 -1442 4795 -1386
rect 4927 -1442 4989 -1386
rect 4737 -1464 4989 -1442
rect 6805 -1384 7057 -1364
rect 6805 -1440 6863 -1384
rect 6995 -1440 7057 -1384
rect 6805 -1462 7057 -1440
rect 8874 -1384 9126 -1364
rect 8874 -1440 8932 -1384
rect 9064 -1440 9126 -1384
rect 8874 -1462 9126 -1440
rect 10942 -1382 11194 -1362
rect 10942 -1438 11000 -1382
rect 11132 -1438 11194 -1382
rect 10942 -1460 11194 -1438
rect 13011 -1384 13263 -1364
rect 13011 -1440 13069 -1384
rect 13201 -1440 13263 -1384
rect 13011 -1462 13263 -1440
rect 15079 -1382 15331 -1362
rect 15079 -1438 15137 -1382
rect 15269 -1438 15331 -1382
rect 15079 -1460 15331 -1438
<< nsubdiff >>
rect 584 874 984 926
rect 584 830 708 874
rect 830 830 984 874
rect 584 782 984 830
rect 2652 876 3052 928
rect 2652 832 2776 876
rect 2898 832 3052 876
rect 2652 784 3052 832
rect 4721 874 5121 926
rect 4721 830 4845 874
rect 4967 830 5121 874
rect 4721 782 5121 830
rect 6789 876 7189 928
rect 6789 832 6913 876
rect 7035 832 7189 876
rect 6789 784 7189 832
rect 8858 876 9258 928
rect 8858 832 8982 876
rect 9104 832 9258 876
rect 8858 784 9258 832
rect 10926 878 11326 930
rect 10926 834 11050 878
rect 11172 834 11326 878
rect 10926 786 11326 834
rect 12995 876 13395 928
rect 12995 832 13119 876
rect 13241 832 13395 876
rect 12995 784 13395 832
rect 15063 878 15463 930
rect 15063 834 15187 878
rect 15309 834 15463 878
rect 15063 786 15463 834
<< psubdiffcont >>
rect 658 -1442 790 -1386
rect 2726 -1440 2858 -1384
rect 4795 -1442 4927 -1386
rect 6863 -1440 6995 -1384
rect 8932 -1440 9064 -1384
rect 11000 -1438 11132 -1382
rect 13069 -1440 13201 -1384
rect 15137 -1438 15269 -1382
<< nsubdiffcont >>
rect 708 830 830 874
rect 2776 832 2898 876
rect 4845 830 4967 874
rect 6913 832 7035 876
rect 8982 832 9104 876
rect 11050 834 11172 878
rect 13119 832 13241 876
rect 15187 834 15309 878
<< poly >>
rect 453 630 749 681
rect 453 615 513 630
rect 571 615 631 630
rect 689 615 749 630
rect 807 615 867 641
rect 925 615 985 641
rect 1043 615 1103 641
rect 2521 632 2817 683
rect 2521 617 2581 632
rect 2639 617 2699 632
rect 2757 617 2817 632
rect 2875 617 2935 643
rect 2993 617 3053 643
rect 3111 617 3171 643
rect 4590 630 4886 681
rect -31 415 29 441
rect 87 415 147 441
rect 205 415 265 441
rect 1290 432 1586 483
rect 1290 415 1350 432
rect 1408 415 1468 432
rect 1526 415 1586 432
rect 2037 417 2097 443
rect 2155 417 2215 443
rect 2273 417 2333 443
rect 4590 615 4650 630
rect 4708 615 4768 630
rect 4826 615 4886 630
rect 4944 615 5004 641
rect 5062 615 5122 641
rect 5180 615 5240 641
rect 6658 632 6954 683
rect 6658 617 6718 632
rect 6776 617 6836 632
rect 6894 617 6954 632
rect 7012 617 7072 643
rect 7130 617 7190 643
rect 7248 617 7308 643
rect 8727 632 9023 683
rect 8727 617 8787 632
rect 8845 617 8905 632
rect 8963 617 9023 632
rect 9081 617 9141 643
rect 9199 617 9259 643
rect 9317 617 9377 643
rect 10795 634 11091 685
rect 10795 619 10855 634
rect 10913 619 10973 634
rect 11031 619 11091 634
rect 11149 619 11209 645
rect 11267 619 11327 645
rect 11385 619 11445 645
rect 12864 632 13160 683
rect 3358 434 3654 485
rect 3358 417 3418 434
rect 3476 417 3536 434
rect 3594 417 3654 434
rect 4106 415 4166 441
rect 4224 415 4284 441
rect 4342 415 4402 441
rect -31 198 29 215
rect 87 198 147 215
rect 205 198 265 215
rect 453 198 513 215
rect -31 147 513 198
rect 571 189 631 215
rect 689 189 749 215
rect 807 196 867 215
rect 925 196 985 215
rect 1043 196 1103 215
rect 1290 196 1350 215
rect 1408 196 1468 215
rect 94 -132 154 147
rect 807 145 1350 196
rect 1392 189 1468 196
rect 1526 189 1586 215
rect 2037 200 2097 217
rect 2155 200 2215 217
rect 2273 200 2333 217
rect 2521 200 2581 217
rect 1392 145 1467 189
rect 2037 149 2581 200
rect 2639 191 2699 217
rect 2757 191 2817 217
rect 2875 198 2935 217
rect 2993 198 3053 217
rect 3111 198 3171 217
rect 3358 198 3418 217
rect 3476 198 3536 217
rect 1392 58 1452 145
rect 1324 48 1452 58
rect 1324 14 1340 48
rect 1374 14 1452 48
rect 396 -55 692 5
rect 396 -78 456 -55
rect 514 -78 574 -55
rect 632 -78 692 -55
rect 750 -54 1046 6
rect 1324 4 1452 14
rect 750 -78 810 -54
rect 868 -78 928 -54
rect 986 -78 1046 -54
rect -70 -146 154 -132
rect -70 -180 -54 -146
rect -20 -180 154 -146
rect -70 -192 154 -180
rect 94 -705 154 -192
rect 396 -504 456 -478
rect 364 -645 431 -638
rect 514 -645 574 -478
rect 632 -504 692 -478
rect 750 -504 810 -478
rect 364 -654 574 -645
rect 364 -688 380 -654
rect 414 -688 574 -654
rect 364 -704 574 -688
rect 94 -721 245 -705
rect 94 -755 195 -721
rect 229 -755 245 -721
rect 94 -771 245 -755
rect 94 -810 154 -771
rect 514 -810 574 -704
rect 868 -645 928 -478
rect 986 -504 1046 -478
rect 1011 -645 1078 -638
rect 868 -654 1078 -645
rect 868 -688 1028 -654
rect 1062 -688 1078 -654
rect 868 -704 1078 -688
rect 630 -738 696 -722
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 630 -788 696 -772
rect 748 -737 814 -722
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 748 -787 814 -771
rect 632 -810 692 -788
rect 750 -810 810 -787
rect 868 -810 928 -704
rect 1392 -706 1452 4
rect 2162 -130 2222 149
rect 2875 147 3418 198
rect 3460 191 3536 198
rect 3594 191 3654 217
rect 5427 432 5723 483
rect 5427 415 5487 432
rect 5545 415 5605 432
rect 5663 415 5723 432
rect 6174 417 6234 443
rect 6292 417 6352 443
rect 6410 417 6470 443
rect 7495 434 7791 485
rect 7495 417 7555 434
rect 7613 417 7673 434
rect 7731 417 7791 434
rect 8243 417 8303 443
rect 8361 417 8421 443
rect 8479 417 8539 443
rect 9564 434 9860 485
rect 9564 417 9624 434
rect 9682 417 9742 434
rect 9800 417 9860 434
rect 10311 419 10371 445
rect 10429 419 10489 445
rect 10547 419 10607 445
rect 12864 617 12924 632
rect 12982 617 13042 632
rect 13100 617 13160 632
rect 13218 617 13278 643
rect 13336 617 13396 643
rect 13454 617 13514 643
rect 14932 634 15228 685
rect 14932 619 14992 634
rect 15050 619 15110 634
rect 15168 619 15228 634
rect 15286 619 15346 645
rect 15404 619 15464 645
rect 15522 619 15582 645
rect 11632 436 11928 487
rect 11632 419 11692 436
rect 11750 419 11810 436
rect 11868 419 11928 436
rect 12380 417 12440 443
rect 12498 417 12558 443
rect 12616 417 12676 443
rect 4106 198 4166 215
rect 4224 198 4284 215
rect 4342 198 4402 215
rect 4590 198 4650 215
rect 3460 147 3535 191
rect 4106 147 4650 198
rect 4708 189 4768 215
rect 4826 189 4886 215
rect 4944 196 5004 215
rect 5062 196 5122 215
rect 5180 196 5240 215
rect 5427 196 5487 215
rect 5545 196 5605 215
rect 3460 60 3520 147
rect 3392 50 3520 60
rect 3392 16 3408 50
rect 3442 16 3520 50
rect 2464 -53 2760 7
rect 2464 -76 2524 -53
rect 2582 -76 2642 -53
rect 2700 -76 2760 -53
rect 2818 -52 3114 8
rect 3392 6 3520 16
rect 2818 -76 2878 -52
rect 2936 -76 2996 -52
rect 3054 -76 3114 -52
rect 1998 -144 2222 -130
rect 1998 -178 2014 -144
rect 2048 -178 2222 -144
rect 1998 -190 2222 -178
rect 1302 -722 1452 -706
rect 1302 -756 1318 -722
rect 1352 -756 1452 -722
rect 1302 -772 1452 -756
rect 1392 -810 1452 -772
rect 2162 -703 2222 -190
rect 2464 -502 2524 -476
rect 2432 -643 2499 -636
rect 2582 -643 2642 -476
rect 2700 -502 2760 -476
rect 2818 -502 2878 -476
rect 2432 -652 2642 -643
rect 2432 -686 2448 -652
rect 2482 -686 2642 -652
rect 2432 -702 2642 -686
rect 2162 -719 2313 -703
rect 2162 -753 2263 -719
rect 2297 -753 2313 -719
rect 2162 -769 2313 -753
rect 2162 -808 2222 -769
rect 2582 -808 2642 -702
rect 2936 -643 2996 -476
rect 3054 -502 3114 -476
rect 3079 -643 3146 -636
rect 2936 -652 3146 -643
rect 2936 -686 3096 -652
rect 3130 -686 3146 -652
rect 2936 -702 3146 -686
rect 2698 -736 2764 -720
rect 2698 -770 2714 -736
rect 2748 -770 2764 -736
rect 2698 -786 2764 -770
rect 2816 -735 2882 -720
rect 2816 -769 2832 -735
rect 2866 -769 2882 -735
rect 2816 -785 2882 -769
rect 2700 -808 2760 -786
rect 2818 -808 2878 -785
rect 2936 -808 2996 -702
rect 3460 -704 3520 6
rect 4231 -132 4291 147
rect 4944 145 5487 196
rect 5529 189 5605 196
rect 5663 189 5723 215
rect 6174 200 6234 217
rect 6292 200 6352 217
rect 6410 200 6470 217
rect 6658 200 6718 217
rect 5529 145 5604 189
rect 6174 149 6718 200
rect 6776 191 6836 217
rect 6894 191 6954 217
rect 7012 198 7072 217
rect 7130 198 7190 217
rect 7248 198 7308 217
rect 7495 198 7555 217
rect 7613 198 7673 217
rect 5529 58 5589 145
rect 5461 48 5589 58
rect 5461 14 5477 48
rect 5511 14 5589 48
rect 4533 -55 4829 5
rect 4533 -78 4593 -55
rect 4651 -78 4711 -55
rect 4769 -78 4829 -55
rect 4887 -54 5183 6
rect 5461 4 5589 14
rect 4887 -78 4947 -54
rect 5005 -78 5065 -54
rect 5123 -78 5183 -54
rect 4067 -146 4291 -132
rect 4067 -180 4083 -146
rect 4117 -180 4291 -146
rect 4067 -192 4291 -180
rect 3370 -720 3520 -704
rect 3370 -754 3386 -720
rect 3420 -754 3520 -720
rect 3370 -770 3520 -754
rect 3460 -808 3520 -770
rect 4231 -705 4291 -192
rect 4533 -504 4593 -478
rect 4501 -645 4568 -638
rect 4651 -645 4711 -478
rect 4769 -504 4829 -478
rect 4887 -504 4947 -478
rect 4501 -654 4711 -645
rect 4501 -688 4517 -654
rect 4551 -688 4711 -654
rect 4501 -704 4711 -688
rect 4231 -721 4382 -705
rect 4231 -755 4332 -721
rect 4366 -755 4382 -721
rect 4231 -771 4382 -755
rect 94 -1036 154 -1010
rect 1392 -1036 1452 -1010
rect 2162 -1034 2222 -1008
rect 4231 -810 4291 -771
rect 4651 -810 4711 -704
rect 5005 -645 5065 -478
rect 5123 -504 5183 -478
rect 5148 -645 5215 -638
rect 5005 -654 5215 -645
rect 5005 -688 5165 -654
rect 5199 -688 5215 -654
rect 5005 -704 5215 -688
rect 4767 -738 4833 -722
rect 4767 -772 4783 -738
rect 4817 -772 4833 -738
rect 4767 -788 4833 -772
rect 4885 -737 4951 -722
rect 4885 -771 4901 -737
rect 4935 -771 4951 -737
rect 4885 -787 4951 -771
rect 4769 -810 4829 -788
rect 4887 -810 4947 -787
rect 5005 -810 5065 -704
rect 5529 -706 5589 4
rect 6299 -130 6359 149
rect 7012 147 7555 198
rect 7597 191 7673 198
rect 7731 191 7791 217
rect 8243 200 8303 217
rect 8361 200 8421 217
rect 8479 200 8539 217
rect 8727 200 8787 217
rect 7597 147 7672 191
rect 8243 149 8787 200
rect 8845 191 8905 217
rect 8963 191 9023 217
rect 9081 198 9141 217
rect 9199 198 9259 217
rect 9317 198 9377 217
rect 9564 198 9624 217
rect 9682 198 9742 217
rect 7597 60 7657 147
rect 7529 50 7657 60
rect 7529 16 7545 50
rect 7579 16 7657 50
rect 6601 -53 6897 7
rect 6601 -76 6661 -53
rect 6719 -76 6779 -53
rect 6837 -76 6897 -53
rect 6955 -52 7251 8
rect 7529 6 7657 16
rect 6955 -76 7015 -52
rect 7073 -76 7133 -52
rect 7191 -76 7251 -52
rect 6135 -144 6359 -130
rect 6135 -178 6151 -144
rect 6185 -178 6359 -144
rect 6135 -190 6359 -178
rect 5439 -722 5589 -706
rect 5439 -756 5455 -722
rect 5489 -756 5589 -722
rect 5439 -772 5589 -756
rect 5529 -810 5589 -772
rect 6299 -703 6359 -190
rect 6601 -502 6661 -476
rect 6569 -643 6636 -636
rect 6719 -643 6779 -476
rect 6837 -502 6897 -476
rect 6955 -502 7015 -476
rect 6569 -652 6779 -643
rect 6569 -686 6585 -652
rect 6619 -686 6779 -652
rect 6569 -702 6779 -686
rect 6299 -719 6450 -703
rect 6299 -753 6400 -719
rect 6434 -753 6450 -719
rect 6299 -769 6450 -753
rect 6299 -808 6359 -769
rect 6719 -808 6779 -702
rect 7073 -643 7133 -476
rect 7191 -502 7251 -476
rect 7216 -643 7283 -636
rect 7073 -652 7283 -643
rect 7073 -686 7233 -652
rect 7267 -686 7283 -652
rect 7073 -702 7283 -686
rect 6835 -736 6901 -720
rect 6835 -770 6851 -736
rect 6885 -770 6901 -736
rect 6835 -786 6901 -770
rect 6953 -735 7019 -720
rect 6953 -769 6969 -735
rect 7003 -769 7019 -735
rect 6953 -785 7019 -769
rect 6837 -808 6897 -786
rect 6955 -808 7015 -785
rect 7073 -808 7133 -702
rect 7597 -704 7657 6
rect 8368 -130 8428 149
rect 9081 147 9624 198
rect 9666 191 9742 198
rect 9800 191 9860 217
rect 10311 202 10371 219
rect 10429 202 10489 219
rect 10547 202 10607 219
rect 10795 202 10855 219
rect 9666 147 9741 191
rect 10311 151 10855 202
rect 10913 193 10973 219
rect 11031 193 11091 219
rect 11149 200 11209 219
rect 11267 200 11327 219
rect 11385 200 11445 219
rect 11632 200 11692 219
rect 11750 200 11810 219
rect 9666 60 9726 147
rect 9598 50 9726 60
rect 9598 16 9614 50
rect 9648 16 9726 50
rect 8670 -53 8966 7
rect 8670 -76 8730 -53
rect 8788 -76 8848 -53
rect 8906 -76 8966 -53
rect 9024 -52 9320 8
rect 9598 6 9726 16
rect 9024 -76 9084 -52
rect 9142 -76 9202 -52
rect 9260 -76 9320 -52
rect 8204 -144 8428 -130
rect 8204 -178 8220 -144
rect 8254 -178 8428 -144
rect 8204 -190 8428 -178
rect 7507 -720 7657 -704
rect 7507 -754 7523 -720
rect 7557 -754 7657 -720
rect 7507 -770 7657 -754
rect 7597 -808 7657 -770
rect 8368 -703 8428 -190
rect 8670 -502 8730 -476
rect 8638 -643 8705 -636
rect 8788 -643 8848 -476
rect 8906 -502 8966 -476
rect 9024 -502 9084 -476
rect 8638 -652 8848 -643
rect 8638 -686 8654 -652
rect 8688 -686 8848 -652
rect 8638 -702 8848 -686
rect 8368 -719 8519 -703
rect 8368 -753 8469 -719
rect 8503 -753 8519 -719
rect 8368 -769 8519 -753
rect 8368 -808 8428 -769
rect 8788 -808 8848 -702
rect 9142 -643 9202 -476
rect 9260 -502 9320 -476
rect 9285 -643 9352 -636
rect 9142 -652 9352 -643
rect 9142 -686 9302 -652
rect 9336 -686 9352 -652
rect 9142 -702 9352 -686
rect 8904 -736 8970 -720
rect 8904 -770 8920 -736
rect 8954 -770 8970 -736
rect 8904 -786 8970 -770
rect 9022 -735 9088 -720
rect 9022 -769 9038 -735
rect 9072 -769 9088 -735
rect 9022 -785 9088 -769
rect 8906 -808 8966 -786
rect 9024 -808 9084 -785
rect 9142 -808 9202 -702
rect 9666 -704 9726 6
rect 10436 -128 10496 151
rect 11149 149 11692 200
rect 11734 193 11810 200
rect 11868 193 11928 219
rect 13701 434 13997 485
rect 13701 417 13761 434
rect 13819 417 13879 434
rect 13937 417 13997 434
rect 14448 419 14508 445
rect 14566 419 14626 445
rect 14684 419 14744 445
rect 15769 436 16065 487
rect 15769 419 15829 436
rect 15887 419 15947 436
rect 16005 419 16065 436
rect 12380 200 12440 217
rect 12498 200 12558 217
rect 12616 200 12676 217
rect 12864 200 12924 217
rect 11734 149 11809 193
rect 12380 149 12924 200
rect 12982 191 13042 217
rect 13100 191 13160 217
rect 13218 198 13278 217
rect 13336 198 13396 217
rect 13454 198 13514 217
rect 13701 198 13761 217
rect 13819 198 13879 217
rect 11734 62 11794 149
rect 11666 52 11794 62
rect 11666 18 11682 52
rect 11716 18 11794 52
rect 10738 -51 11034 9
rect 10738 -74 10798 -51
rect 10856 -74 10916 -51
rect 10974 -74 11034 -51
rect 11092 -50 11388 10
rect 11666 8 11794 18
rect 11092 -74 11152 -50
rect 11210 -74 11270 -50
rect 11328 -74 11388 -50
rect 10272 -142 10496 -128
rect 10272 -176 10288 -142
rect 10322 -176 10496 -142
rect 10272 -188 10496 -176
rect 9576 -720 9726 -704
rect 9576 -754 9592 -720
rect 9626 -754 9726 -720
rect 9576 -770 9726 -754
rect 9666 -808 9726 -770
rect 10436 -701 10496 -188
rect 10738 -500 10798 -474
rect 10706 -641 10773 -634
rect 10856 -641 10916 -474
rect 10974 -500 11034 -474
rect 11092 -500 11152 -474
rect 10706 -650 10916 -641
rect 10706 -684 10722 -650
rect 10756 -684 10916 -650
rect 10706 -700 10916 -684
rect 10436 -717 10587 -701
rect 10436 -751 10537 -717
rect 10571 -751 10587 -717
rect 10436 -767 10587 -751
rect 10436 -806 10496 -767
rect 10856 -806 10916 -700
rect 11210 -641 11270 -474
rect 11328 -500 11388 -474
rect 11353 -641 11420 -634
rect 11210 -650 11420 -641
rect 11210 -684 11370 -650
rect 11404 -684 11420 -650
rect 11210 -700 11420 -684
rect 10972 -734 11038 -718
rect 10972 -768 10988 -734
rect 11022 -768 11038 -734
rect 10972 -784 11038 -768
rect 11090 -733 11156 -718
rect 11090 -767 11106 -733
rect 11140 -767 11156 -733
rect 11090 -783 11156 -767
rect 10974 -806 11034 -784
rect 11092 -806 11152 -783
rect 11210 -806 11270 -700
rect 11734 -702 11794 8
rect 12505 -130 12565 149
rect 13218 147 13761 198
rect 13803 191 13879 198
rect 13937 191 13997 217
rect 14448 202 14508 219
rect 14566 202 14626 219
rect 14684 202 14744 219
rect 14932 202 14992 219
rect 13803 147 13878 191
rect 14448 151 14992 202
rect 15050 193 15110 219
rect 15168 193 15228 219
rect 15286 200 15346 219
rect 15404 200 15464 219
rect 15522 200 15582 219
rect 15769 200 15829 219
rect 15887 200 15947 219
rect 13803 60 13863 147
rect 13735 50 13863 60
rect 13735 16 13751 50
rect 13785 16 13863 50
rect 12807 -53 13103 7
rect 12807 -76 12867 -53
rect 12925 -76 12985 -53
rect 13043 -76 13103 -53
rect 13161 -52 13457 8
rect 13735 6 13863 16
rect 13161 -76 13221 -52
rect 13279 -76 13339 -52
rect 13397 -76 13457 -52
rect 12341 -144 12565 -130
rect 12341 -178 12357 -144
rect 12391 -178 12565 -144
rect 12341 -190 12565 -178
rect 11644 -718 11794 -702
rect 11644 -752 11660 -718
rect 11694 -752 11794 -718
rect 11644 -768 11794 -752
rect 11734 -806 11794 -768
rect 12505 -703 12565 -190
rect 12807 -502 12867 -476
rect 12775 -643 12842 -636
rect 12925 -643 12985 -476
rect 13043 -502 13103 -476
rect 13161 -502 13221 -476
rect 12775 -652 12985 -643
rect 12775 -686 12791 -652
rect 12825 -686 12985 -652
rect 12775 -702 12985 -686
rect 12505 -719 12656 -703
rect 12505 -753 12606 -719
rect 12640 -753 12656 -719
rect 12505 -769 12656 -753
rect 3460 -1034 3520 -1008
rect 4231 -1036 4291 -1010
rect 514 -1236 574 -1210
rect 632 -1236 692 -1210
rect 750 -1236 810 -1210
rect 868 -1236 928 -1210
rect 2582 -1234 2642 -1208
rect 2700 -1234 2760 -1208
rect 2818 -1234 2878 -1208
rect 2936 -1234 2996 -1208
rect 5529 -1036 5589 -1010
rect 6299 -1034 6359 -1008
rect 7597 -1034 7657 -1008
rect 8368 -1034 8428 -1008
rect 9666 -1034 9726 -1008
rect 10436 -1032 10496 -1006
rect 12505 -808 12565 -769
rect 12925 -808 12985 -702
rect 13279 -643 13339 -476
rect 13397 -502 13457 -476
rect 13422 -643 13489 -636
rect 13279 -652 13489 -643
rect 13279 -686 13439 -652
rect 13473 -686 13489 -652
rect 13279 -702 13489 -686
rect 13041 -736 13107 -720
rect 13041 -770 13057 -736
rect 13091 -770 13107 -736
rect 13041 -786 13107 -770
rect 13159 -735 13225 -720
rect 13159 -769 13175 -735
rect 13209 -769 13225 -735
rect 13159 -785 13225 -769
rect 13043 -808 13103 -786
rect 13161 -808 13221 -785
rect 13279 -808 13339 -702
rect 13803 -704 13863 6
rect 14573 -128 14633 151
rect 15286 149 15829 200
rect 15871 193 15947 200
rect 16005 193 16065 219
rect 15871 149 15946 193
rect 15871 62 15931 149
rect 15803 52 15931 62
rect 15803 18 15819 52
rect 15853 18 15931 52
rect 14875 -51 15171 9
rect 14875 -74 14935 -51
rect 14993 -74 15053 -51
rect 15111 -74 15171 -51
rect 15229 -50 15525 10
rect 15803 8 15931 18
rect 15229 -74 15289 -50
rect 15347 -74 15407 -50
rect 15465 -74 15525 -50
rect 14409 -142 14633 -128
rect 14409 -176 14425 -142
rect 14459 -176 14633 -142
rect 14409 -188 14633 -176
rect 13713 -720 13863 -704
rect 13713 -754 13729 -720
rect 13763 -754 13863 -720
rect 13713 -770 13863 -754
rect 13803 -808 13863 -770
rect 14573 -701 14633 -188
rect 14875 -500 14935 -474
rect 14843 -641 14910 -634
rect 14993 -641 15053 -474
rect 15111 -500 15171 -474
rect 15229 -500 15289 -474
rect 14843 -650 15053 -641
rect 14843 -684 14859 -650
rect 14893 -684 15053 -650
rect 14843 -700 15053 -684
rect 14573 -717 14724 -701
rect 14573 -751 14674 -717
rect 14708 -751 14724 -717
rect 14573 -767 14724 -751
rect 14573 -806 14633 -767
rect 14993 -806 15053 -700
rect 15347 -641 15407 -474
rect 15465 -500 15525 -474
rect 15490 -641 15557 -634
rect 15347 -650 15557 -641
rect 15347 -684 15507 -650
rect 15541 -684 15557 -650
rect 15347 -700 15557 -684
rect 15109 -734 15175 -718
rect 15109 -768 15125 -734
rect 15159 -768 15175 -734
rect 15109 -784 15175 -768
rect 15227 -733 15293 -718
rect 15227 -767 15243 -733
rect 15277 -767 15293 -733
rect 15227 -783 15293 -767
rect 15111 -806 15171 -784
rect 15229 -806 15289 -783
rect 15347 -806 15407 -700
rect 15871 -702 15931 8
rect 15781 -718 15931 -702
rect 15781 -752 15797 -718
rect 15831 -752 15931 -718
rect 15781 -768 15931 -752
rect 15871 -806 15931 -768
rect 11734 -1032 11794 -1006
rect 12505 -1034 12565 -1008
rect 4651 -1236 4711 -1210
rect 4769 -1236 4829 -1210
rect 4887 -1236 4947 -1210
rect 5005 -1236 5065 -1210
rect 6719 -1234 6779 -1208
rect 6837 -1234 6897 -1208
rect 6955 -1234 7015 -1208
rect 7073 -1234 7133 -1208
rect 8788 -1234 8848 -1208
rect 8906 -1234 8966 -1208
rect 9024 -1234 9084 -1208
rect 9142 -1234 9202 -1208
rect 10856 -1232 10916 -1206
rect 10974 -1232 11034 -1206
rect 11092 -1232 11152 -1206
rect 11210 -1232 11270 -1206
rect 13803 -1034 13863 -1008
rect 14573 -1032 14633 -1006
rect 15871 -1032 15931 -1006
rect 12925 -1234 12985 -1208
rect 13043 -1234 13103 -1208
rect 13161 -1234 13221 -1208
rect 13279 -1234 13339 -1208
rect 14993 -1232 15053 -1206
rect 15111 -1232 15171 -1206
rect 15229 -1232 15289 -1206
rect 15347 -1232 15407 -1206
<< polycont >>
rect 1340 14 1374 48
rect -54 -180 -20 -146
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1028 -688 1062 -654
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 3408 16 3442 50
rect 2014 -178 2048 -144
rect 1318 -756 1352 -722
rect 2448 -686 2482 -652
rect 2263 -753 2297 -719
rect 3096 -686 3130 -652
rect 2714 -770 2748 -736
rect 2832 -769 2866 -735
rect 5477 14 5511 48
rect 4083 -180 4117 -146
rect 3386 -754 3420 -720
rect 4517 -688 4551 -654
rect 4332 -755 4366 -721
rect 5165 -688 5199 -654
rect 4783 -772 4817 -738
rect 4901 -771 4935 -737
rect 7545 16 7579 50
rect 6151 -178 6185 -144
rect 5455 -756 5489 -722
rect 6585 -686 6619 -652
rect 6400 -753 6434 -719
rect 7233 -686 7267 -652
rect 6851 -770 6885 -736
rect 6969 -769 7003 -735
rect 9614 16 9648 50
rect 8220 -178 8254 -144
rect 7523 -754 7557 -720
rect 8654 -686 8688 -652
rect 8469 -753 8503 -719
rect 9302 -686 9336 -652
rect 8920 -770 8954 -736
rect 9038 -769 9072 -735
rect 11682 18 11716 52
rect 10288 -176 10322 -142
rect 9592 -754 9626 -720
rect 10722 -684 10756 -650
rect 10537 -751 10571 -717
rect 11370 -684 11404 -650
rect 10988 -768 11022 -734
rect 11106 -767 11140 -733
rect 13751 16 13785 50
rect 12357 -178 12391 -144
rect 11660 -752 11694 -718
rect 12791 -686 12825 -652
rect 12606 -753 12640 -719
rect 13439 -686 13473 -652
rect 13057 -770 13091 -736
rect 13175 -769 13209 -735
rect 15819 18 15853 52
rect 14425 -176 14459 -142
rect 13729 -754 13763 -720
rect 14859 -684 14893 -650
rect 14674 -751 14708 -717
rect 15507 -684 15541 -650
rect 15125 -768 15159 -734
rect 15243 -767 15277 -733
rect 15797 -752 15831 -718
<< locali >>
rect 674 874 876 894
rect 674 830 708 874
rect 830 830 876 874
rect 674 820 760 830
rect 798 820 876 830
rect 674 802 876 820
rect 2742 876 2944 896
rect 2742 832 2776 876
rect 2898 832 2944 876
rect 2742 822 2828 832
rect 2866 822 2944 832
rect 2742 804 2944 822
rect 4811 874 5013 894
rect 4811 830 4845 874
rect 4967 830 5013 874
rect 4811 820 4897 830
rect 4935 820 5013 830
rect 4811 802 5013 820
rect 6879 876 7081 896
rect 6879 832 6913 876
rect 7035 832 7081 876
rect 6879 822 6965 832
rect 7003 822 7081 832
rect 6879 804 7081 822
rect 8948 876 9150 896
rect 8948 832 8982 876
rect 9104 832 9150 876
rect 8948 822 9034 832
rect 9072 822 9150 832
rect 8948 804 9150 822
rect 11016 878 11218 898
rect 11016 834 11050 878
rect 11172 834 11218 878
rect 11016 824 11102 834
rect 11140 824 11218 834
rect 11016 806 11218 824
rect 13085 876 13287 896
rect 13085 832 13119 876
rect 13241 832 13287 876
rect 13085 822 13171 832
rect 13209 822 13287 832
rect 13085 804 13287 822
rect 15153 878 15355 898
rect 15153 834 15187 878
rect 15309 834 15355 878
rect 15153 824 15239 834
rect 15277 824 15355 834
rect 15153 806 15355 824
rect 761 656 1031 691
rect 407 603 441 619
rect -77 457 193 492
rect -77 403 -43 457
rect -77 211 -43 227
rect 41 403 75 419
rect 41 211 75 227
rect 159 403 193 457
rect 159 211 193 227
rect 277 403 311 419
rect 277 211 311 227
rect 407 211 441 227
rect 525 603 559 619
rect 525 211 559 227
rect 643 603 677 619
rect 643 211 677 227
rect 761 603 795 656
rect 761 211 795 227
rect 879 603 913 619
rect 879 211 913 227
rect 997 603 1031 656
rect 2829 658 3099 693
rect 997 211 1031 227
rect 1115 603 1149 619
rect 2475 605 2509 621
rect 1991 459 2261 494
rect 1115 211 1149 227
rect 1244 403 1278 419
rect 1244 211 1278 227
rect 1362 403 1396 419
rect 1362 211 1396 227
rect 1480 403 1514 419
rect 1480 211 1514 227
rect 1598 403 1632 419
rect 1598 211 1632 227
rect 1991 405 2025 459
rect 1991 213 2025 229
rect 2109 405 2143 421
rect 2109 213 2143 229
rect 2227 405 2261 459
rect 2227 213 2261 229
rect 2345 405 2379 421
rect 2345 213 2379 229
rect 2475 213 2509 229
rect 2593 605 2627 621
rect 2593 213 2627 229
rect 2711 605 2745 621
rect 2711 213 2745 229
rect 2829 605 2863 658
rect 2829 213 2863 229
rect 2947 605 2981 621
rect 2947 213 2981 229
rect 3065 605 3099 658
rect 4898 656 5168 691
rect 3065 213 3099 229
rect 3183 605 3217 621
rect 4544 603 4578 619
rect 4060 457 4330 492
rect 3183 213 3217 229
rect 3312 405 3346 421
rect 3312 213 3346 229
rect 3430 405 3464 421
rect 3430 213 3464 229
rect 3548 405 3582 421
rect 3548 213 3582 229
rect 3666 405 3700 421
rect 3666 213 3700 229
rect 4060 403 4094 457
rect 4060 211 4094 227
rect 4178 403 4212 419
rect 4178 211 4212 227
rect 4296 403 4330 457
rect 4296 211 4330 227
rect 4414 403 4448 419
rect 4414 211 4448 227
rect 4544 211 4578 227
rect 4662 603 4696 619
rect 4662 211 4696 227
rect 4780 603 4814 619
rect 4780 211 4814 227
rect 4898 603 4932 656
rect 4898 211 4932 227
rect 5016 603 5050 619
rect 5016 211 5050 227
rect 5134 603 5168 656
rect 6966 658 7236 693
rect 5134 211 5168 227
rect 5252 603 5286 619
rect 6612 605 6646 621
rect 6128 459 6398 494
rect 5252 211 5286 227
rect 5381 403 5415 419
rect 5381 211 5415 227
rect 5499 403 5533 419
rect 5499 211 5533 227
rect 5617 403 5651 419
rect 5617 211 5651 227
rect 5735 403 5769 419
rect 5735 211 5769 227
rect 6128 405 6162 459
rect 6128 213 6162 229
rect 6246 405 6280 421
rect 6246 213 6280 229
rect 6364 405 6398 459
rect 6364 213 6398 229
rect 6482 405 6516 421
rect 6482 213 6516 229
rect 6612 213 6646 229
rect 6730 605 6764 621
rect 6730 213 6764 229
rect 6848 605 6882 621
rect 6848 213 6882 229
rect 6966 605 7000 658
rect 6966 213 7000 229
rect 7084 605 7118 621
rect 7084 213 7118 229
rect 7202 605 7236 658
rect 9035 658 9305 693
rect 7202 213 7236 229
rect 7320 605 7354 621
rect 8681 605 8715 621
rect 8197 459 8467 494
rect 7320 213 7354 229
rect 7449 405 7483 421
rect 7449 213 7483 229
rect 7567 405 7601 421
rect 7567 213 7601 229
rect 7685 405 7719 421
rect 7685 213 7719 229
rect 7803 405 7837 421
rect 7803 213 7837 229
rect 8197 405 8231 459
rect 8197 213 8231 229
rect 8315 405 8349 421
rect 8315 213 8349 229
rect 8433 405 8467 459
rect 8433 213 8467 229
rect 8551 405 8585 421
rect 8551 213 8585 229
rect 8681 213 8715 229
rect 8799 605 8833 621
rect 8799 213 8833 229
rect 8917 605 8951 621
rect 8917 213 8951 229
rect 9035 605 9069 658
rect 9035 213 9069 229
rect 9153 605 9187 621
rect 9153 213 9187 229
rect 9271 605 9305 658
rect 11103 660 11373 695
rect 9271 213 9305 229
rect 9389 605 9423 621
rect 10749 607 10783 623
rect 10265 461 10535 496
rect 9389 213 9423 229
rect 9518 405 9552 421
rect 9518 213 9552 229
rect 9636 405 9670 421
rect 9636 213 9670 229
rect 9754 405 9788 421
rect 9754 213 9788 229
rect 9872 405 9906 421
rect 9872 213 9906 229
rect 10265 407 10299 461
rect 10265 215 10299 231
rect 10383 407 10417 423
rect 10383 215 10417 231
rect 10501 407 10535 461
rect 10501 215 10535 231
rect 10619 407 10653 423
rect 10619 215 10653 231
rect 10749 215 10783 231
rect 10867 607 10901 623
rect 10867 215 10901 231
rect 10985 607 11019 623
rect 10985 215 11019 231
rect 11103 607 11137 660
rect 11103 215 11137 231
rect 11221 607 11255 623
rect 11221 215 11255 231
rect 11339 607 11373 660
rect 13172 658 13442 693
rect 11339 215 11373 231
rect 11457 607 11491 623
rect 12818 605 12852 621
rect 12334 459 12604 494
rect 11457 215 11491 231
rect 11586 407 11620 423
rect 11586 215 11620 231
rect 11704 407 11738 423
rect 11704 215 11738 231
rect 11822 407 11856 423
rect 11822 215 11856 231
rect 11940 407 11974 423
rect 11940 215 11974 231
rect 12334 405 12368 459
rect 12334 213 12368 229
rect 12452 405 12486 421
rect 12452 213 12486 229
rect 12570 405 12604 459
rect 12570 213 12604 229
rect 12688 405 12722 421
rect 12688 213 12722 229
rect 12818 213 12852 229
rect 12936 605 12970 621
rect 12936 213 12970 229
rect 13054 605 13088 621
rect 13054 213 13088 229
rect 13172 605 13206 658
rect 13172 213 13206 229
rect 13290 605 13324 621
rect 13290 213 13324 229
rect 13408 605 13442 658
rect 15240 660 15510 695
rect 13408 213 13442 229
rect 13526 605 13560 621
rect 14886 607 14920 623
rect 14402 461 14672 496
rect 13526 213 13560 229
rect 13655 405 13689 421
rect 13655 213 13689 229
rect 13773 405 13807 421
rect 13773 213 13807 229
rect 13891 405 13925 421
rect 13891 213 13925 229
rect 14009 405 14043 421
rect 14009 213 14043 229
rect 14402 407 14436 461
rect 14402 215 14436 231
rect 14520 407 14554 423
rect 14520 215 14554 231
rect 14638 407 14672 461
rect 14638 215 14672 231
rect 14756 407 14790 423
rect 14756 215 14790 231
rect 14886 215 14920 231
rect 15004 607 15038 623
rect 15004 215 15038 231
rect 15122 607 15156 623
rect 15122 215 15156 231
rect 15240 607 15274 660
rect 15240 215 15274 231
rect 15358 607 15392 623
rect 15358 215 15392 231
rect 15476 607 15510 660
rect 15476 215 15510 231
rect 15594 607 15628 623
rect 15594 215 15628 231
rect 15723 407 15757 423
rect 15723 215 15757 231
rect 15841 407 15875 423
rect 15841 215 15875 231
rect 15959 407 15993 423
rect 15959 215 15993 231
rect 16077 407 16111 423
rect 16077 215 16111 231
rect 1324 14 1330 48
rect 1384 14 1390 48
rect 3392 16 3398 50
rect 3452 16 3458 50
rect 5461 14 5467 48
rect 5521 14 5527 48
rect 7529 16 7535 50
rect 7589 16 7595 50
rect 9598 16 9604 50
rect 9658 16 9664 50
rect 11666 18 11672 52
rect 11726 18 11732 52
rect 13735 16 13741 50
rect 13795 16 13801 50
rect 15803 18 15809 52
rect 15863 18 15869 52
rect 350 -90 384 -74
rect 468 -90 502 -74
rect 350 -482 384 -466
rect 467 -466 468 -419
rect 586 -90 620 -74
rect 502 -466 503 -419
rect 467 -524 503 -466
rect 704 -90 738 -74
rect 586 -482 620 -466
rect 702 -466 704 -419
rect 702 -524 738 -466
rect 822 -90 856 -74
rect 822 -482 856 -466
rect 940 -90 974 -74
rect 1058 -90 1092 -74
rect 974 -466 976 -420
rect 940 -524 976 -466
rect 2418 -88 2452 -72
rect 1058 -482 1092 -466
rect 2536 -88 2570 -72
rect 2418 -480 2452 -464
rect 2535 -464 2536 -417
rect 2654 -88 2688 -72
rect 2570 -464 2571 -417
rect 467 -564 1562 -524
rect 486 -565 1562 -564
rect 364 -654 431 -638
rect 364 -688 380 -654
rect 414 -688 431 -654
rect 364 -704 431 -688
rect 195 -721 229 -705
rect 195 -771 229 -755
rect 541 -806 575 -565
rect 2535 -522 2571 -464
rect 2772 -88 2806 -72
rect 2654 -480 2688 -464
rect 2770 -464 2772 -417
rect 2770 -522 2806 -464
rect 2890 -88 2924 -72
rect 2890 -480 2924 -464
rect 3008 -88 3042 -72
rect 3126 -88 3160 -72
rect 3042 -464 3044 -418
rect 3008 -522 3044 -464
rect 4487 -90 4521 -74
rect 3126 -480 3160 -464
rect 4605 -90 4639 -74
rect 4487 -482 4521 -466
rect 4604 -466 4605 -419
rect 4723 -90 4757 -74
rect 4639 -466 4640 -419
rect 2535 -562 3630 -522
rect 2554 -563 3630 -562
rect 1011 -654 1078 -638
rect 1011 -688 1028 -654
rect 1062 -688 1078 -654
rect 1011 -704 1078 -688
rect 2432 -652 2499 -636
rect 2432 -686 2448 -652
rect 2482 -686 2499 -652
rect 2432 -702 2499 -686
rect 1318 -722 1352 -706
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 1318 -772 1352 -756
rect 2263 -719 2297 -703
rect 2263 -769 2297 -753
rect 2609 -804 2643 -563
rect 4604 -524 4640 -466
rect 4841 -90 4875 -74
rect 4723 -482 4757 -466
rect 4839 -466 4841 -419
rect 4839 -524 4875 -466
rect 4959 -90 4993 -74
rect 4959 -482 4993 -466
rect 5077 -90 5111 -74
rect 5195 -90 5229 -74
rect 5111 -466 5113 -420
rect 5077 -524 5113 -466
rect 6555 -88 6589 -72
rect 5195 -482 5229 -466
rect 6673 -88 6707 -72
rect 6555 -480 6589 -464
rect 6672 -464 6673 -417
rect 6791 -88 6825 -72
rect 6707 -464 6708 -417
rect 4604 -564 5699 -524
rect 4623 -565 5699 -564
rect 3079 -652 3146 -636
rect 3079 -686 3096 -652
rect 3130 -686 3146 -652
rect 3079 -702 3146 -686
rect 4501 -654 4568 -638
rect 4501 -688 4517 -654
rect 4551 -688 4568 -654
rect 4501 -704 4568 -688
rect 3386 -720 3420 -704
rect 2698 -770 2714 -736
rect 2748 -770 2764 -736
rect 2816 -769 2832 -735
rect 2866 -769 2882 -735
rect 3386 -770 3420 -754
rect 4332 -721 4366 -705
rect 4332 -771 4366 -755
rect 48 -822 82 -806
rect 48 -1014 82 -998
rect 166 -822 200 -806
rect 166 -1014 200 -998
rect 468 -822 502 -806
rect 541 -822 620 -806
rect 541 -852 586 -822
rect 468 -1265 503 -1198
rect 586 -1214 620 -1198
rect 704 -822 738 -806
rect 704 -1214 738 -1198
rect 822 -822 856 -806
rect 940 -822 974 -806
rect 1346 -822 1380 -806
rect 1346 -1014 1380 -998
rect 1464 -822 1498 -806
rect 1464 -1014 1498 -998
rect 2116 -820 2150 -804
rect 2116 -1012 2150 -996
rect 2234 -820 2268 -804
rect 2234 -1012 2268 -996
rect 2536 -820 2570 -804
rect 822 -1214 856 -1198
rect 939 -1265 974 -1198
rect 468 -1300 974 -1265
rect 2609 -820 2688 -804
rect 2609 -850 2654 -820
rect 2536 -1263 2571 -1196
rect 2654 -1212 2688 -1196
rect 2772 -820 2806 -804
rect 2772 -1212 2806 -1196
rect 2890 -820 2924 -804
rect 3008 -820 3042 -804
rect 3414 -820 3448 -804
rect 3414 -1012 3448 -996
rect 3532 -820 3566 -804
rect 4678 -806 4712 -565
rect 6672 -522 6708 -464
rect 6909 -88 6943 -72
rect 6791 -480 6825 -464
rect 6907 -464 6909 -417
rect 6907 -522 6943 -464
rect 7027 -88 7061 -72
rect 7027 -480 7061 -464
rect 7145 -88 7179 -72
rect 7263 -88 7297 -72
rect 7179 -464 7181 -418
rect 7145 -522 7181 -464
rect 8624 -88 8658 -72
rect 7263 -480 7297 -464
rect 8742 -88 8776 -72
rect 8624 -480 8658 -464
rect 8741 -464 8742 -417
rect 8860 -88 8894 -72
rect 8776 -464 8777 -417
rect 6672 -562 7767 -522
rect 6691 -563 7767 -562
rect 5148 -654 5215 -638
rect 5148 -688 5165 -654
rect 5199 -688 5215 -654
rect 5148 -704 5215 -688
rect 6569 -652 6636 -636
rect 6569 -686 6585 -652
rect 6619 -686 6636 -652
rect 6569 -702 6636 -686
rect 5455 -722 5489 -706
rect 4767 -772 4783 -738
rect 4817 -772 4833 -738
rect 4885 -771 4901 -737
rect 4935 -771 4951 -737
rect 5455 -772 5489 -756
rect 6400 -719 6434 -703
rect 6400 -769 6434 -753
rect 6746 -804 6780 -563
rect 8741 -522 8777 -464
rect 8978 -88 9012 -72
rect 8860 -480 8894 -464
rect 8976 -464 8978 -417
rect 8976 -522 9012 -464
rect 9096 -88 9130 -72
rect 9096 -480 9130 -464
rect 9214 -88 9248 -72
rect 9332 -88 9366 -72
rect 9248 -464 9250 -418
rect 9214 -522 9250 -464
rect 10692 -86 10726 -70
rect 9332 -480 9366 -464
rect 10810 -86 10844 -70
rect 10692 -478 10726 -462
rect 10809 -462 10810 -415
rect 10928 -86 10962 -70
rect 10844 -462 10845 -415
rect 8741 -562 9836 -522
rect 8760 -563 9836 -562
rect 7216 -652 7283 -636
rect 7216 -686 7233 -652
rect 7267 -686 7283 -652
rect 7216 -702 7283 -686
rect 8638 -652 8705 -636
rect 8638 -686 8654 -652
rect 8688 -686 8705 -652
rect 8638 -702 8705 -686
rect 7523 -720 7557 -704
rect 6835 -770 6851 -736
rect 6885 -770 6901 -736
rect 6953 -769 6969 -735
rect 7003 -769 7019 -735
rect 7523 -770 7557 -754
rect 8469 -719 8503 -703
rect 8469 -769 8503 -753
rect 8815 -804 8849 -563
rect 10809 -520 10845 -462
rect 11046 -86 11080 -70
rect 10928 -478 10962 -462
rect 11044 -462 11046 -415
rect 11044 -520 11080 -462
rect 11164 -86 11198 -70
rect 11164 -478 11198 -462
rect 11282 -86 11316 -70
rect 11400 -86 11434 -70
rect 11316 -462 11318 -416
rect 11282 -520 11318 -462
rect 12761 -88 12795 -72
rect 11400 -478 11434 -462
rect 12879 -88 12913 -72
rect 12761 -480 12795 -464
rect 12878 -464 12879 -417
rect 12997 -88 13031 -72
rect 12913 -464 12914 -417
rect 10809 -560 11904 -520
rect 10828 -561 11904 -560
rect 9285 -652 9352 -636
rect 9285 -686 9302 -652
rect 9336 -686 9352 -652
rect 9285 -702 9352 -686
rect 10706 -650 10773 -634
rect 10706 -684 10722 -650
rect 10756 -684 10773 -650
rect 10706 -700 10773 -684
rect 9592 -720 9626 -704
rect 8904 -770 8920 -736
rect 8954 -770 8970 -736
rect 9022 -769 9038 -735
rect 9072 -769 9088 -735
rect 9592 -770 9626 -754
rect 10537 -717 10571 -701
rect 10537 -767 10571 -751
rect 10883 -802 10917 -561
rect 12878 -522 12914 -464
rect 13115 -88 13149 -72
rect 12997 -480 13031 -464
rect 13113 -464 13115 -417
rect 13113 -522 13149 -464
rect 13233 -88 13267 -72
rect 13233 -480 13267 -464
rect 13351 -88 13385 -72
rect 13469 -88 13503 -72
rect 13385 -464 13387 -418
rect 13351 -522 13387 -464
rect 14829 -86 14863 -70
rect 13469 -480 13503 -464
rect 14947 -86 14981 -70
rect 14829 -478 14863 -462
rect 14946 -462 14947 -415
rect 15065 -86 15099 -70
rect 14981 -462 14982 -415
rect 12878 -562 13973 -522
rect 12897 -563 13973 -562
rect 11353 -650 11420 -634
rect 11353 -684 11370 -650
rect 11404 -684 11420 -650
rect 11353 -700 11420 -684
rect 12775 -652 12842 -636
rect 12775 -686 12791 -652
rect 12825 -686 12842 -652
rect 12775 -702 12842 -686
rect 11660 -718 11694 -702
rect 10972 -768 10988 -734
rect 11022 -768 11038 -734
rect 11090 -767 11106 -733
rect 11140 -767 11156 -733
rect 11660 -768 11694 -752
rect 12606 -719 12640 -703
rect 12606 -769 12640 -753
rect 3532 -1012 3566 -996
rect 4185 -822 4219 -806
rect 4185 -1014 4219 -998
rect 4303 -822 4337 -806
rect 4303 -1014 4337 -998
rect 4605 -822 4639 -806
rect 2890 -1212 2924 -1196
rect 3007 -1263 3042 -1196
rect 2536 -1298 3042 -1263
rect 4678 -822 4757 -806
rect 4678 -852 4723 -822
rect 4605 -1265 4640 -1198
rect 4723 -1214 4757 -1198
rect 4841 -822 4875 -806
rect 4841 -1214 4875 -1198
rect 4959 -822 4993 -806
rect 5077 -822 5111 -806
rect 5483 -822 5517 -806
rect 5483 -1014 5517 -998
rect 5601 -822 5635 -806
rect 5601 -1014 5635 -998
rect 6253 -820 6287 -804
rect 6253 -1012 6287 -996
rect 6371 -820 6405 -804
rect 6371 -1012 6405 -996
rect 6673 -820 6707 -804
rect 4959 -1214 4993 -1198
rect 5076 -1265 5111 -1198
rect 4605 -1300 5111 -1265
rect 6746 -820 6825 -804
rect 6746 -850 6791 -820
rect 6673 -1263 6708 -1196
rect 6791 -1212 6825 -1196
rect 6909 -820 6943 -804
rect 6909 -1212 6943 -1196
rect 7027 -820 7061 -804
rect 7145 -820 7179 -804
rect 7551 -820 7585 -804
rect 7551 -1012 7585 -996
rect 7669 -820 7703 -804
rect 7669 -1012 7703 -996
rect 8322 -820 8356 -804
rect 8322 -1012 8356 -996
rect 8440 -820 8474 -804
rect 8440 -1012 8474 -996
rect 8742 -820 8776 -804
rect 7027 -1212 7061 -1196
rect 7144 -1263 7179 -1196
rect 6673 -1298 7179 -1263
rect 8815 -820 8894 -804
rect 8815 -850 8860 -820
rect 8742 -1263 8777 -1196
rect 8860 -1212 8894 -1196
rect 8978 -820 9012 -804
rect 8978 -1212 9012 -1196
rect 9096 -820 9130 -804
rect 9214 -820 9248 -804
rect 9620 -820 9654 -804
rect 9620 -1012 9654 -996
rect 9738 -820 9772 -804
rect 9738 -1012 9772 -996
rect 10390 -818 10424 -802
rect 10390 -1010 10424 -994
rect 10508 -818 10542 -802
rect 10508 -1010 10542 -994
rect 10810 -818 10844 -802
rect 9096 -1212 9130 -1196
rect 9213 -1263 9248 -1196
rect 8742 -1298 9248 -1263
rect 10883 -818 10962 -802
rect 10883 -848 10928 -818
rect 10810 -1261 10845 -1194
rect 10928 -1210 10962 -1194
rect 11046 -818 11080 -802
rect 11046 -1210 11080 -1194
rect 11164 -818 11198 -802
rect 11282 -818 11316 -802
rect 11688 -818 11722 -802
rect 11688 -1010 11722 -994
rect 11806 -818 11840 -802
rect 12952 -804 12986 -563
rect 14946 -520 14982 -462
rect 15183 -86 15217 -70
rect 15065 -478 15099 -462
rect 15181 -462 15183 -415
rect 15181 -520 15217 -462
rect 15301 -86 15335 -70
rect 15301 -478 15335 -462
rect 15419 -86 15453 -70
rect 15537 -86 15571 -70
rect 15453 -462 15455 -416
rect 15419 -520 15455 -462
rect 15537 -478 15571 -462
rect 14946 -560 16041 -520
rect 14965 -561 16041 -560
rect 13422 -652 13489 -636
rect 13422 -686 13439 -652
rect 13473 -686 13489 -652
rect 13422 -702 13489 -686
rect 14843 -650 14910 -634
rect 14843 -684 14859 -650
rect 14893 -684 14910 -650
rect 14843 -700 14910 -684
rect 13729 -720 13763 -704
rect 13041 -770 13057 -736
rect 13091 -770 13107 -736
rect 13159 -769 13175 -735
rect 13209 -769 13225 -735
rect 13729 -770 13763 -754
rect 14674 -717 14708 -701
rect 14674 -767 14708 -751
rect 15020 -802 15054 -561
rect 15490 -650 15557 -634
rect 15490 -684 15507 -650
rect 15541 -684 15557 -650
rect 15490 -700 15557 -684
rect 15797 -718 15831 -702
rect 15109 -768 15125 -734
rect 15159 -768 15175 -734
rect 15227 -767 15243 -733
rect 15277 -767 15293 -733
rect 15797 -768 15831 -752
rect 11806 -1010 11840 -994
rect 12459 -820 12493 -804
rect 12459 -1012 12493 -996
rect 12577 -820 12611 -804
rect 12577 -1012 12611 -996
rect 12879 -820 12913 -804
rect 11164 -1210 11198 -1194
rect 11281 -1261 11316 -1194
rect 10810 -1296 11316 -1261
rect 12952 -820 13031 -804
rect 12952 -850 12997 -820
rect 12879 -1263 12914 -1196
rect 12997 -1212 13031 -1196
rect 13115 -820 13149 -804
rect 13115 -1212 13149 -1196
rect 13233 -820 13267 -804
rect 13351 -820 13385 -804
rect 13757 -820 13791 -804
rect 13757 -1012 13791 -996
rect 13875 -820 13909 -804
rect 13875 -1012 13909 -996
rect 14527 -818 14561 -802
rect 14527 -1010 14561 -994
rect 14645 -818 14679 -802
rect 14645 -1010 14679 -994
rect 14947 -818 14981 -802
rect 13233 -1212 13267 -1196
rect 13350 -1263 13385 -1196
rect 12879 -1298 13385 -1263
rect 15020 -818 15099 -802
rect 15020 -848 15065 -818
rect 14947 -1261 14982 -1194
rect 15065 -1210 15099 -1194
rect 15183 -818 15217 -802
rect 15183 -1210 15217 -1194
rect 15301 -818 15335 -802
rect 15419 -818 15453 -802
rect 15825 -818 15859 -802
rect 15825 -1010 15859 -994
rect 15943 -818 15977 -802
rect 15943 -1010 15977 -994
rect 15301 -1210 15335 -1194
rect 15418 -1261 15453 -1194
rect 14947 -1296 15453 -1261
rect 642 -1386 698 -1370
rect 748 -1386 806 -1370
rect 642 -1442 658 -1386
rect 790 -1442 806 -1386
rect 642 -1458 806 -1442
rect 2710 -1384 2766 -1368
rect 2816 -1384 2874 -1368
rect 2710 -1440 2726 -1384
rect 2858 -1440 2874 -1384
rect 2710 -1456 2874 -1440
rect 4779 -1386 4835 -1370
rect 4885 -1386 4943 -1370
rect 4779 -1442 4795 -1386
rect 4927 -1442 4943 -1386
rect 4779 -1458 4943 -1442
rect 6847 -1384 6903 -1368
rect 6953 -1384 7011 -1368
rect 6847 -1440 6863 -1384
rect 6995 -1440 7011 -1384
rect 6847 -1456 7011 -1440
rect 8916 -1384 8972 -1368
rect 9022 -1384 9080 -1368
rect 8916 -1440 8932 -1384
rect 9064 -1440 9080 -1384
rect 8916 -1456 9080 -1440
rect 10984 -1382 11040 -1366
rect 11090 -1382 11148 -1366
rect 10984 -1438 11000 -1382
rect 11132 -1438 11148 -1382
rect 10984 -1454 11148 -1438
rect 13053 -1384 13109 -1368
rect 13159 -1384 13217 -1368
rect 13053 -1440 13069 -1384
rect 13201 -1440 13217 -1384
rect 13053 -1456 13217 -1440
rect 15121 -1382 15177 -1366
rect 15227 -1382 15285 -1366
rect 15121 -1438 15137 -1382
rect 15269 -1438 15285 -1382
rect 15121 -1454 15285 -1438
<< viali >>
rect 760 830 798 858
rect 760 820 798 830
rect 2828 832 2866 860
rect 2828 822 2866 832
rect 4897 830 4935 858
rect 4897 820 4935 830
rect 6965 832 7003 860
rect 6965 822 7003 832
rect 9034 832 9072 860
rect 9034 822 9072 832
rect 11102 834 11140 862
rect 11102 824 11140 834
rect 13171 832 13209 860
rect 13171 822 13209 832
rect 15239 834 15277 862
rect 15239 824 15277 834
rect -77 227 -43 403
rect 41 227 75 403
rect 159 227 193 403
rect 277 227 311 403
rect 407 227 441 603
rect 525 227 559 603
rect 643 227 677 603
rect 761 227 795 603
rect 879 227 913 603
rect 997 227 1031 603
rect 1115 227 1149 603
rect 1244 227 1278 403
rect 1362 227 1396 403
rect 1480 227 1514 403
rect 1598 227 1632 403
rect 1991 229 2025 405
rect 2109 229 2143 405
rect 2227 229 2261 405
rect 2345 229 2379 405
rect 2475 229 2509 605
rect 2593 229 2627 605
rect 2711 229 2745 605
rect 2829 229 2863 605
rect 2947 229 2981 605
rect 3065 229 3099 605
rect 3183 229 3217 605
rect 3312 229 3346 405
rect 3430 229 3464 405
rect 3548 229 3582 405
rect 3666 229 3700 405
rect 4060 227 4094 403
rect 4178 227 4212 403
rect 4296 227 4330 403
rect 4414 227 4448 403
rect 4544 227 4578 603
rect 4662 227 4696 603
rect 4780 227 4814 603
rect 4898 227 4932 603
rect 5016 227 5050 603
rect 5134 227 5168 603
rect 5252 227 5286 603
rect 5381 227 5415 403
rect 5499 227 5533 403
rect 5617 227 5651 403
rect 5735 227 5769 403
rect 6128 229 6162 405
rect 6246 229 6280 405
rect 6364 229 6398 405
rect 6482 229 6516 405
rect 6612 229 6646 605
rect 6730 229 6764 605
rect 6848 229 6882 605
rect 6966 229 7000 605
rect 7084 229 7118 605
rect 7202 229 7236 605
rect 7320 229 7354 605
rect 7449 229 7483 405
rect 7567 229 7601 405
rect 7685 229 7719 405
rect 7803 229 7837 405
rect 8197 229 8231 405
rect 8315 229 8349 405
rect 8433 229 8467 405
rect 8551 229 8585 405
rect 8681 229 8715 605
rect 8799 229 8833 605
rect 8917 229 8951 605
rect 9035 229 9069 605
rect 9153 229 9187 605
rect 9271 229 9305 605
rect 9389 229 9423 605
rect 9518 229 9552 405
rect 9636 229 9670 405
rect 9754 229 9788 405
rect 9872 229 9906 405
rect 10265 231 10299 407
rect 10383 231 10417 407
rect 10501 231 10535 407
rect 10619 231 10653 407
rect 10749 231 10783 607
rect 10867 231 10901 607
rect 10985 231 11019 607
rect 11103 231 11137 607
rect 11221 231 11255 607
rect 11339 231 11373 607
rect 11457 231 11491 607
rect 11586 231 11620 407
rect 11704 231 11738 407
rect 11822 231 11856 407
rect 11940 231 11974 407
rect 12334 229 12368 405
rect 12452 229 12486 405
rect 12570 229 12604 405
rect 12688 229 12722 405
rect 12818 229 12852 605
rect 12936 229 12970 605
rect 13054 229 13088 605
rect 13172 229 13206 605
rect 13290 229 13324 605
rect 13408 229 13442 605
rect 13526 229 13560 605
rect 13655 229 13689 405
rect 13773 229 13807 405
rect 13891 229 13925 405
rect 14009 229 14043 405
rect 14402 231 14436 407
rect 14520 231 14554 407
rect 14638 231 14672 407
rect 14756 231 14790 407
rect 14886 231 14920 607
rect 15004 231 15038 607
rect 15122 231 15156 607
rect 15240 231 15274 607
rect 15358 231 15392 607
rect 15476 231 15510 607
rect 15594 231 15628 607
rect 15723 231 15757 407
rect 15841 231 15875 407
rect 15959 231 15993 407
rect 16077 231 16111 407
rect 1330 48 1384 58
rect 3398 50 3452 60
rect 1330 14 1340 48
rect 1340 14 1374 48
rect 1374 14 1384 48
rect 3398 16 3408 50
rect 3408 16 3442 50
rect 3442 16 3452 50
rect 5467 48 5521 58
rect 7535 50 7589 60
rect 9604 50 9658 60
rect 11672 52 11726 62
rect 1330 4 1384 14
rect 3398 6 3452 16
rect 5467 14 5477 48
rect 5477 14 5511 48
rect 5511 14 5521 48
rect 7535 16 7545 50
rect 7545 16 7579 50
rect 7579 16 7589 50
rect 9604 16 9614 50
rect 9614 16 9648 50
rect 9648 16 9658 50
rect 11672 18 11682 52
rect 11682 18 11716 52
rect 11716 18 11726 52
rect 13741 50 13795 60
rect 15809 52 15863 62
rect 5467 4 5521 14
rect 7535 6 7589 16
rect 9604 6 9658 16
rect 11672 8 11726 18
rect 13741 16 13751 50
rect 13751 16 13785 50
rect 13785 16 13795 50
rect 15809 18 15819 52
rect 15819 18 15853 52
rect 15853 18 15863 52
rect 13741 6 13795 16
rect 15809 8 15863 18
rect -70 -146 -4 -132
rect -70 -180 -54 -146
rect -54 -180 -20 -146
rect -20 -180 -4 -146
rect -70 -192 -4 -180
rect 350 -466 384 -90
rect 468 -466 502 -90
rect 586 -466 620 -90
rect 704 -466 738 -90
rect 822 -466 856 -90
rect 940 -466 974 -90
rect 1058 -466 1092 -90
rect 1998 -144 2064 -130
rect 1998 -178 2014 -144
rect 2014 -178 2048 -144
rect 2048 -178 2064 -144
rect 1998 -190 2064 -178
rect 2418 -464 2452 -88
rect 2536 -464 2570 -88
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1562 -596 1664 -494
rect 2654 -464 2688 -88
rect 2772 -464 2806 -88
rect 2890 -464 2924 -88
rect 3008 -464 3042 -88
rect 3126 -464 3160 -88
rect 4067 -146 4133 -132
rect 4067 -180 4083 -146
rect 4083 -180 4117 -146
rect 4117 -180 4133 -146
rect 4067 -192 4133 -180
rect 4487 -466 4521 -90
rect 4605 -466 4639 -90
rect 1028 -688 1062 -654
rect 2448 -686 2482 -652
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 1318 -756 1352 -722
rect 2263 -753 2297 -719
rect 3630 -594 3732 -492
rect 4723 -466 4757 -90
rect 4841 -466 4875 -90
rect 4959 -466 4993 -90
rect 5077 -466 5111 -90
rect 5195 -466 5229 -90
rect 6135 -144 6201 -130
rect 6135 -178 6151 -144
rect 6151 -178 6185 -144
rect 6185 -178 6201 -144
rect 6135 -190 6201 -178
rect 6555 -464 6589 -88
rect 6673 -464 6707 -88
rect 3096 -686 3130 -652
rect 4517 -688 4551 -654
rect 2714 -770 2748 -736
rect 2832 -769 2866 -735
rect 3386 -754 3420 -720
rect 4332 -755 4366 -721
rect 48 -998 82 -822
rect 166 -998 200 -822
rect 468 -1198 502 -822
rect 586 -1198 620 -822
rect 704 -1198 738 -822
rect 822 -1198 856 -822
rect 940 -1198 974 -822
rect 1346 -998 1380 -822
rect 1464 -998 1498 -822
rect 2116 -996 2150 -820
rect 2234 -996 2268 -820
rect 2536 -1196 2570 -820
rect 2654 -1196 2688 -820
rect 2772 -1196 2806 -820
rect 2890 -1196 2924 -820
rect 3008 -1196 3042 -820
rect 3414 -996 3448 -820
rect 5699 -596 5801 -494
rect 6791 -464 6825 -88
rect 6909 -464 6943 -88
rect 7027 -464 7061 -88
rect 7145 -464 7179 -88
rect 7263 -464 7297 -88
rect 8204 -144 8270 -130
rect 8204 -178 8220 -144
rect 8220 -178 8254 -144
rect 8254 -178 8270 -144
rect 8204 -190 8270 -178
rect 8624 -464 8658 -88
rect 8742 -464 8776 -88
rect 5165 -688 5199 -654
rect 6585 -686 6619 -652
rect 4783 -772 4817 -738
rect 4901 -771 4935 -737
rect 5455 -756 5489 -722
rect 6400 -753 6434 -719
rect 7767 -594 7869 -492
rect 8860 -464 8894 -88
rect 8978 -464 9012 -88
rect 9096 -464 9130 -88
rect 9214 -464 9248 -88
rect 9332 -464 9366 -88
rect 10272 -142 10338 -128
rect 10272 -176 10288 -142
rect 10288 -176 10322 -142
rect 10322 -176 10338 -142
rect 10272 -188 10338 -176
rect 10692 -462 10726 -86
rect 10810 -462 10844 -86
rect 7233 -686 7267 -652
rect 8654 -686 8688 -652
rect 6851 -770 6885 -736
rect 6969 -769 7003 -735
rect 7523 -754 7557 -720
rect 8469 -753 8503 -719
rect 9836 -594 9938 -492
rect 10928 -462 10962 -86
rect 11046 -462 11080 -86
rect 11164 -462 11198 -86
rect 11282 -462 11316 -86
rect 11400 -462 11434 -86
rect 12341 -144 12407 -130
rect 12341 -178 12357 -144
rect 12357 -178 12391 -144
rect 12391 -178 12407 -144
rect 12341 -190 12407 -178
rect 12761 -464 12795 -88
rect 12879 -464 12913 -88
rect 9302 -686 9336 -652
rect 10722 -684 10756 -650
rect 8920 -770 8954 -736
rect 9038 -769 9072 -735
rect 9592 -754 9626 -720
rect 10537 -751 10571 -717
rect 11904 -592 12006 -490
rect 12997 -464 13031 -88
rect 13115 -464 13149 -88
rect 13233 -464 13267 -88
rect 13351 -464 13385 -88
rect 13469 -464 13503 -88
rect 14409 -142 14475 -128
rect 14409 -176 14425 -142
rect 14425 -176 14459 -142
rect 14459 -176 14475 -142
rect 14409 -188 14475 -176
rect 14829 -462 14863 -86
rect 14947 -462 14981 -86
rect 11370 -684 11404 -650
rect 12791 -686 12825 -652
rect 10988 -768 11022 -734
rect 11106 -767 11140 -733
rect 11660 -752 11694 -718
rect 12606 -753 12640 -719
rect 3532 -996 3566 -820
rect 4185 -998 4219 -822
rect 4303 -998 4337 -822
rect 4605 -1198 4639 -822
rect 4723 -1198 4757 -822
rect 4841 -1198 4875 -822
rect 4959 -1198 4993 -822
rect 5077 -1198 5111 -822
rect 5483 -998 5517 -822
rect 5601 -998 5635 -822
rect 6253 -996 6287 -820
rect 6371 -996 6405 -820
rect 6673 -1196 6707 -820
rect 6791 -1196 6825 -820
rect 6909 -1196 6943 -820
rect 7027 -1196 7061 -820
rect 7145 -1196 7179 -820
rect 7551 -996 7585 -820
rect 7669 -996 7703 -820
rect 8322 -996 8356 -820
rect 8440 -996 8474 -820
rect 8742 -1196 8776 -820
rect 8860 -1196 8894 -820
rect 8978 -1196 9012 -820
rect 9096 -1196 9130 -820
rect 9214 -1196 9248 -820
rect 9620 -996 9654 -820
rect 9738 -996 9772 -820
rect 10390 -994 10424 -818
rect 10508 -994 10542 -818
rect 10810 -1194 10844 -818
rect 10928 -1194 10962 -818
rect 11046 -1194 11080 -818
rect 11164 -1194 11198 -818
rect 11282 -1194 11316 -818
rect 11688 -994 11722 -818
rect 13973 -594 14075 -492
rect 15065 -462 15099 -86
rect 15183 -462 15217 -86
rect 15301 -462 15335 -86
rect 15419 -462 15453 -86
rect 15537 -462 15571 -86
rect 13439 -686 13473 -652
rect 14859 -684 14893 -650
rect 13057 -770 13091 -736
rect 13175 -769 13209 -735
rect 13729 -754 13763 -720
rect 14674 -751 14708 -717
rect 16041 -592 16143 -490
rect 15507 -684 15541 -650
rect 15125 -768 15159 -734
rect 15243 -767 15277 -733
rect 15797 -752 15831 -718
rect 11806 -994 11840 -818
rect 12459 -996 12493 -820
rect 12577 -996 12611 -820
rect 12879 -1196 12913 -820
rect 12997 -1196 13031 -820
rect 13115 -1196 13149 -820
rect 13233 -1196 13267 -820
rect 13351 -1196 13385 -820
rect 13757 -996 13791 -820
rect 13875 -996 13909 -820
rect 14527 -994 14561 -818
rect 14645 -994 14679 -818
rect 14947 -1194 14981 -818
rect 15065 -1194 15099 -818
rect 15183 -1194 15217 -818
rect 15301 -1194 15335 -818
rect 15419 -1194 15453 -818
rect 15825 -994 15859 -818
rect 15943 -994 15977 -818
rect 698 -1386 748 -1364
rect 698 -1406 748 -1386
rect 2766 -1384 2816 -1362
rect 2766 -1404 2816 -1384
rect 4835 -1386 4885 -1364
rect 4835 -1406 4885 -1386
rect 6903 -1384 6953 -1362
rect 6903 -1404 6953 -1384
rect 8972 -1384 9022 -1362
rect 8972 -1404 9022 -1384
rect 11040 -1382 11090 -1360
rect 11040 -1402 11090 -1382
rect 13109 -1384 13159 -1362
rect 13109 -1404 13159 -1384
rect 15177 -1382 15227 -1360
rect 15177 -1402 15227 -1382
<< metal1 >>
rect 740 844 750 866
rect 712 812 750 844
rect 804 844 814 866
rect 2808 846 2818 868
rect 804 812 846 844
rect 712 761 846 812
rect 2780 814 2818 846
rect 2872 846 2882 868
rect 2872 814 2914 846
rect 4877 844 4887 866
rect 2780 763 2914 814
rect 4849 812 4887 844
rect 4941 844 4951 866
rect 6945 846 6955 868
rect 4941 812 4983 844
rect 41 718 1514 761
rect 41 415 75 718
rect 407 615 441 718
rect 643 615 677 718
rect 879 615 913 718
rect 1115 615 1149 718
rect 401 603 447 615
rect -83 403 -37 415
rect -83 227 -77 403
rect -43 227 -37 403
rect -83 215 -37 227
rect 35 403 81 415
rect 35 227 41 403
rect 75 227 81 403
rect 35 215 81 227
rect 153 403 199 415
rect 153 227 159 403
rect 193 227 199 403
rect 153 215 199 227
rect 271 403 317 415
rect 401 403 407 603
rect 271 227 277 403
rect 311 227 407 403
rect 441 227 447 603
rect 271 215 317 227
rect 401 215 447 227
rect 519 603 565 615
rect 519 227 525 603
rect 559 227 565 603
rect 519 215 565 227
rect 637 603 683 615
rect 637 227 643 603
rect 677 227 683 603
rect 637 215 683 227
rect 755 603 801 615
rect 755 227 761 603
rect 795 227 801 603
rect 755 215 801 227
rect 873 603 919 615
rect 873 227 879 603
rect 913 227 919 603
rect 873 215 919 227
rect 991 603 1037 615
rect 991 227 997 603
rect 1031 227 1037 603
rect 991 215 1037 227
rect 1109 603 1155 615
rect 1109 227 1115 603
rect 1149 403 1155 603
rect 1480 415 1514 718
rect 2109 720 3582 763
rect 4849 761 4983 812
rect 6917 814 6955 846
rect 7009 846 7019 868
rect 9014 846 9024 868
rect 7009 814 7051 846
rect 6917 763 7051 814
rect 8986 814 9024 846
rect 9078 846 9088 868
rect 11082 848 11092 870
rect 9078 814 9120 846
rect 8986 763 9120 814
rect 11054 816 11092 848
rect 11146 848 11156 870
rect 11146 816 11188 848
rect 13151 846 13161 868
rect 11054 765 11188 816
rect 13123 814 13161 846
rect 13215 846 13225 868
rect 15219 848 15229 870
rect 13215 814 13257 846
rect 2109 417 2143 720
rect 2475 617 2509 720
rect 2711 617 2745 720
rect 2947 617 2981 720
rect 3183 617 3217 720
rect 2469 605 2515 617
rect 1238 403 1284 415
rect 1149 227 1244 403
rect 1278 227 1284 403
rect 1109 215 1155 227
rect 1238 215 1284 227
rect 1356 403 1402 415
rect 1356 227 1362 403
rect 1396 227 1402 403
rect 1356 215 1402 227
rect 1474 403 1520 415
rect 1474 227 1480 403
rect 1514 227 1520 403
rect 1474 215 1520 227
rect 1592 403 1638 415
rect 1592 227 1598 403
rect 1632 227 1638 403
rect 1592 215 1638 227
rect 1985 405 2031 417
rect 1985 229 1991 405
rect 2025 229 2031 405
rect 1985 217 2031 229
rect 2103 405 2149 417
rect 2103 229 2109 405
rect 2143 229 2149 405
rect 2103 217 2149 229
rect 2221 405 2267 417
rect 2221 229 2227 405
rect 2261 229 2267 405
rect 2221 217 2267 229
rect 2339 405 2385 417
rect 2469 405 2475 605
rect 2339 229 2345 405
rect 2379 229 2475 405
rect 2509 229 2515 605
rect 2339 217 2385 229
rect 2469 217 2515 229
rect 2587 605 2633 617
rect 2587 229 2593 605
rect 2627 229 2633 605
rect 2587 217 2633 229
rect 2705 605 2751 617
rect 2705 229 2711 605
rect 2745 229 2751 605
rect 2705 217 2751 229
rect 2823 605 2869 617
rect 2823 229 2829 605
rect 2863 229 2869 605
rect 2823 217 2869 229
rect 2941 605 2987 617
rect 2941 229 2947 605
rect 2981 229 2987 605
rect 2941 217 2987 229
rect 3059 605 3105 617
rect 3059 229 3065 605
rect 3099 229 3105 605
rect 3059 217 3105 229
rect 3177 605 3223 617
rect 3177 229 3183 605
rect 3217 405 3223 605
rect 3548 417 3582 720
rect 4178 718 5651 761
rect 3306 405 3352 417
rect 3217 229 3312 405
rect 3346 229 3352 405
rect 3177 217 3223 229
rect 3306 217 3352 229
rect 3424 405 3470 417
rect 3424 229 3430 405
rect 3464 229 3470 405
rect 3424 217 3470 229
rect 3542 405 3588 417
rect 3542 229 3548 405
rect 3582 229 3588 405
rect 3542 217 3588 229
rect 3660 405 3706 417
rect 4178 415 4212 718
rect 4544 615 4578 718
rect 4780 615 4814 718
rect 5016 615 5050 718
rect 5252 615 5286 718
rect 4538 603 4584 615
rect 3660 229 3666 405
rect 3700 229 3706 405
rect 3660 217 3706 229
rect 4054 403 4100 415
rect 4054 227 4060 403
rect 4094 227 4100 403
rect -77 181 -43 215
rect 525 181 559 215
rect 761 181 795 215
rect -77 146 82 181
rect 525 146 795 181
rect 1362 181 1396 215
rect 1598 181 1632 215
rect 1362 146 1632 181
rect 1991 183 2025 217
rect 2593 183 2627 217
rect 2829 183 2863 217
rect 1991 148 2150 183
rect 2593 148 2863 183
rect 3430 183 3464 217
rect 3666 183 3700 217
rect 4054 215 4100 227
rect 4172 403 4218 415
rect 4172 227 4178 403
rect 4212 227 4218 403
rect 4172 215 4218 227
rect 4290 403 4336 415
rect 4290 227 4296 403
rect 4330 227 4336 403
rect 4290 215 4336 227
rect 4408 403 4454 415
rect 4538 403 4544 603
rect 4408 227 4414 403
rect 4448 227 4544 403
rect 4578 227 4584 603
rect 4408 215 4454 227
rect 4538 215 4584 227
rect 4656 603 4702 615
rect 4656 227 4662 603
rect 4696 227 4702 603
rect 4656 215 4702 227
rect 4774 603 4820 615
rect 4774 227 4780 603
rect 4814 227 4820 603
rect 4774 215 4820 227
rect 4892 603 4938 615
rect 4892 227 4898 603
rect 4932 227 4938 603
rect 4892 215 4938 227
rect 5010 603 5056 615
rect 5010 227 5016 603
rect 5050 227 5056 603
rect 5010 215 5056 227
rect 5128 603 5174 615
rect 5128 227 5134 603
rect 5168 227 5174 603
rect 5128 215 5174 227
rect 5246 603 5292 615
rect 5246 227 5252 603
rect 5286 403 5292 603
rect 5617 415 5651 718
rect 6246 720 7719 763
rect 6246 417 6280 720
rect 6612 617 6646 720
rect 6848 617 6882 720
rect 7084 617 7118 720
rect 7320 617 7354 720
rect 6606 605 6652 617
rect 5375 403 5421 415
rect 5286 227 5381 403
rect 5415 227 5421 403
rect 5246 215 5292 227
rect 5375 215 5421 227
rect 5493 403 5539 415
rect 5493 227 5499 403
rect 5533 227 5539 403
rect 5493 215 5539 227
rect 5611 403 5657 415
rect 5611 227 5617 403
rect 5651 227 5657 403
rect 5611 215 5657 227
rect 5729 403 5775 415
rect 5729 227 5735 403
rect 5769 227 5775 403
rect 5729 215 5775 227
rect 6122 405 6168 417
rect 6122 229 6128 405
rect 6162 229 6168 405
rect 6122 217 6168 229
rect 6240 405 6286 417
rect 6240 229 6246 405
rect 6280 229 6286 405
rect 6240 217 6286 229
rect 6358 405 6404 417
rect 6358 229 6364 405
rect 6398 229 6404 405
rect 6358 217 6404 229
rect 6476 405 6522 417
rect 6606 405 6612 605
rect 6476 229 6482 405
rect 6516 229 6612 405
rect 6646 229 6652 605
rect 6476 217 6522 229
rect 6606 217 6652 229
rect 6724 605 6770 617
rect 6724 229 6730 605
rect 6764 229 6770 605
rect 6724 217 6770 229
rect 6842 605 6888 617
rect 6842 229 6848 605
rect 6882 229 6888 605
rect 6842 217 6888 229
rect 6960 605 7006 617
rect 6960 229 6966 605
rect 7000 229 7006 605
rect 6960 217 7006 229
rect 7078 605 7124 617
rect 7078 229 7084 605
rect 7118 229 7124 605
rect 7078 217 7124 229
rect 7196 605 7242 617
rect 7196 229 7202 605
rect 7236 229 7242 605
rect 7196 217 7242 229
rect 7314 605 7360 617
rect 7314 229 7320 605
rect 7354 405 7360 605
rect 7685 417 7719 720
rect 8315 720 9788 763
rect 8315 417 8349 720
rect 8681 617 8715 720
rect 8917 617 8951 720
rect 9153 617 9187 720
rect 9389 617 9423 720
rect 8675 605 8721 617
rect 7443 405 7489 417
rect 7354 229 7449 405
rect 7483 229 7489 405
rect 7314 217 7360 229
rect 7443 217 7489 229
rect 7561 405 7607 417
rect 7561 229 7567 405
rect 7601 229 7607 405
rect 7561 217 7607 229
rect 7679 405 7725 417
rect 7679 229 7685 405
rect 7719 229 7725 405
rect 7679 217 7725 229
rect 7797 405 7843 417
rect 7797 229 7803 405
rect 7837 229 7843 405
rect 7797 217 7843 229
rect 8191 405 8237 417
rect 8191 229 8197 405
rect 8231 229 8237 405
rect 8191 217 8237 229
rect 8309 405 8355 417
rect 8309 229 8315 405
rect 8349 229 8355 405
rect 8309 217 8355 229
rect 8427 405 8473 417
rect 8427 229 8433 405
rect 8467 229 8473 405
rect 8427 217 8473 229
rect 8545 405 8591 417
rect 8675 405 8681 605
rect 8545 229 8551 405
rect 8585 229 8681 405
rect 8715 229 8721 605
rect 8545 217 8591 229
rect 8675 217 8721 229
rect 8793 605 8839 617
rect 8793 229 8799 605
rect 8833 229 8839 605
rect 8793 217 8839 229
rect 8911 605 8957 617
rect 8911 229 8917 605
rect 8951 229 8957 605
rect 8911 217 8957 229
rect 9029 605 9075 617
rect 9029 229 9035 605
rect 9069 229 9075 605
rect 9029 217 9075 229
rect 9147 605 9193 617
rect 9147 229 9153 605
rect 9187 229 9193 605
rect 9147 217 9193 229
rect 9265 605 9311 617
rect 9265 229 9271 605
rect 9305 229 9311 605
rect 9265 217 9311 229
rect 9383 605 9429 617
rect 9383 229 9389 605
rect 9423 405 9429 605
rect 9754 417 9788 720
rect 10383 722 11856 765
rect 13123 763 13257 814
rect 15191 816 15229 848
rect 15283 848 15293 870
rect 15283 816 15325 848
rect 15191 765 15325 816
rect 10383 419 10417 722
rect 10749 619 10783 722
rect 10985 619 11019 722
rect 11221 619 11255 722
rect 11457 619 11491 722
rect 10743 607 10789 619
rect 9512 405 9558 417
rect 9423 229 9518 405
rect 9552 229 9558 405
rect 9383 217 9429 229
rect 9512 217 9558 229
rect 9630 405 9676 417
rect 9630 229 9636 405
rect 9670 229 9676 405
rect 9630 217 9676 229
rect 9748 405 9794 417
rect 9748 229 9754 405
rect 9788 229 9794 405
rect 9748 217 9794 229
rect 9866 405 9912 417
rect 9866 229 9872 405
rect 9906 229 9912 405
rect 9866 217 9912 229
rect 10259 407 10305 419
rect 10259 231 10265 407
rect 10299 231 10305 407
rect 10259 219 10305 231
rect 10377 407 10423 419
rect 10377 231 10383 407
rect 10417 231 10423 407
rect 10377 219 10423 231
rect 10495 407 10541 419
rect 10495 231 10501 407
rect 10535 231 10541 407
rect 10495 219 10541 231
rect 10613 407 10659 419
rect 10743 407 10749 607
rect 10613 231 10619 407
rect 10653 231 10749 407
rect 10783 231 10789 607
rect 10613 219 10659 231
rect 10743 219 10789 231
rect 10861 607 10907 619
rect 10861 231 10867 607
rect 10901 231 10907 607
rect 10861 219 10907 231
rect 10979 607 11025 619
rect 10979 231 10985 607
rect 11019 231 11025 607
rect 10979 219 11025 231
rect 11097 607 11143 619
rect 11097 231 11103 607
rect 11137 231 11143 607
rect 11097 219 11143 231
rect 11215 607 11261 619
rect 11215 231 11221 607
rect 11255 231 11261 607
rect 11215 219 11261 231
rect 11333 607 11379 619
rect 11333 231 11339 607
rect 11373 231 11379 607
rect 11333 219 11379 231
rect 11451 607 11497 619
rect 11451 231 11457 607
rect 11491 407 11497 607
rect 11822 419 11856 722
rect 12452 720 13925 763
rect 11580 407 11626 419
rect 11491 231 11586 407
rect 11620 231 11626 407
rect 11451 219 11497 231
rect 11580 219 11626 231
rect 11698 407 11744 419
rect 11698 231 11704 407
rect 11738 231 11744 407
rect 11698 219 11744 231
rect 11816 407 11862 419
rect 11816 231 11822 407
rect 11856 231 11862 407
rect 11816 219 11862 231
rect 11934 407 11980 419
rect 12452 417 12486 720
rect 12818 617 12852 720
rect 13054 617 13088 720
rect 13290 617 13324 720
rect 13526 617 13560 720
rect 12812 605 12858 617
rect 11934 231 11940 407
rect 11974 231 11980 407
rect 11934 219 11980 231
rect 12328 405 12374 417
rect 12328 229 12334 405
rect 12368 229 12374 405
rect 3430 148 3700 183
rect 4060 181 4094 215
rect 4662 181 4696 215
rect 4898 181 4932 215
rect -132 -2 -58 64
rect 8 -2 18 64
rect -132 -132 8 -126
rect -132 -192 -70 -132
rect -4 -192 8 -132
rect -132 -198 8 -192
rect 48 -638 82 146
rect 761 84 795 146
rect 350 46 1092 84
rect 350 -78 384 46
rect 586 -78 620 46
rect 822 -78 856 46
rect 1058 -78 1092 46
rect 1318 58 1396 64
rect 1318 4 1330 58
rect 1384 4 1396 58
rect 1318 -2 1396 4
rect 344 -90 390 -78
rect 344 -466 350 -90
rect 384 -466 390 -90
rect 344 -478 390 -466
rect 462 -90 508 -78
rect 462 -466 468 -90
rect 502 -466 508 -90
rect 462 -478 508 -466
rect 580 -90 626 -78
rect 580 -466 586 -90
rect 620 -466 626 -90
rect 580 -478 626 -466
rect 698 -90 744 -78
rect 698 -466 704 -90
rect 738 -466 744 -90
rect 698 -478 744 -466
rect 816 -90 862 -78
rect 816 -466 822 -90
rect 856 -466 862 -90
rect 816 -478 862 -466
rect 934 -90 980 -78
rect 934 -466 940 -90
rect 974 -466 980 -90
rect 934 -478 980 -466
rect 1052 -90 1098 -78
rect 1052 -466 1058 -90
rect 1092 -466 1098 -90
rect 1052 -478 1098 -466
rect 1464 -637 1498 146
rect 1936 0 2010 66
rect 2076 0 2086 66
rect 1936 -130 2076 -124
rect 1936 -190 1998 -130
rect 2064 -190 2076 -130
rect 1936 -196 2076 -190
rect 1550 -494 1676 -488
rect 1550 -596 1562 -494
rect 1664 -596 1676 -494
rect 1550 -602 1676 -596
rect 1191 -638 1498 -637
rect 48 -643 364 -638
rect 1078 -643 1498 -638
rect 48 -654 431 -643
rect 48 -681 380 -654
rect 48 -810 82 -681
rect 364 -688 380 -681
rect 414 -688 431 -654
rect 364 -694 431 -688
rect 1011 -654 1498 -643
rect 1011 -688 1028 -654
rect 1062 -681 1498 -654
rect 1062 -688 1078 -681
rect 1191 -682 1498 -681
rect 1011 -694 1078 -688
rect 189 -721 245 -709
rect 189 -755 195 -721
rect 229 -722 245 -721
rect 1302 -722 1358 -710
rect 229 -738 696 -722
rect 229 -755 646 -738
rect 189 -771 646 -755
rect 630 -772 646 -771
rect 680 -772 696 -738
rect 630 -779 696 -772
rect 748 -737 1318 -722
rect 748 -771 764 -737
rect 798 -756 1318 -737
rect 1352 -756 1358 -722
rect 798 -771 1358 -756
rect 748 -781 815 -771
rect 1302 -772 1358 -771
rect 1464 -810 1498 -682
rect 2116 -636 2150 148
rect 2829 86 2863 148
rect 2418 48 3160 86
rect 2418 -76 2452 48
rect 2654 -76 2688 48
rect 2890 -76 2924 48
rect 3126 -76 3160 48
rect 3386 60 3464 66
rect 3386 6 3398 60
rect 3452 6 3464 60
rect 3386 0 3464 6
rect 2412 -88 2458 -76
rect 2412 -464 2418 -88
rect 2452 -464 2458 -88
rect 2412 -476 2458 -464
rect 2530 -88 2576 -76
rect 2530 -464 2536 -88
rect 2570 -464 2576 -88
rect 2530 -476 2576 -464
rect 2648 -88 2694 -76
rect 2648 -464 2654 -88
rect 2688 -464 2694 -88
rect 2648 -476 2694 -464
rect 2766 -88 2812 -76
rect 2766 -464 2772 -88
rect 2806 -464 2812 -88
rect 2766 -476 2812 -464
rect 2884 -88 2930 -76
rect 2884 -464 2890 -88
rect 2924 -464 2930 -88
rect 2884 -476 2930 -464
rect 3002 -88 3048 -76
rect 3002 -464 3008 -88
rect 3042 -464 3048 -88
rect 3002 -476 3048 -464
rect 3120 -88 3166 -76
rect 3120 -464 3126 -88
rect 3160 -464 3166 -88
rect 3120 -476 3166 -464
rect 3532 -635 3566 148
rect 4060 146 4219 181
rect 4662 146 4932 181
rect 5499 181 5533 215
rect 5735 181 5769 215
rect 5499 146 5769 181
rect 6128 183 6162 217
rect 6730 183 6764 217
rect 6966 183 7000 217
rect 6128 148 6287 183
rect 6730 148 7000 183
rect 7567 183 7601 217
rect 7803 183 7837 217
rect 7567 148 7837 183
rect 8197 183 8231 217
rect 8799 183 8833 217
rect 9035 183 9069 217
rect 8197 148 8356 183
rect 8799 148 9069 183
rect 9636 183 9670 217
rect 9872 183 9906 217
rect 9636 148 9906 183
rect 10265 185 10299 219
rect 10867 185 10901 219
rect 11103 185 11137 219
rect 10265 150 10424 185
rect 10867 150 11137 185
rect 11704 185 11738 219
rect 11940 185 11974 219
rect 12328 217 12374 229
rect 12446 405 12492 417
rect 12446 229 12452 405
rect 12486 229 12492 405
rect 12446 217 12492 229
rect 12564 405 12610 417
rect 12564 229 12570 405
rect 12604 229 12610 405
rect 12564 217 12610 229
rect 12682 405 12728 417
rect 12812 405 12818 605
rect 12682 229 12688 405
rect 12722 229 12818 405
rect 12852 229 12858 605
rect 12682 217 12728 229
rect 12812 217 12858 229
rect 12930 605 12976 617
rect 12930 229 12936 605
rect 12970 229 12976 605
rect 12930 217 12976 229
rect 13048 605 13094 617
rect 13048 229 13054 605
rect 13088 229 13094 605
rect 13048 217 13094 229
rect 13166 605 13212 617
rect 13166 229 13172 605
rect 13206 229 13212 605
rect 13166 217 13212 229
rect 13284 605 13330 617
rect 13284 229 13290 605
rect 13324 229 13330 605
rect 13284 217 13330 229
rect 13402 605 13448 617
rect 13402 229 13408 605
rect 13442 229 13448 605
rect 13402 217 13448 229
rect 13520 605 13566 617
rect 13520 229 13526 605
rect 13560 405 13566 605
rect 13891 417 13925 720
rect 14520 722 15993 765
rect 14520 419 14554 722
rect 14886 619 14920 722
rect 15122 619 15156 722
rect 15358 619 15392 722
rect 15594 619 15628 722
rect 14880 607 14926 619
rect 13649 405 13695 417
rect 13560 229 13655 405
rect 13689 229 13695 405
rect 13520 217 13566 229
rect 13649 217 13695 229
rect 13767 405 13813 417
rect 13767 229 13773 405
rect 13807 229 13813 405
rect 13767 217 13813 229
rect 13885 405 13931 417
rect 13885 229 13891 405
rect 13925 229 13931 405
rect 13885 217 13931 229
rect 14003 405 14049 417
rect 14003 229 14009 405
rect 14043 229 14049 405
rect 14003 217 14049 229
rect 14396 407 14442 419
rect 14396 231 14402 407
rect 14436 231 14442 407
rect 14396 219 14442 231
rect 14514 407 14560 419
rect 14514 231 14520 407
rect 14554 231 14560 407
rect 14514 219 14560 231
rect 14632 407 14678 419
rect 14632 231 14638 407
rect 14672 231 14678 407
rect 14632 219 14678 231
rect 14750 407 14796 419
rect 14880 407 14886 607
rect 14750 231 14756 407
rect 14790 231 14886 407
rect 14920 231 14926 607
rect 14750 219 14796 231
rect 14880 219 14926 231
rect 14998 607 15044 619
rect 14998 231 15004 607
rect 15038 231 15044 607
rect 14998 219 15044 231
rect 15116 607 15162 619
rect 15116 231 15122 607
rect 15156 231 15162 607
rect 15116 219 15162 231
rect 15234 607 15280 619
rect 15234 231 15240 607
rect 15274 231 15280 607
rect 15234 219 15280 231
rect 15352 607 15398 619
rect 15352 231 15358 607
rect 15392 231 15398 607
rect 15352 219 15398 231
rect 15470 607 15516 619
rect 15470 231 15476 607
rect 15510 231 15516 607
rect 15470 219 15516 231
rect 15588 607 15634 619
rect 15588 231 15594 607
rect 15628 407 15634 607
rect 15959 419 15993 722
rect 15717 407 15763 419
rect 15628 231 15723 407
rect 15757 231 15763 407
rect 15588 219 15634 231
rect 15717 219 15763 231
rect 15835 407 15881 419
rect 15835 231 15841 407
rect 15875 231 15881 407
rect 15835 219 15881 231
rect 15953 407 15999 419
rect 15953 231 15959 407
rect 15993 231 15999 407
rect 15953 219 15999 231
rect 16071 407 16117 419
rect 16071 231 16077 407
rect 16111 231 16117 407
rect 16071 219 16117 231
rect 11704 150 11974 185
rect 12334 183 12368 217
rect 12936 183 12970 217
rect 13172 183 13206 217
rect 4005 -2 4079 64
rect 4145 -2 4155 64
rect 4005 -132 4145 -126
rect 4005 -192 4067 -132
rect 4133 -192 4145 -132
rect 4005 -198 4145 -192
rect 3618 -492 3744 -486
rect 3618 -594 3630 -492
rect 3732 -594 3744 -492
rect 3618 -600 3744 -594
rect 3259 -636 3566 -635
rect 2116 -641 2432 -636
rect 3146 -641 3566 -636
rect 2116 -652 2499 -641
rect 2116 -679 2448 -652
rect 2116 -808 2150 -679
rect 2432 -686 2448 -679
rect 2482 -686 2499 -652
rect 2432 -692 2499 -686
rect 3079 -652 3566 -641
rect 3079 -686 3096 -652
rect 3130 -679 3566 -652
rect 3130 -686 3146 -679
rect 3259 -680 3566 -679
rect 3079 -692 3146 -686
rect 2257 -719 2313 -707
rect 2257 -753 2263 -719
rect 2297 -720 2313 -719
rect 3370 -720 3426 -708
rect 2297 -736 2764 -720
rect 2297 -753 2714 -736
rect 2257 -769 2714 -753
rect 2698 -770 2714 -769
rect 2748 -770 2764 -736
rect 2698 -777 2764 -770
rect 2816 -735 3386 -720
rect 2816 -769 2832 -735
rect 2866 -754 3386 -735
rect 3420 -754 3426 -720
rect 2866 -769 3426 -754
rect 2816 -779 2883 -769
rect 3370 -770 3426 -769
rect 3532 -808 3566 -680
rect 4185 -638 4219 146
rect 4898 84 4932 146
rect 4487 46 5229 84
rect 4487 -78 4521 46
rect 4723 -78 4757 46
rect 4959 -78 4993 46
rect 5195 -78 5229 46
rect 5455 58 5533 64
rect 5455 4 5467 58
rect 5521 4 5533 58
rect 5455 -2 5533 4
rect 4481 -90 4527 -78
rect 4481 -466 4487 -90
rect 4521 -466 4527 -90
rect 4481 -478 4527 -466
rect 4599 -90 4645 -78
rect 4599 -466 4605 -90
rect 4639 -466 4645 -90
rect 4599 -478 4645 -466
rect 4717 -90 4763 -78
rect 4717 -466 4723 -90
rect 4757 -466 4763 -90
rect 4717 -478 4763 -466
rect 4835 -90 4881 -78
rect 4835 -466 4841 -90
rect 4875 -466 4881 -90
rect 4835 -478 4881 -466
rect 4953 -90 4999 -78
rect 4953 -466 4959 -90
rect 4993 -466 4999 -90
rect 4953 -478 4999 -466
rect 5071 -90 5117 -78
rect 5071 -466 5077 -90
rect 5111 -466 5117 -90
rect 5071 -478 5117 -466
rect 5189 -90 5235 -78
rect 5189 -466 5195 -90
rect 5229 -466 5235 -90
rect 5189 -478 5235 -466
rect 5601 -637 5635 146
rect 6073 0 6147 66
rect 6213 0 6223 66
rect 6073 -130 6213 -124
rect 6073 -190 6135 -130
rect 6201 -190 6213 -130
rect 6073 -196 6213 -190
rect 5687 -494 5813 -488
rect 5687 -596 5699 -494
rect 5801 -596 5813 -494
rect 5687 -602 5813 -596
rect 5328 -638 5635 -637
rect 4185 -643 4501 -638
rect 5215 -643 5635 -638
rect 4185 -654 4568 -643
rect 4185 -681 4517 -654
rect 42 -822 88 -810
rect 42 -998 48 -822
rect 82 -998 88 -822
rect 42 -1010 88 -998
rect 160 -822 206 -810
rect 160 -998 166 -822
rect 200 -998 206 -822
rect 160 -1010 206 -998
rect 462 -822 508 -810
rect 165 -1304 199 -1010
rect 462 -1198 468 -822
rect 502 -1198 508 -822
rect 462 -1210 508 -1198
rect 580 -822 626 -810
rect 580 -1198 586 -822
rect 620 -1198 626 -822
rect 580 -1210 626 -1198
rect 698 -822 744 -810
rect 698 -1198 704 -822
rect 738 -1198 744 -822
rect 698 -1210 744 -1198
rect 816 -822 862 -810
rect 816 -1198 822 -822
rect 856 -1198 862 -822
rect 816 -1210 862 -1198
rect 934 -822 980 -810
rect 934 -1198 940 -822
rect 974 -1198 980 -822
rect 1340 -822 1386 -810
rect 1340 -998 1346 -822
rect 1380 -998 1386 -822
rect 1340 -1010 1386 -998
rect 1458 -822 1504 -810
rect 1458 -998 1464 -822
rect 1498 -998 1504 -822
rect 1458 -1010 1504 -998
rect 2110 -820 2156 -808
rect 2110 -996 2116 -820
rect 2150 -996 2156 -820
rect 2110 -1008 2156 -996
rect 2228 -820 2274 -808
rect 2228 -996 2234 -820
rect 2268 -996 2274 -820
rect 2228 -1008 2274 -996
rect 2530 -820 2576 -808
rect 934 -1210 980 -1198
rect 822 -1304 856 -1210
rect 1346 -1304 1379 -1010
rect 165 -1336 1379 -1304
rect 2233 -1302 2267 -1008
rect 2530 -1196 2536 -820
rect 2570 -1196 2576 -820
rect 2530 -1208 2576 -1196
rect 2648 -820 2694 -808
rect 2648 -1196 2654 -820
rect 2688 -1196 2694 -820
rect 2648 -1208 2694 -1196
rect 2766 -820 2812 -808
rect 2766 -1196 2772 -820
rect 2806 -1196 2812 -820
rect 2766 -1208 2812 -1196
rect 2884 -820 2930 -808
rect 2884 -1196 2890 -820
rect 2924 -1196 2930 -820
rect 2884 -1208 2930 -1196
rect 3002 -820 3048 -808
rect 3002 -1196 3008 -820
rect 3042 -1196 3048 -820
rect 3408 -820 3454 -808
rect 3408 -996 3414 -820
rect 3448 -996 3454 -820
rect 3408 -1008 3454 -996
rect 3526 -820 3572 -808
rect 4185 -810 4219 -681
rect 4501 -688 4517 -681
rect 4551 -688 4568 -654
rect 4501 -694 4568 -688
rect 5148 -654 5635 -643
rect 5148 -688 5165 -654
rect 5199 -681 5635 -654
rect 5199 -688 5215 -681
rect 5328 -682 5635 -681
rect 5148 -694 5215 -688
rect 4326 -721 4382 -709
rect 4326 -755 4332 -721
rect 4366 -722 4382 -721
rect 5439 -722 5495 -710
rect 4366 -738 4833 -722
rect 4366 -755 4783 -738
rect 4326 -771 4783 -755
rect 4767 -772 4783 -771
rect 4817 -772 4833 -738
rect 4767 -779 4833 -772
rect 4885 -737 5455 -722
rect 4885 -771 4901 -737
rect 4935 -756 5455 -737
rect 5489 -756 5495 -722
rect 4935 -771 5495 -756
rect 4885 -781 4952 -771
rect 5439 -772 5495 -771
rect 5601 -810 5635 -682
rect 6253 -636 6287 148
rect 6966 86 7000 148
rect 6555 48 7297 86
rect 6555 -76 6589 48
rect 6791 -76 6825 48
rect 7027 -76 7061 48
rect 7263 -76 7297 48
rect 7523 60 7601 66
rect 7523 6 7535 60
rect 7589 6 7601 60
rect 7523 0 7601 6
rect 6549 -88 6595 -76
rect 6549 -464 6555 -88
rect 6589 -464 6595 -88
rect 6549 -476 6595 -464
rect 6667 -88 6713 -76
rect 6667 -464 6673 -88
rect 6707 -464 6713 -88
rect 6667 -476 6713 -464
rect 6785 -88 6831 -76
rect 6785 -464 6791 -88
rect 6825 -464 6831 -88
rect 6785 -476 6831 -464
rect 6903 -88 6949 -76
rect 6903 -464 6909 -88
rect 6943 -464 6949 -88
rect 6903 -476 6949 -464
rect 7021 -88 7067 -76
rect 7021 -464 7027 -88
rect 7061 -464 7067 -88
rect 7021 -476 7067 -464
rect 7139 -88 7185 -76
rect 7139 -464 7145 -88
rect 7179 -464 7185 -88
rect 7139 -476 7185 -464
rect 7257 -88 7303 -76
rect 7257 -464 7263 -88
rect 7297 -464 7303 -88
rect 7257 -476 7303 -464
rect 7669 -635 7703 148
rect 8142 0 8216 66
rect 8282 0 8292 66
rect 8142 -130 8282 -124
rect 8142 -190 8204 -130
rect 8270 -190 8282 -130
rect 8142 -196 8282 -190
rect 7755 -492 7881 -486
rect 7755 -594 7767 -492
rect 7869 -594 7881 -492
rect 7755 -600 7881 -594
rect 7396 -636 7703 -635
rect 6253 -641 6569 -636
rect 7283 -641 7703 -636
rect 6253 -652 6636 -641
rect 6253 -679 6585 -652
rect 6253 -808 6287 -679
rect 6569 -686 6585 -679
rect 6619 -686 6636 -652
rect 6569 -692 6636 -686
rect 7216 -652 7703 -641
rect 7216 -686 7233 -652
rect 7267 -679 7703 -652
rect 7267 -686 7283 -679
rect 7396 -680 7703 -679
rect 7216 -692 7283 -686
rect 6394 -719 6450 -707
rect 6394 -753 6400 -719
rect 6434 -720 6450 -719
rect 7507 -720 7563 -708
rect 6434 -736 6901 -720
rect 6434 -753 6851 -736
rect 6394 -769 6851 -753
rect 6835 -770 6851 -769
rect 6885 -770 6901 -736
rect 6835 -777 6901 -770
rect 6953 -735 7523 -720
rect 6953 -769 6969 -735
rect 7003 -754 7523 -735
rect 7557 -754 7563 -720
rect 7003 -769 7563 -754
rect 6953 -779 7020 -769
rect 7507 -770 7563 -769
rect 7669 -808 7703 -680
rect 8322 -636 8356 148
rect 9035 86 9069 148
rect 8624 48 9366 86
rect 8624 -76 8658 48
rect 8860 -76 8894 48
rect 9096 -76 9130 48
rect 9332 -76 9366 48
rect 9592 60 9670 66
rect 9592 6 9604 60
rect 9658 6 9670 60
rect 9592 0 9670 6
rect 8618 -88 8664 -76
rect 8618 -464 8624 -88
rect 8658 -464 8664 -88
rect 8618 -476 8664 -464
rect 8736 -88 8782 -76
rect 8736 -464 8742 -88
rect 8776 -464 8782 -88
rect 8736 -476 8782 -464
rect 8854 -88 8900 -76
rect 8854 -464 8860 -88
rect 8894 -464 8900 -88
rect 8854 -476 8900 -464
rect 8972 -88 9018 -76
rect 8972 -464 8978 -88
rect 9012 -464 9018 -88
rect 8972 -476 9018 -464
rect 9090 -88 9136 -76
rect 9090 -464 9096 -88
rect 9130 -464 9136 -88
rect 9090 -476 9136 -464
rect 9208 -88 9254 -76
rect 9208 -464 9214 -88
rect 9248 -464 9254 -88
rect 9208 -476 9254 -464
rect 9326 -88 9372 -76
rect 9326 -464 9332 -88
rect 9366 -464 9372 -88
rect 9326 -476 9372 -464
rect 9738 -635 9772 148
rect 10210 2 10284 68
rect 10350 2 10360 68
rect 10210 -128 10350 -122
rect 10210 -188 10272 -128
rect 10338 -188 10350 -128
rect 10210 -194 10350 -188
rect 9824 -492 9950 -486
rect 9824 -594 9836 -492
rect 9938 -594 9950 -492
rect 9824 -600 9950 -594
rect 9465 -636 9772 -635
rect 8322 -641 8638 -636
rect 9352 -641 9772 -636
rect 8322 -652 8705 -641
rect 8322 -679 8654 -652
rect 8322 -808 8356 -679
rect 8638 -686 8654 -679
rect 8688 -686 8705 -652
rect 8638 -692 8705 -686
rect 9285 -652 9772 -641
rect 9285 -686 9302 -652
rect 9336 -679 9772 -652
rect 9336 -686 9352 -679
rect 9465 -680 9772 -679
rect 9285 -692 9352 -686
rect 8463 -719 8519 -707
rect 8463 -753 8469 -719
rect 8503 -720 8519 -719
rect 9576 -720 9632 -708
rect 8503 -736 8970 -720
rect 8503 -753 8920 -736
rect 8463 -769 8920 -753
rect 8904 -770 8920 -769
rect 8954 -770 8970 -736
rect 8904 -777 8970 -770
rect 9022 -735 9592 -720
rect 9022 -769 9038 -735
rect 9072 -754 9592 -735
rect 9626 -754 9632 -720
rect 9072 -769 9632 -754
rect 9022 -779 9089 -769
rect 9576 -770 9632 -769
rect 9738 -808 9772 -680
rect 10390 -634 10424 150
rect 11103 88 11137 150
rect 10692 50 11434 88
rect 10692 -74 10726 50
rect 10928 -74 10962 50
rect 11164 -74 11198 50
rect 11400 -74 11434 50
rect 11660 62 11738 68
rect 11660 8 11672 62
rect 11726 8 11738 62
rect 11660 2 11738 8
rect 10686 -86 10732 -74
rect 10686 -462 10692 -86
rect 10726 -462 10732 -86
rect 10686 -474 10732 -462
rect 10804 -86 10850 -74
rect 10804 -462 10810 -86
rect 10844 -462 10850 -86
rect 10804 -474 10850 -462
rect 10922 -86 10968 -74
rect 10922 -462 10928 -86
rect 10962 -462 10968 -86
rect 10922 -474 10968 -462
rect 11040 -86 11086 -74
rect 11040 -462 11046 -86
rect 11080 -462 11086 -86
rect 11040 -474 11086 -462
rect 11158 -86 11204 -74
rect 11158 -462 11164 -86
rect 11198 -462 11204 -86
rect 11158 -474 11204 -462
rect 11276 -86 11322 -74
rect 11276 -462 11282 -86
rect 11316 -462 11322 -86
rect 11276 -474 11322 -462
rect 11394 -86 11440 -74
rect 11394 -462 11400 -86
rect 11434 -462 11440 -86
rect 11394 -474 11440 -462
rect 11806 -633 11840 150
rect 12334 148 12493 183
rect 12936 148 13206 183
rect 13773 183 13807 217
rect 14009 183 14043 217
rect 13773 148 14043 183
rect 14402 185 14436 219
rect 15004 185 15038 219
rect 15240 185 15274 219
rect 14402 150 14561 185
rect 15004 150 15274 185
rect 15841 185 15875 219
rect 16077 185 16111 219
rect 15841 150 16111 185
rect 12279 0 12353 66
rect 12419 0 12429 66
rect 12279 -130 12419 -124
rect 12279 -190 12341 -130
rect 12407 -190 12419 -130
rect 12279 -196 12419 -190
rect 11892 -490 12018 -484
rect 11892 -592 11904 -490
rect 12006 -592 12018 -490
rect 11892 -598 12018 -592
rect 11533 -634 11840 -633
rect 10390 -639 10706 -634
rect 11420 -639 11840 -634
rect 10390 -650 10773 -639
rect 10390 -677 10722 -650
rect 10390 -806 10424 -677
rect 10706 -684 10722 -677
rect 10756 -684 10773 -650
rect 10706 -690 10773 -684
rect 11353 -650 11840 -639
rect 11353 -684 11370 -650
rect 11404 -677 11840 -650
rect 11404 -684 11420 -677
rect 11533 -678 11840 -677
rect 11353 -690 11420 -684
rect 10531 -717 10587 -705
rect 10531 -751 10537 -717
rect 10571 -718 10587 -717
rect 11644 -718 11700 -706
rect 10571 -734 11038 -718
rect 10571 -751 10988 -734
rect 10531 -767 10988 -751
rect 10972 -768 10988 -767
rect 11022 -768 11038 -734
rect 10972 -775 11038 -768
rect 11090 -733 11660 -718
rect 11090 -767 11106 -733
rect 11140 -752 11660 -733
rect 11694 -752 11700 -718
rect 11140 -767 11700 -752
rect 11090 -777 11157 -767
rect 11644 -768 11700 -767
rect 11806 -806 11840 -678
rect 12459 -636 12493 148
rect 13172 86 13206 148
rect 12761 48 13503 86
rect 12761 -76 12795 48
rect 12997 -76 13031 48
rect 13233 -76 13267 48
rect 13469 -76 13503 48
rect 13729 60 13807 66
rect 13729 6 13741 60
rect 13795 6 13807 60
rect 13729 0 13807 6
rect 12755 -88 12801 -76
rect 12755 -464 12761 -88
rect 12795 -464 12801 -88
rect 12755 -476 12801 -464
rect 12873 -88 12919 -76
rect 12873 -464 12879 -88
rect 12913 -464 12919 -88
rect 12873 -476 12919 -464
rect 12991 -88 13037 -76
rect 12991 -464 12997 -88
rect 13031 -464 13037 -88
rect 12991 -476 13037 -464
rect 13109 -88 13155 -76
rect 13109 -464 13115 -88
rect 13149 -464 13155 -88
rect 13109 -476 13155 -464
rect 13227 -88 13273 -76
rect 13227 -464 13233 -88
rect 13267 -464 13273 -88
rect 13227 -476 13273 -464
rect 13345 -88 13391 -76
rect 13345 -464 13351 -88
rect 13385 -464 13391 -88
rect 13345 -476 13391 -464
rect 13463 -88 13509 -76
rect 13463 -464 13469 -88
rect 13503 -464 13509 -88
rect 13463 -476 13509 -464
rect 13875 -635 13909 148
rect 14347 2 14421 68
rect 14487 2 14497 68
rect 14347 -128 14487 -122
rect 14347 -188 14409 -128
rect 14475 -188 14487 -128
rect 14347 -194 14487 -188
rect 13961 -492 14087 -486
rect 13961 -594 13973 -492
rect 14075 -594 14087 -492
rect 13961 -600 14087 -594
rect 13602 -636 13909 -635
rect 12459 -641 12775 -636
rect 13489 -641 13909 -636
rect 12459 -652 12842 -641
rect 12459 -679 12791 -652
rect 3526 -996 3532 -820
rect 3566 -996 3572 -820
rect 3526 -1008 3572 -996
rect 4179 -822 4225 -810
rect 4179 -998 4185 -822
rect 4219 -998 4225 -822
rect 3002 -1208 3048 -1196
rect 2890 -1302 2924 -1208
rect 3414 -1302 3447 -1008
rect 4179 -1010 4225 -998
rect 4297 -822 4343 -810
rect 4297 -998 4303 -822
rect 4337 -998 4343 -822
rect 4297 -1010 4343 -998
rect 4599 -822 4645 -810
rect 2233 -1334 3447 -1302
rect 4302 -1304 4336 -1010
rect 4599 -1198 4605 -822
rect 4639 -1198 4645 -822
rect 4599 -1210 4645 -1198
rect 4717 -822 4763 -810
rect 4717 -1198 4723 -822
rect 4757 -1198 4763 -822
rect 4717 -1210 4763 -1198
rect 4835 -822 4881 -810
rect 4835 -1198 4841 -822
rect 4875 -1198 4881 -822
rect 4835 -1210 4881 -1198
rect 4953 -822 4999 -810
rect 4953 -1198 4959 -822
rect 4993 -1198 4999 -822
rect 4953 -1210 4999 -1198
rect 5071 -822 5117 -810
rect 5071 -1198 5077 -822
rect 5111 -1198 5117 -822
rect 5477 -822 5523 -810
rect 5477 -998 5483 -822
rect 5517 -998 5523 -822
rect 5477 -1010 5523 -998
rect 5595 -822 5641 -810
rect 5595 -998 5601 -822
rect 5635 -998 5641 -822
rect 5595 -1010 5641 -998
rect 6247 -820 6293 -808
rect 6247 -996 6253 -820
rect 6287 -996 6293 -820
rect 6247 -1008 6293 -996
rect 6365 -820 6411 -808
rect 6365 -996 6371 -820
rect 6405 -996 6411 -820
rect 6365 -1008 6411 -996
rect 6667 -820 6713 -808
rect 5071 -1210 5117 -1198
rect 4959 -1304 4993 -1210
rect 5483 -1304 5516 -1010
rect 658 -1358 790 -1336
rect 658 -1416 692 -1358
rect 754 -1416 790 -1358
rect 658 -1421 790 -1416
rect 2726 -1356 2858 -1334
rect 4302 -1336 5516 -1304
rect 6370 -1302 6404 -1008
rect 6667 -1196 6673 -820
rect 6707 -1196 6713 -820
rect 6667 -1208 6713 -1196
rect 6785 -820 6831 -808
rect 6785 -1196 6791 -820
rect 6825 -1196 6831 -820
rect 6785 -1208 6831 -1196
rect 6903 -820 6949 -808
rect 6903 -1196 6909 -820
rect 6943 -1196 6949 -820
rect 6903 -1208 6949 -1196
rect 7021 -820 7067 -808
rect 7021 -1196 7027 -820
rect 7061 -1196 7067 -820
rect 7021 -1208 7067 -1196
rect 7139 -820 7185 -808
rect 7139 -1196 7145 -820
rect 7179 -1196 7185 -820
rect 7545 -820 7591 -808
rect 7545 -996 7551 -820
rect 7585 -996 7591 -820
rect 7545 -1008 7591 -996
rect 7663 -820 7709 -808
rect 7663 -996 7669 -820
rect 7703 -996 7709 -820
rect 7663 -1008 7709 -996
rect 8316 -820 8362 -808
rect 8316 -996 8322 -820
rect 8356 -996 8362 -820
rect 8316 -1008 8362 -996
rect 8434 -820 8480 -808
rect 8434 -996 8440 -820
rect 8474 -996 8480 -820
rect 8434 -1008 8480 -996
rect 8736 -820 8782 -808
rect 7139 -1208 7185 -1196
rect 7027 -1302 7061 -1208
rect 7551 -1302 7584 -1008
rect 6370 -1334 7584 -1302
rect 8439 -1302 8473 -1008
rect 8736 -1196 8742 -820
rect 8776 -1196 8782 -820
rect 8736 -1208 8782 -1196
rect 8854 -820 8900 -808
rect 8854 -1196 8860 -820
rect 8894 -1196 8900 -820
rect 8854 -1208 8900 -1196
rect 8972 -820 9018 -808
rect 8972 -1196 8978 -820
rect 9012 -1196 9018 -820
rect 8972 -1208 9018 -1196
rect 9090 -820 9136 -808
rect 9090 -1196 9096 -820
rect 9130 -1196 9136 -820
rect 9090 -1208 9136 -1196
rect 9208 -820 9254 -808
rect 9208 -1196 9214 -820
rect 9248 -1196 9254 -820
rect 9614 -820 9660 -808
rect 9614 -996 9620 -820
rect 9654 -996 9660 -820
rect 9614 -1008 9660 -996
rect 9732 -820 9778 -808
rect 9732 -996 9738 -820
rect 9772 -996 9778 -820
rect 9732 -1008 9778 -996
rect 10384 -818 10430 -806
rect 10384 -994 10390 -818
rect 10424 -994 10430 -818
rect 10384 -1006 10430 -994
rect 10502 -818 10548 -806
rect 10502 -994 10508 -818
rect 10542 -994 10548 -818
rect 10502 -1006 10548 -994
rect 10804 -818 10850 -806
rect 9208 -1208 9254 -1196
rect 9096 -1302 9130 -1208
rect 9620 -1302 9653 -1008
rect 8439 -1334 9653 -1302
rect 10507 -1300 10541 -1006
rect 10804 -1194 10810 -818
rect 10844 -1194 10850 -818
rect 10804 -1206 10850 -1194
rect 10922 -818 10968 -806
rect 10922 -1194 10928 -818
rect 10962 -1194 10968 -818
rect 10922 -1206 10968 -1194
rect 11040 -818 11086 -806
rect 11040 -1194 11046 -818
rect 11080 -1194 11086 -818
rect 11040 -1206 11086 -1194
rect 11158 -818 11204 -806
rect 11158 -1194 11164 -818
rect 11198 -1194 11204 -818
rect 11158 -1206 11204 -1194
rect 11276 -818 11322 -806
rect 11276 -1194 11282 -818
rect 11316 -1194 11322 -818
rect 11682 -818 11728 -806
rect 11682 -994 11688 -818
rect 11722 -994 11728 -818
rect 11682 -1006 11728 -994
rect 11800 -818 11846 -806
rect 12459 -808 12493 -679
rect 12775 -686 12791 -679
rect 12825 -686 12842 -652
rect 12775 -692 12842 -686
rect 13422 -652 13909 -641
rect 13422 -686 13439 -652
rect 13473 -679 13909 -652
rect 13473 -686 13489 -679
rect 13602 -680 13909 -679
rect 13422 -692 13489 -686
rect 12600 -719 12656 -707
rect 12600 -753 12606 -719
rect 12640 -720 12656 -719
rect 13713 -720 13769 -708
rect 12640 -736 13107 -720
rect 12640 -753 13057 -736
rect 12600 -769 13057 -753
rect 13041 -770 13057 -769
rect 13091 -770 13107 -736
rect 13041 -777 13107 -770
rect 13159 -735 13729 -720
rect 13159 -769 13175 -735
rect 13209 -754 13729 -735
rect 13763 -754 13769 -720
rect 13209 -769 13769 -754
rect 13159 -779 13226 -769
rect 13713 -770 13769 -769
rect 13875 -808 13909 -680
rect 14527 -634 14561 150
rect 15240 88 15274 150
rect 14829 50 15571 88
rect 14829 -74 14863 50
rect 15065 -74 15099 50
rect 15301 -74 15335 50
rect 15537 -74 15571 50
rect 15797 62 15875 68
rect 15797 8 15809 62
rect 15863 8 15875 62
rect 15797 2 15875 8
rect 14823 -86 14869 -74
rect 14823 -462 14829 -86
rect 14863 -462 14869 -86
rect 14823 -474 14869 -462
rect 14941 -86 14987 -74
rect 14941 -462 14947 -86
rect 14981 -462 14987 -86
rect 14941 -474 14987 -462
rect 15059 -86 15105 -74
rect 15059 -462 15065 -86
rect 15099 -462 15105 -86
rect 15059 -474 15105 -462
rect 15177 -86 15223 -74
rect 15177 -462 15183 -86
rect 15217 -462 15223 -86
rect 15177 -474 15223 -462
rect 15295 -86 15341 -74
rect 15295 -462 15301 -86
rect 15335 -462 15341 -86
rect 15295 -474 15341 -462
rect 15413 -86 15459 -74
rect 15413 -462 15419 -86
rect 15453 -462 15459 -86
rect 15413 -474 15459 -462
rect 15531 -86 15577 -74
rect 15531 -462 15537 -86
rect 15571 -462 15577 -86
rect 15531 -474 15577 -462
rect 15943 -633 15977 150
rect 16029 -490 16155 -484
rect 16029 -592 16041 -490
rect 16143 -592 16155 -490
rect 16029 -598 16155 -592
rect 15670 -634 15977 -633
rect 14527 -639 14843 -634
rect 15557 -639 15977 -634
rect 14527 -650 14910 -639
rect 14527 -677 14859 -650
rect 14527 -806 14561 -677
rect 14843 -684 14859 -677
rect 14893 -684 14910 -650
rect 14843 -690 14910 -684
rect 15490 -650 15977 -639
rect 15490 -684 15507 -650
rect 15541 -677 15977 -650
rect 15541 -684 15557 -677
rect 15670 -678 15977 -677
rect 15490 -690 15557 -684
rect 14668 -717 14724 -705
rect 14668 -751 14674 -717
rect 14708 -718 14724 -717
rect 15781 -718 15837 -706
rect 14708 -734 15175 -718
rect 14708 -751 15125 -734
rect 14668 -767 15125 -751
rect 15109 -768 15125 -767
rect 15159 -768 15175 -734
rect 15109 -775 15175 -768
rect 15227 -733 15797 -718
rect 15227 -767 15243 -733
rect 15277 -752 15797 -733
rect 15831 -752 15837 -718
rect 15277 -767 15837 -752
rect 15227 -777 15294 -767
rect 15781 -768 15837 -767
rect 15943 -806 15977 -678
rect 11800 -994 11806 -818
rect 11840 -994 11846 -818
rect 11800 -1006 11846 -994
rect 12453 -820 12499 -808
rect 12453 -996 12459 -820
rect 12493 -996 12499 -820
rect 11276 -1206 11322 -1194
rect 11164 -1300 11198 -1206
rect 11688 -1300 11721 -1006
rect 12453 -1008 12499 -996
rect 12571 -820 12617 -808
rect 12571 -996 12577 -820
rect 12611 -996 12617 -820
rect 12571 -1008 12617 -996
rect 12873 -820 12919 -808
rect 10507 -1332 11721 -1300
rect 12576 -1302 12610 -1008
rect 12873 -1196 12879 -820
rect 12913 -1196 12919 -820
rect 12873 -1208 12919 -1196
rect 12991 -820 13037 -808
rect 12991 -1196 12997 -820
rect 13031 -1196 13037 -820
rect 12991 -1208 13037 -1196
rect 13109 -820 13155 -808
rect 13109 -1196 13115 -820
rect 13149 -1196 13155 -820
rect 13109 -1208 13155 -1196
rect 13227 -820 13273 -808
rect 13227 -1196 13233 -820
rect 13267 -1196 13273 -820
rect 13227 -1208 13273 -1196
rect 13345 -820 13391 -808
rect 13345 -1196 13351 -820
rect 13385 -1196 13391 -820
rect 13751 -820 13797 -808
rect 13751 -996 13757 -820
rect 13791 -996 13797 -820
rect 13751 -1008 13797 -996
rect 13869 -820 13915 -808
rect 13869 -996 13875 -820
rect 13909 -996 13915 -820
rect 13869 -1008 13915 -996
rect 14521 -818 14567 -806
rect 14521 -994 14527 -818
rect 14561 -994 14567 -818
rect 14521 -1006 14567 -994
rect 14639 -818 14685 -806
rect 14639 -994 14645 -818
rect 14679 -994 14685 -818
rect 14639 -1006 14685 -994
rect 14941 -818 14987 -806
rect 13345 -1208 13391 -1196
rect 13233 -1302 13267 -1208
rect 13757 -1302 13790 -1008
rect 2726 -1414 2760 -1356
rect 2822 -1414 2858 -1356
rect 2726 -1419 2858 -1414
rect 4795 -1358 4927 -1336
rect 4795 -1416 4829 -1358
rect 4891 -1416 4927 -1358
rect 4795 -1421 4927 -1416
rect 6863 -1356 6995 -1334
rect 6863 -1414 6897 -1356
rect 6959 -1414 6995 -1356
rect 6863 -1419 6995 -1414
rect 8932 -1356 9064 -1334
rect 8932 -1414 8966 -1356
rect 9028 -1414 9064 -1356
rect 8932 -1419 9064 -1414
rect 11000 -1354 11132 -1332
rect 12576 -1334 13790 -1302
rect 14644 -1300 14678 -1006
rect 14941 -1194 14947 -818
rect 14981 -1194 14987 -818
rect 14941 -1206 14987 -1194
rect 15059 -818 15105 -806
rect 15059 -1194 15065 -818
rect 15099 -1194 15105 -818
rect 15059 -1206 15105 -1194
rect 15177 -818 15223 -806
rect 15177 -1194 15183 -818
rect 15217 -1194 15223 -818
rect 15177 -1206 15223 -1194
rect 15295 -818 15341 -806
rect 15295 -1194 15301 -818
rect 15335 -1194 15341 -818
rect 15295 -1206 15341 -1194
rect 15413 -818 15459 -806
rect 15413 -1194 15419 -818
rect 15453 -1194 15459 -818
rect 15819 -818 15865 -806
rect 15819 -994 15825 -818
rect 15859 -994 15865 -818
rect 15819 -1006 15865 -994
rect 15937 -818 15983 -806
rect 15937 -994 15943 -818
rect 15977 -994 15983 -818
rect 15937 -1006 15983 -994
rect 15413 -1206 15459 -1194
rect 15301 -1300 15335 -1206
rect 15825 -1300 15858 -1006
rect 14644 -1332 15858 -1300
rect 11000 -1412 11034 -1354
rect 11096 -1412 11132 -1354
rect 11000 -1417 11132 -1412
rect 13069 -1356 13201 -1334
rect 13069 -1414 13103 -1356
rect 13165 -1414 13201 -1356
rect 13069 -1419 13201 -1414
rect 15137 -1354 15269 -1332
rect 15137 -1412 15171 -1354
rect 15233 -1412 15269 -1354
rect 15137 -1417 15269 -1412
<< via1 >>
rect 750 858 804 866
rect 750 820 760 858
rect 760 820 798 858
rect 798 820 804 858
rect 2818 860 2872 868
rect 750 812 804 820
rect 2818 822 2828 860
rect 2828 822 2866 860
rect 2866 822 2872 860
rect 2818 814 2872 822
rect 4887 858 4941 866
rect 4887 820 4897 858
rect 4897 820 4935 858
rect 4935 820 4941 858
rect 6955 860 7009 868
rect 4887 812 4941 820
rect 6955 822 6965 860
rect 6965 822 7003 860
rect 7003 822 7009 860
rect 9024 860 9078 868
rect 6955 814 7009 822
rect 9024 822 9034 860
rect 9034 822 9072 860
rect 9072 822 9078 860
rect 11092 862 11146 870
rect 9024 814 9078 822
rect 11092 824 11102 862
rect 11102 824 11140 862
rect 11140 824 11146 862
rect 11092 816 11146 824
rect 13161 860 13215 868
rect 13161 822 13171 860
rect 13171 822 13209 860
rect 13209 822 13215 860
rect 15229 862 15283 870
rect 13161 814 13215 822
rect 15229 824 15239 862
rect 15239 824 15277 862
rect 15277 824 15283 862
rect 15229 816 15283 824
rect -58 -2 8 64
rect 1330 4 1384 58
rect 2010 0 2076 66
rect 3398 6 3452 60
rect 4079 -2 4145 64
rect 5467 4 5521 58
rect 6147 0 6213 66
rect 7535 6 7589 60
rect 8216 0 8282 66
rect 9604 6 9658 60
rect 10284 2 10350 68
rect 11672 8 11726 62
rect 12353 0 12419 66
rect 13741 6 13795 60
rect 14421 2 14487 68
rect 692 -1364 754 -1358
rect 692 -1406 698 -1364
rect 698 -1406 748 -1364
rect 748 -1406 754 -1364
rect 692 -1416 754 -1406
rect 15809 8 15863 62
rect 2760 -1362 2822 -1356
rect 2760 -1404 2766 -1362
rect 2766 -1404 2816 -1362
rect 2816 -1404 2822 -1362
rect 2760 -1414 2822 -1404
rect 4829 -1364 4891 -1358
rect 4829 -1406 4835 -1364
rect 4835 -1406 4885 -1364
rect 4885 -1406 4891 -1364
rect 4829 -1416 4891 -1406
rect 6897 -1362 6959 -1356
rect 6897 -1404 6903 -1362
rect 6903 -1404 6953 -1362
rect 6953 -1404 6959 -1362
rect 6897 -1414 6959 -1404
rect 8966 -1362 9028 -1356
rect 8966 -1404 8972 -1362
rect 8972 -1404 9022 -1362
rect 9022 -1404 9028 -1362
rect 8966 -1414 9028 -1404
rect 11034 -1360 11096 -1354
rect 11034 -1402 11040 -1360
rect 11040 -1402 11090 -1360
rect 11090 -1402 11096 -1360
rect 11034 -1412 11096 -1402
rect 13103 -1362 13165 -1356
rect 13103 -1404 13109 -1362
rect 13109 -1404 13159 -1362
rect 13159 -1404 13165 -1362
rect 13103 -1414 13165 -1404
rect 15171 -1360 15233 -1354
rect 15171 -1402 15177 -1360
rect 15177 -1402 15227 -1360
rect 15227 -1402 15233 -1360
rect 15171 -1412 15233 -1402
<< metal2 >>
rect 738 874 816 884
rect 738 794 816 804
rect 2806 876 2884 886
rect 2806 796 2884 806
rect 4875 874 4953 884
rect 4875 794 4953 804
rect 6943 876 7021 886
rect 6943 796 7021 806
rect 9012 876 9090 886
rect 9012 796 9090 806
rect 11080 878 11158 888
rect 11080 798 11158 808
rect 13149 876 13227 886
rect 13149 796 13227 806
rect 15217 878 15295 888
rect 15217 798 15295 808
rect -64 -2 -58 64
rect 8 58 1384 64
rect 8 4 1330 58
rect 8 -2 1384 4
rect 2004 0 2010 66
rect 2076 60 3452 66
rect 2076 6 3398 60
rect 2076 0 3452 6
rect 4073 -2 4079 64
rect 4145 58 5521 64
rect 4145 4 5467 58
rect 4145 -2 5521 4
rect 6141 0 6147 66
rect 6213 60 7589 66
rect 6213 6 7535 60
rect 6213 0 7589 6
rect 8210 0 8216 66
rect 8282 60 9658 66
rect 8282 6 9604 60
rect 8282 0 9658 6
rect 10278 2 10284 68
rect 10350 62 11726 68
rect 10350 8 11672 62
rect 10350 2 11726 8
rect 12347 0 12353 66
rect 12419 60 13795 66
rect 12419 6 13741 60
rect 12419 0 13795 6
rect 14415 2 14421 68
rect 14487 62 15863 68
rect 14487 8 15809 62
rect 14487 2 15863 8
rect 686 -1356 758 -1346
rect 686 -1436 758 -1426
rect 2754 -1354 2826 -1344
rect 2754 -1434 2826 -1424
rect 4823 -1356 4895 -1346
rect 4823 -1436 4895 -1426
rect 6891 -1354 6963 -1344
rect 6891 -1434 6963 -1424
rect 8960 -1354 9032 -1344
rect 8960 -1434 9032 -1424
rect 11028 -1352 11100 -1342
rect 11028 -1432 11100 -1422
rect 13097 -1354 13169 -1344
rect 13097 -1434 13169 -1424
rect 15165 -1352 15237 -1342
rect 15165 -1432 15237 -1422
<< via2 >>
rect 738 866 816 874
rect 738 812 750 866
rect 750 812 804 866
rect 804 812 816 866
rect 738 804 816 812
rect 2806 868 2884 876
rect 2806 814 2818 868
rect 2818 814 2872 868
rect 2872 814 2884 868
rect 2806 806 2884 814
rect 4875 866 4953 874
rect 4875 812 4887 866
rect 4887 812 4941 866
rect 4941 812 4953 866
rect 4875 804 4953 812
rect 6943 868 7021 876
rect 6943 814 6955 868
rect 6955 814 7009 868
rect 7009 814 7021 868
rect 6943 806 7021 814
rect 9012 868 9090 876
rect 9012 814 9024 868
rect 9024 814 9078 868
rect 9078 814 9090 868
rect 9012 806 9090 814
rect 11080 870 11158 878
rect 11080 816 11092 870
rect 11092 816 11146 870
rect 11146 816 11158 870
rect 11080 808 11158 816
rect 13149 868 13227 876
rect 13149 814 13161 868
rect 13161 814 13215 868
rect 13215 814 13227 868
rect 13149 806 13227 814
rect 15217 870 15295 878
rect 15217 816 15229 870
rect 15229 816 15283 870
rect 15283 816 15295 870
rect 15217 808 15295 816
rect 686 -1358 758 -1356
rect 686 -1416 692 -1358
rect 692 -1416 754 -1358
rect 754 -1416 758 -1358
rect 686 -1426 758 -1416
rect 2754 -1356 2826 -1354
rect 2754 -1414 2760 -1356
rect 2760 -1414 2822 -1356
rect 2822 -1414 2826 -1356
rect 2754 -1424 2826 -1414
rect 4823 -1358 4895 -1356
rect 4823 -1416 4829 -1358
rect 4829 -1416 4891 -1358
rect 4891 -1416 4895 -1358
rect 4823 -1426 4895 -1416
rect 6891 -1356 6963 -1354
rect 6891 -1414 6897 -1356
rect 6897 -1414 6959 -1356
rect 6959 -1414 6963 -1356
rect 6891 -1424 6963 -1414
rect 8960 -1356 9032 -1354
rect 8960 -1414 8966 -1356
rect 8966 -1414 9028 -1356
rect 9028 -1414 9032 -1356
rect 8960 -1424 9032 -1414
rect 11028 -1354 11100 -1352
rect 11028 -1412 11034 -1354
rect 11034 -1412 11096 -1354
rect 11096 -1412 11100 -1354
rect 11028 -1422 11100 -1412
rect 13097 -1356 13169 -1354
rect 13097 -1414 13103 -1356
rect 13103 -1414 13165 -1356
rect 13165 -1414 13169 -1356
rect 13097 -1424 13169 -1414
rect 15165 -1354 15237 -1352
rect 15165 -1412 15171 -1354
rect 15171 -1412 15233 -1354
rect 15233 -1412 15237 -1354
rect 15165 -1422 15237 -1412
<< metal3 >>
rect 668 876 882 880
rect 668 804 738 876
rect 814 874 882 876
rect 816 804 882 874
rect 2736 878 2950 882
rect 2736 806 2806 878
rect 2882 876 2950 878
rect 2884 806 2950 876
rect 2736 804 2950 806
rect 4805 876 5019 880
rect 4805 804 4875 876
rect 4951 874 5019 876
rect 4953 804 5019 874
rect 6873 878 7087 882
rect 6873 806 6943 878
rect 7019 876 7087 878
rect 7021 806 7087 876
rect 6873 804 7087 806
rect 8942 878 9156 882
rect 8942 806 9012 878
rect 9088 876 9156 878
rect 9090 806 9156 876
rect 11010 880 11224 884
rect 11010 808 11080 880
rect 11156 878 11224 880
rect 11158 808 11224 878
rect 11010 806 11224 808
rect 13079 878 13293 882
rect 13079 806 13149 878
rect 13225 876 13293 878
rect 13227 806 13293 876
rect 15147 880 15361 884
rect 15147 808 15217 880
rect 15293 878 15361 880
rect 15295 808 15361 878
rect 15147 806 15361 808
rect 8942 804 9156 806
rect 668 802 882 804
rect 728 799 826 802
rect 2796 801 2894 804
rect 4805 802 5019 804
rect 4865 799 4963 802
rect 6933 801 7031 804
rect 9002 801 9100 804
rect 11070 803 11168 806
rect 13079 804 13293 806
rect 13139 801 13237 804
rect 15207 803 15305 806
rect 10990 -1338 11142 -1336
rect 15127 -1338 15279 -1336
rect 2716 -1340 2868 -1338
rect 6853 -1340 7005 -1338
rect 8922 -1340 9074 -1338
rect 648 -1342 800 -1340
rect 646 -1346 800 -1342
rect 646 -1434 676 -1346
rect 770 -1434 800 -1346
rect 646 -1440 800 -1434
rect 2714 -1344 2868 -1340
rect 4785 -1342 4937 -1340
rect 2714 -1432 2744 -1344
rect 2838 -1432 2868 -1344
rect 2714 -1438 2868 -1432
rect 648 -1450 800 -1440
rect 2716 -1448 2868 -1438
rect 4783 -1346 4937 -1342
rect 4783 -1434 4813 -1346
rect 4907 -1434 4937 -1346
rect 4783 -1440 4937 -1434
rect 6851 -1344 7005 -1340
rect 6851 -1432 6881 -1344
rect 6975 -1432 7005 -1344
rect 6851 -1438 7005 -1432
rect 8920 -1344 9074 -1340
rect 8920 -1432 8950 -1344
rect 9044 -1432 9074 -1344
rect 8920 -1438 9074 -1432
rect 10988 -1342 11142 -1338
rect 13059 -1340 13211 -1338
rect 10988 -1430 11018 -1342
rect 11112 -1430 11142 -1342
rect 10988 -1436 11142 -1430
rect 4785 -1450 4937 -1440
rect 6853 -1448 7005 -1438
rect 8922 -1448 9074 -1438
rect 10990 -1446 11142 -1436
rect 13057 -1344 13211 -1340
rect 13057 -1432 13087 -1344
rect 13181 -1432 13211 -1344
rect 13057 -1438 13211 -1432
rect 15125 -1342 15279 -1338
rect 15125 -1430 15155 -1342
rect 15249 -1430 15279 -1342
rect 15125 -1436 15279 -1430
rect 13059 -1448 13211 -1438
rect 15127 -1446 15279 -1436
<< via3 >>
rect 738 874 814 876
rect 738 810 814 874
rect 2806 876 2882 878
rect 2806 812 2882 876
rect 4875 874 4951 876
rect 4875 810 4951 874
rect 6943 876 7019 878
rect 6943 812 7019 876
rect 9012 876 9088 878
rect 9012 812 9088 876
rect 11080 878 11156 880
rect 11080 814 11156 878
rect 13149 876 13225 878
rect 13149 812 13225 876
rect 15217 878 15293 880
rect 15217 814 15293 878
rect 676 -1356 770 -1346
rect 676 -1426 686 -1356
rect 686 -1426 758 -1356
rect 758 -1426 770 -1356
rect 676 -1434 770 -1426
rect 2744 -1354 2838 -1344
rect 2744 -1424 2754 -1354
rect 2754 -1424 2826 -1354
rect 2826 -1424 2838 -1354
rect 2744 -1432 2838 -1424
rect 4813 -1356 4907 -1346
rect 4813 -1426 4823 -1356
rect 4823 -1426 4895 -1356
rect 4895 -1426 4907 -1356
rect 4813 -1434 4907 -1426
rect 6881 -1354 6975 -1344
rect 6881 -1424 6891 -1354
rect 6891 -1424 6963 -1354
rect 6963 -1424 6975 -1354
rect 6881 -1432 6975 -1424
rect 8950 -1354 9044 -1344
rect 8950 -1424 8960 -1354
rect 8960 -1424 9032 -1354
rect 9032 -1424 9044 -1354
rect 8950 -1432 9044 -1424
rect 11018 -1352 11112 -1342
rect 11018 -1422 11028 -1352
rect 11028 -1422 11100 -1352
rect 11100 -1422 11112 -1352
rect 11018 -1430 11112 -1422
rect 13087 -1354 13181 -1344
rect 13087 -1424 13097 -1354
rect 13097 -1424 13169 -1354
rect 13169 -1424 13181 -1354
rect 13087 -1432 13181 -1424
rect 15155 -1352 15249 -1342
rect 15155 -1422 15165 -1352
rect 15165 -1422 15237 -1352
rect 15237 -1422 15249 -1352
rect 15155 -1430 15249 -1422
<< metal4 >>
rect -106 880 16132 1012
rect -106 878 11080 880
rect -106 876 2806 878
rect -106 810 738 876
rect 814 812 2806 876
rect 2882 876 6943 878
rect 2882 812 4875 876
rect 814 810 4875 812
rect 4951 812 6943 876
rect 7019 812 9012 878
rect 9088 814 11080 878
rect 11156 878 15217 880
rect 11156 814 13149 878
rect 9088 812 13149 814
rect 13225 814 15217 878
rect 15293 814 16132 880
rect 13225 812 16132 814
rect 4951 810 16132 812
rect -106 768 16132 810
rect 2118 -1340 3482 -1338
rect 6255 -1340 7619 -1338
rect 8324 -1340 9688 -1338
rect 10392 -1340 11756 -1336
rect 12461 -1340 13825 -1338
rect 14529 -1340 16080 -1336
rect -10 -1342 16080 -1340
rect -10 -1344 11018 -1342
rect -10 -1346 2744 -1344
rect -10 -1434 676 -1346
rect 770 -1432 2744 -1346
rect 2838 -1346 6881 -1344
rect 2838 -1432 4813 -1346
rect 770 -1434 4813 -1432
rect 4907 -1432 6881 -1346
rect 6975 -1432 8950 -1344
rect 9044 -1430 11018 -1344
rect 11112 -1344 15155 -1342
rect 11112 -1430 13087 -1344
rect 9044 -1432 13087 -1430
rect 13181 -1430 15155 -1344
rect 15249 -1430 16080 -1342
rect 13181 -1432 16080 -1430
rect 4907 -1434 16080 -1432
rect -10 -1530 16080 -1434
<< labels >>
flabel metal4 7782 -1524 8178 -1430 1 FreeSerif 1120 0 0 0 VSS
port 1 n
flabel metal4 7782 776 8182 898 1 FreeSerif 1120 0 0 0 VDD
port 2 n
flabel metal1 -132 -196 -92 -146 1 FreeSerif 480 0 0 0 A[0]
port 3 n
flabel metal1 1938 -192 1978 -142 1 FreeSerif 480 0 0 0 A[1]
port 4 n
flabel metal1 4008 -194 4048 -144 1 FreeSerif 480 0 0 0 A[2]
port 5 n
flabel metal1 6074 -194 6114 -144 1 FreeSerif 480 0 0 0 A[3]
port 6 n
flabel metal1 8144 -194 8184 -144 1 FreeSerif 480 0 0 0 A[4]
port 7 n
flabel metal1 10212 -192 10252 -142 1 FreeSerif 480 0 0 0 A[5]
port 8 n
flabel metal1 12280 -194 12320 -144 1 FreeSerif 480 0 0 0 A[6]
port 9 n
flabel metal1 14348 -194 14388 -144 1 FreeSerif 480 0 0 0 A[7]
port 10 n
flabel metal1 -130 0 -90 50 1 FreeSerif 480 0 0 0 B[0]
port 11 n
flabel metal1 1938 2 1978 52 1 FreeSerif 480 0 0 0 B[1]
port 12 n
flabel metal1 4008 0 4048 50 1 FreeSerif 480 0 0 0 B[2]
port 13 n
flabel metal1 6074 2 6114 52 1 FreeSerif 480 0 0 0 B[3]
port 14 n
flabel metal1 8144 2 8184 52 1 FreeSerif 480 0 0 0 B[4]
port 15 n
flabel metal1 10212 2 10252 52 1 FreeSerif 480 0 0 0 B[5]
port 16 n
flabel metal1 12280 2 12320 52 1 FreeSerif 480 0 0 0 B[6]
port 17 n
flabel metal1 14350 4 14390 54 1 FreeSerif 480 0 0 0 B[7]
port 18 n
flabel metal1 1570 -570 1676 -510 1 FreeSerif 560 0 0 0 Y[0]
port 19 n
flabel metal1 3632 -568 3738 -508 1 FreeSerif 560 0 0 0 Y[1]
port 20 n
flabel metal1 5702 -568 5808 -508 1 FreeSerif 560 0 0 0 Y[2]
port 21 n
flabel metal1 7762 -572 7868 -512 1 FreeSerif 560 0 0 0 Y[3]
port 22 n
flabel metal1 9844 -564 9950 -504 1 FreeSerif 560 0 0 0 Y[4]
port 23 n
flabel metal1 11910 -562 12016 -502 1 FreeSerif 560 0 0 0 Y[5]
port 24 n
flabel metal1 13978 -568 14084 -508 1 FreeSerif 560 0 0 0 Y[6]
port 25 n
flabel metal1 16044 -562 16150 -502 1 FreeSerif 560 0 0 0 Y[7]
port 26 n
<< end >>
