* NGSPICE file created from logic_inverter_pex.ext - technology: sky130B

.subckt logic_inverter A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2]
+ Y[3] Y[4] Y[5] Y[6] Y[7] VSS VDD
X0 VDD.t35 A[5].t0 Y[5].t3 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1 Y[3].t3 A[3].t0 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2 Y[6].t3 A[6].t0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 VDD.t43 A[0].t0 Y[0].t3 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4 Y[1].t3 A[1].t0 VSS.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 Y[3].t2 A[3].t1 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6 Y[4].t2 A[4].t0 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7 Y[0].t0 A[0].t1 VSS.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8 Y[4].t3 A[4].t1 VSS.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X9 VDD.t25 A[6].t1 Y[6].t2 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10 Y[0].t2 A[0].t2 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X11 Y[0].t1 A[0].t3 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X12 Y[1].t2 A[1].t1 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X13 Y[5].t0 A[5].t1 VSS.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X14 Y[7].t2 A[7].t0 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X15 VDD.t19 A[3].t2 Y[3].t1 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X16 Y[4].t1 A[4].t2 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X17 Y[5].t2 A[5].t2 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X18 Y[5].t1 A[5].t3 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X19 Y[6].t1 A[6].t2 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X20 VDD.t45 A[2].t0 Y[2].t2 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X21 VDD.t29 A[7].t1 Y[7].t1 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X22 Y[1].t1 A[1].t2 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X23 Y[2].t1 A[2].t1 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X24 VDD.t41 A[4].t3 Y[4].t0 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X25 Y[7].t0 A[7].t2 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 VDD.t23 A[1].t3 Y[1].t0 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X27 Y[3].t0 A[3].t3 VSS.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 Y[2].t0 A[2].t2 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X29 Y[2].t3 A[2].t3 VSS.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X30 Y[7].t3 A[7].t3 VSS.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X31 Y[6].t0 A[6].t3 VSS.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 A[5].n0 A[5].t3 185.301
R1 A[5].n0 A[5].t2 185.301
R2 A[5].n1 A[5].t1 140.583
R3 A[5].n0 A[5].t0 107.646
R4 A[5].n1 A[5].n0 61.856
R5 A[5] A[5].n1 13.908
R6 Y[5].n1 Y[5].n0 197.272
R7 Y[5].n1 Y[5].t1 28.568
R8 Y[5].n0 Y[5].t3 28.565
R9 Y[5].n0 Y[5].t2 28.565
R10 Y[5] Y[5].t0 18.14
R11 Y[5] Y[5].n2 0.593
R12 Y[5].n2 Y[5] 0.593
R13 Y[5] Y[5].n1 0.49
R14 Y[5].n2 Y[5] 0.078
R15 Y[5].n2 Y[5] 0.049
R16 Y[5].n2 Y[5] 0.049
R17 VDD.n33 VDD.t16 174.172
R18 VDD.n40 VDD.t46 173.061
R19 VDD.n47 VDD.t2 172.51
R20 VDD.n0 VDD.t8 172.51
R21 VDD.n6 VDD.t30 172.51
R22 VDD.n12 VDD.t10 172.51
R23 VDD.n18 VDD.t4 172.51
R24 VDD.n30 VDD.t12 172.51
R25 VDD.n32 VDD.t20 170.712
R26 VDD.n39 VDD.t36 169.626
R27 VDD.n29 VDD.t6 169.089
R28 VDD.n46 VDD.t14 169.088
R29 VDD.n1 VDD.t38 169.088
R30 VDD.n7 VDD.t32 169.088
R31 VDD.n13 VDD.t0 169.088
R32 VDD.n19 VDD.t26 169.088
R33 VDD.n50 VDD.t15 29.208
R34 VDD.n4 VDD.t39 29.208
R35 VDD.n10 VDD.t33 29.208
R36 VDD.n16 VDD.t1 29.208
R37 VDD.n22 VDD.t27 29.208
R38 VDD.n28 VDD.t7 29.208
R39 VDD.n43 VDD.t37 29.202
R40 VDD.n36 VDD.t21 29.191
R41 VDD.n35 VDD.t17 28.565
R42 VDD.n35 VDD.t23 28.565
R43 VDD.n42 VDD.t47 28.565
R44 VDD.n42 VDD.t45 28.565
R45 VDD.n49 VDD.t3 28.565
R46 VDD.n49 VDD.t19 28.565
R47 VDD.n3 VDD.t9 28.565
R48 VDD.n3 VDD.t41 28.565
R49 VDD.n9 VDD.t31 28.565
R50 VDD.n9 VDD.t35 28.565
R51 VDD.n15 VDD.t11 28.565
R52 VDD.n15 VDD.t25 28.565
R53 VDD.n21 VDD.t5 28.565
R54 VDD.n21 VDD.t29 28.565
R55 VDD.n27 VDD.t13 28.565
R56 VDD.n27 VDD.t43 28.565
R57 VDD.n50 VDD.n49 0.386
R58 VDD.n4 VDD.n3 0.386
R59 VDD.n10 VDD.n9 0.386
R60 VDD.n16 VDD.n15 0.386
R61 VDD.n22 VDD.n21 0.386
R62 VDD.n28 VDD.n27 0.386
R63 VDD.n43 VDD.n42 0.38
R64 VDD.n36 VDD.n35 0.369
R65 VDD.n48 VDD.n47 0.285
R66 VDD.n31 VDD.n30 0.285
R67 VDD.n41 VDD.n40 0.285
R68 VDD.n34 VDD.n33 0.285
R69 VDD.t42 VDD.n29 0.244
R70 VDD.t22 VDD.n32 0.244
R71 VDD.t44 VDD.n39 0.243
R72 VDD.t18 VDD.n46 0.243
R73 VDD.n1 VDD.t40 0.243
R74 VDD.n7 VDD.t34 0.243
R75 VDD.n13 VDD.t24 0.243
R76 VDD.n19 VDD.t28 0.243
R77 VDD.n24 VDD.n23 0.183
R78 VDD.n38 VDD.n31 0.182
R79 VDD.n52 VDD.n45 0.182
R80 VDD.n25 VDD.n24 0.181
R81 VDD.n26 VDD.n25 0.181
R82 VDD.n45 VDD.n38 0.181
R83 VDD VDD.n26 0.098
R84 VDD.n37 VDD.n36 0.079
R85 VDD.n44 VDD.n43 0.079
R86 VDD.n51 VDD.n50 0.079
R87 VDD.n5 VDD.n4 0.079
R88 VDD.n11 VDD.n10 0.079
R89 VDD.n17 VDD.n16 0.079
R90 VDD.n23 VDD.n22 0.079
R91 VDD.n31 VDD.n28 0.078
R92 VDD VDD.n52 0.036
R93 VDD.n33 VDD.t22 0.021
R94 VDD.n40 VDD.t44 0.021
R95 VDD.n47 VDD.t18 0.021
R96 VDD.t40 VDD.n0 0.021
R97 VDD.t34 VDD.n6 0.021
R98 VDD.t24 VDD.n12 0.021
R99 VDD.t28 VDD.n18 0.021
R100 VDD.n30 VDD.t42 0.021
R101 VDD.n48 VDD.n46 0.003
R102 VDD.n2 VDD.n1 0.003
R103 VDD.n8 VDD.n7 0.003
R104 VDD.n14 VDD.n13 0.003
R105 VDD.n20 VDD.n19 0.003
R106 VDD.n41 VDD.n39 0.003
R107 VDD.n34 VDD.n32 0.003
R108 VDD.n31 VDD.n29 0.002
R109 VDD.n38 VDD.n37 0.001
R110 VDD.n37 VDD.n34 0.001
R111 VDD.n45 VDD.n44 0.001
R112 VDD.n44 VDD.n41 0.001
R113 VDD.n52 VDD.n51 0.001
R114 VDD.n51 VDD.n48 0.001
R115 VDD.n26 VDD.n5 0.001
R116 VDD.n5 VDD.n2 0.001
R117 VDD.n25 VDD.n11 0.001
R118 VDD.n11 VDD.n8 0.001
R119 VDD.n24 VDD.n17 0.001
R120 VDD.n17 VDD.n14 0.001
R121 VDD.n23 VDD.n20 0.001
R122 A[3].n0 A[3].t0 185.301
R123 A[3].n0 A[3].t1 185.301
R124 A[3].n1 A[3].t3 140.583
R125 A[3].n0 A[3].t2 107.646
R126 A[3].n1 A[3].n0 61.856
R127 A[3] A[3].n1 13.908
R128 Y[3].n1 Y[3].n0 197.272
R129 Y[3].n1 Y[3].t3 28.568
R130 Y[3].n0 Y[3].t1 28.565
R131 Y[3].n0 Y[3].t2 28.565
R132 Y[3] Y[3].t0 18.14
R133 Y[3] Y[3].n2 0.593
R134 Y[3].n2 Y[3] 0.593
R135 Y[3] Y[3].n1 0.49
R136 Y[3].n2 Y[3] 0.078
R137 Y[3].n2 Y[3] 0.049
R138 Y[3].n2 Y[3] 0.049
R139 A[6].n0 A[6].t2 185.301
R140 A[6].n0 A[6].t0 185.301
R141 A[6].n1 A[6].t3 137.369
R142 A[6].n0 A[6].t1 107.646
R143 A[6].n1 A[6].n0 61.856
R144 A[6] A[6].n1 13.908
R145 Y[6].n1 Y[6].n0 197.272
R146 Y[6].n1 Y[6].t1 28.568
R147 Y[6].n0 Y[6].t2 28.565
R148 Y[6].n0 Y[6].t3 28.565
R149 Y[6] Y[6].t0 18.129
R150 Y[6] Y[6].n2 0.593
R151 Y[6].n2 Y[6] 0.593
R152 Y[6] Y[6].n1 0.49
R153 Y[6].n2 Y[6] 0.078
R154 Y[6].n2 Y[6] 0.049
R155 Y[6].n2 Y[6] 0.049
R156 A[0].n0 A[0].t3 185.301
R157 A[0].n0 A[0].t2 185.301
R158 A[0].n1 A[0].t1 140.583
R159 A[0].n0 A[0].t0 107.646
R160 A[0].n1 A[0].n0 61.856
R161 A[0] A[0].n1 13.908
R162 Y[0].n1 Y[0].n0 197.272
R163 Y[0].n1 Y[0].t1 28.568
R164 Y[0].n0 Y[0].t3 28.565
R165 Y[0].n0 Y[0].t2 28.565
R166 Y[0] Y[0].t0 18.14
R167 Y[0] Y[0].n2 0.593
R168 Y[0].n2 Y[0] 0.593
R169 Y[0] Y[0].n1 0.49
R170 Y[0].n2 Y[0] 0.078
R171 Y[0].n2 Y[0] 0.049
R172 Y[0].n2 Y[0] 0.049
R173 A[1].n0 A[1].t1 190.121
R174 A[1].n0 A[1].t2 190.121
R175 A[1].n1 A[1].t0 137.369
R176 A[1].n0 A[1].t3 112.466
R177 A[1].n1 A[1].n0 61.856
R178 A[1] A[1].n1 13.908
R179 VSS.n0 VSS.t1 18.151
R180 VSS.n3 VSS.t0 18.141
R181 VSS.n3 VSS.t7 17.97
R182 VSS.n0 VSS.t3 17.97
R183 VSS.n4 VSS.t6 17.959
R184 VSS.n5 VSS.t4 17.959
R185 VSS.n2 VSS.t2 17.959
R186 VSS.n1 VSS.t5 17.959
R187 VSS.n5 VSS.n4 0.182
R188 VSS.n1 VSS.n0 0.181
R189 VSS.n2 VSS.n1 0.181
R190 VSS.n4 VSS.n3 0.181
R191 VSS VSS.n2 0.08
R192 VSS VSS.n5 0.052
R193 Y[1].n1 Y[1].n0 192.754
R194 Y[1].n1 Y[1].t2 28.568
R195 Y[1].n0 Y[1].t0 28.565
R196 Y[1].n0 Y[1].t1 28.565
R197 Y[1] Y[1].t3 18.129
R198 Y[1] Y[1].n2 0.593
R199 Y[1].n2 Y[1] 0.593
R200 Y[1] Y[1].n1 0.505
R201 Y[1].n2 Y[1] 0.078
R202 Y[1].n2 Y[1] 0.049
R203 Y[1].n2 Y[1] 0.049
R204 A[4].n0 A[4].t0 185.301
R205 A[4].n0 A[4].t2 185.301
R206 A[4].n1 A[4].t1 140.583
R207 A[4].n0 A[4].t3 107.646
R208 A[4].n1 A[4].n0 61.856
R209 A[4] A[4].n1 13.908
R210 Y[4].n1 Y[4].n0 197.272
R211 Y[4].n1 Y[4].t2 28.568
R212 Y[4].n0 Y[4].t0 28.565
R213 Y[4].n0 Y[4].t1 28.565
R214 Y[4] Y[4].t3 18.14
R215 Y[4] Y[4].n2 0.593
R216 Y[4].n2 Y[4] 0.593
R217 Y[4] Y[4].n1 0.49
R218 Y[4].n2 Y[4] 0.078
R219 Y[4].n2 Y[4] 0.049
R220 Y[4].n2 Y[4] 0.049
R221 A[7].n0 A[7].t2 185.301
R222 A[7].n0 A[7].t0 185.301
R223 A[7].n1 A[7].t3 137.369
R224 A[7].n0 A[7].t1 107.646
R225 A[7].n1 A[7].n0 61.856
R226 A[7] A[7].n1 13.908
R227 Y[7].n1 Y[7].n0 197.272
R228 Y[7].n1 Y[7].t0 28.568
R229 Y[7].n0 Y[7].t1 28.565
R230 Y[7].n0 Y[7].t2 28.565
R231 Y[7] Y[7].t3 18.129
R232 Y[7] Y[7].n2 0.593
R233 Y[7].n2 Y[7] 0.593
R234 Y[7] Y[7].n1 0.49
R235 Y[7].n2 Y[7] 0.078
R236 Y[7].n2 Y[7] 0.049
R237 Y[7].n2 Y[7] 0.049
R238 A[2].n0 A[2].t1 186.908
R239 A[2].n0 A[2].t2 186.908
R240 A[2].n1 A[2].t3 140.583
R241 A[2].n0 A[2].t0 109.253
R242 A[2].n1 A[2].n0 61.856
R243 A[2] A[2].n1 13.908
R244 Y[2].n1 Y[2].n0 195.766
R245 Y[2].n1 Y[2].t1 28.568
R246 Y[2].n0 Y[2].t2 28.565
R247 Y[2].n0 Y[2].t0 28.565
R248 Y[2] Y[2].t3 18.14
R249 Y[2] Y[2].n2 0.593
R250 Y[2].n2 Y[2] 0.593
R251 Y[2] Y[2].n1 0.496
R252 Y[2].n2 Y[2] 0.078
R253 Y[2].n2 Y[2] 0.049
R254 Y[2].n2 Y[2] 0.049
C0 A[5] Y[4] 0.02fF
C1 A[4] Y[5] 0.01fF
C2 A[4] Y[4] 0.06fF
C3 A[3] Y[5] 0.00fF
C4 A[5] Y[3] 0.00fF
C5 A[6] A[7] 0.01fF
C6 A[5] A[7] 0.00fF
C7 A[3] Y[4] 0.01fF
C8 A[4] Y[3] 0.02fF
C9 Y[4] Y[2] 0.00fF
C10 A[5] A[6] 0.01fF
C11 A[3] Y[3] 0.06fF
C12 Y[4] A[2] 0.00fF
C13 Y[3] Y[2] 0.02fF
C14 A[4] A[6] 0.00fF
C15 Y[3] A[2] 0.01fF
C16 A[4] A[5] 0.01fF
C17 Y[7] VDD 0.90fF
C18 Y[3] Y[1] 0.00fF
C19 A[3] A[5] 0.00fF
C20 Y[6] VDD 0.96fF
C21 A[3] A[4] 0.01fF
C22 Y[3] A[1] 0.00fF
C23 A[4] Y[2] 0.00fF
C24 Y[5] VDD 0.97fF
C25 A[4] A[2] 0.00fF
C26 A[3] Y[2] 0.02fF
C27 Y[4] VDD 0.97fF
C28 A[3] A[2] 0.01fF
C29 Y[3] VDD 0.97fF
C30 A[2] Y[2] 0.06fF
C31 A[7] VDD 0.20fF
C32 A[3] Y[1] 0.00fF
C33 Y[1] Y[2] 0.02fF
C34 A[6] VDD 0.21fF
C35 Y[1] A[2] 0.02fF
C36 Y[0] Y[2] 0.00fF
C37 A[5] VDD 0.21fF
C38 A[3] A[1] 0.00fF
C39 Y[0] A[2] 0.00fF
C40 A[1] Y[2] 0.01fF
C41 A[4] VDD 0.21fF
C42 A[1] A[2] 0.01fF
C43 A[0] Y[2] 0.00fF
C44 Y[0] Y[1] 0.02fF
C45 A[3] VDD 0.21fF
C46 A[1] Y[1] 0.06fF
C47 VDD Y[2] 0.96fF
C48 A[0] A[2] 0.00fF
C49 A[0] Y[1] 0.01fF
C50 VDD A[2] 0.21fF
C51 A[1] Y[0] 0.02fF
C52 VDD Y[1] 0.97fF
C53 A[0] Y[0] 0.07fF
C54 A[0] A[1] 0.01fF
C55 VDD Y[0] 0.96fF
C56 VDD A[1] 0.21fF
C57 VDD A[0] 0.20fF
C58 Y[6] Y[7] 0.02fF
C59 Y[5] Y[7] 0.00fF
C60 Y[5] Y[6] 0.02fF
C61 Y[4] Y[6] 0.00fF
C62 Y[4] Y[5] 0.02fF
C63 A[7] Y[7] 0.06fF
C64 A[6] Y[7] 0.01fF
C65 A[7] Y[6] 0.02fF
C66 Y[3] Y[5] 0.00fF
C67 A[7] Y[5] 0.00fF
C68 A[5] Y[7] 0.00fF
C69 Y[3] Y[4] 0.02fF
C70 A[6] Y[6] 0.06fF
C71 A[6] Y[5] 0.02fF
C72 A[5] Y[6] 0.01fF
C73 A[4] Y[6] 0.00fF
C74 A[5] Y[5] 0.06fF
C75 A[6] Y[4] 0.00fF
.ends

