magic
tech sky130B
magscale 1 2
timestamp 1735941024
<< nwell >>
rect 1455 4932 1742 4933
rect 2602 4932 2837 4933
rect -1027 4878 -787 4879
rect -1030 4645 -787 4878
rect -1030 4463 -786 4645
rect 1452 4535 1742 4932
rect 2429 4539 2911 4932
rect -1468 4139 -276 4463
rect 857 4068 1742 4535
rect 857 4015 1743 4068
rect 1999 4015 2911 4539
rect 857 4011 1744 4015
rect 1286 3726 1744 4011
rect 2429 3756 2911 4015
rect 1286 3428 1770 3726
rect 2428 3432 2912 3756
rect -1013 3228 -773 3229
rect -1016 2995 -773 3228
rect -1016 2813 -772 2995
rect -1454 2489 -262 2813
rect 2698 2396 2926 2886
rect 9 2196 1332 2396
rect 2392 2196 3230 2396
rect 9 1872 3713 2196
rect -1018 1624 -778 1625
rect -1021 1391 -778 1624
rect -1021 1209 -777 1391
rect -1459 885 -267 1209
rect 437 1179 1275 1872
rect 2335 1179 3173 1872
<< nmos >>
rect -1137 3564 -1077 3964
rect -1019 3564 -959 3964
rect -784 3764 -724 3964
rect 861 3490 921 3690
rect 979 3490 1039 3690
rect 1097 3490 1157 3690
rect 2003 3494 2063 3694
rect 2121 3494 2181 3694
rect 2239 3494 2299 3694
rect -1123 1914 -1063 2314
rect -1005 1914 -945 2314
rect -770 2114 -710 2314
rect -1128 310 -1068 710
rect -1010 310 -950 710
rect -775 510 -715 710
rect 229 709 289 909
rect 649 509 709 909
rect 767 509 827 909
rect 885 509 945 909
rect 1003 509 1063 909
rect 1527 709 1587 909
rect 2127 709 2187 909
rect 2547 509 2607 909
rect 2665 509 2725 909
rect 2783 509 2843 909
rect 2901 509 2961 909
rect 3425 709 3485 909
<< pmos >>
rect -1374 4201 -1314 4401
rect -1256 4201 -1196 4401
rect -1138 4201 -1078 4401
rect -1020 4201 -960 4401
rect -902 4201 -842 4401
rect -784 4201 -724 4401
rect -666 4201 -606 4401
rect -548 4201 -488 4401
rect -430 4201 -370 4401
rect 951 4073 1011 4473
rect 1069 4073 1129 4473
rect 1187 4073 1247 4473
rect 1305 4073 1365 4473
rect 1423 4073 1483 4473
rect 1541 4073 1601 4473
rect 2093 4077 2153 4477
rect 2211 4077 2271 4477
rect 2329 4077 2389 4477
rect 2447 4077 2507 4477
rect 2565 4077 2625 4477
rect 2683 4077 2743 4477
rect 1380 3490 1440 3690
rect 1498 3490 1558 3690
rect 1616 3490 1676 3690
rect 2522 3494 2582 3694
rect 2640 3494 2700 3694
rect 2758 3494 2818 3694
rect -1360 2551 -1300 2751
rect -1242 2551 -1182 2751
rect -1124 2551 -1064 2751
rect -1006 2551 -946 2751
rect -888 2551 -828 2751
rect -770 2551 -710 2751
rect -652 2551 -592 2751
rect -534 2551 -474 2751
rect -416 2551 -356 2751
rect 104 1934 164 2134
rect 222 1934 282 2134
rect 340 1934 400 2134
rect 588 1934 648 2334
rect 706 1934 766 2334
rect 824 1934 884 2334
rect 942 1934 1002 2334
rect 1060 1934 1120 2334
rect 1178 1934 1238 2334
rect 1425 1934 1485 2134
rect 1543 1934 1603 2134
rect 1661 1934 1721 2134
rect 2002 1934 2062 2134
rect 2120 1934 2180 2134
rect 2238 1934 2298 2134
rect 2486 1934 2546 2334
rect 2604 1934 2664 2334
rect 2722 1934 2782 2334
rect 2840 1934 2900 2334
rect 2958 1934 3018 2334
rect 3076 1934 3136 2334
rect 3323 1934 3383 2134
rect 3441 1934 3501 2134
rect 3559 1934 3619 2134
rect -1365 947 -1305 1147
rect -1247 947 -1187 1147
rect -1129 947 -1069 1147
rect -1011 947 -951 1147
rect -893 947 -833 1147
rect -775 947 -715 1147
rect -657 947 -597 1147
rect -539 947 -479 1147
rect -421 947 -361 1147
rect 531 1241 591 1641
rect 649 1241 709 1641
rect 767 1241 827 1641
rect 885 1241 945 1641
rect 1003 1241 1063 1641
rect 1121 1241 1181 1641
rect 2429 1241 2489 1641
rect 2547 1241 2607 1641
rect 2665 1241 2725 1641
rect 2783 1241 2843 1641
rect 2901 1241 2961 1641
rect 3019 1241 3079 1641
<< ndiff >>
rect -1195 3952 -1137 3964
rect -1195 3576 -1183 3952
rect -1149 3576 -1137 3952
rect -1195 3564 -1137 3576
rect -1077 3952 -1019 3964
rect -1077 3576 -1065 3952
rect -1031 3576 -1019 3952
rect -1077 3564 -1019 3576
rect -959 3952 -901 3964
rect -959 3576 -947 3952
rect -913 3576 -901 3952
rect -842 3952 -784 3964
rect -842 3776 -830 3952
rect -796 3776 -784 3952
rect -842 3764 -784 3776
rect -724 3952 -666 3964
rect -724 3776 -712 3952
rect -678 3776 -666 3952
rect -724 3764 -666 3776
rect 803 3678 861 3690
rect -959 3564 -901 3576
rect 803 3502 815 3678
rect 849 3502 861 3678
rect 803 3490 861 3502
rect 921 3678 979 3690
rect 921 3502 933 3678
rect 967 3502 979 3678
rect 921 3490 979 3502
rect 1039 3678 1097 3690
rect 1039 3502 1051 3678
rect 1085 3502 1097 3678
rect 1039 3490 1097 3502
rect 1157 3678 1215 3690
rect 1157 3502 1169 3678
rect 1203 3502 1215 3678
rect 1157 3490 1215 3502
rect 1945 3682 2003 3694
rect 1945 3506 1957 3682
rect 1991 3506 2003 3682
rect 1945 3494 2003 3506
rect 2063 3682 2121 3694
rect 2063 3506 2075 3682
rect 2109 3506 2121 3682
rect 2063 3494 2121 3506
rect 2181 3682 2239 3694
rect 2181 3506 2193 3682
rect 2227 3506 2239 3682
rect 2181 3494 2239 3506
rect 2299 3682 2357 3694
rect 2299 3506 2311 3682
rect 2345 3506 2357 3682
rect 2299 3494 2357 3506
rect -1181 2302 -1123 2314
rect -1181 1926 -1169 2302
rect -1135 1926 -1123 2302
rect -1181 1914 -1123 1926
rect -1063 2302 -1005 2314
rect -1063 1926 -1051 2302
rect -1017 1926 -1005 2302
rect -1063 1914 -1005 1926
rect -945 2302 -887 2314
rect -945 1926 -933 2302
rect -899 1926 -887 2302
rect -828 2302 -770 2314
rect -828 2126 -816 2302
rect -782 2126 -770 2302
rect -828 2114 -770 2126
rect -710 2302 -652 2314
rect -710 2126 -698 2302
rect -664 2126 -652 2302
rect -710 2114 -652 2126
rect -945 1914 -887 1926
rect 171 897 229 909
rect 171 721 183 897
rect 217 721 229 897
rect -1186 698 -1128 710
rect -1186 322 -1174 698
rect -1140 322 -1128 698
rect -1186 310 -1128 322
rect -1068 698 -1010 710
rect -1068 322 -1056 698
rect -1022 322 -1010 698
rect -1068 310 -1010 322
rect -950 698 -892 710
rect -950 322 -938 698
rect -904 322 -892 698
rect -833 698 -775 710
rect -833 522 -821 698
rect -787 522 -775 698
rect -833 510 -775 522
rect -715 698 -657 710
rect 171 709 229 721
rect 289 897 347 909
rect 289 721 301 897
rect 335 721 347 897
rect 289 709 347 721
rect 591 897 649 909
rect -715 522 -703 698
rect -669 522 -657 698
rect -715 510 -657 522
rect 591 521 603 897
rect 637 521 649 897
rect 591 509 649 521
rect 709 897 767 909
rect 709 521 721 897
rect 755 521 767 897
rect 709 509 767 521
rect 827 897 885 909
rect 827 521 839 897
rect 873 521 885 897
rect 827 509 885 521
rect 945 897 1003 909
rect 945 521 957 897
rect 991 521 1003 897
rect 945 509 1003 521
rect 1063 897 1121 909
rect 1063 521 1075 897
rect 1109 521 1121 897
rect 1469 897 1527 909
rect 1469 721 1481 897
rect 1515 721 1527 897
rect 1469 709 1527 721
rect 1587 897 1645 909
rect 1587 721 1599 897
rect 1633 721 1645 897
rect 1587 709 1645 721
rect 2069 897 2127 909
rect 2069 721 2081 897
rect 2115 721 2127 897
rect 2069 709 2127 721
rect 2187 897 2245 909
rect 2187 721 2199 897
rect 2233 721 2245 897
rect 2187 709 2245 721
rect 2489 897 2547 909
rect 1063 509 1121 521
rect 2489 521 2501 897
rect 2535 521 2547 897
rect 2489 509 2547 521
rect 2607 897 2665 909
rect 2607 521 2619 897
rect 2653 521 2665 897
rect 2607 509 2665 521
rect 2725 897 2783 909
rect 2725 521 2737 897
rect 2771 521 2783 897
rect 2725 509 2783 521
rect 2843 897 2901 909
rect 2843 521 2855 897
rect 2889 521 2901 897
rect 2843 509 2901 521
rect 2961 897 3019 909
rect 2961 521 2973 897
rect 3007 521 3019 897
rect 3367 897 3425 909
rect 3367 721 3379 897
rect 3413 721 3425 897
rect 3367 709 3425 721
rect 3485 897 3543 909
rect 3485 721 3497 897
rect 3531 721 3543 897
rect 3485 709 3543 721
rect 2961 509 3019 521
rect -950 310 -892 322
<< pdiff >>
rect 893 4461 951 4473
rect -1432 4389 -1374 4401
rect -1432 4213 -1420 4389
rect -1386 4213 -1374 4389
rect -1432 4201 -1374 4213
rect -1314 4389 -1256 4401
rect -1314 4213 -1302 4389
rect -1268 4213 -1256 4389
rect -1314 4201 -1256 4213
rect -1196 4389 -1138 4401
rect -1196 4213 -1184 4389
rect -1150 4213 -1138 4389
rect -1196 4201 -1138 4213
rect -1078 4389 -1020 4401
rect -1078 4213 -1066 4389
rect -1032 4213 -1020 4389
rect -1078 4201 -1020 4213
rect -960 4389 -902 4401
rect -960 4213 -948 4389
rect -914 4213 -902 4389
rect -960 4201 -902 4213
rect -842 4389 -784 4401
rect -842 4213 -830 4389
rect -796 4213 -784 4389
rect -842 4201 -784 4213
rect -724 4389 -666 4401
rect -724 4213 -712 4389
rect -678 4213 -666 4389
rect -724 4201 -666 4213
rect -606 4389 -548 4401
rect -606 4213 -594 4389
rect -560 4213 -548 4389
rect -606 4201 -548 4213
rect -488 4389 -430 4401
rect -488 4213 -476 4389
rect -442 4213 -430 4389
rect -488 4201 -430 4213
rect -370 4389 -312 4401
rect -370 4213 -358 4389
rect -324 4213 -312 4389
rect -370 4201 -312 4213
rect 893 4085 905 4461
rect 939 4085 951 4461
rect 893 4073 951 4085
rect 1011 4461 1069 4473
rect 1011 4085 1023 4461
rect 1057 4085 1069 4461
rect 1011 4073 1069 4085
rect 1129 4461 1187 4473
rect 1129 4085 1141 4461
rect 1175 4085 1187 4461
rect 1129 4073 1187 4085
rect 1247 4461 1305 4473
rect 1247 4085 1259 4461
rect 1293 4085 1305 4461
rect 1247 4073 1305 4085
rect 1365 4461 1423 4473
rect 1365 4085 1377 4461
rect 1411 4085 1423 4461
rect 1365 4073 1423 4085
rect 1483 4461 1541 4473
rect 1483 4085 1495 4461
rect 1529 4085 1541 4461
rect 1483 4073 1541 4085
rect 1601 4461 1659 4473
rect 1601 4085 1613 4461
rect 1647 4085 1659 4461
rect 1601 4073 1659 4085
rect 2035 4465 2093 4477
rect 2035 4089 2047 4465
rect 2081 4089 2093 4465
rect 2035 4077 2093 4089
rect 2153 4465 2211 4477
rect 2153 4089 2165 4465
rect 2199 4089 2211 4465
rect 2153 4077 2211 4089
rect 2271 4465 2329 4477
rect 2271 4089 2283 4465
rect 2317 4089 2329 4465
rect 2271 4077 2329 4089
rect 2389 4465 2447 4477
rect 2389 4089 2401 4465
rect 2435 4089 2447 4465
rect 2389 4077 2447 4089
rect 2507 4465 2565 4477
rect 2507 4089 2519 4465
rect 2553 4089 2565 4465
rect 2507 4077 2565 4089
rect 2625 4465 2683 4477
rect 2625 4089 2637 4465
rect 2671 4089 2683 4465
rect 2625 4077 2683 4089
rect 2743 4465 2801 4477
rect 2743 4089 2755 4465
rect 2789 4089 2801 4465
rect 2743 4077 2801 4089
rect 1322 3678 1380 3690
rect 1322 3502 1334 3678
rect 1368 3502 1380 3678
rect 1322 3490 1380 3502
rect 1440 3678 1498 3690
rect 1440 3502 1452 3678
rect 1486 3502 1498 3678
rect 1440 3490 1498 3502
rect 1558 3678 1616 3690
rect 1558 3502 1570 3678
rect 1604 3502 1616 3678
rect 1558 3490 1616 3502
rect 1676 3678 1734 3690
rect 1676 3502 1688 3678
rect 1722 3502 1734 3678
rect 1676 3490 1734 3502
rect 2464 3682 2522 3694
rect 2464 3506 2476 3682
rect 2510 3506 2522 3682
rect 2464 3494 2522 3506
rect 2582 3682 2640 3694
rect 2582 3506 2594 3682
rect 2628 3506 2640 3682
rect 2582 3494 2640 3506
rect 2700 3682 2758 3694
rect 2700 3506 2712 3682
rect 2746 3506 2758 3682
rect 2700 3494 2758 3506
rect 2818 3682 2876 3694
rect 2818 3506 2830 3682
rect 2864 3506 2876 3682
rect 2818 3494 2876 3506
rect -1418 2739 -1360 2751
rect -1418 2563 -1406 2739
rect -1372 2563 -1360 2739
rect -1418 2551 -1360 2563
rect -1300 2739 -1242 2751
rect -1300 2563 -1288 2739
rect -1254 2563 -1242 2739
rect -1300 2551 -1242 2563
rect -1182 2739 -1124 2751
rect -1182 2563 -1170 2739
rect -1136 2563 -1124 2739
rect -1182 2551 -1124 2563
rect -1064 2739 -1006 2751
rect -1064 2563 -1052 2739
rect -1018 2563 -1006 2739
rect -1064 2551 -1006 2563
rect -946 2739 -888 2751
rect -946 2563 -934 2739
rect -900 2563 -888 2739
rect -946 2551 -888 2563
rect -828 2739 -770 2751
rect -828 2563 -816 2739
rect -782 2563 -770 2739
rect -828 2551 -770 2563
rect -710 2739 -652 2751
rect -710 2563 -698 2739
rect -664 2563 -652 2739
rect -710 2551 -652 2563
rect -592 2739 -534 2751
rect -592 2563 -580 2739
rect -546 2563 -534 2739
rect -592 2551 -534 2563
rect -474 2739 -416 2751
rect -474 2563 -462 2739
rect -428 2563 -416 2739
rect -474 2551 -416 2563
rect -356 2739 -298 2751
rect -356 2563 -344 2739
rect -310 2563 -298 2739
rect -356 2551 -298 2563
rect 530 2322 588 2334
rect 46 2122 104 2134
rect 46 1946 58 2122
rect 92 1946 104 2122
rect 46 1934 104 1946
rect 164 2122 222 2134
rect 164 1946 176 2122
rect 210 1946 222 2122
rect 164 1934 222 1946
rect 282 2122 340 2134
rect 282 1946 294 2122
rect 328 1946 340 2122
rect 282 1934 340 1946
rect 400 2122 458 2134
rect 400 1946 412 2122
rect 446 1946 458 2122
rect 400 1934 458 1946
rect 530 1946 542 2322
rect 576 1946 588 2322
rect 530 1934 588 1946
rect 648 2322 706 2334
rect 648 1946 660 2322
rect 694 1946 706 2322
rect 648 1934 706 1946
rect 766 2322 824 2334
rect 766 1946 778 2322
rect 812 1946 824 2322
rect 766 1934 824 1946
rect 884 2322 942 2334
rect 884 1946 896 2322
rect 930 1946 942 2322
rect 884 1934 942 1946
rect 1002 2322 1060 2334
rect 1002 1946 1014 2322
rect 1048 1946 1060 2322
rect 1002 1934 1060 1946
rect 1120 2322 1178 2334
rect 1120 1946 1132 2322
rect 1166 1946 1178 2322
rect 1120 1934 1178 1946
rect 1238 2322 1296 2334
rect 1238 1946 1250 2322
rect 1284 1946 1296 2322
rect 2428 2322 2486 2334
rect 1238 1934 1296 1946
rect 1367 2122 1425 2134
rect 1367 1946 1379 2122
rect 1413 1946 1425 2122
rect 1367 1934 1425 1946
rect 1485 2122 1543 2134
rect 1485 1946 1497 2122
rect 1531 1946 1543 2122
rect 1485 1934 1543 1946
rect 1603 2122 1661 2134
rect 1603 1946 1615 2122
rect 1649 1946 1661 2122
rect 1603 1934 1661 1946
rect 1721 2122 1779 2134
rect 1721 1946 1733 2122
rect 1767 1946 1779 2122
rect 1721 1934 1779 1946
rect 1944 2122 2002 2134
rect 1944 1946 1956 2122
rect 1990 1946 2002 2122
rect 1944 1934 2002 1946
rect 2062 2122 2120 2134
rect 2062 1946 2074 2122
rect 2108 1946 2120 2122
rect 2062 1934 2120 1946
rect 2180 2122 2238 2134
rect 2180 1946 2192 2122
rect 2226 1946 2238 2122
rect 2180 1934 2238 1946
rect 2298 2122 2356 2134
rect 2298 1946 2310 2122
rect 2344 1946 2356 2122
rect 2298 1934 2356 1946
rect 2428 1946 2440 2322
rect 2474 1946 2486 2322
rect 2428 1934 2486 1946
rect 2546 2322 2604 2334
rect 2546 1946 2558 2322
rect 2592 1946 2604 2322
rect 2546 1934 2604 1946
rect 2664 2322 2722 2334
rect 2664 1946 2676 2322
rect 2710 1946 2722 2322
rect 2664 1934 2722 1946
rect 2782 2322 2840 2334
rect 2782 1946 2794 2322
rect 2828 1946 2840 2322
rect 2782 1934 2840 1946
rect 2900 2322 2958 2334
rect 2900 1946 2912 2322
rect 2946 1946 2958 2322
rect 2900 1934 2958 1946
rect 3018 2322 3076 2334
rect 3018 1946 3030 2322
rect 3064 1946 3076 2322
rect 3018 1934 3076 1946
rect 3136 2322 3194 2334
rect 3136 1946 3148 2322
rect 3182 1946 3194 2322
rect 3136 1934 3194 1946
rect 3265 2122 3323 2134
rect 3265 1946 3277 2122
rect 3311 1946 3323 2122
rect 3265 1934 3323 1946
rect 3383 2122 3441 2134
rect 3383 1946 3395 2122
rect 3429 1946 3441 2122
rect 3383 1934 3441 1946
rect 3501 2122 3559 2134
rect 3501 1946 3513 2122
rect 3547 1946 3559 2122
rect 3501 1934 3559 1946
rect 3619 2122 3677 2134
rect 3619 1946 3631 2122
rect 3665 1946 3677 2122
rect 3619 1934 3677 1946
rect -1423 1135 -1365 1147
rect -1423 959 -1411 1135
rect -1377 959 -1365 1135
rect -1423 947 -1365 959
rect -1305 1135 -1247 1147
rect -1305 959 -1293 1135
rect -1259 959 -1247 1135
rect -1305 947 -1247 959
rect -1187 1135 -1129 1147
rect -1187 959 -1175 1135
rect -1141 959 -1129 1135
rect -1187 947 -1129 959
rect -1069 1135 -1011 1147
rect -1069 959 -1057 1135
rect -1023 959 -1011 1135
rect -1069 947 -1011 959
rect -951 1135 -893 1147
rect -951 959 -939 1135
rect -905 959 -893 1135
rect -951 947 -893 959
rect -833 1135 -775 1147
rect -833 959 -821 1135
rect -787 959 -775 1135
rect -833 947 -775 959
rect -715 1135 -657 1147
rect -715 959 -703 1135
rect -669 959 -657 1135
rect -715 947 -657 959
rect -597 1135 -539 1147
rect -597 959 -585 1135
rect -551 959 -539 1135
rect -597 947 -539 959
rect -479 1135 -421 1147
rect -479 959 -467 1135
rect -433 959 -421 1135
rect -479 947 -421 959
rect -361 1135 -303 1147
rect -361 959 -349 1135
rect -315 959 -303 1135
rect -361 947 -303 959
rect 473 1629 531 1641
rect 473 1253 485 1629
rect 519 1253 531 1629
rect 473 1241 531 1253
rect 591 1629 649 1641
rect 591 1253 603 1629
rect 637 1253 649 1629
rect 591 1241 649 1253
rect 709 1629 767 1641
rect 709 1253 721 1629
rect 755 1253 767 1629
rect 709 1241 767 1253
rect 827 1629 885 1641
rect 827 1253 839 1629
rect 873 1253 885 1629
rect 827 1241 885 1253
rect 945 1629 1003 1641
rect 945 1253 957 1629
rect 991 1253 1003 1629
rect 945 1241 1003 1253
rect 1063 1629 1121 1641
rect 1063 1253 1075 1629
rect 1109 1253 1121 1629
rect 1063 1241 1121 1253
rect 1181 1629 1239 1641
rect 1181 1253 1193 1629
rect 1227 1253 1239 1629
rect 1181 1241 1239 1253
rect 2371 1629 2429 1641
rect 2371 1253 2383 1629
rect 2417 1253 2429 1629
rect 2371 1241 2429 1253
rect 2489 1629 2547 1641
rect 2489 1253 2501 1629
rect 2535 1253 2547 1629
rect 2489 1241 2547 1253
rect 2607 1629 2665 1641
rect 2607 1253 2619 1629
rect 2653 1253 2665 1629
rect 2607 1241 2665 1253
rect 2725 1629 2783 1641
rect 2725 1253 2737 1629
rect 2771 1253 2783 1629
rect 2725 1241 2783 1253
rect 2843 1629 2901 1641
rect 2843 1253 2855 1629
rect 2889 1253 2901 1629
rect 2843 1241 2901 1253
rect 2961 1629 3019 1641
rect 2961 1253 2973 1629
rect 3007 1253 3019 1629
rect 2961 1241 3019 1253
rect 3079 1629 3137 1641
rect 3079 1253 3091 1629
rect 3125 1253 3137 1629
rect 3079 1241 3137 1253
<< ndiffc >>
rect -1183 3576 -1149 3952
rect -1065 3576 -1031 3952
rect -947 3576 -913 3952
rect -830 3776 -796 3952
rect -712 3776 -678 3952
rect 815 3502 849 3678
rect 933 3502 967 3678
rect 1051 3502 1085 3678
rect 1169 3502 1203 3678
rect 1957 3506 1991 3682
rect 2075 3506 2109 3682
rect 2193 3506 2227 3682
rect 2311 3506 2345 3682
rect -1169 1926 -1135 2302
rect -1051 1926 -1017 2302
rect -933 1926 -899 2302
rect -816 2126 -782 2302
rect -698 2126 -664 2302
rect 183 721 217 897
rect -1174 322 -1140 698
rect -1056 322 -1022 698
rect -938 322 -904 698
rect -821 522 -787 698
rect 301 721 335 897
rect -703 522 -669 698
rect 603 521 637 897
rect 721 521 755 897
rect 839 521 873 897
rect 957 521 991 897
rect 1075 521 1109 897
rect 1481 721 1515 897
rect 1599 721 1633 897
rect 2081 721 2115 897
rect 2199 721 2233 897
rect 2501 521 2535 897
rect 2619 521 2653 897
rect 2737 521 2771 897
rect 2855 521 2889 897
rect 2973 521 3007 897
rect 3379 721 3413 897
rect 3497 721 3531 897
<< pdiffc >>
rect -1420 4213 -1386 4389
rect -1302 4213 -1268 4389
rect -1184 4213 -1150 4389
rect -1066 4213 -1032 4389
rect -948 4213 -914 4389
rect -830 4213 -796 4389
rect -712 4213 -678 4389
rect -594 4213 -560 4389
rect -476 4213 -442 4389
rect -358 4213 -324 4389
rect 905 4085 939 4461
rect 1023 4085 1057 4461
rect 1141 4085 1175 4461
rect 1259 4085 1293 4461
rect 1377 4085 1411 4461
rect 1495 4085 1529 4461
rect 1613 4085 1647 4461
rect 2047 4089 2081 4465
rect 2165 4089 2199 4465
rect 2283 4089 2317 4465
rect 2401 4089 2435 4465
rect 2519 4089 2553 4465
rect 2637 4089 2671 4465
rect 2755 4089 2789 4465
rect 1334 3502 1368 3678
rect 1452 3502 1486 3678
rect 1570 3502 1604 3678
rect 1688 3502 1722 3678
rect 2476 3506 2510 3682
rect 2594 3506 2628 3682
rect 2712 3506 2746 3682
rect 2830 3506 2864 3682
rect -1406 2563 -1372 2739
rect -1288 2563 -1254 2739
rect -1170 2563 -1136 2739
rect -1052 2563 -1018 2739
rect -934 2563 -900 2739
rect -816 2563 -782 2739
rect -698 2563 -664 2739
rect -580 2563 -546 2739
rect -462 2563 -428 2739
rect -344 2563 -310 2739
rect 58 1946 92 2122
rect 176 1946 210 2122
rect 294 1946 328 2122
rect 412 1946 446 2122
rect 542 1946 576 2322
rect 660 1946 694 2322
rect 778 1946 812 2322
rect 896 1946 930 2322
rect 1014 1946 1048 2322
rect 1132 1946 1166 2322
rect 1250 1946 1284 2322
rect 1379 1946 1413 2122
rect 1497 1946 1531 2122
rect 1615 1946 1649 2122
rect 1733 1946 1767 2122
rect 1956 1946 1990 2122
rect 2074 1946 2108 2122
rect 2192 1946 2226 2122
rect 2310 1946 2344 2122
rect 2440 1946 2474 2322
rect 2558 1946 2592 2322
rect 2676 1946 2710 2322
rect 2794 1946 2828 2322
rect 2912 1946 2946 2322
rect 3030 1946 3064 2322
rect 3148 1946 3182 2322
rect 3277 1946 3311 2122
rect 3395 1946 3429 2122
rect 3513 1946 3547 2122
rect 3631 1946 3665 2122
rect -1411 959 -1377 1135
rect -1293 959 -1259 1135
rect -1175 959 -1141 1135
rect -1057 959 -1023 1135
rect -939 959 -905 1135
rect -821 959 -787 1135
rect -703 959 -669 1135
rect -585 959 -551 1135
rect -467 959 -433 1135
rect -349 959 -315 1135
rect 485 1253 519 1629
rect 603 1253 637 1629
rect 721 1253 755 1629
rect 839 1253 873 1629
rect 957 1253 991 1629
rect 1075 1253 1109 1629
rect 1193 1253 1227 1629
rect 2383 1253 2417 1629
rect 2501 1253 2535 1629
rect 2619 1253 2653 1629
rect 2737 1253 2771 1629
rect 2855 1253 2889 1629
rect 2973 1253 3007 1629
rect 3091 1253 3125 1629
<< psubdiff >>
rect -659 3626 -425 3660
rect -659 3536 -613 3626
rect -450 3536 -425 3626
rect -659 3505 -425 3536
rect 838 3255 993 3301
rect 838 3092 869 3255
rect 959 3092 993 3255
rect 838 3067 993 3092
rect 1980 3253 2135 3299
rect 1980 3090 2011 3253
rect 2101 3090 2135 3253
rect 1980 3065 2135 3090
rect -645 1976 -411 2010
rect -645 1886 -599 1976
rect -436 1886 -411 1976
rect -645 1855 -411 1886
rect -650 372 -416 406
rect -650 282 -604 372
rect -441 282 -416 372
rect -650 251 -416 282
rect 782 212 937 258
rect 782 49 813 212
rect 903 49 937 212
rect 782 24 937 49
<< nsubdiff >>
rect 1493 4857 1646 4897
rect -989 4803 -836 4843
rect -989 4654 -946 4803
rect -879 4654 -836 4803
rect -989 4585 -836 4654
rect 1493 4708 1536 4857
rect 1603 4708 1646 4857
rect 1493 4639 1646 4708
rect 2640 4857 2793 4897
rect 2640 4708 2683 4857
rect 2750 4708 2793 4857
rect 2640 4639 2793 4708
rect -975 3153 -822 3193
rect -975 3004 -932 3153
rect -865 3004 -822 3153
rect -975 2935 -822 3004
rect 2736 2810 2889 2850
rect 2736 2661 2779 2810
rect 2846 2661 2889 2810
rect 2736 2592 2889 2661
rect -980 1549 -827 1589
rect -980 1400 -937 1549
rect -870 1400 -827 1549
rect -980 1331 -827 1400
<< psubdiffcont >>
rect -613 3536 -450 3626
rect 869 3092 959 3255
rect 2011 3090 2101 3253
rect -599 1886 -436 1976
rect -604 282 -441 372
rect 813 49 903 212
<< nsubdiffcont >>
rect -946 4654 -879 4803
rect 1536 4708 1603 4857
rect 2683 4708 2750 4857
rect -932 3004 -865 3153
rect 2779 2661 2846 2810
rect -937 1400 -870 1549
<< poly >>
rect 774 4637 840 4653
rect 1904 4643 1970 4659
rect 774 4603 790 4637
rect 824 4630 840 4637
rect 824 4603 1349 4630
rect 774 4587 1349 4603
rect 1904 4609 1920 4643
rect 1954 4634 1970 4643
rect 1954 4609 2491 4634
rect 1904 4591 2491 4609
rect 1305 4535 1349 4587
rect 2447 4539 2491 4591
rect 774 4519 1247 4535
rect 774 4485 790 4519
rect 824 4494 1247 4519
rect 824 4493 1011 4494
rect 824 4485 840 4493
rect 774 4469 840 4485
rect 951 4473 1011 4493
rect 1069 4473 1129 4494
rect 1187 4473 1247 4494
rect 1305 4494 1601 4535
rect 1305 4473 1365 4494
rect 1423 4473 1483 4494
rect 1541 4473 1601 4494
rect 1904 4523 2389 4539
rect 1904 4489 1920 4523
rect 1954 4498 2389 4523
rect 1954 4497 2153 4498
rect 1954 4489 1970 4497
rect 1904 4473 1970 4489
rect 2093 4477 2153 4497
rect 2211 4477 2271 4498
rect 2329 4477 2389 4498
rect 2447 4498 2743 4539
rect 2447 4477 2507 4498
rect 2565 4477 2625 4498
rect 2683 4477 2743 4498
rect -1374 4422 -1078 4458
rect -1374 4401 -1314 4422
rect -1256 4401 -1196 4422
rect -1138 4401 -1078 4422
rect -1020 4421 -724 4457
rect -1020 4401 -960 4421
rect -902 4401 -842 4421
rect -784 4401 -724 4421
rect -666 4421 -370 4457
rect -666 4401 -606 4421
rect -548 4401 -488 4421
rect -430 4401 -370 4421
rect -1374 4175 -1314 4201
rect -1256 4175 -1196 4201
rect -1138 4175 -1078 4201
rect -1020 4181 -960 4201
rect -1020 4175 -959 4181
rect -902 4175 -842 4201
rect -784 4175 -724 4201
rect -1137 3990 -1079 4175
rect -1137 3964 -1077 3990
rect -1019 3964 -959 4175
rect -666 4169 -606 4201
rect -548 4175 -488 4201
rect -430 4175 -370 4201
rect -669 4153 -603 4169
rect -669 4119 -653 4153
rect -619 4119 -603 4153
rect -669 4103 -603 4119
rect 951 4056 1011 4073
rect -787 4036 -721 4052
rect -787 4002 -771 4036
rect -737 4002 -721 4036
rect -787 3986 -721 4002
rect -784 3964 -724 3986
rect 951 3967 1012 4056
rect 1069 4047 1129 4073
rect 1187 4047 1247 4073
rect 861 3914 1012 3967
rect -784 3738 -724 3764
rect 861 3690 921 3914
rect 1305 3872 1365 4073
rect 1423 4047 1483 4073
rect 1541 4047 1601 4073
rect 2093 4060 2153 4077
rect 2093 3971 2154 4060
rect 2211 4051 2271 4077
rect 2329 4051 2389 4077
rect 979 3821 1365 3872
rect 2003 3918 2154 3971
rect 979 3690 1039 3821
rect 1094 3763 1160 3779
rect 1094 3729 1110 3763
rect 1144 3729 1160 3763
rect 1094 3713 1160 3729
rect 1097 3690 1157 3713
rect 1380 3690 1440 3716
rect 1498 3690 1558 3716
rect 1616 3690 1676 3716
rect 2003 3694 2063 3918
rect 2447 3876 2507 4077
rect 2565 4051 2625 4077
rect 2683 4051 2743 4077
rect 2121 3825 2507 3876
rect 2121 3694 2181 3825
rect 2236 3767 2302 3783
rect 2236 3733 2252 3767
rect 2286 3733 2302 3767
rect 2236 3717 2302 3733
rect 2239 3694 2299 3717
rect 2522 3694 2582 3720
rect 2640 3694 2700 3720
rect 2758 3694 2818 3720
rect -1137 3542 -1077 3564
rect -1019 3542 -959 3564
rect -1140 3526 -1074 3542
rect -1140 3492 -1124 3526
rect -1090 3492 -1074 3526
rect -1140 3476 -1074 3492
rect -1022 3526 -956 3542
rect -1022 3492 -1006 3526
rect -972 3492 -956 3526
rect -1022 3476 -956 3492
rect 861 3464 921 3490
rect 979 3464 1039 3490
rect 1097 3458 1157 3490
rect 1380 3458 1440 3490
rect 1498 3458 1558 3490
rect 1616 3458 1676 3490
rect 2003 3468 2063 3494
rect 2121 3468 2181 3494
rect 1097 3417 1676 3458
rect 2239 3462 2299 3494
rect 2522 3462 2582 3494
rect 2640 3462 2700 3494
rect 2758 3462 2818 3494
rect 2239 3421 2818 3462
rect -1360 2772 -1064 2808
rect -1360 2751 -1300 2772
rect -1242 2751 -1182 2772
rect -1124 2751 -1064 2772
rect -1006 2771 -710 2807
rect -1006 2751 -946 2771
rect -888 2751 -828 2771
rect -770 2751 -710 2771
rect -652 2771 -356 2807
rect -652 2751 -592 2771
rect -534 2751 -474 2771
rect -416 2751 -356 2771
rect -1360 2525 -1300 2551
rect -1242 2525 -1182 2551
rect -1124 2525 -1064 2551
rect -1006 2531 -946 2551
rect -1006 2525 -945 2531
rect -888 2525 -828 2551
rect -770 2525 -710 2551
rect -1123 2340 -1065 2525
rect -1123 2314 -1063 2340
rect -1005 2314 -945 2525
rect -652 2519 -592 2551
rect -534 2525 -474 2551
rect -416 2525 -356 2551
rect -655 2503 -589 2519
rect -655 2469 -639 2503
rect -605 2469 -589 2503
rect -655 2453 -589 2469
rect -773 2386 -707 2402
rect -773 2352 -757 2386
rect -723 2352 -707 2386
rect -773 2336 -707 2352
rect 588 2349 884 2400
rect -770 2314 -710 2336
rect 588 2334 648 2349
rect 706 2334 766 2349
rect 824 2334 884 2349
rect 942 2334 1002 2360
rect 1060 2334 1120 2360
rect 1178 2334 1238 2360
rect 2486 2349 2782 2400
rect 2486 2334 2546 2349
rect 2604 2334 2664 2349
rect 2722 2334 2782 2349
rect 2840 2334 2900 2360
rect 2958 2334 3018 2360
rect 3076 2334 3136 2360
rect 104 2134 164 2160
rect 222 2134 282 2160
rect 340 2134 400 2160
rect -770 2088 -710 2114
rect -1123 1892 -1063 1914
rect -1005 1898 -945 1914
rect -1126 1876 -1060 1892
rect -1126 1842 -1110 1876
rect -1076 1842 -1060 1876
rect -1126 1826 -1060 1842
rect -1011 1876 -937 1898
rect -1011 1842 -992 1876
rect -958 1842 -937 1876
rect 1425 2151 1721 2202
rect 1425 2134 1485 2151
rect 1543 2134 1603 2151
rect 1661 2134 1721 2151
rect 2002 2134 2062 2160
rect 2120 2134 2180 2160
rect 2238 2134 2298 2160
rect 3323 2151 3619 2202
rect 3323 2134 3383 2151
rect 3441 2134 3501 2151
rect 3559 2134 3619 2151
rect 104 1917 164 1934
rect 222 1917 282 1934
rect 340 1917 400 1934
rect 588 1917 648 1934
rect 104 1866 648 1917
rect 706 1908 766 1934
rect 824 1908 884 1934
rect 942 1915 1002 1934
rect 1060 1915 1120 1934
rect 1178 1915 1238 1934
rect 1425 1915 1485 1934
rect 1543 1915 1603 1934
rect -1011 1785 -937 1842
rect 229 1785 289 1866
rect 942 1864 1485 1915
rect 1527 1908 1603 1915
rect 1661 1908 1721 1934
rect 2002 1917 2062 1934
rect 2120 1917 2180 1934
rect 2238 1917 2298 1934
rect 2486 1917 2546 1934
rect 1527 1864 1602 1908
rect 2002 1866 2546 1917
rect 2604 1908 2664 1934
rect 2722 1908 2782 1934
rect 2840 1915 2900 1934
rect 2958 1915 3018 1934
rect 3076 1915 3136 1934
rect 3323 1915 3383 1934
rect 3441 1915 3501 1934
rect -1011 1760 289 1785
rect -1012 1712 289 1760
rect 1527 1744 1587 1864
rect -1365 1168 -1069 1204
rect -1365 1147 -1305 1168
rect -1247 1147 -1187 1168
rect -1129 1147 -1069 1168
rect -1011 1167 -715 1203
rect -1011 1147 -951 1167
rect -893 1147 -833 1167
rect -775 1147 -715 1167
rect -657 1167 -361 1203
rect -657 1147 -597 1167
rect -539 1147 -479 1167
rect -421 1147 -361 1167
rect 229 1014 289 1712
rect 531 1664 827 1724
rect 531 1641 591 1664
rect 649 1641 709 1664
rect 767 1641 827 1664
rect 885 1665 1181 1725
rect 1526 1724 1587 1744
rect 885 1641 945 1665
rect 1003 1641 1063 1665
rect 1121 1641 1181 1665
rect 1507 1708 1587 1724
rect 1507 1674 1522 1708
rect 1556 1674 1587 1708
rect 1507 1658 1587 1674
rect 1526 1635 1587 1658
rect 1527 1489 1587 1635
rect 1526 1316 1587 1489
rect 531 1215 591 1241
rect 499 1074 566 1081
rect 649 1074 709 1241
rect 767 1215 827 1241
rect 885 1215 945 1241
rect 499 1065 709 1074
rect 499 1031 515 1065
rect 549 1031 709 1065
rect 499 1015 709 1031
rect 229 998 380 1014
rect 229 964 330 998
rect 364 964 380 998
rect 229 948 380 964
rect -1365 921 -1305 947
rect -1247 921 -1187 947
rect -1129 921 -1069 947
rect -1011 927 -951 947
rect -1011 921 -950 927
rect -893 921 -833 947
rect -775 921 -715 947
rect -1128 736 -1070 921
rect -1128 710 -1068 736
rect -1010 710 -950 921
rect -657 915 -597 947
rect -539 921 -479 947
rect -421 921 -361 947
rect -660 899 -594 915
rect 229 909 289 948
rect 649 909 709 1015
rect 1003 1074 1063 1241
rect 1121 1215 1181 1241
rect 1146 1074 1213 1081
rect 1003 1065 1213 1074
rect 1003 1031 1163 1065
rect 1197 1031 1213 1065
rect 1003 1015 1213 1031
rect 765 981 831 997
rect 765 947 781 981
rect 815 947 831 981
rect 765 931 831 947
rect 883 982 949 997
rect 883 948 899 982
rect 933 948 949 982
rect 883 932 949 948
rect 767 909 827 931
rect 885 909 945 932
rect 1003 909 1063 1015
rect 1527 1013 1587 1316
rect 1437 997 1587 1013
rect 1437 963 1453 997
rect 1487 963 1587 997
rect 1437 947 1587 963
rect 1527 909 1587 947
rect 2127 1208 2187 1866
rect 2840 1864 3383 1915
rect 3425 1908 3501 1915
rect 3559 1908 3619 1934
rect 3425 1864 3500 1908
rect 2429 1664 2725 1724
rect 2429 1641 2489 1664
rect 2547 1641 2607 1664
rect 2665 1641 2725 1664
rect 2783 1665 3079 1725
rect 2783 1641 2843 1665
rect 2901 1641 2961 1665
rect 3019 1641 3079 1665
rect 3425 1711 3485 1864
rect 3425 1687 3679 1711
rect 3425 1653 3629 1687
rect 3663 1653 3679 1687
rect 3425 1637 3679 1653
rect 2429 1215 2489 1241
rect 2127 1192 2194 1208
rect 2127 1158 2143 1192
rect 2177 1158 2194 1192
rect 2127 1142 2194 1158
rect 2127 1014 2187 1142
rect 2397 1074 2464 1081
rect 2547 1074 2607 1241
rect 2665 1215 2725 1241
rect 2783 1215 2843 1241
rect 2397 1065 2607 1074
rect 2397 1031 2413 1065
rect 2447 1031 2607 1065
rect 2397 1015 2607 1031
rect 2127 998 2278 1014
rect 2127 964 2228 998
rect 2262 964 2278 998
rect 2127 948 2278 964
rect 2127 909 2187 948
rect 2547 909 2607 1015
rect 2901 1074 2961 1241
rect 3019 1215 3079 1241
rect 3042 1075 3109 1082
rect 3036 1074 3109 1075
rect 2901 1066 3109 1074
rect 2901 1032 3059 1066
rect 3093 1032 3109 1066
rect 2901 1016 3109 1032
rect 2901 1015 3098 1016
rect 2663 981 2729 997
rect 2663 947 2679 981
rect 2713 947 2729 981
rect 2663 931 2729 947
rect 2781 982 2847 997
rect 2781 948 2797 982
rect 2831 948 2847 982
rect 2781 932 2847 948
rect 2665 909 2725 931
rect 2783 909 2843 932
rect 2901 909 2961 1015
rect 3425 1013 3485 1637
rect 3335 997 3485 1013
rect 3335 963 3351 997
rect 3385 963 3485 997
rect 3335 947 3485 963
rect 3425 909 3485 947
rect -660 865 -644 899
rect -610 865 -594 899
rect -660 849 -594 865
rect -778 782 -712 798
rect -778 748 -762 782
rect -728 748 -712 782
rect -778 732 -712 748
rect -775 710 -715 732
rect 229 683 289 709
rect -775 484 -715 510
rect 1527 683 1587 709
rect 2127 683 2187 709
rect 3425 683 3485 709
rect 649 483 709 509
rect 767 483 827 509
rect 885 483 945 509
rect 1003 483 1063 509
rect 2547 483 2607 509
rect 2665 483 2725 509
rect 2783 483 2843 509
rect 2901 483 2961 509
rect -1128 288 -1068 310
rect -1010 288 -950 310
rect -1131 272 -1065 288
rect -1131 238 -1115 272
rect -1081 238 -1065 272
rect -1131 222 -1065 238
rect -1013 272 -947 288
rect -1013 238 -997 272
rect -963 238 -947 272
rect -1013 222 -947 238
<< polycont >>
rect 790 4603 824 4637
rect 1920 4609 1954 4643
rect 790 4485 824 4519
rect 1920 4489 1954 4523
rect -653 4119 -619 4153
rect -771 4002 -737 4036
rect 1110 3729 1144 3763
rect 2252 3733 2286 3767
rect -1124 3492 -1090 3526
rect -1006 3492 -972 3526
rect -639 2469 -605 2503
rect -757 2352 -723 2386
rect -1110 1842 -1076 1876
rect -992 1842 -958 1876
rect 1522 1674 1556 1708
rect 515 1031 549 1065
rect 330 964 364 998
rect 1163 1031 1197 1065
rect 781 947 815 981
rect 899 948 933 982
rect 1453 963 1487 997
rect 3629 1653 3663 1687
rect 2143 1158 2177 1192
rect 2413 1031 2447 1065
rect 2228 964 2262 998
rect 3059 1032 3093 1066
rect 2679 947 2713 981
rect 2797 948 2831 982
rect 3351 963 3385 997
rect -644 865 -610 899
rect -762 748 -728 782
rect -1115 238 -1081 272
rect -997 238 -963 272
<< locali >>
rect -1025 4803 -802 4879
rect -1025 4654 -946 4803
rect -879 4654 -802 4803
rect -1025 4548 -802 4654
rect 1457 4857 1680 4933
rect 1457 4708 1536 4857
rect 1603 4708 1680 4857
rect 790 4637 824 4653
rect 790 4587 824 4603
rect 1457 4602 1680 4708
rect 2604 4857 2827 4933
rect 2604 4708 2683 4857
rect 2750 4708 2827 4857
rect 1920 4643 1954 4659
rect 1920 4593 1954 4609
rect 2604 4602 2827 4708
rect 790 4519 824 4535
rect -594 4439 -324 4473
rect 790 4469 824 4485
rect 1920 4523 1954 4539
rect -1420 4389 -1386 4405
rect -1420 4197 -1386 4213
rect -1302 4389 -1268 4405
rect -1302 4197 -1268 4213
rect -1184 4389 -1150 4405
rect -1184 4197 -1150 4213
rect -1066 4389 -1032 4405
rect -1066 4197 -1032 4213
rect -948 4389 -914 4405
rect -948 4197 -914 4213
rect -830 4389 -796 4405
rect -830 4197 -796 4213
rect -712 4389 -678 4405
rect -712 4197 -678 4213
rect -594 4389 -560 4439
rect -594 4197 -560 4213
rect -476 4389 -442 4405
rect -476 4197 -442 4213
rect -358 4389 -324 4439
rect -358 4197 -324 4213
rect 905 4461 939 4477
rect -669 4119 -653 4153
rect -619 4119 -603 4153
rect 905 4069 939 4085
rect 1023 4461 1057 4477
rect 1023 4069 1057 4085
rect 1141 4461 1175 4477
rect 1141 4069 1175 4085
rect 1259 4461 1293 4477
rect 1259 4069 1293 4085
rect 1377 4461 1411 4477
rect 1377 4069 1411 4085
rect 1495 4461 1529 4477
rect 1495 4069 1529 4085
rect 1613 4461 1647 4477
rect 1920 4473 1954 4489
rect 1613 4069 1647 4085
rect 2047 4465 2081 4481
rect 2047 4073 2081 4089
rect 2165 4465 2199 4481
rect 2165 4073 2199 4089
rect 2283 4465 2317 4481
rect 2283 4073 2317 4089
rect 2401 4465 2435 4481
rect 2401 4073 2435 4089
rect 2519 4465 2553 4481
rect 2519 4073 2553 4089
rect 2637 4465 2671 4481
rect 2637 4073 2671 4089
rect 2755 4465 2789 4481
rect 2755 4073 2789 4089
rect -787 4002 -771 4036
rect -737 4002 -721 4036
rect -1183 3952 -1149 3968
rect -1183 3560 -1149 3576
rect -1065 3952 -1031 3968
rect -1065 3560 -1031 3576
rect -947 3952 -913 3968
rect -830 3952 -796 3968
rect -830 3760 -796 3776
rect -712 3952 -678 3968
rect -712 3760 -678 3776
rect 1094 3729 1110 3763
rect 1144 3729 1160 3763
rect 2236 3733 2252 3767
rect 2286 3733 2302 3767
rect 815 3678 849 3694
rect -947 3560 -913 3576
rect -660 3626 -411 3669
rect -660 3536 -613 3626
rect -450 3536 -411 3626
rect -1140 3492 -1124 3526
rect -1090 3492 -1074 3526
rect -1022 3492 -1006 3526
rect -972 3492 -956 3526
rect -660 3497 -411 3536
rect 815 3486 849 3502
rect 933 3678 967 3694
rect 933 3486 967 3502
rect 1051 3678 1085 3694
rect 1051 3486 1085 3502
rect 1169 3678 1203 3694
rect 1169 3486 1203 3502
rect 1334 3678 1368 3694
rect 1334 3486 1368 3502
rect 1452 3678 1486 3694
rect 1452 3486 1486 3502
rect 1570 3678 1604 3694
rect 1570 3486 1604 3502
rect 1688 3678 1722 3694
rect 1688 3486 1722 3502
rect 1957 3682 1991 3698
rect 1957 3490 1991 3506
rect 2075 3682 2109 3698
rect 2075 3490 2109 3506
rect 2193 3682 2227 3698
rect 2193 3490 2227 3506
rect 2311 3682 2345 3698
rect 2311 3490 2345 3506
rect 2476 3682 2510 3698
rect 2476 3490 2510 3506
rect 2594 3682 2628 3698
rect 2594 3490 2628 3506
rect 2712 3682 2746 3698
rect 2712 3490 2746 3506
rect 2830 3682 2864 3698
rect 2830 3490 2864 3506
rect 830 3255 1002 3302
rect -1011 3153 -788 3229
rect -1011 3004 -932 3153
rect -865 3004 -788 3153
rect 830 3092 869 3255
rect 959 3092 1002 3255
rect 830 3053 1002 3092
rect 1972 3253 2144 3300
rect 1972 3090 2011 3253
rect 2101 3090 2144 3253
rect 1972 3051 2144 3090
rect -1011 2898 -788 3004
rect -580 2789 -310 2823
rect -1406 2739 -1372 2755
rect -1406 2547 -1372 2563
rect -1288 2739 -1254 2755
rect -1288 2547 -1254 2563
rect -1170 2739 -1136 2755
rect -1170 2547 -1136 2563
rect -1052 2739 -1018 2755
rect -1052 2547 -1018 2563
rect -934 2739 -900 2755
rect -934 2547 -900 2563
rect -816 2739 -782 2755
rect -816 2547 -782 2563
rect -698 2739 -664 2755
rect -698 2547 -664 2563
rect -580 2739 -546 2789
rect -580 2547 -546 2563
rect -462 2739 -428 2755
rect -462 2547 -428 2563
rect -344 2739 -310 2789
rect -344 2547 -310 2563
rect 2700 2810 2925 2886
rect 2700 2661 2779 2810
rect 2846 2661 2925 2810
rect 2700 2555 2925 2661
rect -655 2469 -639 2503
rect -605 2469 -589 2503
rect -773 2352 -757 2386
rect -723 2352 -707 2386
rect 896 2375 1166 2410
rect 542 2322 576 2338
rect -1169 2302 -1135 2318
rect -1169 1910 -1135 1926
rect -1051 2302 -1017 2318
rect -1051 1910 -1017 1926
rect -933 2302 -899 2318
rect -816 2302 -782 2318
rect -816 2110 -782 2126
rect -698 2302 -664 2318
rect -698 2110 -664 2126
rect 58 2176 328 2211
rect 58 2122 92 2176
rect -933 1910 -899 1926
rect -646 1976 -397 2019
rect -646 1886 -599 1976
rect -436 1886 -397 1976
rect 58 1930 92 1946
rect 176 2122 210 2138
rect 176 1930 210 1946
rect 294 2122 328 2176
rect 294 1930 328 1946
rect 412 2122 446 2138
rect 412 1930 446 1946
rect 542 1930 576 1946
rect 660 2322 694 2338
rect 660 1930 694 1946
rect 778 2322 812 2338
rect 778 1930 812 1946
rect 896 2322 930 2375
rect 896 1930 930 1946
rect 1014 2322 1048 2338
rect 1014 1930 1048 1946
rect 1132 2322 1166 2375
rect 2794 2375 3064 2410
rect 1132 1930 1166 1946
rect 1250 2322 1284 2338
rect 2440 2322 2474 2338
rect 1956 2176 2226 2211
rect 1250 1930 1284 1946
rect 1379 2122 1413 2138
rect 1379 1930 1413 1946
rect 1497 2122 1531 2138
rect 1497 1930 1531 1946
rect 1615 2122 1649 2138
rect 1615 1930 1649 1946
rect 1733 2122 1767 2138
rect 1733 1930 1767 1946
rect 1956 2122 1990 2176
rect 1956 1930 1990 1946
rect 2074 2122 2108 2138
rect 2074 1930 2108 1946
rect 2192 2122 2226 2176
rect 2192 1930 2226 1946
rect 2310 2122 2344 2138
rect 2310 1930 2344 1946
rect 2440 1930 2474 1946
rect 2558 2322 2592 2338
rect 2558 1930 2592 1946
rect 2676 2322 2710 2338
rect 2676 1930 2710 1946
rect 2794 2322 2828 2375
rect 2794 1930 2828 1946
rect 2912 2322 2946 2338
rect 2912 1930 2946 1946
rect 3030 2322 3064 2375
rect 3030 1930 3064 1946
rect 3148 2322 3182 2338
rect 3148 1930 3182 1946
rect 3277 2122 3311 2138
rect 3277 1930 3311 1946
rect 3395 2122 3429 2138
rect 3395 1930 3429 1946
rect 3513 2122 3547 2138
rect 3513 1930 3547 1946
rect 3631 2122 3665 2138
rect 3631 1930 3665 1946
rect -1126 1842 -1110 1876
rect -1076 1842 -1060 1876
rect -1008 1842 -992 1876
rect -958 1842 -942 1876
rect -646 1847 -397 1886
rect 1522 1708 1556 1724
rect 1522 1658 1556 1674
rect 3612 1687 3679 1703
rect 3612 1653 3629 1687
rect 3663 1653 3679 1687
rect 485 1629 519 1645
rect -1016 1549 -793 1625
rect -1016 1400 -937 1549
rect -870 1400 -793 1549
rect -1016 1294 -793 1400
rect 603 1629 637 1645
rect 485 1237 519 1253
rect 602 1253 603 1300
rect 721 1629 755 1645
rect 637 1253 638 1300
rect -585 1185 -315 1219
rect -1411 1135 -1377 1151
rect -1411 943 -1377 959
rect -1293 1135 -1259 1151
rect -1293 943 -1259 959
rect -1175 1135 -1141 1151
rect -1175 943 -1141 959
rect -1057 1135 -1023 1151
rect -1057 943 -1023 959
rect -939 1135 -905 1151
rect -939 943 -905 959
rect -821 1135 -787 1151
rect -821 943 -787 959
rect -703 1135 -669 1151
rect -703 943 -669 959
rect -585 1135 -551 1185
rect -585 943 -551 959
rect -467 1135 -433 1151
rect -467 943 -433 959
rect -349 1135 -315 1185
rect 602 1195 638 1253
rect 839 1629 873 1645
rect 721 1237 755 1253
rect 837 1253 839 1300
rect 837 1195 873 1253
rect 957 1629 991 1645
rect 957 1237 991 1253
rect 1075 1629 1109 1645
rect 1193 1629 1227 1645
rect 1109 1253 1111 1299
rect 1075 1195 1111 1253
rect 1193 1237 1227 1253
rect 2383 1629 2417 1645
rect 2501 1629 2535 1645
rect 2383 1237 2417 1253
rect 2500 1253 2501 1300
rect 2619 1629 2653 1645
rect 2535 1253 2536 1300
rect 1698 1195 2195 1213
rect 602 1192 2195 1195
rect 602 1158 2143 1192
rect 2177 1158 2195 1192
rect 602 1155 2195 1158
rect 2500 1195 2536 1253
rect 2737 1629 2771 1645
rect 2619 1237 2653 1253
rect 2735 1253 2737 1300
rect 2735 1195 2771 1253
rect 2855 1629 2889 1645
rect 2855 1237 2889 1253
rect 2973 1629 3007 1645
rect 3091 1629 3125 1645
rect 3612 1637 3679 1653
rect 3007 1253 3009 1299
rect 2973 1195 3009 1253
rect 3091 1237 3125 1253
rect 3596 1224 3696 1225
rect 3596 1195 3752 1224
rect 2500 1155 3752 1195
rect 621 1154 2195 1155
rect 2519 1154 3752 1155
rect 499 1065 566 1081
rect 499 1031 515 1065
rect 549 1031 566 1065
rect 499 1015 566 1031
rect -349 943 -315 959
rect 330 998 364 1014
rect 330 948 364 964
rect 676 913 710 1154
rect 1698 1137 2195 1154
rect 1146 1065 1213 1081
rect 1146 1031 1163 1065
rect 1197 1031 1213 1065
rect 1146 1015 1213 1031
rect 2397 1065 2464 1081
rect 2397 1031 2413 1065
rect 2447 1031 2464 1065
rect 2397 1015 2464 1031
rect 1453 997 1487 1013
rect 765 947 781 981
rect 815 947 831 981
rect 883 948 899 982
rect 933 948 949 982
rect 1453 947 1487 963
rect 2228 998 2262 1014
rect 2228 948 2262 964
rect 2574 913 2608 1154
rect 3596 1126 3752 1154
rect 3596 1125 3696 1126
rect 3042 1066 3109 1082
rect 3042 1032 3059 1066
rect 3093 1032 3109 1066
rect 3042 1016 3109 1032
rect 3351 997 3385 1013
rect 2663 947 2679 981
rect 2713 947 2729 981
rect 2781 948 2797 982
rect 2831 948 2847 982
rect 3351 947 3385 963
rect -660 865 -644 899
rect -610 865 -594 899
rect 183 897 217 913
rect -778 748 -762 782
rect -728 748 -712 782
rect -1174 698 -1140 714
rect -1174 306 -1140 322
rect -1056 698 -1022 714
rect -1056 306 -1022 322
rect -938 698 -904 714
rect -821 698 -787 714
rect -821 506 -787 522
rect -703 698 -669 714
rect 183 705 217 721
rect 301 897 335 913
rect 301 705 335 721
rect 603 897 637 913
rect -703 506 -669 522
rect 676 897 755 913
rect 676 867 721 897
rect 603 454 638 521
rect 721 505 755 521
rect 839 897 873 913
rect 839 505 873 521
rect 957 897 991 913
rect 1075 897 1109 913
rect 1481 897 1515 913
rect 1481 705 1515 721
rect 1599 897 1633 913
rect 1599 705 1633 721
rect 2081 897 2115 913
rect 2081 705 2115 721
rect 2199 897 2233 913
rect 2199 705 2233 721
rect 2501 897 2535 913
rect 957 505 991 521
rect 1074 454 1109 521
rect 603 419 1109 454
rect 2574 897 2653 913
rect 2574 867 2619 897
rect 2501 454 2536 521
rect 2619 505 2653 521
rect 2737 897 2771 913
rect 2737 505 2771 521
rect 2855 897 2889 913
rect 2973 897 3007 913
rect 3379 897 3413 913
rect 3379 705 3413 721
rect 3497 897 3531 913
rect 3497 705 3531 721
rect 2855 505 2889 521
rect 2972 454 3007 521
rect 2501 419 3007 454
rect -938 306 -904 322
rect -651 372 -402 415
rect -651 282 -604 372
rect -441 282 -402 372
rect -1131 238 -1115 272
rect -1081 238 -1065 272
rect -1013 238 -997 272
rect -963 238 -947 272
rect -651 243 -402 282
rect 774 212 946 259
rect 774 49 813 212
rect 903 49 946 212
rect 774 9 946 49
<< viali >>
rect 790 4603 824 4637
rect 1920 4609 1954 4643
rect 790 4485 824 4519
rect 1920 4489 1954 4523
rect -1420 4213 -1386 4389
rect -1302 4213 -1268 4389
rect -1184 4213 -1150 4389
rect -1066 4213 -1032 4389
rect -948 4213 -914 4389
rect -830 4213 -796 4389
rect -712 4213 -678 4389
rect -594 4213 -560 4389
rect -476 4213 -442 4389
rect -358 4213 -324 4389
rect -653 4119 -619 4153
rect 905 4085 939 4461
rect 1023 4085 1057 4461
rect 1141 4085 1175 4461
rect 1259 4085 1293 4461
rect 1377 4085 1411 4461
rect 1495 4085 1529 4461
rect 1613 4085 1647 4461
rect 2047 4089 2081 4465
rect 2165 4089 2199 4465
rect 2283 4089 2317 4465
rect 2401 4089 2435 4465
rect 2519 4089 2553 4465
rect 2637 4089 2671 4465
rect 2755 4089 2789 4465
rect -771 4002 -737 4036
rect -1183 3576 -1149 3952
rect -1065 3576 -1031 3952
rect -947 3576 -913 3952
rect -830 3776 -796 3952
rect -712 3776 -678 3952
rect 1110 3729 1144 3763
rect 2252 3733 2286 3767
rect -1124 3492 -1090 3526
rect -1006 3492 -972 3526
rect 815 3502 849 3678
rect 933 3502 967 3678
rect 1051 3502 1085 3678
rect 1169 3502 1203 3678
rect 1334 3502 1368 3678
rect 1452 3502 1486 3678
rect 1570 3502 1604 3678
rect 1688 3502 1722 3678
rect 1957 3506 1991 3682
rect 2075 3506 2109 3682
rect 2193 3506 2227 3682
rect 2311 3506 2345 3682
rect 2476 3506 2510 3682
rect 2594 3506 2628 3682
rect 2712 3506 2746 3682
rect 2830 3506 2864 3682
rect -1406 2563 -1372 2739
rect -1288 2563 -1254 2739
rect -1170 2563 -1136 2739
rect -1052 2563 -1018 2739
rect -934 2563 -900 2739
rect -816 2563 -782 2739
rect -698 2563 -664 2739
rect -580 2563 -546 2739
rect -462 2563 -428 2739
rect -344 2563 -310 2739
rect -639 2469 -605 2503
rect -757 2352 -723 2386
rect -1169 1926 -1135 2302
rect -1051 1926 -1017 2302
rect -933 1926 -899 2302
rect -816 2126 -782 2302
rect -698 2126 -664 2302
rect 58 1946 92 2122
rect 176 1946 210 2122
rect 294 1946 328 2122
rect 412 1946 446 2122
rect 542 1946 576 2322
rect 660 1946 694 2322
rect 778 1946 812 2322
rect 896 1946 930 2322
rect 1014 1946 1048 2322
rect 1132 1946 1166 2322
rect 1250 1946 1284 2322
rect 1379 1946 1413 2122
rect 1497 1946 1531 2122
rect 1615 1946 1649 2122
rect 1733 1946 1767 2122
rect 1956 1946 1990 2122
rect 2074 1946 2108 2122
rect 2192 1946 2226 2122
rect 2310 1946 2344 2122
rect 2440 1946 2474 2322
rect 2558 1946 2592 2322
rect 2676 1946 2710 2322
rect 2794 1946 2828 2322
rect 2912 1946 2946 2322
rect 3030 1946 3064 2322
rect 3148 1946 3182 2322
rect 3277 1946 3311 2122
rect 3395 1946 3429 2122
rect 3513 1946 3547 2122
rect 3631 1946 3665 2122
rect -1110 1842 -1076 1876
rect -992 1842 -958 1876
rect 1522 1674 1556 1708
rect 3629 1653 3663 1687
rect 485 1253 519 1629
rect 603 1253 637 1629
rect -1411 959 -1377 1135
rect -1293 959 -1259 1135
rect -1175 959 -1141 1135
rect -1057 959 -1023 1135
rect -939 959 -905 1135
rect -821 959 -787 1135
rect -703 959 -669 1135
rect -585 959 -551 1135
rect -467 959 -433 1135
rect 721 1253 755 1629
rect 839 1253 873 1629
rect 957 1253 991 1629
rect 1075 1253 1109 1629
rect 1193 1253 1227 1629
rect 2383 1253 2417 1629
rect 2501 1253 2535 1629
rect 2619 1253 2653 1629
rect 2737 1253 2771 1629
rect 2855 1253 2889 1629
rect 2973 1253 3007 1629
rect 3091 1253 3125 1629
rect -349 959 -315 1135
rect 515 1031 549 1065
rect 330 964 364 998
rect 1163 1031 1197 1065
rect 2413 1031 2447 1065
rect 781 947 815 981
rect 899 948 933 982
rect 1453 963 1487 997
rect 2228 964 2262 998
rect 3752 1126 3884 1224
rect 3059 1032 3093 1066
rect 2679 947 2713 981
rect 2797 948 2831 982
rect 3351 963 3385 997
rect -644 865 -610 899
rect -762 748 -728 782
rect 183 721 217 897
rect -1174 322 -1140 698
rect -1056 322 -1022 698
rect -938 322 -904 698
rect -821 522 -787 698
rect 301 721 335 897
rect -703 522 -669 698
rect 603 521 637 897
rect 721 521 755 897
rect 839 521 873 897
rect 957 521 991 897
rect 1075 521 1109 897
rect 1481 721 1515 897
rect 1599 721 1633 897
rect 2081 721 2115 897
rect 2199 721 2233 897
rect 2501 521 2535 897
rect 2619 521 2653 897
rect 2737 521 2771 897
rect 2855 521 2889 897
rect 2973 521 3007 897
rect 3379 721 3413 897
rect 3497 721 3531 897
rect -1115 238 -1081 272
rect -997 238 -963 272
<< metal1 >>
rect -1023 4687 -803 4707
rect -1023 4579 -979 4687
rect -847 4579 -803 4687
rect 774 4645 830 4653
rect -1023 4537 -803 4579
rect -152 4637 830 4645
rect -152 4603 790 4637
rect 824 4603 830 4637
rect 1493 4633 1503 4741
rect 1635 4678 1645 4741
rect 1635 4667 1647 4678
rect 1635 4633 1648 4667
rect 1904 4657 1960 4659
rect -152 4587 830 4603
rect 1503 4595 1648 4633
rect -152 4586 827 4587
rect -1419 4507 -442 4537
rect -1419 4401 -1387 4507
rect -1183 4401 -1151 4507
rect -947 4401 -915 4507
rect -711 4401 -679 4507
rect -476 4401 -442 4507
rect -1426 4389 -1380 4401
rect -1426 4213 -1420 4389
rect -1386 4213 -1380 4389
rect -1426 4201 -1380 4213
rect -1308 4389 -1262 4401
rect -1308 4213 -1302 4389
rect -1268 4213 -1262 4389
rect -1308 4201 -1262 4213
rect -1190 4389 -1144 4401
rect -1190 4213 -1184 4389
rect -1150 4213 -1144 4389
rect -1190 4201 -1144 4213
rect -1072 4389 -1026 4401
rect -1072 4213 -1066 4389
rect -1032 4213 -1026 4389
rect -1072 4201 -1026 4213
rect -954 4389 -908 4401
rect -954 4213 -948 4389
rect -914 4213 -908 4389
rect -954 4201 -908 4213
rect -836 4389 -790 4401
rect -836 4213 -830 4389
rect -796 4213 -790 4389
rect -836 4201 -790 4213
rect -718 4389 -672 4401
rect -718 4213 -712 4389
rect -678 4213 -672 4389
rect -718 4201 -672 4213
rect -600 4389 -554 4401
rect -600 4213 -594 4389
rect -560 4213 -554 4389
rect -600 4201 -554 4213
rect -482 4389 -436 4401
rect -482 4213 -476 4389
rect -442 4213 -436 4389
rect -482 4201 -436 4213
rect -364 4389 -318 4401
rect -364 4213 -358 4389
rect -324 4213 -318 4389
rect -364 4201 -318 4213
rect -1303 4107 -1267 4201
rect -1067 4107 -1031 4201
rect -831 4108 -795 4201
rect -669 4153 -603 4160
rect -669 4119 -653 4153
rect -619 4119 -603 4153
rect -669 4108 -603 4119
rect -831 4107 -603 4108
rect -1303 4078 -603 4107
rect -1303 4077 -721 4078
rect -1183 3964 -1149 4077
rect -787 4036 -721 4077
rect -787 4002 -771 4036
rect -737 4002 -721 4036
rect -787 3995 -721 4002
rect -359 3996 -324 4201
rect -152 3996 -85 4586
rect 1607 4563 1648 4595
rect 1894 4591 1904 4657
rect 1960 4591 1970 4657
rect 2640 4633 2650 4741
rect 2782 4678 2792 4741
rect 2782 4667 2794 4678
rect 2782 4633 2795 4667
rect 2650 4595 2795 4633
rect 2754 4567 2795 4595
rect 1023 4535 1293 4563
rect 764 4469 774 4535
rect 840 4469 850 4535
rect 1023 4473 1057 4535
rect 1259 4473 1293 4535
rect 1377 4535 1648 4563
rect 2165 4539 2435 4567
rect 1377 4473 1411 4535
rect 1613 4473 1648 4535
rect 1789 4523 1960 4539
rect 1789 4489 1920 4523
rect 1954 4489 1960 4523
rect 1789 4473 1960 4489
rect 2165 4477 2199 4539
rect 2401 4477 2435 4539
rect 2519 4539 2795 4567
rect 2519 4477 2553 4539
rect 2755 4477 2795 4539
rect 899 4461 945 4473
rect 899 4085 905 4461
rect 939 4085 945 4461
rect 899 4073 945 4085
rect 1017 4461 1063 4473
rect 1017 4085 1023 4461
rect 1057 4085 1063 4461
rect 1017 4073 1063 4085
rect 1135 4461 1181 4473
rect 1135 4085 1141 4461
rect 1175 4085 1181 4461
rect 1135 4073 1181 4085
rect 1253 4461 1299 4473
rect 1253 4085 1259 4461
rect 1293 4085 1299 4461
rect 1253 4073 1299 4085
rect 1371 4461 1417 4473
rect 1371 4085 1377 4461
rect 1411 4085 1417 4461
rect 1371 4073 1417 4085
rect 1489 4461 1535 4473
rect 1489 4085 1495 4461
rect 1529 4085 1535 4461
rect 1489 4073 1535 4085
rect 1607 4461 1653 4473
rect 1607 4085 1613 4461
rect 1647 4085 1653 4461
rect 1607 4073 1653 4085
rect -359 3968 -85 3996
rect -713 3964 -85 3968
rect -1189 3952 -1143 3964
rect -2361 3559 -2072 3734
rect -1189 3576 -1183 3952
rect -1149 3576 -1143 3952
rect -1189 3564 -1143 3576
rect -1071 3952 -1025 3964
rect -1071 3576 -1065 3952
rect -1031 3576 -1025 3952
rect -1071 3564 -1025 3576
rect -953 3952 -907 3964
rect -953 3576 -947 3952
rect -913 3600 -907 3952
rect -836 3952 -790 3964
rect -836 3776 -830 3952
rect -796 3776 -790 3952
rect -836 3764 -790 3776
rect -718 3952 -85 3964
rect -718 3776 -712 3952
rect -678 3939 -85 3952
rect 905 4031 939 4073
rect 1141 4031 1175 4073
rect 905 4003 1175 4031
rect 1259 4032 1293 4073
rect 1495 4032 1529 4073
rect 1259 4003 1529 4032
rect 905 3955 939 4003
rect -678 3776 -672 3939
rect 905 3925 968 3955
rect -718 3764 -672 3776
rect 933 3833 968 3925
rect 933 3797 1160 3833
rect 1430 3822 1440 3919
rect 1539 3822 1549 3919
rect 1613 3890 1647 4073
rect 1613 3836 1722 3890
rect -830 3648 -795 3764
rect 933 3690 968 3797
rect 1094 3763 1160 3797
rect 1094 3729 1110 3763
rect 1144 3729 1160 3763
rect 1441 3821 1538 3822
rect 1441 3754 1498 3821
rect 1094 3723 1160 3729
rect 1335 3718 1604 3754
rect 1335 3690 1368 3718
rect 1571 3690 1604 3718
rect 1688 3690 1722 3836
rect 809 3678 855 3690
rect -699 3648 -591 3658
rect -830 3600 -699 3648
rect -913 3576 -699 3600
rect -953 3564 -699 3576
rect -947 3560 -699 3564
rect -2361 3532 -1311 3559
rect -2361 3526 -1074 3532
rect -2361 3492 -1124 3526
rect -1090 3492 -1074 3526
rect -2361 3476 -1074 3492
rect -1022 3526 -956 3532
rect -1022 3492 -1006 3526
rect -972 3492 -956 3526
rect -773 3516 -699 3560
rect -699 3506 -591 3516
rect -2361 3460 -1311 3476
rect -2361 3459 -1374 3460
rect -2361 3455 -1839 3459
rect -2361 3454 -2072 3455
rect -2344 3044 -2055 3206
rect -2344 2938 -2207 3044
rect -2095 3031 -2055 3044
rect -2095 2938 -2053 3031
rect -2344 2927 -2053 2938
rect -2344 2926 -2055 2927
rect -2344 1932 -2056 2094
rect -2344 1826 -2208 1932
rect -2096 1930 -2056 1932
rect -2090 1919 -2056 1930
rect -2344 1824 -2202 1826
rect -2090 1824 -2055 1919
rect -2344 1815 -2055 1824
rect -2344 1814 -2056 1815
rect -2344 1813 -2088 1814
rect -1932 1561 -1839 3455
rect -1776 3396 -1310 3418
rect -1022 3396 -956 3492
rect 809 3502 815 3678
rect 849 3502 855 3678
rect 809 3490 855 3502
rect 927 3678 973 3690
rect 927 3502 933 3678
rect 967 3502 973 3678
rect 927 3490 973 3502
rect 1045 3678 1091 3690
rect 1045 3502 1051 3678
rect 1085 3502 1091 3678
rect 1045 3490 1091 3502
rect 1163 3678 1209 3690
rect 1163 3502 1169 3678
rect 1203 3623 1209 3678
rect 1328 3678 1374 3690
rect 1328 3623 1334 3678
rect 1203 3535 1334 3623
rect 1203 3502 1209 3535
rect 1163 3490 1209 3502
rect 1328 3502 1334 3535
rect 1368 3502 1374 3678
rect 1328 3490 1374 3502
rect 1446 3678 1492 3690
rect 1446 3502 1452 3678
rect 1486 3502 1492 3678
rect 1446 3490 1492 3502
rect 1564 3678 1610 3690
rect 1564 3502 1570 3678
rect 1604 3502 1610 3678
rect 1564 3490 1610 3502
rect 1682 3678 1728 3690
rect 1682 3502 1688 3678
rect 1722 3502 1728 3678
rect 1682 3490 1728 3502
rect 815 3451 849 3490
rect 1051 3451 1085 3490
rect 815 3416 1085 3451
rect 1452 3452 1485 3490
rect 1688 3452 1721 3490
rect 1452 3416 1721 3452
rect -1776 3348 -956 3396
rect 849 3415 1085 3416
rect -1776 3317 -1310 3348
rect 849 3341 981 3415
rect -1776 3061 -1671 3317
rect 839 3233 849 3341
rect 981 3233 991 3341
rect -1776 2955 -1713 3061
rect -1601 2955 -1591 3061
rect -1009 3037 -789 3057
rect -1776 2944 -1627 2955
rect -1776 1767 -1671 2944
rect -1009 2929 -965 3037
rect -833 2929 -789 3037
rect -1009 2887 -789 2929
rect 1789 2902 1851 4473
rect 2041 4465 2087 4477
rect 2041 4089 2047 4465
rect 2081 4089 2087 4465
rect 2041 4077 2087 4089
rect 2159 4465 2205 4477
rect 2159 4089 2165 4465
rect 2199 4089 2205 4465
rect 2159 4077 2205 4089
rect 2277 4465 2323 4477
rect 2277 4089 2283 4465
rect 2317 4089 2323 4465
rect 2277 4077 2323 4089
rect 2395 4465 2441 4477
rect 2395 4089 2401 4465
rect 2435 4089 2441 4465
rect 2395 4077 2441 4089
rect 2513 4465 2559 4477
rect 2513 4089 2519 4465
rect 2553 4089 2559 4465
rect 2513 4077 2559 4089
rect 2631 4465 2677 4477
rect 2631 4089 2637 4465
rect 2671 4089 2677 4465
rect 2631 4077 2677 4089
rect 2749 4465 2795 4477
rect 2749 4089 2755 4465
rect 2789 4089 2795 4465
rect 2749 4077 2795 4089
rect 2047 4035 2081 4077
rect 2283 4035 2317 4077
rect 2047 4007 2317 4035
rect 2401 4036 2435 4077
rect 2637 4036 2671 4077
rect 2401 4007 2671 4036
rect 2047 3959 2081 4007
rect 2047 3929 2110 3959
rect 2075 3837 2110 3929
rect 2582 3899 2682 3920
rect 2582 3845 2596 3899
rect 2661 3845 2682 3899
rect 2582 3840 2682 3845
rect 2755 3894 2789 4077
rect 2755 3840 2864 3894
rect 2075 3801 2302 3837
rect 2075 3694 2110 3801
rect 2236 3767 2302 3801
rect 2236 3733 2252 3767
rect 2286 3733 2302 3767
rect 2583 3825 2680 3840
rect 2583 3758 2640 3825
rect 2236 3727 2302 3733
rect 2477 3722 2746 3758
rect 2477 3694 2510 3722
rect 2713 3694 2746 3722
rect 2830 3694 2864 3840
rect 3681 3833 3691 3908
rect 3759 3833 3859 3908
rect 3708 3832 3859 3833
rect 1951 3682 1997 3694
rect 1951 3506 1957 3682
rect 1991 3506 1997 3682
rect 1951 3494 1997 3506
rect 2069 3682 2115 3694
rect 2069 3506 2075 3682
rect 2109 3506 2115 3682
rect 2069 3494 2115 3506
rect 2187 3682 2233 3694
rect 2187 3506 2193 3682
rect 2227 3506 2233 3682
rect 2187 3494 2233 3506
rect 2305 3682 2351 3694
rect 2305 3506 2311 3682
rect 2345 3627 2351 3682
rect 2470 3682 2516 3694
rect 2470 3627 2476 3682
rect 2345 3539 2476 3627
rect 2345 3506 2351 3539
rect 2305 3494 2351 3506
rect 2470 3506 2476 3539
rect 2510 3506 2516 3682
rect 2470 3494 2516 3506
rect 2588 3682 2634 3694
rect 2588 3506 2594 3682
rect 2628 3506 2634 3682
rect 2588 3494 2634 3506
rect 2706 3682 2752 3694
rect 2706 3506 2712 3682
rect 2746 3506 2752 3682
rect 2706 3494 2752 3506
rect 2824 3682 2870 3694
rect 2824 3506 2830 3682
rect 2864 3506 2870 3682
rect 2824 3494 2870 3506
rect 1957 3455 1991 3494
rect 2193 3455 2227 3494
rect 1957 3419 2227 3455
rect 2594 3456 2627 3494
rect 2830 3456 2863 3494
rect 2594 3420 2863 3456
rect 1957 3418 2123 3419
rect 1991 3339 2123 3418
rect 1981 3231 1991 3339
rect 2123 3231 2133 3339
rect -1405 2857 -428 2887
rect 1789 2885 1852 2902
rect 1714 2881 1852 2885
rect -1405 2751 -1373 2857
rect -1169 2751 -1137 2857
rect -933 2751 -901 2857
rect -697 2751 -665 2857
rect -462 2751 -428 2857
rect -118 2847 1852 2881
rect -120 2818 1852 2847
rect -120 2802 -74 2818
rect 1714 2816 1852 2818
rect -1412 2739 -1366 2751
rect -1412 2563 -1406 2739
rect -1372 2563 -1366 2739
rect -1412 2551 -1366 2563
rect -1294 2739 -1248 2751
rect -1294 2563 -1288 2739
rect -1254 2563 -1248 2739
rect -1294 2551 -1248 2563
rect -1176 2739 -1130 2751
rect -1176 2563 -1170 2739
rect -1136 2563 -1130 2739
rect -1176 2551 -1130 2563
rect -1058 2739 -1012 2751
rect -1058 2563 -1052 2739
rect -1018 2563 -1012 2739
rect -1058 2551 -1012 2563
rect -940 2739 -894 2751
rect -940 2563 -934 2739
rect -900 2563 -894 2739
rect -940 2551 -894 2563
rect -822 2739 -776 2751
rect -822 2563 -816 2739
rect -782 2563 -776 2739
rect -822 2551 -776 2563
rect -704 2739 -658 2751
rect -704 2563 -698 2739
rect -664 2563 -658 2739
rect -704 2551 -658 2563
rect -586 2739 -540 2751
rect -586 2563 -580 2739
rect -546 2563 -540 2739
rect -586 2551 -540 2563
rect -468 2739 -422 2751
rect -468 2563 -462 2739
rect -428 2563 -422 2739
rect -468 2551 -422 2563
rect -350 2739 -304 2751
rect -350 2563 -344 2739
rect -310 2563 -304 2739
rect -350 2551 -304 2563
rect -1289 2457 -1253 2551
rect -1053 2457 -1017 2551
rect -817 2458 -781 2551
rect -655 2503 -589 2510
rect -655 2469 -639 2503
rect -605 2469 -589 2503
rect -655 2458 -589 2469
rect -817 2457 -589 2458
rect -1289 2428 -589 2457
rect -1289 2427 -707 2428
rect -1169 2314 -1135 2427
rect -773 2386 -707 2427
rect -773 2352 -757 2386
rect -723 2352 -707 2386
rect -773 2345 -707 2352
rect -345 2333 -310 2551
rect -121 2350 -74 2802
rect 838 2586 848 2694
rect 980 2586 990 2694
rect 2736 2586 2746 2694
rect 2878 2586 2888 2694
rect 848 2546 980 2586
rect 2746 2546 2878 2586
rect 847 2480 980 2546
rect 2745 2480 2878 2546
rect 176 2437 1649 2480
rect -121 2334 -75 2350
rect -156 2333 -75 2334
rect -345 2318 -75 2333
rect -699 2314 -75 2318
rect -1175 2302 -1129 2314
rect -1440 1824 -1430 1942
rect -1312 1910 -1302 1942
rect -1175 1926 -1169 2302
rect -1135 1926 -1129 2302
rect -1175 1914 -1129 1926
rect -1057 2302 -1011 2314
rect -1057 1926 -1051 2302
rect -1017 1926 -1011 2302
rect -1057 1914 -1011 1926
rect -939 2302 -893 2314
rect -939 1926 -933 2302
rect -899 1950 -893 2302
rect -822 2302 -776 2314
rect -822 2126 -816 2302
rect -782 2126 -776 2302
rect -822 2114 -776 2126
rect -704 2302 -75 2314
rect -704 2126 -698 2302
rect -664 2290 -75 2302
rect -664 2289 -422 2290
rect -664 2126 -658 2289
rect -156 2288 -75 2290
rect 176 2134 210 2437
rect 542 2334 576 2437
rect 778 2334 812 2437
rect 1014 2334 1048 2437
rect 1250 2334 1284 2437
rect 536 2322 582 2334
rect -704 2114 -658 2126
rect 52 2122 98 2134
rect -816 1998 -781 2114
rect -685 1998 -577 2008
rect -816 1950 -685 1998
rect -899 1926 -685 1950
rect -939 1914 -685 1926
rect -933 1910 -685 1914
rect -1312 1882 -1297 1910
rect -1312 1876 -1060 1882
rect -1312 1842 -1110 1876
rect -1076 1842 -1060 1876
rect -1312 1826 -1060 1842
rect -1008 1876 -942 1882
rect -1008 1842 -992 1876
rect -958 1842 -942 1876
rect -759 1866 -685 1910
rect 52 1946 58 2122
rect 92 1946 98 2122
rect 52 1934 98 1946
rect 170 2122 216 2134
rect 170 1946 176 2122
rect 210 1946 216 2122
rect 170 1934 216 1946
rect 288 2122 334 2134
rect 288 1946 294 2122
rect 328 1946 334 2122
rect 288 1934 334 1946
rect 406 2122 452 2134
rect 536 2122 542 2322
rect 406 1946 412 2122
rect 446 1946 542 2122
rect 576 1946 582 2322
rect 406 1934 452 1946
rect 536 1934 582 1946
rect 654 2322 700 2334
rect 654 1946 660 2322
rect 694 1946 700 2322
rect 654 1934 700 1946
rect 772 2322 818 2334
rect 772 1946 778 2322
rect 812 1946 818 2322
rect 772 1934 818 1946
rect 890 2322 936 2334
rect 890 1946 896 2322
rect 930 1946 936 2322
rect 890 1934 936 1946
rect 1008 2322 1054 2334
rect 1008 1946 1014 2322
rect 1048 1946 1054 2322
rect 1008 1934 1054 1946
rect 1126 2322 1172 2334
rect 1126 1946 1132 2322
rect 1166 1946 1172 2322
rect 1126 1934 1172 1946
rect 1244 2322 1290 2334
rect 1244 1946 1250 2322
rect 1284 2122 1290 2322
rect 1615 2134 1649 2437
rect 2074 2437 3547 2480
rect 2074 2134 2108 2437
rect 2440 2334 2474 2437
rect 2676 2334 2710 2437
rect 2912 2334 2946 2437
rect 3148 2334 3182 2437
rect 2434 2322 2480 2334
rect 1373 2122 1419 2134
rect 1284 1946 1379 2122
rect 1413 1946 1419 2122
rect 1244 1934 1290 1946
rect 1373 1934 1419 1946
rect 1491 2122 1537 2134
rect 1491 1946 1497 2122
rect 1531 1946 1537 2122
rect 1491 1934 1537 1946
rect 1609 2122 1655 2134
rect 1609 1946 1615 2122
rect 1649 1946 1655 2122
rect 1609 1934 1655 1946
rect 1727 2122 1773 2134
rect 1727 1946 1733 2122
rect 1767 1946 1773 2122
rect 1727 1934 1773 1946
rect 1950 2122 1996 2134
rect 1950 1946 1956 2122
rect 1990 1946 1996 2122
rect 1950 1934 1996 1946
rect 2068 2122 2114 2134
rect 2068 1946 2074 2122
rect 2108 1946 2114 2122
rect 2068 1934 2114 1946
rect 2186 2122 2232 2134
rect 2186 1946 2192 2122
rect 2226 1946 2232 2122
rect 2186 1934 2232 1946
rect 2304 2122 2350 2134
rect 2434 2122 2440 2322
rect 2304 1946 2310 2122
rect 2344 1946 2440 2122
rect 2474 1946 2480 2322
rect 2304 1934 2350 1946
rect 2434 1934 2480 1946
rect 2552 2322 2598 2334
rect 2552 1946 2558 2322
rect 2592 1946 2598 2322
rect 2552 1934 2598 1946
rect 2670 2322 2716 2334
rect 2670 1946 2676 2322
rect 2710 1946 2716 2322
rect 2670 1934 2716 1946
rect 2788 2322 2834 2334
rect 2788 1946 2794 2322
rect 2828 1946 2834 2322
rect 2788 1934 2834 1946
rect 2906 2322 2952 2334
rect 2906 1946 2912 2322
rect 2946 1946 2952 2322
rect 2906 1934 2952 1946
rect 3024 2322 3070 2334
rect 3024 1946 3030 2322
rect 3064 1946 3070 2322
rect 3024 1934 3070 1946
rect 3142 2322 3188 2334
rect 3142 1946 3148 2322
rect 3182 2122 3188 2322
rect 3513 2134 3547 2437
rect 3271 2122 3317 2134
rect 3182 1946 3277 2122
rect 3311 1946 3317 2122
rect 3142 1934 3188 1946
rect 3271 1934 3317 1946
rect 3389 2122 3435 2134
rect 3389 1946 3395 2122
rect 3429 1946 3435 2122
rect 3389 1934 3435 1946
rect 3507 2122 3553 2134
rect 3507 1946 3513 2122
rect 3547 1946 3553 2122
rect 3507 1934 3553 1946
rect 3625 2122 3671 2134
rect 3625 1946 3631 2122
rect 3665 1946 3671 2122
rect 3625 1934 3671 1946
rect -685 1856 -577 1866
rect 58 1900 92 1934
rect 660 1900 694 1934
rect 896 1900 930 1934
rect 58 1865 217 1900
rect 660 1865 930 1900
rect 1497 1900 1531 1934
rect 1733 1900 1767 1934
rect 1497 1865 1767 1900
rect 1956 1900 1990 1934
rect 2558 1900 2592 1934
rect 2794 1900 2828 1934
rect 1956 1865 2115 1900
rect 2558 1865 2828 1900
rect 3395 1900 3429 1934
rect 3631 1900 3665 1934
rect 3395 1865 3665 1900
rect -1312 1824 -1297 1826
rect -1397 1810 -1297 1824
rect -1397 1767 -1297 1768
rect -1776 1746 -1297 1767
rect -1008 1746 -942 1842
rect -1776 1698 -942 1746
rect -1776 1669 -1297 1698
rect -1776 1667 -1671 1669
rect -1397 1668 -1297 1669
rect -1943 1482 -1933 1561
rect -1840 1482 -1830 1561
rect -1932 308 -1839 1482
rect -1014 1433 -794 1453
rect -1014 1325 -970 1433
rect -838 1325 -794 1433
rect -1014 1283 -794 1325
rect -1410 1253 -433 1283
rect -1410 1147 -1378 1253
rect -1174 1147 -1142 1253
rect -938 1147 -906 1253
rect -702 1147 -670 1253
rect -467 1147 -433 1253
rect -1417 1135 -1371 1147
rect -1417 959 -1411 1135
rect -1377 959 -1371 1135
rect -1417 947 -1371 959
rect -1299 1135 -1253 1147
rect -1299 959 -1293 1135
rect -1259 959 -1253 1135
rect -1299 947 -1253 959
rect -1181 1135 -1135 1147
rect -1181 959 -1175 1135
rect -1141 959 -1135 1135
rect -1181 947 -1135 959
rect -1063 1135 -1017 1147
rect -1063 959 -1057 1135
rect -1023 959 -1017 1135
rect -1063 947 -1017 959
rect -945 1135 -899 1147
rect -945 959 -939 1135
rect -905 959 -899 1135
rect -945 947 -899 959
rect -827 1135 -781 1147
rect -827 959 -821 1135
rect -787 959 -781 1135
rect -827 947 -781 959
rect -709 1135 -663 1147
rect -709 959 -703 1135
rect -669 959 -663 1135
rect -709 947 -663 959
rect -591 1135 -545 1147
rect -591 959 -585 1135
rect -551 959 -545 1135
rect -591 947 -545 959
rect -473 1135 -427 1147
rect -473 959 -467 1135
rect -433 959 -427 1135
rect -473 947 -427 959
rect -355 1135 -309 1147
rect -355 959 -349 1135
rect -315 959 -309 1135
rect -355 947 -309 959
rect 183 1081 217 1865
rect 896 1803 930 1865
rect 485 1765 1227 1803
rect 485 1641 519 1765
rect 721 1641 755 1765
rect 957 1641 991 1765
rect 1193 1641 1227 1765
rect 1483 1658 1493 1724
rect 1556 1658 1566 1724
rect 479 1629 525 1641
rect 479 1253 485 1629
rect 519 1253 525 1629
rect 479 1241 525 1253
rect 597 1629 643 1641
rect 597 1253 603 1629
rect 637 1253 643 1629
rect 597 1241 643 1253
rect 715 1629 761 1641
rect 715 1253 721 1629
rect 755 1253 761 1629
rect 715 1241 761 1253
rect 833 1629 879 1641
rect 833 1253 839 1629
rect 873 1253 879 1629
rect 833 1241 879 1253
rect 951 1629 997 1641
rect 951 1253 957 1629
rect 991 1253 997 1629
rect 951 1241 997 1253
rect 1069 1629 1115 1641
rect 1069 1253 1075 1629
rect 1109 1253 1115 1629
rect 1069 1241 1115 1253
rect 1187 1629 1233 1641
rect 1187 1253 1193 1629
rect 1227 1253 1233 1629
rect 1187 1241 1233 1253
rect 1599 1082 1633 1865
rect 1326 1081 1633 1082
rect 183 1076 499 1081
rect 1213 1076 1633 1081
rect 183 1065 566 1076
rect 183 1038 515 1065
rect -1294 853 -1258 947
rect -1058 853 -1022 947
rect -822 854 -786 947
rect -660 899 -594 906
rect -660 865 -644 899
rect -610 865 -594 899
rect -660 854 -594 865
rect -822 853 -594 854
rect -1294 824 -594 853
rect -1294 823 -712 824
rect -1174 710 -1140 823
rect -778 782 -712 823
rect -778 748 -762 782
rect -728 748 -712 782
rect -778 741 -712 748
rect -350 714 -315 947
rect 183 909 217 1038
rect 499 1031 515 1038
rect 549 1031 566 1065
rect 499 1025 566 1031
rect 1146 1065 1633 1076
rect 1146 1031 1163 1065
rect 1197 1038 1633 1065
rect 1197 1031 1213 1038
rect 1326 1037 1633 1038
rect 1146 1025 1213 1031
rect 324 998 380 1010
rect 324 964 330 998
rect 364 997 380 998
rect 1437 997 1493 1009
rect 364 981 831 997
rect 364 964 781 981
rect 324 948 781 964
rect 765 947 781 948
rect 815 947 831 981
rect 765 940 831 947
rect 883 982 1453 997
rect 883 948 899 982
rect 933 963 1453 982
rect 1487 963 1493 997
rect 933 948 1493 963
rect 883 938 950 948
rect 1437 947 1493 948
rect 1599 909 1633 1037
rect 2081 1081 2115 1865
rect 2794 1803 2828 1865
rect 2383 1765 3125 1803
rect 2383 1641 2417 1765
rect 2619 1641 2653 1765
rect 2855 1641 2889 1765
rect 3091 1641 3125 1765
rect 2377 1629 2423 1641
rect 2377 1253 2383 1629
rect 2417 1253 2423 1629
rect 2377 1241 2423 1253
rect 2495 1629 2541 1641
rect 2495 1253 2501 1629
rect 2535 1253 2541 1629
rect 2495 1241 2541 1253
rect 2613 1629 2659 1641
rect 2613 1253 2619 1629
rect 2653 1253 2659 1629
rect 2613 1241 2659 1253
rect 2731 1629 2777 1641
rect 2731 1253 2737 1629
rect 2771 1253 2777 1629
rect 2731 1241 2777 1253
rect 2849 1629 2895 1641
rect 2849 1253 2855 1629
rect 2889 1253 2895 1629
rect 2849 1241 2895 1253
rect 2967 1629 3013 1641
rect 2967 1253 2973 1629
rect 3007 1253 3013 1629
rect 2967 1241 3013 1253
rect 3085 1629 3131 1641
rect 3085 1253 3091 1629
rect 3125 1253 3131 1629
rect 3085 1241 3131 1253
rect 3497 1082 3531 1865
rect 3109 1081 3178 1082
rect 3224 1081 3531 1082
rect 2081 1076 2397 1081
rect 3109 1077 3531 1081
rect 2081 1065 2464 1076
rect 2081 1038 2413 1065
rect 2081 909 2115 1038
rect 2397 1031 2413 1038
rect 2447 1031 2464 1065
rect 2397 1025 2464 1031
rect 3042 1066 3531 1077
rect 3042 1032 3059 1066
rect 3093 1038 3531 1066
rect 3093 1032 3109 1038
rect 3224 1037 3531 1038
rect 3042 1026 3109 1032
rect 2222 998 2278 1010
rect 2222 964 2228 998
rect 2262 997 2278 998
rect 3335 997 3391 1009
rect 2262 981 2729 997
rect 2262 964 2679 981
rect 2222 948 2679 964
rect 2663 947 2679 948
rect 2713 947 2729 981
rect 2663 940 2729 947
rect 2781 982 3351 997
rect 2781 948 2797 982
rect 2831 963 3351 982
rect 3385 963 3391 997
rect 2831 948 3391 963
rect 2781 938 2848 948
rect 3335 947 3391 948
rect 3497 909 3531 1037
rect 3612 1687 3679 1711
rect 3612 1653 3629 1687
rect 3663 1653 3679 1687
rect -704 710 -315 714
rect -1180 698 -1134 710
rect -1180 322 -1174 698
rect -1140 322 -1134 698
rect -1180 310 -1134 322
rect -1062 698 -1016 710
rect -1062 322 -1056 698
rect -1022 322 -1016 698
rect -1062 310 -1016 322
rect -944 698 -898 710
rect -944 322 -938 698
rect -904 346 -898 698
rect -827 698 -781 710
rect -827 522 -821 698
rect -787 522 -781 698
rect -827 510 -781 522
rect -709 698 -315 710
rect 177 897 223 909
rect 177 721 183 897
rect 217 721 223 897
rect 177 709 223 721
rect 295 897 341 909
rect 295 721 301 897
rect 335 721 341 897
rect 295 709 341 721
rect 597 897 643 909
rect -709 522 -703 698
rect -669 685 -315 698
rect -669 522 -663 685
rect -393 682 -315 685
rect -393 630 -383 682
rect -320 630 -310 682
rect -388 624 -315 630
rect -709 510 -663 522
rect -821 394 -786 510
rect 300 415 334 709
rect 597 521 603 897
rect 637 521 643 897
rect 597 509 643 521
rect 715 897 761 909
rect 715 521 721 897
rect 755 521 761 897
rect 715 509 761 521
rect 833 897 879 909
rect 833 521 839 897
rect 873 521 879 897
rect 833 509 879 521
rect 951 897 997 909
rect 951 521 957 897
rect 991 521 997 897
rect 951 509 997 521
rect 1069 897 1115 909
rect 1069 521 1075 897
rect 1109 521 1115 897
rect 1475 897 1521 909
rect 1475 721 1481 897
rect 1515 721 1521 897
rect 1475 709 1521 721
rect 1593 897 1639 909
rect 1593 721 1599 897
rect 1633 721 1639 897
rect 1593 709 1639 721
rect 2075 897 2121 909
rect 2075 721 2081 897
rect 2115 721 2121 897
rect 2075 709 2121 721
rect 2193 897 2239 909
rect 2193 721 2199 897
rect 2233 721 2239 897
rect 2193 709 2239 721
rect 2495 897 2541 909
rect 1069 509 1115 521
rect 957 415 991 509
rect 1481 415 1514 709
rect -690 394 -582 404
rect -821 346 -690 394
rect -904 322 -690 346
rect -944 310 -690 322
rect -1932 306 -1347 308
rect -938 306 -690 310
rect -1932 278 -1302 306
rect -1932 272 -1065 278
rect -1932 238 -1115 272
rect -1081 238 -1065 272
rect -1932 222 -1065 238
rect -1013 272 -947 278
rect -1013 238 -997 272
rect -963 238 -947 272
rect -764 262 -690 306
rect 300 383 1514 415
rect 2198 415 2232 709
rect 2495 521 2501 897
rect 2535 521 2541 897
rect 2495 509 2541 521
rect 2613 897 2659 909
rect 2613 521 2619 897
rect 2653 521 2659 897
rect 2613 509 2659 521
rect 2731 897 2777 909
rect 2731 521 2737 897
rect 2771 521 2777 897
rect 2731 509 2777 521
rect 2849 897 2895 909
rect 2849 521 2855 897
rect 2889 521 2895 897
rect 2849 509 2895 521
rect 2967 897 3013 909
rect 2967 521 2973 897
rect 3007 521 3013 897
rect 3373 897 3419 909
rect 3373 721 3379 897
rect 3413 721 3419 897
rect 3373 709 3419 721
rect 3491 897 3537 909
rect 3491 721 3497 897
rect 3531 721 3537 897
rect 3491 709 3537 721
rect 2967 509 3013 521
rect 2855 415 2889 509
rect 3379 415 3412 709
rect 2198 383 3412 415
rect 793 298 925 383
rect 2691 298 2823 383
rect -690 252 -582 262
rect -1932 206 -1302 222
rect -1932 202 -1347 206
rect -1932 201 -1831 202
rect -1402 153 -1302 164
rect -1438 47 -1428 153
rect -1316 142 -1302 153
rect -1013 142 -947 238
rect 783 190 793 298
rect 925 190 935 298
rect 2681 190 2691 298
rect 2823 190 2833 298
rect 3612 270 3679 1653
rect 3740 1224 3896 1230
rect 3740 1126 3752 1224
rect 3884 1126 3896 1224
rect 3740 1120 3896 1126
rect -1316 94 -947 142
rect -1316 64 -1302 94
rect -1316 47 -1306 64
rect -1014 -9 -948 94
rect 3612 -9 3678 270
rect -1016 -89 3678 -9
<< via1 >>
rect -979 4579 -847 4687
rect 1503 4633 1635 4741
rect 1904 4643 1960 4657
rect 1904 4609 1920 4643
rect 1920 4609 1954 4643
rect 1954 4609 1960 4643
rect 1904 4591 1960 4609
rect 2650 4633 2782 4741
rect 774 4519 840 4535
rect 774 4485 790 4519
rect 790 4485 824 4519
rect 824 4485 840 4519
rect 774 4469 840 4485
rect 1440 3822 1539 3919
rect -699 3516 -591 3648
rect -2207 2938 -2095 3044
rect -2208 1930 -2096 1932
rect -2208 1826 -2090 1930
rect -2202 1824 -2090 1826
rect 849 3233 981 3341
rect -1713 2955 -1601 3061
rect -965 2929 -833 3037
rect 2596 3845 2661 3899
rect 3691 3833 3759 3908
rect 1991 3231 2123 3339
rect 848 2586 980 2694
rect 2746 2586 2878 2694
rect -1430 1824 -1312 1942
rect -685 1866 -577 1998
rect -1933 1482 -1840 1561
rect -970 1325 -838 1433
rect 1493 1708 1556 1724
rect 1493 1674 1522 1708
rect 1522 1674 1556 1708
rect 1493 1658 1556 1674
rect -383 630 -320 682
rect -690 262 -582 394
rect -1428 47 -1316 153
rect 793 190 925 298
rect 2691 190 2823 298
<< metal2 >>
rect 1492 4752 1645 4762
rect -990 4698 -837 4708
rect 2639 4752 2792 4762
rect 1904 4657 1960 4667
rect 1492 4613 1645 4623
rect -990 4559 -837 4569
rect 1779 4591 1904 4653
rect 1960 4591 1961 4653
rect 2639 4613 2792 4623
rect 774 4542 840 4545
rect -152 4535 840 4542
rect -152 4469 774 4535
rect -719 3506 -709 3659
rect -580 3506 -570 3659
rect -2219 3071 -2052 3072
rect -1712 3071 -1596 3072
rect -2219 3061 -1596 3071
rect -2219 3044 -1713 3061
rect -2219 2938 -2207 3044
rect -2095 2955 -1713 3044
rect -1601 2955 -1596 3061
rect -2095 2938 -1596 2955
rect -2219 2929 -1596 2938
rect -976 3048 -823 3058
rect -976 2909 -823 2919
rect -2220 1950 -2055 1960
rect -2220 1949 -2052 1950
rect -1430 1949 -1312 1952
rect -2220 1942 -1312 1949
rect -2220 1932 -1430 1942
rect -2220 1826 -2208 1932
rect -2096 1930 -1430 1932
rect -2220 1824 -2202 1826
rect -2090 1824 -1430 1930
rect -705 1856 -695 2009
rect -566 1856 -556 2009
rect -2220 1817 -1312 1824
rect -2214 1815 -1312 1817
rect -2177 1814 -1312 1815
rect -1943 1570 -1828 1580
rect -1943 1463 -1828 1473
rect -1433 163 -1317 1814
rect -981 1444 -828 1454
rect -981 1305 -828 1315
rect -383 686 -320 692
rect -152 686 -84 4469
rect 774 4459 840 4469
rect 1779 3930 1839 4591
rect 1904 4581 1960 4591
rect 1701 3929 1839 3930
rect 1439 3919 1839 3929
rect 1439 3822 1440 3919
rect 1539 3822 1839 3919
rect 2596 3908 2661 3909
rect 3691 3908 3759 3918
rect 2595 3899 3691 3908
rect 2595 3845 2596 3899
rect 2661 3845 3691 3899
rect 2595 3834 3691 3845
rect 3691 3823 3759 3833
rect 1439 3814 1839 3822
rect 1439 3810 1748 3814
rect 839 3351 992 3361
rect 839 3212 992 3222
rect 1981 3349 2134 3359
rect 1981 3210 2134 3220
rect 837 2705 990 2715
rect 837 2566 990 2576
rect 2735 2705 2888 2715
rect 2735 2566 2888 2576
rect 1478 1734 1556 1744
rect 1478 1638 1556 1648
rect -388 682 -84 686
rect -388 630 -383 682
rect -320 630 -84 682
rect -388 624 -84 630
rect -383 620 -320 624
rect -710 252 -700 405
rect -571 252 -561 405
rect 783 308 936 318
rect 783 169 936 179
rect 2681 308 2834 318
rect 2681 169 2834 179
rect -1433 153 -1316 163
rect -1433 47 -1428 153
rect -1433 37 -1316 47
rect -1433 36 -1317 37
<< via2 >>
rect 1492 4741 1645 4752
rect -990 4687 -837 4698
rect -990 4579 -979 4687
rect -979 4579 -847 4687
rect -847 4579 -837 4687
rect 1492 4633 1503 4741
rect 1503 4633 1635 4741
rect 1635 4633 1645 4741
rect 2639 4741 2792 4752
rect 1492 4623 1645 4633
rect -990 4569 -837 4579
rect 2639 4633 2650 4741
rect 2650 4633 2782 4741
rect 2782 4633 2792 4741
rect 2639 4623 2792 4633
rect -709 3648 -580 3659
rect -709 3516 -699 3648
rect -699 3516 -591 3648
rect -591 3516 -580 3648
rect -709 3506 -580 3516
rect -976 3037 -823 3048
rect -976 2929 -965 3037
rect -965 2929 -833 3037
rect -833 2929 -823 3037
rect -976 2919 -823 2929
rect -695 1998 -566 2009
rect -695 1866 -685 1998
rect -685 1866 -577 1998
rect -577 1866 -566 1998
rect -695 1856 -566 1866
rect -1943 1561 -1828 1570
rect -1943 1482 -1933 1561
rect -1933 1482 -1840 1561
rect -1840 1482 -1828 1561
rect -1943 1473 -1828 1482
rect -981 1433 -828 1444
rect -981 1325 -970 1433
rect -970 1325 -838 1433
rect -838 1325 -828 1433
rect -981 1315 -828 1325
rect 839 3341 992 3351
rect 839 3233 849 3341
rect 849 3233 981 3341
rect 981 3233 992 3341
rect 839 3222 992 3233
rect 1981 3339 2134 3349
rect 1981 3231 1991 3339
rect 1991 3231 2123 3339
rect 2123 3231 2134 3339
rect 1981 3220 2134 3231
rect 837 2694 990 2705
rect 837 2586 848 2694
rect 848 2586 980 2694
rect 980 2586 990 2694
rect 837 2576 990 2586
rect 2735 2694 2888 2705
rect 2735 2586 2746 2694
rect 2746 2586 2878 2694
rect 2878 2586 2888 2694
rect 2735 2576 2888 2586
rect 1478 1724 1556 1734
rect 1478 1658 1493 1724
rect 1493 1658 1556 1724
rect 1478 1648 1556 1658
rect -700 394 -571 405
rect -700 262 -690 394
rect -690 262 -582 394
rect -582 262 -571 394
rect -700 252 -571 262
rect 783 298 936 308
rect 783 190 793 298
rect 793 190 925 298
rect 925 190 936 298
rect 783 179 936 190
rect 2681 298 2834 308
rect 2681 190 2691 298
rect 2691 190 2823 298
rect 2823 190 2834 298
rect 2681 179 2834 190
<< metal3 >>
rect -1022 4550 -1012 4729
rect -813 4550 -803 4729
rect 1460 4604 1470 4783
rect 1669 4604 1679 4783
rect 2607 4604 2617 4783
rect 2816 4604 2826 4783
rect -728 3681 -549 3691
rect -728 3473 -549 3482
rect 806 3191 815 3370
rect 1014 3191 1024 3370
rect 1948 3189 1957 3368
rect 2156 3189 2166 3368
rect -1008 2900 -998 3079
rect -799 2900 -789 3079
rect 805 2557 815 2736
rect 1014 2557 1024 2736
rect 2703 2557 2713 2736
rect 2912 2557 2922 2736
rect -714 2031 -535 2041
rect -714 1823 -535 1832
rect -1932 1738 -1840 1739
rect 1466 1738 1570 1740
rect -1932 1734 1570 1738
rect -1932 1648 1478 1734
rect 1556 1648 1570 1734
rect -1932 1635 1570 1648
rect -1932 1575 -1840 1635
rect -1953 1570 -1818 1575
rect -1953 1473 -1943 1570
rect -1828 1473 -1818 1570
rect -1953 1468 -1818 1473
rect -1013 1296 -1003 1475
rect -804 1296 -794 1475
rect -719 427 -540 437
rect -719 219 -540 228
rect 749 148 759 327
rect 958 148 968 327
rect 2647 148 2657 327
rect 2856 148 2866 327
<< via3 >>
rect -1012 4698 -813 4729
rect -1012 4569 -990 4698
rect -990 4569 -837 4698
rect -837 4569 -813 4698
rect -1012 4550 -813 4569
rect 1470 4752 1669 4783
rect 1470 4623 1492 4752
rect 1492 4623 1645 4752
rect 1645 4623 1669 4752
rect 1470 4604 1669 4623
rect 2617 4752 2816 4783
rect 2617 4623 2639 4752
rect 2639 4623 2792 4752
rect 2792 4623 2816 4752
rect 2617 4604 2816 4623
rect -728 3659 -549 3681
rect -728 3506 -709 3659
rect -709 3506 -580 3659
rect -580 3506 -549 3659
rect -728 3482 -549 3506
rect 815 3351 1014 3370
rect 815 3222 839 3351
rect 839 3222 992 3351
rect 992 3222 1014 3351
rect 815 3191 1014 3222
rect 1957 3349 2156 3368
rect 1957 3220 1981 3349
rect 1981 3220 2134 3349
rect 2134 3220 2156 3349
rect 1957 3189 2156 3220
rect -998 3048 -799 3079
rect -998 2919 -976 3048
rect -976 2919 -823 3048
rect -823 2919 -799 3048
rect -998 2900 -799 2919
rect 815 2705 1014 2736
rect 815 2576 837 2705
rect 837 2576 990 2705
rect 990 2576 1014 2705
rect 815 2557 1014 2576
rect 2713 2705 2912 2736
rect 2713 2576 2735 2705
rect 2735 2576 2888 2705
rect 2888 2576 2912 2705
rect 2713 2557 2912 2576
rect -714 2009 -535 2031
rect -714 1856 -695 2009
rect -695 1856 -566 2009
rect -566 1856 -535 2009
rect -714 1832 -535 1856
rect -1003 1444 -804 1475
rect -1003 1315 -981 1444
rect -981 1315 -828 1444
rect -828 1315 -804 1444
rect -1003 1296 -804 1315
rect -719 405 -540 427
rect -719 252 -700 405
rect -700 252 -571 405
rect -571 252 -540 405
rect -719 228 -540 252
rect 759 308 958 327
rect 759 179 783 308
rect 783 179 936 308
rect 936 179 958 308
rect 759 148 958 179
rect 2657 308 2856 327
rect 2657 179 2681 308
rect 2681 179 2834 308
rect 2834 179 2856 308
rect 2657 148 2856 179
<< metal4 >>
rect -1034 4889 3399 5054
rect -1033 4783 3395 4889
rect -1033 4729 1470 4783
rect -1033 4550 -1012 4729
rect -813 4604 1470 4729
rect 1669 4604 2617 4783
rect 2816 4604 3395 4783
rect -813 4550 3395 4604
rect -1033 4344 3395 4550
rect -1553 3079 -658 3293
rect -1553 2900 -998 3079
rect -799 2911 -658 3079
rect -799 2906 -313 2911
rect 1565 2906 1912 2909
rect 2779 2906 3395 4344
rect -799 2900 3395 2906
rect -1553 2736 3395 2900
rect -1553 2557 815 2736
rect 1014 2557 2713 2736
rect 2912 2557 3395 2736
rect -1553 2401 3395 2557
rect -1553 1671 -1383 2401
rect 2779 2396 3395 2401
rect -1553 1475 -285 1671
rect -1553 1296 -1003 1475
rect -804 1296 -285 1475
rect -1553 1027 -285 1296
rect 735 327 980 330
rect 735 309 759 327
rect 958 309 980 327
rect 2633 327 2878 330
rect 2633 309 2657 327
rect 2856 309 2878 327
rect 631 5 655 242
rect 1165 5 2501 191
rect 631 0 2998 5
rect 1019 -2 2690 0
<< via4 >>
rect -787 3681 -277 3759
rect -787 3482 -728 3681
rect -728 3482 -549 3681
rect -549 3482 -277 3681
rect -787 3455 -277 3482
rect 781 3370 1085 3521
rect 781 3191 815 3370
rect 815 3191 1014 3370
rect 1014 3191 1085 3370
rect 781 3011 1085 3191
rect 1915 3368 2219 3531
rect 1915 3189 1957 3368
rect 1957 3189 2156 3368
rect 2156 3189 2219 3368
rect 1915 3021 2219 3189
rect -793 2031 -283 2099
rect -793 1832 -714 2031
rect -714 1832 -535 2031
rect -535 1832 -283 2031
rect -793 1795 -283 1832
rect -794 427 -284 494
rect -794 228 -719 427
rect -719 228 -540 427
rect -540 228 -284 427
rect -794 190 -284 228
rect 655 148 759 309
rect 759 148 958 309
rect 958 148 1165 309
rect 655 5 1165 148
rect 2501 148 2657 309
rect 2657 148 2856 309
rect 2856 148 3011 309
rect 2501 5 3011 148
<< metal5 >>
rect -938 3759 3036 3923
rect -938 3455 -787 3759
rect -277 3531 3036 3759
rect -277 3521 1915 3531
rect -277 3455 781 3521
rect -938 3011 781 3455
rect 1085 3021 1915 3521
rect 2219 3021 3036 3531
rect 1085 3011 3036 3021
rect -938 2099 3036 3011
rect -938 1795 -793 2099
rect -283 1795 3036 2099
rect -938 494 3036 1795
rect -938 190 -794 494
rect -284 309 3036 494
rect -284 190 655 309
rect -938 5 655 190
rect 1165 5 2501 309
rect 3011 5 3036 309
rect -938 -464 3036 5
<< labels >>
flabel metal4 -326 4738 1080 5035 1 FreeSans 1200 0 0 0 VDD
port 1 n
flabel metal5 -332 -431 1079 -151 1 FreeSans 1200 0 0 0 VSS
port 2 n
flabel metal1 -2345 3479 -2095 3706 1 FreeSans 400 0 0 0 A
port 3 n
flabel metal1 -2327 2944 -2075 3182 1 FreeSans 400 0 0 0 B
port 4 n
flabel metal1 -2332 1830 -2070 2075 1 FreeSans 240 0 0 0 carry_in
port 5 n
flabel metal1 3722 3839 3846 3900 1 FreeSans 240 0 0 0 carry_out
port 6 n
flabel viali 3752 1126 3884 1224 1 FreeSans 400 0 0 0 Y
port 7 n
<< end >>
