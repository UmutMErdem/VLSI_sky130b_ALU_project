magic
tech sky130B
magscale 1 2
timestamp 1736091534
<< nwell >>
rect 3806 5396 4093 5397
rect 4953 5396 5188 5397
rect 1324 5342 1564 5343
rect 1321 5109 1564 5342
rect 1321 4927 1565 5109
rect 3803 4999 4093 5396
rect 4780 5003 5262 5396
rect 10319 5393 10606 5394
rect 11466 5393 11701 5394
rect 7837 5339 8077 5340
rect 883 4603 2075 4927
rect 3208 4532 4093 4999
rect 3208 4479 4094 4532
rect 4350 4479 5262 5003
rect 7834 5106 8077 5339
rect 7834 4924 8078 5106
rect 10316 4996 10606 5393
rect 11293 5000 11775 5393
rect 23411 5392 23698 5393
rect 24558 5392 24793 5393
rect 16853 5388 17140 5389
rect 18000 5388 18235 5389
rect 14371 5334 14611 5335
rect 7396 4600 8588 4924
rect 3208 4475 4095 4479
rect 3637 4190 4095 4475
rect 4780 4220 5262 4479
rect 9721 4529 10606 4996
rect 9721 4476 10607 4529
rect 10863 4476 11775 5000
rect 14368 5101 14611 5334
rect 14368 4919 14612 5101
rect 16850 4991 17140 5388
rect 17827 4995 18309 5388
rect 20929 5338 21169 5339
rect 13930 4595 15122 4919
rect 9721 4472 10608 4476
rect 3637 3892 4121 4190
rect 4779 3896 5263 4220
rect 10150 4187 10608 4472
rect 11293 4217 11775 4476
rect 16255 4524 17140 4991
rect 16255 4471 17141 4524
rect 17397 4471 18309 4995
rect 20926 5105 21169 5338
rect 20926 4923 21170 5105
rect 23408 4995 23698 5392
rect 24385 4999 24867 5392
rect 20488 4599 21680 4923
rect 22813 4528 23698 4995
rect 22813 4475 23699 4528
rect 23955 4475 24867 4999
rect 22813 4471 23700 4475
rect 16255 4467 17142 4471
rect 10150 3889 10634 4187
rect 11292 3893 11776 4217
rect 16684 4182 17142 4467
rect 17827 4212 18309 4471
rect 16684 3884 17168 4182
rect 17826 3888 18310 4212
rect 23242 4186 23700 4471
rect 24385 4216 24867 4475
rect 23242 3888 23726 4186
rect 24384 3892 24868 4216
rect 1338 3692 1578 3693
rect 1335 3459 1578 3692
rect 7851 3689 8091 3690
rect 1335 3277 1579 3459
rect 7848 3456 8091 3689
rect 20943 3688 21183 3689
rect 14385 3684 14625 3685
rect 897 2953 2089 3277
rect 5049 2860 5277 3350
rect 7848 3274 8092 3456
rect 14382 3451 14625 3684
rect 20940 3455 21183 3688
rect 7410 2950 8602 3274
rect 2360 2660 3683 2860
rect 4743 2660 5581 2860
rect 11562 2857 11790 3347
rect 14382 3269 14626 3451
rect 13944 2945 15136 3269
rect 2360 2336 6064 2660
rect 8873 2657 10196 2857
rect 11256 2657 12094 2857
rect 18096 2852 18324 3342
rect 20940 3273 21184 3455
rect 20502 2949 21694 3273
rect 24654 2856 24882 3346
rect 1333 2088 1573 2089
rect 1330 1855 1573 2088
rect 1330 1673 1574 1855
rect 892 1349 2084 1673
rect 2788 1643 3626 2336
rect 4686 1643 5524 2336
rect 8873 2333 12577 2657
rect 15407 2652 16730 2852
rect 17790 2652 18628 2852
rect 21965 2656 23288 2856
rect 24348 2656 25186 2856
rect 7846 2085 8086 2086
rect 7843 1852 8086 2085
rect 7843 1670 8087 1852
rect 7405 1346 8597 1670
rect 9301 1640 10139 2333
rect 11199 1640 12037 2333
rect 15407 2328 19111 2652
rect 21965 2332 25669 2656
rect 14380 2080 14620 2081
rect 14377 1847 14620 2080
rect 14377 1665 14621 1847
rect 13939 1341 15131 1665
rect 15835 1635 16673 2328
rect 17733 1635 18571 2328
rect 20938 2084 21178 2085
rect 20935 1851 21178 2084
rect 20935 1669 21179 1851
rect 20497 1345 21689 1669
rect 22393 1639 23231 2332
rect 24291 1639 25129 2332
rect 20499 -208 20734 -207
rect 21594 -208 21881 -207
rect 13986 -211 14221 -210
rect 15081 -211 15368 -210
rect 894 -212 1129 -211
rect 1989 -212 2276 -211
rect 820 -605 1302 -212
rect 820 -1129 1732 -605
rect 1989 -609 2279 -212
rect 7452 -216 7687 -215
rect 8547 -216 8834 -215
rect 4518 -266 4758 -265
rect 4518 -499 4761 -266
rect 1989 -1076 2874 -609
rect 4517 -681 4761 -499
rect 7378 -609 7860 -216
rect 4007 -1005 5199 -681
rect 1988 -1129 2874 -1076
rect 820 -1388 1302 -1129
rect 1987 -1133 2874 -1129
rect 7378 -1133 8290 -609
rect 8547 -613 8837 -216
rect 11076 -270 11316 -269
rect 11076 -503 11319 -270
rect 8547 -1080 9432 -613
rect 11075 -685 11319 -503
rect 13912 -604 14394 -211
rect 10565 -1009 11757 -685
rect 8546 -1133 9432 -1080
rect 819 -1712 1303 -1388
rect 1987 -1418 2445 -1133
rect 7378 -1392 7860 -1133
rect 8545 -1137 9432 -1133
rect 13912 -1128 14824 -604
rect 15081 -608 15371 -211
rect 17610 -265 17850 -264
rect 17610 -498 17853 -265
rect 15081 -1075 15966 -608
rect 17609 -680 17853 -498
rect 20425 -601 20907 -208
rect 17099 -1004 18291 -680
rect 15080 -1128 15966 -1075
rect 1961 -1716 2445 -1418
rect 7377 -1716 7861 -1392
rect 8545 -1422 9003 -1137
rect 13912 -1387 14394 -1128
rect 15079 -1132 15966 -1128
rect 20425 -1125 21337 -601
rect 21594 -605 21884 -208
rect 24123 -262 24363 -261
rect 24123 -495 24366 -262
rect 21594 -1072 22479 -605
rect 24122 -677 24366 -495
rect 23612 -1001 24804 -677
rect 21593 -1125 22479 -1072
rect 8519 -1720 9003 -1422
rect 13911 -1711 14395 -1387
rect 15079 -1417 15537 -1132
rect 20425 -1384 20907 -1125
rect 21592 -1129 22479 -1125
rect 15053 -1715 15537 -1417
rect 20424 -1708 20908 -1384
rect 21592 -1414 22050 -1129
rect 21566 -1712 22050 -1414
rect 24109 -1912 24349 -1911
rect 17596 -1915 17836 -1914
rect 4504 -1916 4744 -1915
rect 4504 -2149 4747 -1916
rect 805 -2748 1033 -2258
rect 4503 -2331 4747 -2149
rect 11062 -1920 11302 -1919
rect 11062 -2153 11305 -1920
rect 17596 -2148 17839 -1915
rect 24109 -2145 24352 -1912
rect 3993 -2655 5185 -2331
rect 501 -2948 1339 -2748
rect 2399 -2948 3722 -2748
rect 7363 -2752 7591 -2262
rect 11061 -2335 11305 -2153
rect 10551 -2659 11743 -2335
rect 13897 -2747 14125 -2257
rect 17595 -2330 17839 -2148
rect 17085 -2654 18277 -2330
rect 20410 -2744 20638 -2254
rect 24108 -2327 24352 -2145
rect 23598 -2651 24790 -2327
rect 18 -3272 3722 -2948
rect 7059 -2952 7897 -2752
rect 8957 -2952 10280 -2752
rect 13593 -2947 14431 -2747
rect 15491 -2947 16814 -2747
rect 20106 -2944 20944 -2744
rect 22004 -2944 23327 -2744
rect 558 -3965 1396 -3272
rect 2456 -3965 3294 -3272
rect 6576 -3276 10280 -2952
rect 13110 -3271 16814 -2947
rect 19623 -3268 23327 -2944
rect 4509 -3520 4749 -3519
rect 4509 -3753 4752 -3520
rect 4508 -3935 4752 -3753
rect 3998 -4259 5190 -3935
rect 7116 -3969 7954 -3276
rect 9014 -3969 9852 -3276
rect 11067 -3524 11307 -3523
rect 11067 -3757 11310 -3524
rect 11066 -3939 11310 -3757
rect 10556 -4263 11748 -3939
rect 13650 -3964 14488 -3271
rect 15548 -3964 16386 -3271
rect 17601 -3519 17841 -3518
rect 17601 -3752 17844 -3519
rect 17600 -3934 17844 -3752
rect 17090 -4258 18282 -3934
rect 20163 -3961 21001 -3268
rect 22061 -3961 22899 -3268
rect 24114 -3516 24354 -3515
rect 24114 -3749 24357 -3516
rect 24113 -3931 24357 -3749
rect 23603 -4255 24795 -3931
<< nmos >>
rect 1214 4028 1274 4428
rect 1332 4028 1392 4428
rect 1567 4228 1627 4428
rect 3212 3954 3272 4154
rect 3330 3954 3390 4154
rect 3448 3954 3508 4154
rect 4354 3958 4414 4158
rect 4472 3958 4532 4158
rect 4590 3958 4650 4158
rect 7727 4025 7787 4425
rect 7845 4025 7905 4425
rect 8080 4225 8140 4425
rect 9725 3951 9785 4151
rect 9843 3951 9903 4151
rect 9961 3951 10021 4151
rect 10867 3955 10927 4155
rect 10985 3955 11045 4155
rect 11103 3955 11163 4155
rect 14261 4020 14321 4420
rect 14379 4020 14439 4420
rect 14614 4220 14674 4420
rect 16259 3946 16319 4146
rect 16377 3946 16437 4146
rect 16495 3946 16555 4146
rect 17401 3950 17461 4150
rect 17519 3950 17579 4150
rect 17637 3950 17697 4150
rect 20819 4024 20879 4424
rect 20937 4024 20997 4424
rect 21172 4224 21232 4424
rect 22817 3950 22877 4150
rect 22935 3950 22995 4150
rect 23053 3950 23113 4150
rect 23959 3954 24019 4154
rect 24077 3954 24137 4154
rect 24195 3954 24255 4154
rect 1228 2378 1288 2778
rect 1346 2378 1406 2778
rect 1581 2578 1641 2778
rect 7741 2375 7801 2775
rect 7859 2375 7919 2775
rect 8094 2575 8154 2775
rect 1223 774 1283 1174
rect 1341 774 1401 1174
rect 1576 974 1636 1174
rect 2580 1173 2640 1373
rect 3000 973 3060 1373
rect 3118 973 3178 1373
rect 3236 973 3296 1373
rect 3354 973 3414 1373
rect 3878 1173 3938 1373
rect 4478 1173 4538 1373
rect 4898 973 4958 1373
rect 5016 973 5076 1373
rect 5134 973 5194 1373
rect 5252 973 5312 1373
rect 5776 1173 5836 1373
rect 14275 2370 14335 2770
rect 14393 2370 14453 2770
rect 14628 2570 14688 2770
rect 7736 771 7796 1171
rect 7854 771 7914 1171
rect 8089 971 8149 1171
rect 9093 1170 9153 1370
rect 9513 970 9573 1370
rect 9631 970 9691 1370
rect 9749 970 9809 1370
rect 9867 970 9927 1370
rect 10391 1170 10451 1370
rect 10991 1170 11051 1370
rect 11411 970 11471 1370
rect 11529 970 11589 1370
rect 11647 970 11707 1370
rect 11765 970 11825 1370
rect 12289 1170 12349 1370
rect 20833 2374 20893 2774
rect 20951 2374 21011 2774
rect 21186 2574 21246 2774
rect 14270 766 14330 1166
rect 14388 766 14448 1166
rect 14623 966 14683 1166
rect 15627 1165 15687 1365
rect 16047 965 16107 1365
rect 16165 965 16225 1365
rect 16283 965 16343 1365
rect 16401 965 16461 1365
rect 16925 1165 16985 1365
rect 17525 1165 17585 1365
rect 17945 965 18005 1365
rect 18063 965 18123 1365
rect 18181 965 18241 1365
rect 18299 965 18359 1365
rect 18823 1165 18883 1365
rect 20828 770 20888 1170
rect 20946 770 21006 1170
rect 21181 970 21241 1170
rect 22185 1169 22245 1369
rect 22605 969 22665 1369
rect 22723 969 22783 1369
rect 22841 969 22901 1369
rect 22959 969 23019 1369
rect 23483 1169 23543 1369
rect 24083 1169 24143 1369
rect 24503 969 24563 1369
rect 24621 969 24681 1369
rect 24739 969 24799 1369
rect 24857 969 24917 1369
rect 25381 1169 25441 1369
rect 1432 -1650 1492 -1450
rect 1550 -1650 1610 -1450
rect 1668 -1650 1728 -1450
rect 4455 -1380 4515 -1180
rect 2574 -1654 2634 -1454
rect 2692 -1654 2752 -1454
rect 2810 -1654 2870 -1454
rect 4690 -1580 4750 -1180
rect 4808 -1580 4868 -1180
rect 7990 -1654 8050 -1454
rect 8108 -1654 8168 -1454
rect 8226 -1654 8286 -1454
rect 11013 -1384 11073 -1184
rect 9132 -1658 9192 -1458
rect 9250 -1658 9310 -1458
rect 9368 -1658 9428 -1458
rect 11248 -1584 11308 -1184
rect 11366 -1584 11426 -1184
rect 14524 -1649 14584 -1449
rect 14642 -1649 14702 -1449
rect 14760 -1649 14820 -1449
rect 17547 -1379 17607 -1179
rect 15666 -1653 15726 -1453
rect 15784 -1653 15844 -1453
rect 15902 -1653 15962 -1453
rect 17782 -1579 17842 -1179
rect 17900 -1579 17960 -1179
rect 21037 -1646 21097 -1446
rect 21155 -1646 21215 -1446
rect 21273 -1646 21333 -1446
rect 24060 -1376 24120 -1176
rect 22179 -1650 22239 -1450
rect 22297 -1650 22357 -1450
rect 22415 -1650 22475 -1450
rect 24295 -1576 24355 -1176
rect 24413 -1576 24473 -1176
rect 4441 -3030 4501 -2830
rect 4676 -3230 4736 -2830
rect 4794 -3230 4854 -2830
rect 10999 -3034 11059 -2834
rect 246 -4435 306 -4235
rect 770 -4635 830 -4235
rect 888 -4635 948 -4235
rect 1006 -4635 1066 -4235
rect 1124 -4635 1184 -4235
rect 1544 -4435 1604 -4235
rect 2144 -4435 2204 -4235
rect 2668 -4635 2728 -4235
rect 2786 -4635 2846 -4235
rect 2904 -4635 2964 -4235
rect 3022 -4635 3082 -4235
rect 3442 -4435 3502 -4235
rect 11234 -3234 11294 -2834
rect 11352 -3234 11412 -2834
rect 17533 -3029 17593 -2829
rect 4446 -4634 4506 -4434
rect 4681 -4834 4741 -4434
rect 4799 -4834 4859 -4434
rect 6804 -4439 6864 -4239
rect 7328 -4639 7388 -4239
rect 7446 -4639 7506 -4239
rect 7564 -4639 7624 -4239
rect 7682 -4639 7742 -4239
rect 8102 -4439 8162 -4239
rect 8702 -4439 8762 -4239
rect 9226 -4639 9286 -4239
rect 9344 -4639 9404 -4239
rect 9462 -4639 9522 -4239
rect 9580 -4639 9640 -4239
rect 10000 -4439 10060 -4239
rect 17768 -3229 17828 -2829
rect 17886 -3229 17946 -2829
rect 24046 -3026 24106 -2826
rect 13338 -4434 13398 -4234
rect 11004 -4638 11064 -4438
rect 11239 -4838 11299 -4438
rect 11357 -4838 11417 -4438
rect 13862 -4634 13922 -4234
rect 13980 -4634 14040 -4234
rect 14098 -4634 14158 -4234
rect 14216 -4634 14276 -4234
rect 14636 -4434 14696 -4234
rect 15236 -4434 15296 -4234
rect 15760 -4634 15820 -4234
rect 15878 -4634 15938 -4234
rect 15996 -4634 16056 -4234
rect 16114 -4634 16174 -4234
rect 16534 -4434 16594 -4234
rect 24281 -3226 24341 -2826
rect 24399 -3226 24459 -2826
rect 19851 -4431 19911 -4231
rect 17538 -4633 17598 -4433
rect 17773 -4833 17833 -4433
rect 17891 -4833 17951 -4433
rect 20375 -4631 20435 -4231
rect 20493 -4631 20553 -4231
rect 20611 -4631 20671 -4231
rect 20729 -4631 20789 -4231
rect 21149 -4431 21209 -4231
rect 21749 -4431 21809 -4231
rect 22273 -4631 22333 -4231
rect 22391 -4631 22451 -4231
rect 22509 -4631 22569 -4231
rect 22627 -4631 22687 -4231
rect 23047 -4431 23107 -4231
rect 24051 -4630 24111 -4430
rect 24286 -4830 24346 -4430
rect 24404 -4830 24464 -4430
<< pmos >>
rect 977 4665 1037 4865
rect 1095 4665 1155 4865
rect 1213 4665 1273 4865
rect 1331 4665 1391 4865
rect 1449 4665 1509 4865
rect 1567 4665 1627 4865
rect 1685 4665 1745 4865
rect 1803 4665 1863 4865
rect 1921 4665 1981 4865
rect 3302 4537 3362 4937
rect 3420 4537 3480 4937
rect 3538 4537 3598 4937
rect 3656 4537 3716 4937
rect 3774 4537 3834 4937
rect 3892 4537 3952 4937
rect 4444 4541 4504 4941
rect 4562 4541 4622 4941
rect 4680 4541 4740 4941
rect 4798 4541 4858 4941
rect 4916 4541 4976 4941
rect 5034 4541 5094 4941
rect 7490 4662 7550 4862
rect 7608 4662 7668 4862
rect 7726 4662 7786 4862
rect 7844 4662 7904 4862
rect 7962 4662 8022 4862
rect 8080 4662 8140 4862
rect 8198 4662 8258 4862
rect 8316 4662 8376 4862
rect 8434 4662 8494 4862
rect 9815 4534 9875 4934
rect 9933 4534 9993 4934
rect 10051 4534 10111 4934
rect 10169 4534 10229 4934
rect 10287 4534 10347 4934
rect 10405 4534 10465 4934
rect 10957 4538 11017 4938
rect 11075 4538 11135 4938
rect 11193 4538 11253 4938
rect 11311 4538 11371 4938
rect 11429 4538 11489 4938
rect 11547 4538 11607 4938
rect 14024 4657 14084 4857
rect 14142 4657 14202 4857
rect 14260 4657 14320 4857
rect 14378 4657 14438 4857
rect 14496 4657 14556 4857
rect 14614 4657 14674 4857
rect 14732 4657 14792 4857
rect 14850 4657 14910 4857
rect 14968 4657 15028 4857
rect 3731 3954 3791 4154
rect 3849 3954 3909 4154
rect 3967 3954 4027 4154
rect 4873 3958 4933 4158
rect 4991 3958 5051 4158
rect 5109 3958 5169 4158
rect 16349 4529 16409 4929
rect 16467 4529 16527 4929
rect 16585 4529 16645 4929
rect 16703 4529 16763 4929
rect 16821 4529 16881 4929
rect 16939 4529 16999 4929
rect 17491 4533 17551 4933
rect 17609 4533 17669 4933
rect 17727 4533 17787 4933
rect 17845 4533 17905 4933
rect 17963 4533 18023 4933
rect 18081 4533 18141 4933
rect 20582 4661 20642 4861
rect 20700 4661 20760 4861
rect 20818 4661 20878 4861
rect 20936 4661 20996 4861
rect 21054 4661 21114 4861
rect 21172 4661 21232 4861
rect 21290 4661 21350 4861
rect 21408 4661 21468 4861
rect 21526 4661 21586 4861
rect 10244 3951 10304 4151
rect 10362 3951 10422 4151
rect 10480 3951 10540 4151
rect 11386 3955 11446 4155
rect 11504 3955 11564 4155
rect 11622 3955 11682 4155
rect 22907 4533 22967 4933
rect 23025 4533 23085 4933
rect 23143 4533 23203 4933
rect 23261 4533 23321 4933
rect 23379 4533 23439 4933
rect 23497 4533 23557 4933
rect 24049 4537 24109 4937
rect 24167 4537 24227 4937
rect 24285 4537 24345 4937
rect 24403 4537 24463 4937
rect 24521 4537 24581 4937
rect 24639 4537 24699 4937
rect 16778 3946 16838 4146
rect 16896 3946 16956 4146
rect 17014 3946 17074 4146
rect 17920 3950 17980 4150
rect 18038 3950 18098 4150
rect 18156 3950 18216 4150
rect 23336 3950 23396 4150
rect 23454 3950 23514 4150
rect 23572 3950 23632 4150
rect 24478 3954 24538 4154
rect 24596 3954 24656 4154
rect 24714 3954 24774 4154
rect 991 3015 1051 3215
rect 1109 3015 1169 3215
rect 1227 3015 1287 3215
rect 1345 3015 1405 3215
rect 1463 3015 1523 3215
rect 1581 3015 1641 3215
rect 1699 3015 1759 3215
rect 1817 3015 1877 3215
rect 1935 3015 1995 3215
rect 7504 3012 7564 3212
rect 7622 3012 7682 3212
rect 7740 3012 7800 3212
rect 7858 3012 7918 3212
rect 7976 3012 8036 3212
rect 8094 3012 8154 3212
rect 8212 3012 8272 3212
rect 8330 3012 8390 3212
rect 8448 3012 8508 3212
rect 2455 2398 2515 2598
rect 2573 2398 2633 2598
rect 2691 2398 2751 2598
rect 2939 2398 2999 2798
rect 3057 2398 3117 2798
rect 3175 2398 3235 2798
rect 3293 2398 3353 2798
rect 3411 2398 3471 2798
rect 3529 2398 3589 2798
rect 3776 2398 3836 2598
rect 3894 2398 3954 2598
rect 4012 2398 4072 2598
rect 4353 2398 4413 2598
rect 4471 2398 4531 2598
rect 4589 2398 4649 2598
rect 4837 2398 4897 2798
rect 4955 2398 5015 2798
rect 5073 2398 5133 2798
rect 5191 2398 5251 2798
rect 5309 2398 5369 2798
rect 5427 2398 5487 2798
rect 14038 3007 14098 3207
rect 14156 3007 14216 3207
rect 14274 3007 14334 3207
rect 14392 3007 14452 3207
rect 14510 3007 14570 3207
rect 14628 3007 14688 3207
rect 14746 3007 14806 3207
rect 14864 3007 14924 3207
rect 14982 3007 15042 3207
rect 20596 3011 20656 3211
rect 20714 3011 20774 3211
rect 20832 3011 20892 3211
rect 20950 3011 21010 3211
rect 21068 3011 21128 3211
rect 21186 3011 21246 3211
rect 21304 3011 21364 3211
rect 21422 3011 21482 3211
rect 21540 3011 21600 3211
rect 5674 2398 5734 2598
rect 5792 2398 5852 2598
rect 5910 2398 5970 2598
rect 986 1411 1046 1611
rect 1104 1411 1164 1611
rect 1222 1411 1282 1611
rect 1340 1411 1400 1611
rect 1458 1411 1518 1611
rect 1576 1411 1636 1611
rect 1694 1411 1754 1611
rect 1812 1411 1872 1611
rect 1930 1411 1990 1611
rect 2882 1705 2942 2105
rect 3000 1705 3060 2105
rect 3118 1705 3178 2105
rect 3236 1705 3296 2105
rect 3354 1705 3414 2105
rect 3472 1705 3532 2105
rect 8968 2395 9028 2595
rect 9086 2395 9146 2595
rect 9204 2395 9264 2595
rect 9452 2395 9512 2795
rect 9570 2395 9630 2795
rect 9688 2395 9748 2795
rect 9806 2395 9866 2795
rect 9924 2395 9984 2795
rect 10042 2395 10102 2795
rect 10289 2395 10349 2595
rect 10407 2395 10467 2595
rect 10525 2395 10585 2595
rect 10866 2395 10926 2595
rect 10984 2395 11044 2595
rect 11102 2395 11162 2595
rect 11350 2395 11410 2795
rect 11468 2395 11528 2795
rect 11586 2395 11646 2795
rect 11704 2395 11764 2795
rect 11822 2395 11882 2795
rect 11940 2395 12000 2795
rect 12187 2395 12247 2595
rect 12305 2395 12365 2595
rect 12423 2395 12483 2595
rect 4780 1705 4840 2105
rect 4898 1705 4958 2105
rect 5016 1705 5076 2105
rect 5134 1705 5194 2105
rect 5252 1705 5312 2105
rect 5370 1705 5430 2105
rect 7499 1408 7559 1608
rect 7617 1408 7677 1608
rect 7735 1408 7795 1608
rect 7853 1408 7913 1608
rect 7971 1408 8031 1608
rect 8089 1408 8149 1608
rect 8207 1408 8267 1608
rect 8325 1408 8385 1608
rect 8443 1408 8503 1608
rect 9395 1702 9455 2102
rect 9513 1702 9573 2102
rect 9631 1702 9691 2102
rect 9749 1702 9809 2102
rect 9867 1702 9927 2102
rect 9985 1702 10045 2102
rect 15502 2390 15562 2590
rect 15620 2390 15680 2590
rect 15738 2390 15798 2590
rect 15986 2390 16046 2790
rect 16104 2390 16164 2790
rect 16222 2390 16282 2790
rect 16340 2390 16400 2790
rect 16458 2390 16518 2790
rect 16576 2390 16636 2790
rect 16823 2390 16883 2590
rect 16941 2390 17001 2590
rect 17059 2390 17119 2590
rect 17400 2390 17460 2590
rect 17518 2390 17578 2590
rect 17636 2390 17696 2590
rect 17884 2390 17944 2790
rect 18002 2390 18062 2790
rect 18120 2390 18180 2790
rect 18238 2390 18298 2790
rect 18356 2390 18416 2790
rect 18474 2390 18534 2790
rect 18721 2390 18781 2590
rect 18839 2390 18899 2590
rect 18957 2390 19017 2590
rect 11293 1702 11353 2102
rect 11411 1702 11471 2102
rect 11529 1702 11589 2102
rect 11647 1702 11707 2102
rect 11765 1702 11825 2102
rect 11883 1702 11943 2102
rect 14033 1403 14093 1603
rect 14151 1403 14211 1603
rect 14269 1403 14329 1603
rect 14387 1403 14447 1603
rect 14505 1403 14565 1603
rect 14623 1403 14683 1603
rect 14741 1403 14801 1603
rect 14859 1403 14919 1603
rect 14977 1403 15037 1603
rect 15929 1697 15989 2097
rect 16047 1697 16107 2097
rect 16165 1697 16225 2097
rect 16283 1697 16343 2097
rect 16401 1697 16461 2097
rect 16519 1697 16579 2097
rect 22060 2394 22120 2594
rect 22178 2394 22238 2594
rect 22296 2394 22356 2594
rect 22544 2394 22604 2794
rect 22662 2394 22722 2794
rect 22780 2394 22840 2794
rect 22898 2394 22958 2794
rect 23016 2394 23076 2794
rect 23134 2394 23194 2794
rect 23381 2394 23441 2594
rect 23499 2394 23559 2594
rect 23617 2394 23677 2594
rect 23958 2394 24018 2594
rect 24076 2394 24136 2594
rect 24194 2394 24254 2594
rect 24442 2394 24502 2794
rect 24560 2394 24620 2794
rect 24678 2394 24738 2794
rect 24796 2394 24856 2794
rect 24914 2394 24974 2794
rect 25032 2394 25092 2794
rect 25279 2394 25339 2594
rect 25397 2394 25457 2594
rect 25515 2394 25575 2594
rect 17827 1697 17887 2097
rect 17945 1697 18005 2097
rect 18063 1697 18123 2097
rect 18181 1697 18241 2097
rect 18299 1697 18359 2097
rect 18417 1697 18477 2097
rect 20591 1407 20651 1607
rect 20709 1407 20769 1607
rect 20827 1407 20887 1607
rect 20945 1407 21005 1607
rect 21063 1407 21123 1607
rect 21181 1407 21241 1607
rect 21299 1407 21359 1607
rect 21417 1407 21477 1607
rect 21535 1407 21595 1607
rect 22487 1701 22547 2101
rect 22605 1701 22665 2101
rect 22723 1701 22783 2101
rect 22841 1701 22901 2101
rect 22959 1701 23019 2101
rect 23077 1701 23137 2101
rect 24385 1701 24445 2101
rect 24503 1701 24563 2101
rect 24621 1701 24681 2101
rect 24739 1701 24799 2101
rect 24857 1701 24917 2101
rect 24975 1701 25035 2101
rect 988 -1067 1048 -667
rect 1106 -1067 1166 -667
rect 1224 -1067 1284 -667
rect 1342 -1067 1402 -667
rect 1460 -1067 1520 -667
rect 1578 -1067 1638 -667
rect 2130 -1071 2190 -671
rect 2248 -1071 2308 -671
rect 2366 -1071 2426 -671
rect 2484 -1071 2544 -671
rect 2602 -1071 2662 -671
rect 2720 -1071 2780 -671
rect 4101 -943 4161 -743
rect 4219 -943 4279 -743
rect 4337 -943 4397 -743
rect 4455 -943 4515 -743
rect 4573 -943 4633 -743
rect 4691 -943 4751 -743
rect 4809 -943 4869 -743
rect 4927 -943 4987 -743
rect 5045 -943 5105 -743
rect 7546 -1071 7606 -671
rect 7664 -1071 7724 -671
rect 7782 -1071 7842 -671
rect 7900 -1071 7960 -671
rect 8018 -1071 8078 -671
rect 8136 -1071 8196 -671
rect 913 -1650 973 -1450
rect 1031 -1650 1091 -1450
rect 1149 -1650 1209 -1450
rect 2055 -1654 2115 -1454
rect 2173 -1654 2233 -1454
rect 2291 -1654 2351 -1454
rect 8688 -1075 8748 -675
rect 8806 -1075 8866 -675
rect 8924 -1075 8984 -675
rect 9042 -1075 9102 -675
rect 9160 -1075 9220 -675
rect 9278 -1075 9338 -675
rect 10659 -947 10719 -747
rect 10777 -947 10837 -747
rect 10895 -947 10955 -747
rect 11013 -947 11073 -747
rect 11131 -947 11191 -747
rect 11249 -947 11309 -747
rect 11367 -947 11427 -747
rect 11485 -947 11545 -747
rect 11603 -947 11663 -747
rect 14080 -1066 14140 -666
rect 14198 -1066 14258 -666
rect 14316 -1066 14376 -666
rect 14434 -1066 14494 -666
rect 14552 -1066 14612 -666
rect 14670 -1066 14730 -666
rect 7471 -1654 7531 -1454
rect 7589 -1654 7649 -1454
rect 7707 -1654 7767 -1454
rect 8613 -1658 8673 -1458
rect 8731 -1658 8791 -1458
rect 8849 -1658 8909 -1458
rect 15222 -1070 15282 -670
rect 15340 -1070 15400 -670
rect 15458 -1070 15518 -670
rect 15576 -1070 15636 -670
rect 15694 -1070 15754 -670
rect 15812 -1070 15872 -670
rect 17193 -942 17253 -742
rect 17311 -942 17371 -742
rect 17429 -942 17489 -742
rect 17547 -942 17607 -742
rect 17665 -942 17725 -742
rect 17783 -942 17843 -742
rect 17901 -942 17961 -742
rect 18019 -942 18079 -742
rect 18137 -942 18197 -742
rect 20593 -1063 20653 -663
rect 20711 -1063 20771 -663
rect 20829 -1063 20889 -663
rect 20947 -1063 21007 -663
rect 21065 -1063 21125 -663
rect 21183 -1063 21243 -663
rect 14005 -1649 14065 -1449
rect 14123 -1649 14183 -1449
rect 14241 -1649 14301 -1449
rect 15147 -1653 15207 -1453
rect 15265 -1653 15325 -1453
rect 15383 -1653 15443 -1453
rect 21735 -1067 21795 -667
rect 21853 -1067 21913 -667
rect 21971 -1067 22031 -667
rect 22089 -1067 22149 -667
rect 22207 -1067 22267 -667
rect 22325 -1067 22385 -667
rect 23706 -939 23766 -739
rect 23824 -939 23884 -739
rect 23942 -939 24002 -739
rect 24060 -939 24120 -739
rect 24178 -939 24238 -739
rect 24296 -939 24356 -739
rect 24414 -939 24474 -739
rect 24532 -939 24592 -739
rect 24650 -939 24710 -739
rect 20518 -1646 20578 -1446
rect 20636 -1646 20696 -1446
rect 20754 -1646 20814 -1446
rect 21660 -1650 21720 -1450
rect 21778 -1650 21838 -1450
rect 21896 -1650 21956 -1450
rect 4087 -2593 4147 -2393
rect 4205 -2593 4265 -2393
rect 4323 -2593 4383 -2393
rect 4441 -2593 4501 -2393
rect 4559 -2593 4619 -2393
rect 4677 -2593 4737 -2393
rect 4795 -2593 4855 -2393
rect 4913 -2593 4973 -2393
rect 5031 -2593 5091 -2393
rect 10645 -2597 10705 -2397
rect 10763 -2597 10823 -2397
rect 10881 -2597 10941 -2397
rect 10999 -2597 11059 -2397
rect 11117 -2597 11177 -2397
rect 11235 -2597 11295 -2397
rect 11353 -2597 11413 -2397
rect 11471 -2597 11531 -2397
rect 11589 -2597 11649 -2397
rect 17179 -2592 17239 -2392
rect 17297 -2592 17357 -2392
rect 17415 -2592 17475 -2392
rect 17533 -2592 17593 -2392
rect 17651 -2592 17711 -2392
rect 17769 -2592 17829 -2392
rect 17887 -2592 17947 -2392
rect 18005 -2592 18065 -2392
rect 18123 -2592 18183 -2392
rect 23692 -2589 23752 -2389
rect 23810 -2589 23870 -2389
rect 23928 -2589 23988 -2389
rect 24046 -2589 24106 -2389
rect 24164 -2589 24224 -2389
rect 24282 -2589 24342 -2389
rect 24400 -2589 24460 -2389
rect 24518 -2589 24578 -2389
rect 24636 -2589 24696 -2389
rect 112 -3210 172 -3010
rect 230 -3210 290 -3010
rect 348 -3210 408 -3010
rect 595 -3210 655 -2810
rect 713 -3210 773 -2810
rect 831 -3210 891 -2810
rect 949 -3210 1009 -2810
rect 1067 -3210 1127 -2810
rect 1185 -3210 1245 -2810
rect 1433 -3210 1493 -3010
rect 1551 -3210 1611 -3010
rect 1669 -3210 1729 -3010
rect 2010 -3210 2070 -3010
rect 2128 -3210 2188 -3010
rect 2246 -3210 2306 -3010
rect 2493 -3210 2553 -2810
rect 2611 -3210 2671 -2810
rect 2729 -3210 2789 -2810
rect 2847 -3210 2907 -2810
rect 2965 -3210 3025 -2810
rect 3083 -3210 3143 -2810
rect 3331 -3210 3391 -3010
rect 3449 -3210 3509 -3010
rect 3567 -3210 3627 -3010
rect 652 -3903 712 -3503
rect 770 -3903 830 -3503
rect 888 -3903 948 -3503
rect 1006 -3903 1066 -3503
rect 1124 -3903 1184 -3503
rect 1242 -3903 1302 -3503
rect 6670 -3214 6730 -3014
rect 6788 -3214 6848 -3014
rect 6906 -3214 6966 -3014
rect 7153 -3214 7213 -2814
rect 7271 -3214 7331 -2814
rect 7389 -3214 7449 -2814
rect 7507 -3214 7567 -2814
rect 7625 -3214 7685 -2814
rect 7743 -3214 7803 -2814
rect 7991 -3214 8051 -3014
rect 8109 -3214 8169 -3014
rect 8227 -3214 8287 -3014
rect 8568 -3214 8628 -3014
rect 8686 -3214 8746 -3014
rect 8804 -3214 8864 -3014
rect 9051 -3214 9111 -2814
rect 9169 -3214 9229 -2814
rect 9287 -3214 9347 -2814
rect 9405 -3214 9465 -2814
rect 9523 -3214 9583 -2814
rect 9641 -3214 9701 -2814
rect 9889 -3214 9949 -3014
rect 10007 -3214 10067 -3014
rect 10125 -3214 10185 -3014
rect 2550 -3903 2610 -3503
rect 2668 -3903 2728 -3503
rect 2786 -3903 2846 -3503
rect 2904 -3903 2964 -3503
rect 3022 -3903 3082 -3503
rect 3140 -3903 3200 -3503
rect 4092 -4197 4152 -3997
rect 4210 -4197 4270 -3997
rect 4328 -4197 4388 -3997
rect 4446 -4197 4506 -3997
rect 4564 -4197 4624 -3997
rect 4682 -4197 4742 -3997
rect 4800 -4197 4860 -3997
rect 4918 -4197 4978 -3997
rect 5036 -4197 5096 -3997
rect 7210 -3907 7270 -3507
rect 7328 -3907 7388 -3507
rect 7446 -3907 7506 -3507
rect 7564 -3907 7624 -3507
rect 7682 -3907 7742 -3507
rect 7800 -3907 7860 -3507
rect 13204 -3209 13264 -3009
rect 13322 -3209 13382 -3009
rect 13440 -3209 13500 -3009
rect 13687 -3209 13747 -2809
rect 13805 -3209 13865 -2809
rect 13923 -3209 13983 -2809
rect 14041 -3209 14101 -2809
rect 14159 -3209 14219 -2809
rect 14277 -3209 14337 -2809
rect 14525 -3209 14585 -3009
rect 14643 -3209 14703 -3009
rect 14761 -3209 14821 -3009
rect 15102 -3209 15162 -3009
rect 15220 -3209 15280 -3009
rect 15338 -3209 15398 -3009
rect 15585 -3209 15645 -2809
rect 15703 -3209 15763 -2809
rect 15821 -3209 15881 -2809
rect 15939 -3209 15999 -2809
rect 16057 -3209 16117 -2809
rect 16175 -3209 16235 -2809
rect 16423 -3209 16483 -3009
rect 16541 -3209 16601 -3009
rect 16659 -3209 16719 -3009
rect 9108 -3907 9168 -3507
rect 9226 -3907 9286 -3507
rect 9344 -3907 9404 -3507
rect 9462 -3907 9522 -3507
rect 9580 -3907 9640 -3507
rect 9698 -3907 9758 -3507
rect 10650 -4201 10710 -4001
rect 10768 -4201 10828 -4001
rect 10886 -4201 10946 -4001
rect 11004 -4201 11064 -4001
rect 11122 -4201 11182 -4001
rect 11240 -4201 11300 -4001
rect 11358 -4201 11418 -4001
rect 11476 -4201 11536 -4001
rect 11594 -4201 11654 -4001
rect 13744 -3902 13804 -3502
rect 13862 -3902 13922 -3502
rect 13980 -3902 14040 -3502
rect 14098 -3902 14158 -3502
rect 14216 -3902 14276 -3502
rect 14334 -3902 14394 -3502
rect 19717 -3206 19777 -3006
rect 19835 -3206 19895 -3006
rect 19953 -3206 20013 -3006
rect 20200 -3206 20260 -2806
rect 20318 -3206 20378 -2806
rect 20436 -3206 20496 -2806
rect 20554 -3206 20614 -2806
rect 20672 -3206 20732 -2806
rect 20790 -3206 20850 -2806
rect 21038 -3206 21098 -3006
rect 21156 -3206 21216 -3006
rect 21274 -3206 21334 -3006
rect 21615 -3206 21675 -3006
rect 21733 -3206 21793 -3006
rect 21851 -3206 21911 -3006
rect 22098 -3206 22158 -2806
rect 22216 -3206 22276 -2806
rect 22334 -3206 22394 -2806
rect 22452 -3206 22512 -2806
rect 22570 -3206 22630 -2806
rect 22688 -3206 22748 -2806
rect 22936 -3206 22996 -3006
rect 23054 -3206 23114 -3006
rect 23172 -3206 23232 -3006
rect 15642 -3902 15702 -3502
rect 15760 -3902 15820 -3502
rect 15878 -3902 15938 -3502
rect 15996 -3902 16056 -3502
rect 16114 -3902 16174 -3502
rect 16232 -3902 16292 -3502
rect 17184 -4196 17244 -3996
rect 17302 -4196 17362 -3996
rect 17420 -4196 17480 -3996
rect 17538 -4196 17598 -3996
rect 17656 -4196 17716 -3996
rect 17774 -4196 17834 -3996
rect 17892 -4196 17952 -3996
rect 18010 -4196 18070 -3996
rect 18128 -4196 18188 -3996
rect 20257 -3899 20317 -3499
rect 20375 -3899 20435 -3499
rect 20493 -3899 20553 -3499
rect 20611 -3899 20671 -3499
rect 20729 -3899 20789 -3499
rect 20847 -3899 20907 -3499
rect 22155 -3899 22215 -3499
rect 22273 -3899 22333 -3499
rect 22391 -3899 22451 -3499
rect 22509 -3899 22569 -3499
rect 22627 -3899 22687 -3499
rect 22745 -3899 22805 -3499
rect 23697 -4193 23757 -3993
rect 23815 -4193 23875 -3993
rect 23933 -4193 23993 -3993
rect 24051 -4193 24111 -3993
rect 24169 -4193 24229 -3993
rect 24287 -4193 24347 -3993
rect 24405 -4193 24465 -3993
rect 24523 -4193 24583 -3993
rect 24641 -4193 24701 -3993
<< ndiff >>
rect 1156 4416 1214 4428
rect 1156 4040 1168 4416
rect 1202 4040 1214 4416
rect 1156 4028 1214 4040
rect 1274 4416 1332 4428
rect 1274 4040 1286 4416
rect 1320 4040 1332 4416
rect 1274 4028 1332 4040
rect 1392 4416 1450 4428
rect 1392 4040 1404 4416
rect 1438 4040 1450 4416
rect 1509 4416 1567 4428
rect 1509 4240 1521 4416
rect 1555 4240 1567 4416
rect 1509 4228 1567 4240
rect 1627 4416 1685 4428
rect 1627 4240 1639 4416
rect 1673 4240 1685 4416
rect 1627 4228 1685 4240
rect 7669 4413 7727 4425
rect 3154 4142 3212 4154
rect 1392 4028 1450 4040
rect 3154 3966 3166 4142
rect 3200 3966 3212 4142
rect 3154 3954 3212 3966
rect 3272 4142 3330 4154
rect 3272 3966 3284 4142
rect 3318 3966 3330 4142
rect 3272 3954 3330 3966
rect 3390 4142 3448 4154
rect 3390 3966 3402 4142
rect 3436 3966 3448 4142
rect 3390 3954 3448 3966
rect 3508 4142 3566 4154
rect 3508 3966 3520 4142
rect 3554 3966 3566 4142
rect 3508 3954 3566 3966
rect 4296 4146 4354 4158
rect 4296 3970 4308 4146
rect 4342 3970 4354 4146
rect 4296 3958 4354 3970
rect 4414 4146 4472 4158
rect 4414 3970 4426 4146
rect 4460 3970 4472 4146
rect 4414 3958 4472 3970
rect 4532 4146 4590 4158
rect 4532 3970 4544 4146
rect 4578 3970 4590 4146
rect 4532 3958 4590 3970
rect 4650 4146 4708 4158
rect 4650 3970 4662 4146
rect 4696 3970 4708 4146
rect 4650 3958 4708 3970
rect 7669 4037 7681 4413
rect 7715 4037 7727 4413
rect 7669 4025 7727 4037
rect 7787 4413 7845 4425
rect 7787 4037 7799 4413
rect 7833 4037 7845 4413
rect 7787 4025 7845 4037
rect 7905 4413 7963 4425
rect 7905 4037 7917 4413
rect 7951 4037 7963 4413
rect 8022 4413 8080 4425
rect 8022 4237 8034 4413
rect 8068 4237 8080 4413
rect 8022 4225 8080 4237
rect 8140 4413 8198 4425
rect 8140 4237 8152 4413
rect 8186 4237 8198 4413
rect 8140 4225 8198 4237
rect 14203 4408 14261 4420
rect 9667 4139 9725 4151
rect 7905 4025 7963 4037
rect 9667 3963 9679 4139
rect 9713 3963 9725 4139
rect 9667 3951 9725 3963
rect 9785 4139 9843 4151
rect 9785 3963 9797 4139
rect 9831 3963 9843 4139
rect 9785 3951 9843 3963
rect 9903 4139 9961 4151
rect 9903 3963 9915 4139
rect 9949 3963 9961 4139
rect 9903 3951 9961 3963
rect 10021 4139 10079 4151
rect 10021 3963 10033 4139
rect 10067 3963 10079 4139
rect 10021 3951 10079 3963
rect 10809 4143 10867 4155
rect 10809 3967 10821 4143
rect 10855 3967 10867 4143
rect 10809 3955 10867 3967
rect 10927 4143 10985 4155
rect 10927 3967 10939 4143
rect 10973 3967 10985 4143
rect 10927 3955 10985 3967
rect 11045 4143 11103 4155
rect 11045 3967 11057 4143
rect 11091 3967 11103 4143
rect 11045 3955 11103 3967
rect 11163 4143 11221 4155
rect 11163 3967 11175 4143
rect 11209 3967 11221 4143
rect 11163 3955 11221 3967
rect 14203 4032 14215 4408
rect 14249 4032 14261 4408
rect 14203 4020 14261 4032
rect 14321 4408 14379 4420
rect 14321 4032 14333 4408
rect 14367 4032 14379 4408
rect 14321 4020 14379 4032
rect 14439 4408 14497 4420
rect 14439 4032 14451 4408
rect 14485 4032 14497 4408
rect 14556 4408 14614 4420
rect 14556 4232 14568 4408
rect 14602 4232 14614 4408
rect 14556 4220 14614 4232
rect 14674 4408 14732 4420
rect 14674 4232 14686 4408
rect 14720 4232 14732 4408
rect 14674 4220 14732 4232
rect 20761 4412 20819 4424
rect 16201 4134 16259 4146
rect 14439 4020 14497 4032
rect 16201 3958 16213 4134
rect 16247 3958 16259 4134
rect 16201 3946 16259 3958
rect 16319 4134 16377 4146
rect 16319 3958 16331 4134
rect 16365 3958 16377 4134
rect 16319 3946 16377 3958
rect 16437 4134 16495 4146
rect 16437 3958 16449 4134
rect 16483 3958 16495 4134
rect 16437 3946 16495 3958
rect 16555 4134 16613 4146
rect 16555 3958 16567 4134
rect 16601 3958 16613 4134
rect 16555 3946 16613 3958
rect 17343 4138 17401 4150
rect 17343 3962 17355 4138
rect 17389 3962 17401 4138
rect 17343 3950 17401 3962
rect 17461 4138 17519 4150
rect 17461 3962 17473 4138
rect 17507 3962 17519 4138
rect 17461 3950 17519 3962
rect 17579 4138 17637 4150
rect 17579 3962 17591 4138
rect 17625 3962 17637 4138
rect 17579 3950 17637 3962
rect 17697 4138 17755 4150
rect 17697 3962 17709 4138
rect 17743 3962 17755 4138
rect 17697 3950 17755 3962
rect 20761 4036 20773 4412
rect 20807 4036 20819 4412
rect 20761 4024 20819 4036
rect 20879 4412 20937 4424
rect 20879 4036 20891 4412
rect 20925 4036 20937 4412
rect 20879 4024 20937 4036
rect 20997 4412 21055 4424
rect 20997 4036 21009 4412
rect 21043 4036 21055 4412
rect 21114 4412 21172 4424
rect 21114 4236 21126 4412
rect 21160 4236 21172 4412
rect 21114 4224 21172 4236
rect 21232 4412 21290 4424
rect 21232 4236 21244 4412
rect 21278 4236 21290 4412
rect 21232 4224 21290 4236
rect 22759 4138 22817 4150
rect 20997 4024 21055 4036
rect 22759 3962 22771 4138
rect 22805 3962 22817 4138
rect 22759 3950 22817 3962
rect 22877 4138 22935 4150
rect 22877 3962 22889 4138
rect 22923 3962 22935 4138
rect 22877 3950 22935 3962
rect 22995 4138 23053 4150
rect 22995 3962 23007 4138
rect 23041 3962 23053 4138
rect 22995 3950 23053 3962
rect 23113 4138 23171 4150
rect 23113 3962 23125 4138
rect 23159 3962 23171 4138
rect 23113 3950 23171 3962
rect 23901 4142 23959 4154
rect 23901 3966 23913 4142
rect 23947 3966 23959 4142
rect 23901 3954 23959 3966
rect 24019 4142 24077 4154
rect 24019 3966 24031 4142
rect 24065 3966 24077 4142
rect 24019 3954 24077 3966
rect 24137 4142 24195 4154
rect 24137 3966 24149 4142
rect 24183 3966 24195 4142
rect 24137 3954 24195 3966
rect 24255 4142 24313 4154
rect 24255 3966 24267 4142
rect 24301 3966 24313 4142
rect 24255 3954 24313 3966
rect 1170 2766 1228 2778
rect 1170 2390 1182 2766
rect 1216 2390 1228 2766
rect 1170 2378 1228 2390
rect 1288 2766 1346 2778
rect 1288 2390 1300 2766
rect 1334 2390 1346 2766
rect 1288 2378 1346 2390
rect 1406 2766 1464 2778
rect 1406 2390 1418 2766
rect 1452 2390 1464 2766
rect 1523 2766 1581 2778
rect 1523 2590 1535 2766
rect 1569 2590 1581 2766
rect 1523 2578 1581 2590
rect 1641 2766 1699 2778
rect 1641 2590 1653 2766
rect 1687 2590 1699 2766
rect 1641 2578 1699 2590
rect 1406 2378 1464 2390
rect 7683 2763 7741 2775
rect 7683 2387 7695 2763
rect 7729 2387 7741 2763
rect 7683 2375 7741 2387
rect 7801 2763 7859 2775
rect 7801 2387 7813 2763
rect 7847 2387 7859 2763
rect 7801 2375 7859 2387
rect 7919 2763 7977 2775
rect 7919 2387 7931 2763
rect 7965 2387 7977 2763
rect 8036 2763 8094 2775
rect 8036 2587 8048 2763
rect 8082 2587 8094 2763
rect 8036 2575 8094 2587
rect 8154 2763 8212 2775
rect 8154 2587 8166 2763
rect 8200 2587 8212 2763
rect 8154 2575 8212 2587
rect 7919 2375 7977 2387
rect 14217 2758 14275 2770
rect 2522 1361 2580 1373
rect 2522 1185 2534 1361
rect 2568 1185 2580 1361
rect 1165 1162 1223 1174
rect 1165 786 1177 1162
rect 1211 786 1223 1162
rect 1165 774 1223 786
rect 1283 1162 1341 1174
rect 1283 786 1295 1162
rect 1329 786 1341 1162
rect 1283 774 1341 786
rect 1401 1162 1459 1174
rect 1401 786 1413 1162
rect 1447 786 1459 1162
rect 1518 1162 1576 1174
rect 1518 986 1530 1162
rect 1564 986 1576 1162
rect 1518 974 1576 986
rect 1636 1162 1694 1174
rect 2522 1173 2580 1185
rect 2640 1361 2698 1373
rect 2640 1185 2652 1361
rect 2686 1185 2698 1361
rect 2640 1173 2698 1185
rect 2942 1361 3000 1373
rect 1636 986 1648 1162
rect 1682 986 1694 1162
rect 1636 974 1694 986
rect 2942 985 2954 1361
rect 2988 985 3000 1361
rect 2942 973 3000 985
rect 3060 1361 3118 1373
rect 3060 985 3072 1361
rect 3106 985 3118 1361
rect 3060 973 3118 985
rect 3178 1361 3236 1373
rect 3178 985 3190 1361
rect 3224 985 3236 1361
rect 3178 973 3236 985
rect 3296 1361 3354 1373
rect 3296 985 3308 1361
rect 3342 985 3354 1361
rect 3296 973 3354 985
rect 3414 1361 3472 1373
rect 3414 985 3426 1361
rect 3460 985 3472 1361
rect 3820 1361 3878 1373
rect 3820 1185 3832 1361
rect 3866 1185 3878 1361
rect 3820 1173 3878 1185
rect 3938 1361 3996 1373
rect 3938 1185 3950 1361
rect 3984 1185 3996 1361
rect 3938 1173 3996 1185
rect 4420 1361 4478 1373
rect 4420 1185 4432 1361
rect 4466 1185 4478 1361
rect 4420 1173 4478 1185
rect 4538 1361 4596 1373
rect 4538 1185 4550 1361
rect 4584 1185 4596 1361
rect 4538 1173 4596 1185
rect 4840 1361 4898 1373
rect 3414 973 3472 985
rect 4840 985 4852 1361
rect 4886 985 4898 1361
rect 4840 973 4898 985
rect 4958 1361 5016 1373
rect 4958 985 4970 1361
rect 5004 985 5016 1361
rect 4958 973 5016 985
rect 5076 1361 5134 1373
rect 5076 985 5088 1361
rect 5122 985 5134 1361
rect 5076 973 5134 985
rect 5194 1361 5252 1373
rect 5194 985 5206 1361
rect 5240 985 5252 1361
rect 5194 973 5252 985
rect 5312 1361 5370 1373
rect 5312 985 5324 1361
rect 5358 985 5370 1361
rect 5718 1361 5776 1373
rect 5718 1185 5730 1361
rect 5764 1185 5776 1361
rect 5718 1173 5776 1185
rect 5836 1361 5894 1373
rect 5836 1185 5848 1361
rect 5882 1185 5894 1361
rect 5836 1173 5894 1185
rect 14217 2382 14229 2758
rect 14263 2382 14275 2758
rect 14217 2370 14275 2382
rect 14335 2758 14393 2770
rect 14335 2382 14347 2758
rect 14381 2382 14393 2758
rect 14335 2370 14393 2382
rect 14453 2758 14511 2770
rect 14453 2382 14465 2758
rect 14499 2382 14511 2758
rect 14570 2758 14628 2770
rect 14570 2582 14582 2758
rect 14616 2582 14628 2758
rect 14570 2570 14628 2582
rect 14688 2758 14746 2770
rect 14688 2582 14700 2758
rect 14734 2582 14746 2758
rect 14688 2570 14746 2582
rect 14453 2370 14511 2382
rect 20775 2762 20833 2774
rect 9035 1358 9093 1370
rect 9035 1182 9047 1358
rect 9081 1182 9093 1358
rect 7678 1159 7736 1171
rect 5312 973 5370 985
rect 1401 774 1459 786
rect 7678 783 7690 1159
rect 7724 783 7736 1159
rect 7678 771 7736 783
rect 7796 1159 7854 1171
rect 7796 783 7808 1159
rect 7842 783 7854 1159
rect 7796 771 7854 783
rect 7914 1159 7972 1171
rect 7914 783 7926 1159
rect 7960 783 7972 1159
rect 8031 1159 8089 1171
rect 8031 983 8043 1159
rect 8077 983 8089 1159
rect 8031 971 8089 983
rect 8149 1159 8207 1171
rect 9035 1170 9093 1182
rect 9153 1358 9211 1370
rect 9153 1182 9165 1358
rect 9199 1182 9211 1358
rect 9153 1170 9211 1182
rect 9455 1358 9513 1370
rect 8149 983 8161 1159
rect 8195 983 8207 1159
rect 8149 971 8207 983
rect 9455 982 9467 1358
rect 9501 982 9513 1358
rect 9455 970 9513 982
rect 9573 1358 9631 1370
rect 9573 982 9585 1358
rect 9619 982 9631 1358
rect 9573 970 9631 982
rect 9691 1358 9749 1370
rect 9691 982 9703 1358
rect 9737 982 9749 1358
rect 9691 970 9749 982
rect 9809 1358 9867 1370
rect 9809 982 9821 1358
rect 9855 982 9867 1358
rect 9809 970 9867 982
rect 9927 1358 9985 1370
rect 9927 982 9939 1358
rect 9973 982 9985 1358
rect 10333 1358 10391 1370
rect 10333 1182 10345 1358
rect 10379 1182 10391 1358
rect 10333 1170 10391 1182
rect 10451 1358 10509 1370
rect 10451 1182 10463 1358
rect 10497 1182 10509 1358
rect 10451 1170 10509 1182
rect 10933 1358 10991 1370
rect 10933 1182 10945 1358
rect 10979 1182 10991 1358
rect 10933 1170 10991 1182
rect 11051 1358 11109 1370
rect 11051 1182 11063 1358
rect 11097 1182 11109 1358
rect 11051 1170 11109 1182
rect 11353 1358 11411 1370
rect 9927 970 9985 982
rect 11353 982 11365 1358
rect 11399 982 11411 1358
rect 11353 970 11411 982
rect 11471 1358 11529 1370
rect 11471 982 11483 1358
rect 11517 982 11529 1358
rect 11471 970 11529 982
rect 11589 1358 11647 1370
rect 11589 982 11601 1358
rect 11635 982 11647 1358
rect 11589 970 11647 982
rect 11707 1358 11765 1370
rect 11707 982 11719 1358
rect 11753 982 11765 1358
rect 11707 970 11765 982
rect 11825 1358 11883 1370
rect 11825 982 11837 1358
rect 11871 982 11883 1358
rect 12231 1358 12289 1370
rect 12231 1182 12243 1358
rect 12277 1182 12289 1358
rect 12231 1170 12289 1182
rect 12349 1358 12407 1370
rect 12349 1182 12361 1358
rect 12395 1182 12407 1358
rect 12349 1170 12407 1182
rect 20775 2386 20787 2762
rect 20821 2386 20833 2762
rect 20775 2374 20833 2386
rect 20893 2762 20951 2774
rect 20893 2386 20905 2762
rect 20939 2386 20951 2762
rect 20893 2374 20951 2386
rect 21011 2762 21069 2774
rect 21011 2386 21023 2762
rect 21057 2386 21069 2762
rect 21128 2762 21186 2774
rect 21128 2586 21140 2762
rect 21174 2586 21186 2762
rect 21128 2574 21186 2586
rect 21246 2762 21304 2774
rect 21246 2586 21258 2762
rect 21292 2586 21304 2762
rect 21246 2574 21304 2586
rect 21011 2374 21069 2386
rect 15569 1353 15627 1365
rect 15569 1177 15581 1353
rect 15615 1177 15627 1353
rect 14212 1154 14270 1166
rect 11825 970 11883 982
rect 7914 771 7972 783
rect 14212 778 14224 1154
rect 14258 778 14270 1154
rect 14212 766 14270 778
rect 14330 1154 14388 1166
rect 14330 778 14342 1154
rect 14376 778 14388 1154
rect 14330 766 14388 778
rect 14448 1154 14506 1166
rect 14448 778 14460 1154
rect 14494 778 14506 1154
rect 14565 1154 14623 1166
rect 14565 978 14577 1154
rect 14611 978 14623 1154
rect 14565 966 14623 978
rect 14683 1154 14741 1166
rect 15569 1165 15627 1177
rect 15687 1353 15745 1365
rect 15687 1177 15699 1353
rect 15733 1177 15745 1353
rect 15687 1165 15745 1177
rect 15989 1353 16047 1365
rect 14683 978 14695 1154
rect 14729 978 14741 1154
rect 14683 966 14741 978
rect 15989 977 16001 1353
rect 16035 977 16047 1353
rect 15989 965 16047 977
rect 16107 1353 16165 1365
rect 16107 977 16119 1353
rect 16153 977 16165 1353
rect 16107 965 16165 977
rect 16225 1353 16283 1365
rect 16225 977 16237 1353
rect 16271 977 16283 1353
rect 16225 965 16283 977
rect 16343 1353 16401 1365
rect 16343 977 16355 1353
rect 16389 977 16401 1353
rect 16343 965 16401 977
rect 16461 1353 16519 1365
rect 16461 977 16473 1353
rect 16507 977 16519 1353
rect 16867 1353 16925 1365
rect 16867 1177 16879 1353
rect 16913 1177 16925 1353
rect 16867 1165 16925 1177
rect 16985 1353 17043 1365
rect 16985 1177 16997 1353
rect 17031 1177 17043 1353
rect 16985 1165 17043 1177
rect 17467 1353 17525 1365
rect 17467 1177 17479 1353
rect 17513 1177 17525 1353
rect 17467 1165 17525 1177
rect 17585 1353 17643 1365
rect 17585 1177 17597 1353
rect 17631 1177 17643 1353
rect 17585 1165 17643 1177
rect 17887 1353 17945 1365
rect 16461 965 16519 977
rect 17887 977 17899 1353
rect 17933 977 17945 1353
rect 17887 965 17945 977
rect 18005 1353 18063 1365
rect 18005 977 18017 1353
rect 18051 977 18063 1353
rect 18005 965 18063 977
rect 18123 1353 18181 1365
rect 18123 977 18135 1353
rect 18169 977 18181 1353
rect 18123 965 18181 977
rect 18241 1353 18299 1365
rect 18241 977 18253 1353
rect 18287 977 18299 1353
rect 18241 965 18299 977
rect 18359 1353 18417 1365
rect 18359 977 18371 1353
rect 18405 977 18417 1353
rect 18765 1353 18823 1365
rect 18765 1177 18777 1353
rect 18811 1177 18823 1353
rect 18765 1165 18823 1177
rect 18883 1353 18941 1365
rect 18883 1177 18895 1353
rect 18929 1177 18941 1353
rect 18883 1165 18941 1177
rect 22127 1357 22185 1369
rect 22127 1181 22139 1357
rect 22173 1181 22185 1357
rect 20770 1158 20828 1170
rect 18359 965 18417 977
rect 14448 766 14506 778
rect 20770 782 20782 1158
rect 20816 782 20828 1158
rect 20770 770 20828 782
rect 20888 1158 20946 1170
rect 20888 782 20900 1158
rect 20934 782 20946 1158
rect 20888 770 20946 782
rect 21006 1158 21064 1170
rect 21006 782 21018 1158
rect 21052 782 21064 1158
rect 21123 1158 21181 1170
rect 21123 982 21135 1158
rect 21169 982 21181 1158
rect 21123 970 21181 982
rect 21241 1158 21299 1170
rect 22127 1169 22185 1181
rect 22245 1357 22303 1369
rect 22245 1181 22257 1357
rect 22291 1181 22303 1357
rect 22245 1169 22303 1181
rect 22547 1357 22605 1369
rect 21241 982 21253 1158
rect 21287 982 21299 1158
rect 21241 970 21299 982
rect 22547 981 22559 1357
rect 22593 981 22605 1357
rect 22547 969 22605 981
rect 22665 1357 22723 1369
rect 22665 981 22677 1357
rect 22711 981 22723 1357
rect 22665 969 22723 981
rect 22783 1357 22841 1369
rect 22783 981 22795 1357
rect 22829 981 22841 1357
rect 22783 969 22841 981
rect 22901 1357 22959 1369
rect 22901 981 22913 1357
rect 22947 981 22959 1357
rect 22901 969 22959 981
rect 23019 1357 23077 1369
rect 23019 981 23031 1357
rect 23065 981 23077 1357
rect 23425 1357 23483 1369
rect 23425 1181 23437 1357
rect 23471 1181 23483 1357
rect 23425 1169 23483 1181
rect 23543 1357 23601 1369
rect 23543 1181 23555 1357
rect 23589 1181 23601 1357
rect 23543 1169 23601 1181
rect 24025 1357 24083 1369
rect 24025 1181 24037 1357
rect 24071 1181 24083 1357
rect 24025 1169 24083 1181
rect 24143 1357 24201 1369
rect 24143 1181 24155 1357
rect 24189 1181 24201 1357
rect 24143 1169 24201 1181
rect 24445 1357 24503 1369
rect 23019 969 23077 981
rect 24445 981 24457 1357
rect 24491 981 24503 1357
rect 24445 969 24503 981
rect 24563 1357 24621 1369
rect 24563 981 24575 1357
rect 24609 981 24621 1357
rect 24563 969 24621 981
rect 24681 1357 24739 1369
rect 24681 981 24693 1357
rect 24727 981 24739 1357
rect 24681 969 24739 981
rect 24799 1357 24857 1369
rect 24799 981 24811 1357
rect 24845 981 24857 1357
rect 24799 969 24857 981
rect 24917 1357 24975 1369
rect 24917 981 24929 1357
rect 24963 981 24975 1357
rect 25323 1357 25381 1369
rect 25323 1181 25335 1357
rect 25369 1181 25381 1357
rect 25323 1169 25381 1181
rect 25441 1357 25499 1369
rect 25441 1181 25453 1357
rect 25487 1181 25499 1357
rect 25441 1169 25499 1181
rect 24917 969 24975 981
rect 21006 770 21064 782
rect 1374 -1462 1432 -1450
rect 1374 -1638 1386 -1462
rect 1420 -1638 1432 -1462
rect 1374 -1650 1432 -1638
rect 1492 -1462 1550 -1450
rect 1492 -1638 1504 -1462
rect 1538 -1638 1550 -1462
rect 1492 -1650 1550 -1638
rect 1610 -1462 1668 -1450
rect 1610 -1638 1622 -1462
rect 1656 -1638 1668 -1462
rect 1610 -1650 1668 -1638
rect 1728 -1462 1786 -1450
rect 4397 -1192 4455 -1180
rect 4397 -1368 4409 -1192
rect 4443 -1368 4455 -1192
rect 4397 -1380 4455 -1368
rect 4515 -1192 4573 -1180
rect 4515 -1368 4527 -1192
rect 4561 -1368 4573 -1192
rect 4515 -1380 4573 -1368
rect 4632 -1192 4690 -1180
rect 1728 -1638 1740 -1462
rect 1774 -1638 1786 -1462
rect 1728 -1650 1786 -1638
rect 2516 -1466 2574 -1454
rect 2516 -1642 2528 -1466
rect 2562 -1642 2574 -1466
rect 2516 -1654 2574 -1642
rect 2634 -1466 2692 -1454
rect 2634 -1642 2646 -1466
rect 2680 -1642 2692 -1466
rect 2634 -1654 2692 -1642
rect 2752 -1466 2810 -1454
rect 2752 -1642 2764 -1466
rect 2798 -1642 2810 -1466
rect 2752 -1654 2810 -1642
rect 2870 -1466 2928 -1454
rect 2870 -1642 2882 -1466
rect 2916 -1642 2928 -1466
rect 4632 -1568 4644 -1192
rect 4678 -1568 4690 -1192
rect 4632 -1580 4690 -1568
rect 4750 -1192 4808 -1180
rect 4750 -1568 4762 -1192
rect 4796 -1568 4808 -1192
rect 4750 -1580 4808 -1568
rect 4868 -1192 4926 -1180
rect 4868 -1568 4880 -1192
rect 4914 -1568 4926 -1192
rect 4868 -1580 4926 -1568
rect 2870 -1654 2928 -1642
rect 7932 -1466 7990 -1454
rect 7932 -1642 7944 -1466
rect 7978 -1642 7990 -1466
rect 7932 -1654 7990 -1642
rect 8050 -1466 8108 -1454
rect 8050 -1642 8062 -1466
rect 8096 -1642 8108 -1466
rect 8050 -1654 8108 -1642
rect 8168 -1466 8226 -1454
rect 8168 -1642 8180 -1466
rect 8214 -1642 8226 -1466
rect 8168 -1654 8226 -1642
rect 8286 -1466 8344 -1454
rect 10955 -1196 11013 -1184
rect 10955 -1372 10967 -1196
rect 11001 -1372 11013 -1196
rect 10955 -1384 11013 -1372
rect 11073 -1196 11131 -1184
rect 11073 -1372 11085 -1196
rect 11119 -1372 11131 -1196
rect 11073 -1384 11131 -1372
rect 11190 -1196 11248 -1184
rect 8286 -1642 8298 -1466
rect 8332 -1642 8344 -1466
rect 8286 -1654 8344 -1642
rect 9074 -1470 9132 -1458
rect 9074 -1646 9086 -1470
rect 9120 -1646 9132 -1470
rect 9074 -1658 9132 -1646
rect 9192 -1470 9250 -1458
rect 9192 -1646 9204 -1470
rect 9238 -1646 9250 -1470
rect 9192 -1658 9250 -1646
rect 9310 -1470 9368 -1458
rect 9310 -1646 9322 -1470
rect 9356 -1646 9368 -1470
rect 9310 -1658 9368 -1646
rect 9428 -1470 9486 -1458
rect 9428 -1646 9440 -1470
rect 9474 -1646 9486 -1470
rect 11190 -1572 11202 -1196
rect 11236 -1572 11248 -1196
rect 11190 -1584 11248 -1572
rect 11308 -1196 11366 -1184
rect 11308 -1572 11320 -1196
rect 11354 -1572 11366 -1196
rect 11308 -1584 11366 -1572
rect 11426 -1196 11484 -1184
rect 11426 -1572 11438 -1196
rect 11472 -1572 11484 -1196
rect 11426 -1584 11484 -1572
rect 9428 -1658 9486 -1646
rect 14466 -1461 14524 -1449
rect 14466 -1637 14478 -1461
rect 14512 -1637 14524 -1461
rect 14466 -1649 14524 -1637
rect 14584 -1461 14642 -1449
rect 14584 -1637 14596 -1461
rect 14630 -1637 14642 -1461
rect 14584 -1649 14642 -1637
rect 14702 -1461 14760 -1449
rect 14702 -1637 14714 -1461
rect 14748 -1637 14760 -1461
rect 14702 -1649 14760 -1637
rect 14820 -1461 14878 -1449
rect 17489 -1191 17547 -1179
rect 17489 -1367 17501 -1191
rect 17535 -1367 17547 -1191
rect 17489 -1379 17547 -1367
rect 17607 -1191 17665 -1179
rect 17607 -1367 17619 -1191
rect 17653 -1367 17665 -1191
rect 17607 -1379 17665 -1367
rect 17724 -1191 17782 -1179
rect 14820 -1637 14832 -1461
rect 14866 -1637 14878 -1461
rect 14820 -1649 14878 -1637
rect 15608 -1465 15666 -1453
rect 15608 -1641 15620 -1465
rect 15654 -1641 15666 -1465
rect 15608 -1653 15666 -1641
rect 15726 -1465 15784 -1453
rect 15726 -1641 15738 -1465
rect 15772 -1641 15784 -1465
rect 15726 -1653 15784 -1641
rect 15844 -1465 15902 -1453
rect 15844 -1641 15856 -1465
rect 15890 -1641 15902 -1465
rect 15844 -1653 15902 -1641
rect 15962 -1465 16020 -1453
rect 15962 -1641 15974 -1465
rect 16008 -1641 16020 -1465
rect 17724 -1567 17736 -1191
rect 17770 -1567 17782 -1191
rect 17724 -1579 17782 -1567
rect 17842 -1191 17900 -1179
rect 17842 -1567 17854 -1191
rect 17888 -1567 17900 -1191
rect 17842 -1579 17900 -1567
rect 17960 -1191 18018 -1179
rect 17960 -1567 17972 -1191
rect 18006 -1567 18018 -1191
rect 17960 -1579 18018 -1567
rect 15962 -1653 16020 -1641
rect 20979 -1458 21037 -1446
rect 20979 -1634 20991 -1458
rect 21025 -1634 21037 -1458
rect 20979 -1646 21037 -1634
rect 21097 -1458 21155 -1446
rect 21097 -1634 21109 -1458
rect 21143 -1634 21155 -1458
rect 21097 -1646 21155 -1634
rect 21215 -1458 21273 -1446
rect 21215 -1634 21227 -1458
rect 21261 -1634 21273 -1458
rect 21215 -1646 21273 -1634
rect 21333 -1458 21391 -1446
rect 24002 -1188 24060 -1176
rect 24002 -1364 24014 -1188
rect 24048 -1364 24060 -1188
rect 24002 -1376 24060 -1364
rect 24120 -1188 24178 -1176
rect 24120 -1364 24132 -1188
rect 24166 -1364 24178 -1188
rect 24120 -1376 24178 -1364
rect 24237 -1188 24295 -1176
rect 21333 -1634 21345 -1458
rect 21379 -1634 21391 -1458
rect 21333 -1646 21391 -1634
rect 22121 -1462 22179 -1450
rect 22121 -1638 22133 -1462
rect 22167 -1638 22179 -1462
rect 22121 -1650 22179 -1638
rect 22239 -1462 22297 -1450
rect 22239 -1638 22251 -1462
rect 22285 -1638 22297 -1462
rect 22239 -1650 22297 -1638
rect 22357 -1462 22415 -1450
rect 22357 -1638 22369 -1462
rect 22403 -1638 22415 -1462
rect 22357 -1650 22415 -1638
rect 22475 -1462 22533 -1450
rect 22475 -1638 22487 -1462
rect 22521 -1638 22533 -1462
rect 24237 -1564 24249 -1188
rect 24283 -1564 24295 -1188
rect 24237 -1576 24295 -1564
rect 24355 -1188 24413 -1176
rect 24355 -1564 24367 -1188
rect 24401 -1564 24413 -1188
rect 24355 -1576 24413 -1564
rect 24473 -1188 24531 -1176
rect 24473 -1564 24485 -1188
rect 24519 -1564 24531 -1188
rect 24473 -1576 24531 -1564
rect 22475 -1650 22533 -1638
rect 4383 -2842 4441 -2830
rect 4383 -3018 4395 -2842
rect 4429 -3018 4441 -2842
rect 4383 -3030 4441 -3018
rect 4501 -2842 4559 -2830
rect 4501 -3018 4513 -2842
rect 4547 -3018 4559 -2842
rect 4501 -3030 4559 -3018
rect 4618 -2842 4676 -2830
rect 4618 -3218 4630 -2842
rect 4664 -3218 4676 -2842
rect 4618 -3230 4676 -3218
rect 4736 -2842 4794 -2830
rect 4736 -3218 4748 -2842
rect 4782 -3218 4794 -2842
rect 4736 -3230 4794 -3218
rect 4854 -2842 4912 -2830
rect 4854 -3218 4866 -2842
rect 4900 -3218 4912 -2842
rect 10941 -2846 10999 -2834
rect 10941 -3022 10953 -2846
rect 10987 -3022 10999 -2846
rect 10941 -3034 10999 -3022
rect 11059 -2846 11117 -2834
rect 11059 -3022 11071 -2846
rect 11105 -3022 11117 -2846
rect 11059 -3034 11117 -3022
rect 11176 -2846 11234 -2834
rect 4854 -3230 4912 -3218
rect 188 -4247 246 -4235
rect 188 -4423 200 -4247
rect 234 -4423 246 -4247
rect 188 -4435 246 -4423
rect 306 -4247 364 -4235
rect 306 -4423 318 -4247
rect 352 -4423 364 -4247
rect 306 -4435 364 -4423
rect 712 -4247 770 -4235
rect 712 -4623 724 -4247
rect 758 -4623 770 -4247
rect 712 -4635 770 -4623
rect 830 -4247 888 -4235
rect 830 -4623 842 -4247
rect 876 -4623 888 -4247
rect 830 -4635 888 -4623
rect 948 -4247 1006 -4235
rect 948 -4623 960 -4247
rect 994 -4623 1006 -4247
rect 948 -4635 1006 -4623
rect 1066 -4247 1124 -4235
rect 1066 -4623 1078 -4247
rect 1112 -4623 1124 -4247
rect 1066 -4635 1124 -4623
rect 1184 -4247 1242 -4235
rect 1184 -4623 1196 -4247
rect 1230 -4623 1242 -4247
rect 1486 -4247 1544 -4235
rect 1486 -4423 1498 -4247
rect 1532 -4423 1544 -4247
rect 1486 -4435 1544 -4423
rect 1604 -4247 1662 -4235
rect 1604 -4423 1616 -4247
rect 1650 -4423 1662 -4247
rect 1604 -4435 1662 -4423
rect 2086 -4247 2144 -4235
rect 2086 -4423 2098 -4247
rect 2132 -4423 2144 -4247
rect 2086 -4435 2144 -4423
rect 2204 -4247 2262 -4235
rect 2204 -4423 2216 -4247
rect 2250 -4423 2262 -4247
rect 2204 -4435 2262 -4423
rect 2610 -4247 2668 -4235
rect 1184 -4635 1242 -4623
rect 2610 -4623 2622 -4247
rect 2656 -4623 2668 -4247
rect 2610 -4635 2668 -4623
rect 2728 -4247 2786 -4235
rect 2728 -4623 2740 -4247
rect 2774 -4623 2786 -4247
rect 2728 -4635 2786 -4623
rect 2846 -4247 2904 -4235
rect 2846 -4623 2858 -4247
rect 2892 -4623 2904 -4247
rect 2846 -4635 2904 -4623
rect 2964 -4247 3022 -4235
rect 2964 -4623 2976 -4247
rect 3010 -4623 3022 -4247
rect 2964 -4635 3022 -4623
rect 3082 -4247 3140 -4235
rect 3082 -4623 3094 -4247
rect 3128 -4623 3140 -4247
rect 3384 -4247 3442 -4235
rect 3384 -4423 3396 -4247
rect 3430 -4423 3442 -4247
rect 3384 -4435 3442 -4423
rect 3502 -4247 3560 -4235
rect 3502 -4423 3514 -4247
rect 3548 -4423 3560 -4247
rect 3502 -4435 3560 -4423
rect 11176 -3222 11188 -2846
rect 11222 -3222 11234 -2846
rect 11176 -3234 11234 -3222
rect 11294 -2846 11352 -2834
rect 11294 -3222 11306 -2846
rect 11340 -3222 11352 -2846
rect 11294 -3234 11352 -3222
rect 11412 -2846 11470 -2834
rect 11412 -3222 11424 -2846
rect 11458 -3222 11470 -2846
rect 17475 -2841 17533 -2829
rect 17475 -3017 17487 -2841
rect 17521 -3017 17533 -2841
rect 17475 -3029 17533 -3017
rect 17593 -2841 17651 -2829
rect 17593 -3017 17605 -2841
rect 17639 -3017 17651 -2841
rect 17593 -3029 17651 -3017
rect 17710 -2841 17768 -2829
rect 11412 -3234 11470 -3222
rect 6746 -4251 6804 -4239
rect 6746 -4427 6758 -4251
rect 6792 -4427 6804 -4251
rect 4388 -4446 4446 -4434
rect 3082 -4635 3140 -4623
rect 4388 -4622 4400 -4446
rect 4434 -4622 4446 -4446
rect 4388 -4634 4446 -4622
rect 4506 -4446 4564 -4434
rect 4506 -4622 4518 -4446
rect 4552 -4622 4564 -4446
rect 4506 -4634 4564 -4622
rect 4623 -4446 4681 -4434
rect 4623 -4822 4635 -4446
rect 4669 -4822 4681 -4446
rect 4623 -4834 4681 -4822
rect 4741 -4446 4799 -4434
rect 4741 -4822 4753 -4446
rect 4787 -4822 4799 -4446
rect 4741 -4834 4799 -4822
rect 4859 -4446 4917 -4434
rect 6746 -4439 6804 -4427
rect 6864 -4251 6922 -4239
rect 6864 -4427 6876 -4251
rect 6910 -4427 6922 -4251
rect 6864 -4439 6922 -4427
rect 7270 -4251 7328 -4239
rect 4859 -4822 4871 -4446
rect 4905 -4822 4917 -4446
rect 7270 -4627 7282 -4251
rect 7316 -4627 7328 -4251
rect 7270 -4639 7328 -4627
rect 7388 -4251 7446 -4239
rect 7388 -4627 7400 -4251
rect 7434 -4627 7446 -4251
rect 7388 -4639 7446 -4627
rect 7506 -4251 7564 -4239
rect 7506 -4627 7518 -4251
rect 7552 -4627 7564 -4251
rect 7506 -4639 7564 -4627
rect 7624 -4251 7682 -4239
rect 7624 -4627 7636 -4251
rect 7670 -4627 7682 -4251
rect 7624 -4639 7682 -4627
rect 7742 -4251 7800 -4239
rect 7742 -4627 7754 -4251
rect 7788 -4627 7800 -4251
rect 8044 -4251 8102 -4239
rect 8044 -4427 8056 -4251
rect 8090 -4427 8102 -4251
rect 8044 -4439 8102 -4427
rect 8162 -4251 8220 -4239
rect 8162 -4427 8174 -4251
rect 8208 -4427 8220 -4251
rect 8162 -4439 8220 -4427
rect 8644 -4251 8702 -4239
rect 8644 -4427 8656 -4251
rect 8690 -4427 8702 -4251
rect 8644 -4439 8702 -4427
rect 8762 -4251 8820 -4239
rect 8762 -4427 8774 -4251
rect 8808 -4427 8820 -4251
rect 8762 -4439 8820 -4427
rect 9168 -4251 9226 -4239
rect 7742 -4639 7800 -4627
rect 9168 -4627 9180 -4251
rect 9214 -4627 9226 -4251
rect 9168 -4639 9226 -4627
rect 9286 -4251 9344 -4239
rect 9286 -4627 9298 -4251
rect 9332 -4627 9344 -4251
rect 9286 -4639 9344 -4627
rect 9404 -4251 9462 -4239
rect 9404 -4627 9416 -4251
rect 9450 -4627 9462 -4251
rect 9404 -4639 9462 -4627
rect 9522 -4251 9580 -4239
rect 9522 -4627 9534 -4251
rect 9568 -4627 9580 -4251
rect 9522 -4639 9580 -4627
rect 9640 -4251 9698 -4239
rect 9640 -4627 9652 -4251
rect 9686 -4627 9698 -4251
rect 9942 -4251 10000 -4239
rect 9942 -4427 9954 -4251
rect 9988 -4427 10000 -4251
rect 9942 -4439 10000 -4427
rect 10060 -4251 10118 -4239
rect 10060 -4427 10072 -4251
rect 10106 -4427 10118 -4251
rect 10060 -4439 10118 -4427
rect 17710 -3217 17722 -2841
rect 17756 -3217 17768 -2841
rect 17710 -3229 17768 -3217
rect 17828 -2841 17886 -2829
rect 17828 -3217 17840 -2841
rect 17874 -3217 17886 -2841
rect 17828 -3229 17886 -3217
rect 17946 -2841 18004 -2829
rect 17946 -3217 17958 -2841
rect 17992 -3217 18004 -2841
rect 23988 -2838 24046 -2826
rect 23988 -3014 24000 -2838
rect 24034 -3014 24046 -2838
rect 23988 -3026 24046 -3014
rect 24106 -2838 24164 -2826
rect 24106 -3014 24118 -2838
rect 24152 -3014 24164 -2838
rect 24106 -3026 24164 -3014
rect 24223 -2838 24281 -2826
rect 17946 -3229 18004 -3217
rect 13280 -4246 13338 -4234
rect 13280 -4422 13292 -4246
rect 13326 -4422 13338 -4246
rect 13280 -4434 13338 -4422
rect 13398 -4246 13456 -4234
rect 13398 -4422 13410 -4246
rect 13444 -4422 13456 -4246
rect 13398 -4434 13456 -4422
rect 13804 -4246 13862 -4234
rect 10946 -4450 11004 -4438
rect 9640 -4639 9698 -4627
rect 10946 -4626 10958 -4450
rect 10992 -4626 11004 -4450
rect 10946 -4638 11004 -4626
rect 11064 -4450 11122 -4438
rect 11064 -4626 11076 -4450
rect 11110 -4626 11122 -4450
rect 11064 -4638 11122 -4626
rect 11181 -4450 11239 -4438
rect 4859 -4834 4917 -4822
rect 11181 -4826 11193 -4450
rect 11227 -4826 11239 -4450
rect 11181 -4838 11239 -4826
rect 11299 -4450 11357 -4438
rect 11299 -4826 11311 -4450
rect 11345 -4826 11357 -4450
rect 11299 -4838 11357 -4826
rect 11417 -4450 11475 -4438
rect 11417 -4826 11429 -4450
rect 11463 -4826 11475 -4450
rect 13804 -4622 13816 -4246
rect 13850 -4622 13862 -4246
rect 13804 -4634 13862 -4622
rect 13922 -4246 13980 -4234
rect 13922 -4622 13934 -4246
rect 13968 -4622 13980 -4246
rect 13922 -4634 13980 -4622
rect 14040 -4246 14098 -4234
rect 14040 -4622 14052 -4246
rect 14086 -4622 14098 -4246
rect 14040 -4634 14098 -4622
rect 14158 -4246 14216 -4234
rect 14158 -4622 14170 -4246
rect 14204 -4622 14216 -4246
rect 14158 -4634 14216 -4622
rect 14276 -4246 14334 -4234
rect 14276 -4622 14288 -4246
rect 14322 -4622 14334 -4246
rect 14578 -4246 14636 -4234
rect 14578 -4422 14590 -4246
rect 14624 -4422 14636 -4246
rect 14578 -4434 14636 -4422
rect 14696 -4246 14754 -4234
rect 14696 -4422 14708 -4246
rect 14742 -4422 14754 -4246
rect 14696 -4434 14754 -4422
rect 15178 -4246 15236 -4234
rect 15178 -4422 15190 -4246
rect 15224 -4422 15236 -4246
rect 15178 -4434 15236 -4422
rect 15296 -4246 15354 -4234
rect 15296 -4422 15308 -4246
rect 15342 -4422 15354 -4246
rect 15296 -4434 15354 -4422
rect 15702 -4246 15760 -4234
rect 14276 -4634 14334 -4622
rect 15702 -4622 15714 -4246
rect 15748 -4622 15760 -4246
rect 15702 -4634 15760 -4622
rect 15820 -4246 15878 -4234
rect 15820 -4622 15832 -4246
rect 15866 -4622 15878 -4246
rect 15820 -4634 15878 -4622
rect 15938 -4246 15996 -4234
rect 15938 -4622 15950 -4246
rect 15984 -4622 15996 -4246
rect 15938 -4634 15996 -4622
rect 16056 -4246 16114 -4234
rect 16056 -4622 16068 -4246
rect 16102 -4622 16114 -4246
rect 16056 -4634 16114 -4622
rect 16174 -4246 16232 -4234
rect 16174 -4622 16186 -4246
rect 16220 -4622 16232 -4246
rect 16476 -4246 16534 -4234
rect 16476 -4422 16488 -4246
rect 16522 -4422 16534 -4246
rect 16476 -4434 16534 -4422
rect 16594 -4246 16652 -4234
rect 16594 -4422 16606 -4246
rect 16640 -4422 16652 -4246
rect 16594 -4434 16652 -4422
rect 24223 -3214 24235 -2838
rect 24269 -3214 24281 -2838
rect 24223 -3226 24281 -3214
rect 24341 -2838 24399 -2826
rect 24341 -3214 24353 -2838
rect 24387 -3214 24399 -2838
rect 24341 -3226 24399 -3214
rect 24459 -2838 24517 -2826
rect 24459 -3214 24471 -2838
rect 24505 -3214 24517 -2838
rect 24459 -3226 24517 -3214
rect 19793 -4243 19851 -4231
rect 19793 -4419 19805 -4243
rect 19839 -4419 19851 -4243
rect 19793 -4431 19851 -4419
rect 19911 -4243 19969 -4231
rect 19911 -4419 19923 -4243
rect 19957 -4419 19969 -4243
rect 19911 -4431 19969 -4419
rect 20317 -4243 20375 -4231
rect 17480 -4445 17538 -4433
rect 16174 -4634 16232 -4622
rect 17480 -4621 17492 -4445
rect 17526 -4621 17538 -4445
rect 17480 -4633 17538 -4621
rect 17598 -4445 17656 -4433
rect 17598 -4621 17610 -4445
rect 17644 -4621 17656 -4445
rect 17598 -4633 17656 -4621
rect 17715 -4445 17773 -4433
rect 11417 -4838 11475 -4826
rect 17715 -4821 17727 -4445
rect 17761 -4821 17773 -4445
rect 17715 -4833 17773 -4821
rect 17833 -4445 17891 -4433
rect 17833 -4821 17845 -4445
rect 17879 -4821 17891 -4445
rect 17833 -4833 17891 -4821
rect 17951 -4445 18009 -4433
rect 17951 -4821 17963 -4445
rect 17997 -4821 18009 -4445
rect 20317 -4619 20329 -4243
rect 20363 -4619 20375 -4243
rect 20317 -4631 20375 -4619
rect 20435 -4243 20493 -4231
rect 20435 -4619 20447 -4243
rect 20481 -4619 20493 -4243
rect 20435 -4631 20493 -4619
rect 20553 -4243 20611 -4231
rect 20553 -4619 20565 -4243
rect 20599 -4619 20611 -4243
rect 20553 -4631 20611 -4619
rect 20671 -4243 20729 -4231
rect 20671 -4619 20683 -4243
rect 20717 -4619 20729 -4243
rect 20671 -4631 20729 -4619
rect 20789 -4243 20847 -4231
rect 20789 -4619 20801 -4243
rect 20835 -4619 20847 -4243
rect 21091 -4243 21149 -4231
rect 21091 -4419 21103 -4243
rect 21137 -4419 21149 -4243
rect 21091 -4431 21149 -4419
rect 21209 -4243 21267 -4231
rect 21209 -4419 21221 -4243
rect 21255 -4419 21267 -4243
rect 21209 -4431 21267 -4419
rect 21691 -4243 21749 -4231
rect 21691 -4419 21703 -4243
rect 21737 -4419 21749 -4243
rect 21691 -4431 21749 -4419
rect 21809 -4243 21867 -4231
rect 21809 -4419 21821 -4243
rect 21855 -4419 21867 -4243
rect 21809 -4431 21867 -4419
rect 22215 -4243 22273 -4231
rect 20789 -4631 20847 -4619
rect 22215 -4619 22227 -4243
rect 22261 -4619 22273 -4243
rect 22215 -4631 22273 -4619
rect 22333 -4243 22391 -4231
rect 22333 -4619 22345 -4243
rect 22379 -4619 22391 -4243
rect 22333 -4631 22391 -4619
rect 22451 -4243 22509 -4231
rect 22451 -4619 22463 -4243
rect 22497 -4619 22509 -4243
rect 22451 -4631 22509 -4619
rect 22569 -4243 22627 -4231
rect 22569 -4619 22581 -4243
rect 22615 -4619 22627 -4243
rect 22569 -4631 22627 -4619
rect 22687 -4243 22745 -4231
rect 22687 -4619 22699 -4243
rect 22733 -4619 22745 -4243
rect 22989 -4243 23047 -4231
rect 22989 -4419 23001 -4243
rect 23035 -4419 23047 -4243
rect 22989 -4431 23047 -4419
rect 23107 -4243 23165 -4231
rect 23107 -4419 23119 -4243
rect 23153 -4419 23165 -4243
rect 23107 -4431 23165 -4419
rect 23993 -4442 24051 -4430
rect 22687 -4631 22745 -4619
rect 23993 -4618 24005 -4442
rect 24039 -4618 24051 -4442
rect 23993 -4630 24051 -4618
rect 24111 -4442 24169 -4430
rect 24111 -4618 24123 -4442
rect 24157 -4618 24169 -4442
rect 24111 -4630 24169 -4618
rect 24228 -4442 24286 -4430
rect 17951 -4833 18009 -4821
rect 24228 -4818 24240 -4442
rect 24274 -4818 24286 -4442
rect 24228 -4830 24286 -4818
rect 24346 -4442 24404 -4430
rect 24346 -4818 24358 -4442
rect 24392 -4818 24404 -4442
rect 24346 -4830 24404 -4818
rect 24464 -4442 24522 -4430
rect 24464 -4818 24476 -4442
rect 24510 -4818 24522 -4442
rect 24464 -4830 24522 -4818
<< pdiff >>
rect 3244 4925 3302 4937
rect 919 4853 977 4865
rect 919 4677 931 4853
rect 965 4677 977 4853
rect 919 4665 977 4677
rect 1037 4853 1095 4865
rect 1037 4677 1049 4853
rect 1083 4677 1095 4853
rect 1037 4665 1095 4677
rect 1155 4853 1213 4865
rect 1155 4677 1167 4853
rect 1201 4677 1213 4853
rect 1155 4665 1213 4677
rect 1273 4853 1331 4865
rect 1273 4677 1285 4853
rect 1319 4677 1331 4853
rect 1273 4665 1331 4677
rect 1391 4853 1449 4865
rect 1391 4677 1403 4853
rect 1437 4677 1449 4853
rect 1391 4665 1449 4677
rect 1509 4853 1567 4865
rect 1509 4677 1521 4853
rect 1555 4677 1567 4853
rect 1509 4665 1567 4677
rect 1627 4853 1685 4865
rect 1627 4677 1639 4853
rect 1673 4677 1685 4853
rect 1627 4665 1685 4677
rect 1745 4853 1803 4865
rect 1745 4677 1757 4853
rect 1791 4677 1803 4853
rect 1745 4665 1803 4677
rect 1863 4853 1921 4865
rect 1863 4677 1875 4853
rect 1909 4677 1921 4853
rect 1863 4665 1921 4677
rect 1981 4853 2039 4865
rect 1981 4677 1993 4853
rect 2027 4677 2039 4853
rect 1981 4665 2039 4677
rect 3244 4549 3256 4925
rect 3290 4549 3302 4925
rect 3244 4537 3302 4549
rect 3362 4925 3420 4937
rect 3362 4549 3374 4925
rect 3408 4549 3420 4925
rect 3362 4537 3420 4549
rect 3480 4925 3538 4937
rect 3480 4549 3492 4925
rect 3526 4549 3538 4925
rect 3480 4537 3538 4549
rect 3598 4925 3656 4937
rect 3598 4549 3610 4925
rect 3644 4549 3656 4925
rect 3598 4537 3656 4549
rect 3716 4925 3774 4937
rect 3716 4549 3728 4925
rect 3762 4549 3774 4925
rect 3716 4537 3774 4549
rect 3834 4925 3892 4937
rect 3834 4549 3846 4925
rect 3880 4549 3892 4925
rect 3834 4537 3892 4549
rect 3952 4925 4010 4937
rect 3952 4549 3964 4925
rect 3998 4549 4010 4925
rect 3952 4537 4010 4549
rect 4386 4929 4444 4941
rect 4386 4553 4398 4929
rect 4432 4553 4444 4929
rect 4386 4541 4444 4553
rect 4504 4929 4562 4941
rect 4504 4553 4516 4929
rect 4550 4553 4562 4929
rect 4504 4541 4562 4553
rect 4622 4929 4680 4941
rect 4622 4553 4634 4929
rect 4668 4553 4680 4929
rect 4622 4541 4680 4553
rect 4740 4929 4798 4941
rect 4740 4553 4752 4929
rect 4786 4553 4798 4929
rect 4740 4541 4798 4553
rect 4858 4929 4916 4941
rect 4858 4553 4870 4929
rect 4904 4553 4916 4929
rect 4858 4541 4916 4553
rect 4976 4929 5034 4941
rect 4976 4553 4988 4929
rect 5022 4553 5034 4929
rect 4976 4541 5034 4553
rect 5094 4929 5152 4941
rect 5094 4553 5106 4929
rect 5140 4553 5152 4929
rect 9757 4922 9815 4934
rect 7432 4850 7490 4862
rect 7432 4674 7444 4850
rect 7478 4674 7490 4850
rect 7432 4662 7490 4674
rect 7550 4850 7608 4862
rect 7550 4674 7562 4850
rect 7596 4674 7608 4850
rect 7550 4662 7608 4674
rect 7668 4850 7726 4862
rect 7668 4674 7680 4850
rect 7714 4674 7726 4850
rect 7668 4662 7726 4674
rect 7786 4850 7844 4862
rect 7786 4674 7798 4850
rect 7832 4674 7844 4850
rect 7786 4662 7844 4674
rect 7904 4850 7962 4862
rect 7904 4674 7916 4850
rect 7950 4674 7962 4850
rect 7904 4662 7962 4674
rect 8022 4850 8080 4862
rect 8022 4674 8034 4850
rect 8068 4674 8080 4850
rect 8022 4662 8080 4674
rect 8140 4850 8198 4862
rect 8140 4674 8152 4850
rect 8186 4674 8198 4850
rect 8140 4662 8198 4674
rect 8258 4850 8316 4862
rect 8258 4674 8270 4850
rect 8304 4674 8316 4850
rect 8258 4662 8316 4674
rect 8376 4850 8434 4862
rect 8376 4674 8388 4850
rect 8422 4674 8434 4850
rect 8376 4662 8434 4674
rect 8494 4850 8552 4862
rect 8494 4674 8506 4850
rect 8540 4674 8552 4850
rect 8494 4662 8552 4674
rect 5094 4541 5152 4553
rect 9757 4546 9769 4922
rect 9803 4546 9815 4922
rect 9757 4534 9815 4546
rect 9875 4922 9933 4934
rect 9875 4546 9887 4922
rect 9921 4546 9933 4922
rect 9875 4534 9933 4546
rect 9993 4922 10051 4934
rect 9993 4546 10005 4922
rect 10039 4546 10051 4922
rect 9993 4534 10051 4546
rect 10111 4922 10169 4934
rect 10111 4546 10123 4922
rect 10157 4546 10169 4922
rect 10111 4534 10169 4546
rect 10229 4922 10287 4934
rect 10229 4546 10241 4922
rect 10275 4546 10287 4922
rect 10229 4534 10287 4546
rect 10347 4922 10405 4934
rect 10347 4546 10359 4922
rect 10393 4546 10405 4922
rect 10347 4534 10405 4546
rect 10465 4922 10523 4934
rect 10465 4546 10477 4922
rect 10511 4546 10523 4922
rect 10465 4534 10523 4546
rect 10899 4926 10957 4938
rect 10899 4550 10911 4926
rect 10945 4550 10957 4926
rect 10899 4538 10957 4550
rect 11017 4926 11075 4938
rect 11017 4550 11029 4926
rect 11063 4550 11075 4926
rect 11017 4538 11075 4550
rect 11135 4926 11193 4938
rect 11135 4550 11147 4926
rect 11181 4550 11193 4926
rect 11135 4538 11193 4550
rect 11253 4926 11311 4938
rect 11253 4550 11265 4926
rect 11299 4550 11311 4926
rect 11253 4538 11311 4550
rect 11371 4926 11429 4938
rect 11371 4550 11383 4926
rect 11417 4550 11429 4926
rect 11371 4538 11429 4550
rect 11489 4926 11547 4938
rect 11489 4550 11501 4926
rect 11535 4550 11547 4926
rect 11489 4538 11547 4550
rect 11607 4926 11665 4938
rect 11607 4550 11619 4926
rect 11653 4550 11665 4926
rect 16291 4917 16349 4929
rect 13966 4845 14024 4857
rect 13966 4669 13978 4845
rect 14012 4669 14024 4845
rect 13966 4657 14024 4669
rect 14084 4845 14142 4857
rect 14084 4669 14096 4845
rect 14130 4669 14142 4845
rect 14084 4657 14142 4669
rect 14202 4845 14260 4857
rect 14202 4669 14214 4845
rect 14248 4669 14260 4845
rect 14202 4657 14260 4669
rect 14320 4845 14378 4857
rect 14320 4669 14332 4845
rect 14366 4669 14378 4845
rect 14320 4657 14378 4669
rect 14438 4845 14496 4857
rect 14438 4669 14450 4845
rect 14484 4669 14496 4845
rect 14438 4657 14496 4669
rect 14556 4845 14614 4857
rect 14556 4669 14568 4845
rect 14602 4669 14614 4845
rect 14556 4657 14614 4669
rect 14674 4845 14732 4857
rect 14674 4669 14686 4845
rect 14720 4669 14732 4845
rect 14674 4657 14732 4669
rect 14792 4845 14850 4857
rect 14792 4669 14804 4845
rect 14838 4669 14850 4845
rect 14792 4657 14850 4669
rect 14910 4845 14968 4857
rect 14910 4669 14922 4845
rect 14956 4669 14968 4845
rect 14910 4657 14968 4669
rect 15028 4845 15086 4857
rect 15028 4669 15040 4845
rect 15074 4669 15086 4845
rect 15028 4657 15086 4669
rect 11607 4538 11665 4550
rect 3673 4142 3731 4154
rect 3673 3966 3685 4142
rect 3719 3966 3731 4142
rect 3673 3954 3731 3966
rect 3791 4142 3849 4154
rect 3791 3966 3803 4142
rect 3837 3966 3849 4142
rect 3791 3954 3849 3966
rect 3909 4142 3967 4154
rect 3909 3966 3921 4142
rect 3955 3966 3967 4142
rect 3909 3954 3967 3966
rect 4027 4142 4085 4154
rect 4027 3966 4039 4142
rect 4073 3966 4085 4142
rect 4027 3954 4085 3966
rect 4815 4146 4873 4158
rect 4815 3970 4827 4146
rect 4861 3970 4873 4146
rect 4815 3958 4873 3970
rect 4933 4146 4991 4158
rect 4933 3970 4945 4146
rect 4979 3970 4991 4146
rect 4933 3958 4991 3970
rect 5051 4146 5109 4158
rect 5051 3970 5063 4146
rect 5097 3970 5109 4146
rect 5051 3958 5109 3970
rect 5169 4146 5227 4158
rect 5169 3970 5181 4146
rect 5215 3970 5227 4146
rect 16291 4541 16303 4917
rect 16337 4541 16349 4917
rect 16291 4529 16349 4541
rect 16409 4917 16467 4929
rect 16409 4541 16421 4917
rect 16455 4541 16467 4917
rect 16409 4529 16467 4541
rect 16527 4917 16585 4929
rect 16527 4541 16539 4917
rect 16573 4541 16585 4917
rect 16527 4529 16585 4541
rect 16645 4917 16703 4929
rect 16645 4541 16657 4917
rect 16691 4541 16703 4917
rect 16645 4529 16703 4541
rect 16763 4917 16821 4929
rect 16763 4541 16775 4917
rect 16809 4541 16821 4917
rect 16763 4529 16821 4541
rect 16881 4917 16939 4929
rect 16881 4541 16893 4917
rect 16927 4541 16939 4917
rect 16881 4529 16939 4541
rect 16999 4917 17057 4929
rect 16999 4541 17011 4917
rect 17045 4541 17057 4917
rect 16999 4529 17057 4541
rect 17433 4921 17491 4933
rect 17433 4545 17445 4921
rect 17479 4545 17491 4921
rect 17433 4533 17491 4545
rect 17551 4921 17609 4933
rect 17551 4545 17563 4921
rect 17597 4545 17609 4921
rect 17551 4533 17609 4545
rect 17669 4921 17727 4933
rect 17669 4545 17681 4921
rect 17715 4545 17727 4921
rect 17669 4533 17727 4545
rect 17787 4921 17845 4933
rect 17787 4545 17799 4921
rect 17833 4545 17845 4921
rect 17787 4533 17845 4545
rect 17905 4921 17963 4933
rect 17905 4545 17917 4921
rect 17951 4545 17963 4921
rect 17905 4533 17963 4545
rect 18023 4921 18081 4933
rect 18023 4545 18035 4921
rect 18069 4545 18081 4921
rect 18023 4533 18081 4545
rect 18141 4921 18199 4933
rect 18141 4545 18153 4921
rect 18187 4545 18199 4921
rect 22849 4921 22907 4933
rect 20524 4849 20582 4861
rect 20524 4673 20536 4849
rect 20570 4673 20582 4849
rect 20524 4661 20582 4673
rect 20642 4849 20700 4861
rect 20642 4673 20654 4849
rect 20688 4673 20700 4849
rect 20642 4661 20700 4673
rect 20760 4849 20818 4861
rect 20760 4673 20772 4849
rect 20806 4673 20818 4849
rect 20760 4661 20818 4673
rect 20878 4849 20936 4861
rect 20878 4673 20890 4849
rect 20924 4673 20936 4849
rect 20878 4661 20936 4673
rect 20996 4849 21054 4861
rect 20996 4673 21008 4849
rect 21042 4673 21054 4849
rect 20996 4661 21054 4673
rect 21114 4849 21172 4861
rect 21114 4673 21126 4849
rect 21160 4673 21172 4849
rect 21114 4661 21172 4673
rect 21232 4849 21290 4861
rect 21232 4673 21244 4849
rect 21278 4673 21290 4849
rect 21232 4661 21290 4673
rect 21350 4849 21408 4861
rect 21350 4673 21362 4849
rect 21396 4673 21408 4849
rect 21350 4661 21408 4673
rect 21468 4849 21526 4861
rect 21468 4673 21480 4849
rect 21514 4673 21526 4849
rect 21468 4661 21526 4673
rect 21586 4849 21644 4861
rect 21586 4673 21598 4849
rect 21632 4673 21644 4849
rect 21586 4661 21644 4673
rect 18141 4533 18199 4545
rect 5169 3958 5227 3970
rect 10186 4139 10244 4151
rect 10186 3963 10198 4139
rect 10232 3963 10244 4139
rect 10186 3951 10244 3963
rect 10304 4139 10362 4151
rect 10304 3963 10316 4139
rect 10350 3963 10362 4139
rect 10304 3951 10362 3963
rect 10422 4139 10480 4151
rect 10422 3963 10434 4139
rect 10468 3963 10480 4139
rect 10422 3951 10480 3963
rect 10540 4139 10598 4151
rect 10540 3963 10552 4139
rect 10586 3963 10598 4139
rect 10540 3951 10598 3963
rect 11328 4143 11386 4155
rect 11328 3967 11340 4143
rect 11374 3967 11386 4143
rect 11328 3955 11386 3967
rect 11446 4143 11504 4155
rect 11446 3967 11458 4143
rect 11492 3967 11504 4143
rect 11446 3955 11504 3967
rect 11564 4143 11622 4155
rect 11564 3967 11576 4143
rect 11610 3967 11622 4143
rect 11564 3955 11622 3967
rect 11682 4143 11740 4155
rect 11682 3967 11694 4143
rect 11728 3967 11740 4143
rect 22849 4545 22861 4921
rect 22895 4545 22907 4921
rect 22849 4533 22907 4545
rect 22967 4921 23025 4933
rect 22967 4545 22979 4921
rect 23013 4545 23025 4921
rect 22967 4533 23025 4545
rect 23085 4921 23143 4933
rect 23085 4545 23097 4921
rect 23131 4545 23143 4921
rect 23085 4533 23143 4545
rect 23203 4921 23261 4933
rect 23203 4545 23215 4921
rect 23249 4545 23261 4921
rect 23203 4533 23261 4545
rect 23321 4921 23379 4933
rect 23321 4545 23333 4921
rect 23367 4545 23379 4921
rect 23321 4533 23379 4545
rect 23439 4921 23497 4933
rect 23439 4545 23451 4921
rect 23485 4545 23497 4921
rect 23439 4533 23497 4545
rect 23557 4921 23615 4933
rect 23557 4545 23569 4921
rect 23603 4545 23615 4921
rect 23557 4533 23615 4545
rect 23991 4925 24049 4937
rect 23991 4549 24003 4925
rect 24037 4549 24049 4925
rect 23991 4537 24049 4549
rect 24109 4925 24167 4937
rect 24109 4549 24121 4925
rect 24155 4549 24167 4925
rect 24109 4537 24167 4549
rect 24227 4925 24285 4937
rect 24227 4549 24239 4925
rect 24273 4549 24285 4925
rect 24227 4537 24285 4549
rect 24345 4925 24403 4937
rect 24345 4549 24357 4925
rect 24391 4549 24403 4925
rect 24345 4537 24403 4549
rect 24463 4925 24521 4937
rect 24463 4549 24475 4925
rect 24509 4549 24521 4925
rect 24463 4537 24521 4549
rect 24581 4925 24639 4937
rect 24581 4549 24593 4925
rect 24627 4549 24639 4925
rect 24581 4537 24639 4549
rect 24699 4925 24757 4937
rect 24699 4549 24711 4925
rect 24745 4549 24757 4925
rect 24699 4537 24757 4549
rect 11682 3955 11740 3967
rect 16720 4134 16778 4146
rect 16720 3958 16732 4134
rect 16766 3958 16778 4134
rect 16720 3946 16778 3958
rect 16838 4134 16896 4146
rect 16838 3958 16850 4134
rect 16884 3958 16896 4134
rect 16838 3946 16896 3958
rect 16956 4134 17014 4146
rect 16956 3958 16968 4134
rect 17002 3958 17014 4134
rect 16956 3946 17014 3958
rect 17074 4134 17132 4146
rect 17074 3958 17086 4134
rect 17120 3958 17132 4134
rect 17074 3946 17132 3958
rect 17862 4138 17920 4150
rect 17862 3962 17874 4138
rect 17908 3962 17920 4138
rect 17862 3950 17920 3962
rect 17980 4138 18038 4150
rect 17980 3962 17992 4138
rect 18026 3962 18038 4138
rect 17980 3950 18038 3962
rect 18098 4138 18156 4150
rect 18098 3962 18110 4138
rect 18144 3962 18156 4138
rect 18098 3950 18156 3962
rect 18216 4138 18274 4150
rect 18216 3962 18228 4138
rect 18262 3962 18274 4138
rect 18216 3950 18274 3962
rect 23278 4138 23336 4150
rect 23278 3962 23290 4138
rect 23324 3962 23336 4138
rect 23278 3950 23336 3962
rect 23396 4138 23454 4150
rect 23396 3962 23408 4138
rect 23442 3962 23454 4138
rect 23396 3950 23454 3962
rect 23514 4138 23572 4150
rect 23514 3962 23526 4138
rect 23560 3962 23572 4138
rect 23514 3950 23572 3962
rect 23632 4138 23690 4150
rect 23632 3962 23644 4138
rect 23678 3962 23690 4138
rect 23632 3950 23690 3962
rect 24420 4142 24478 4154
rect 24420 3966 24432 4142
rect 24466 3966 24478 4142
rect 24420 3954 24478 3966
rect 24538 4142 24596 4154
rect 24538 3966 24550 4142
rect 24584 3966 24596 4142
rect 24538 3954 24596 3966
rect 24656 4142 24714 4154
rect 24656 3966 24668 4142
rect 24702 3966 24714 4142
rect 24656 3954 24714 3966
rect 24774 4142 24832 4154
rect 24774 3966 24786 4142
rect 24820 3966 24832 4142
rect 24774 3954 24832 3966
rect 933 3203 991 3215
rect 933 3027 945 3203
rect 979 3027 991 3203
rect 933 3015 991 3027
rect 1051 3203 1109 3215
rect 1051 3027 1063 3203
rect 1097 3027 1109 3203
rect 1051 3015 1109 3027
rect 1169 3203 1227 3215
rect 1169 3027 1181 3203
rect 1215 3027 1227 3203
rect 1169 3015 1227 3027
rect 1287 3203 1345 3215
rect 1287 3027 1299 3203
rect 1333 3027 1345 3203
rect 1287 3015 1345 3027
rect 1405 3203 1463 3215
rect 1405 3027 1417 3203
rect 1451 3027 1463 3203
rect 1405 3015 1463 3027
rect 1523 3203 1581 3215
rect 1523 3027 1535 3203
rect 1569 3027 1581 3203
rect 1523 3015 1581 3027
rect 1641 3203 1699 3215
rect 1641 3027 1653 3203
rect 1687 3027 1699 3203
rect 1641 3015 1699 3027
rect 1759 3203 1817 3215
rect 1759 3027 1771 3203
rect 1805 3027 1817 3203
rect 1759 3015 1817 3027
rect 1877 3203 1935 3215
rect 1877 3027 1889 3203
rect 1923 3027 1935 3203
rect 1877 3015 1935 3027
rect 1995 3203 2053 3215
rect 1995 3027 2007 3203
rect 2041 3027 2053 3203
rect 7446 3200 7504 3212
rect 1995 3015 2053 3027
rect 7446 3024 7458 3200
rect 7492 3024 7504 3200
rect 7446 3012 7504 3024
rect 7564 3200 7622 3212
rect 7564 3024 7576 3200
rect 7610 3024 7622 3200
rect 7564 3012 7622 3024
rect 7682 3200 7740 3212
rect 7682 3024 7694 3200
rect 7728 3024 7740 3200
rect 7682 3012 7740 3024
rect 7800 3200 7858 3212
rect 7800 3024 7812 3200
rect 7846 3024 7858 3200
rect 7800 3012 7858 3024
rect 7918 3200 7976 3212
rect 7918 3024 7930 3200
rect 7964 3024 7976 3200
rect 7918 3012 7976 3024
rect 8036 3200 8094 3212
rect 8036 3024 8048 3200
rect 8082 3024 8094 3200
rect 8036 3012 8094 3024
rect 8154 3200 8212 3212
rect 8154 3024 8166 3200
rect 8200 3024 8212 3200
rect 8154 3012 8212 3024
rect 8272 3200 8330 3212
rect 8272 3024 8284 3200
rect 8318 3024 8330 3200
rect 8272 3012 8330 3024
rect 8390 3200 8448 3212
rect 8390 3024 8402 3200
rect 8436 3024 8448 3200
rect 8390 3012 8448 3024
rect 8508 3200 8566 3212
rect 8508 3024 8520 3200
rect 8554 3024 8566 3200
rect 13980 3195 14038 3207
rect 8508 3012 8566 3024
rect 13980 3019 13992 3195
rect 14026 3019 14038 3195
rect 2881 2786 2939 2798
rect 2397 2586 2455 2598
rect 2397 2410 2409 2586
rect 2443 2410 2455 2586
rect 2397 2398 2455 2410
rect 2515 2586 2573 2598
rect 2515 2410 2527 2586
rect 2561 2410 2573 2586
rect 2515 2398 2573 2410
rect 2633 2586 2691 2598
rect 2633 2410 2645 2586
rect 2679 2410 2691 2586
rect 2633 2398 2691 2410
rect 2751 2586 2809 2598
rect 2751 2410 2763 2586
rect 2797 2410 2809 2586
rect 2751 2398 2809 2410
rect 2881 2410 2893 2786
rect 2927 2410 2939 2786
rect 2881 2398 2939 2410
rect 2999 2786 3057 2798
rect 2999 2410 3011 2786
rect 3045 2410 3057 2786
rect 2999 2398 3057 2410
rect 3117 2786 3175 2798
rect 3117 2410 3129 2786
rect 3163 2410 3175 2786
rect 3117 2398 3175 2410
rect 3235 2786 3293 2798
rect 3235 2410 3247 2786
rect 3281 2410 3293 2786
rect 3235 2398 3293 2410
rect 3353 2786 3411 2798
rect 3353 2410 3365 2786
rect 3399 2410 3411 2786
rect 3353 2398 3411 2410
rect 3471 2786 3529 2798
rect 3471 2410 3483 2786
rect 3517 2410 3529 2786
rect 3471 2398 3529 2410
rect 3589 2786 3647 2798
rect 3589 2410 3601 2786
rect 3635 2410 3647 2786
rect 4779 2786 4837 2798
rect 3589 2398 3647 2410
rect 3718 2586 3776 2598
rect 3718 2410 3730 2586
rect 3764 2410 3776 2586
rect 3718 2398 3776 2410
rect 3836 2586 3894 2598
rect 3836 2410 3848 2586
rect 3882 2410 3894 2586
rect 3836 2398 3894 2410
rect 3954 2586 4012 2598
rect 3954 2410 3966 2586
rect 4000 2410 4012 2586
rect 3954 2398 4012 2410
rect 4072 2586 4130 2598
rect 4072 2410 4084 2586
rect 4118 2410 4130 2586
rect 4072 2398 4130 2410
rect 4295 2586 4353 2598
rect 4295 2410 4307 2586
rect 4341 2410 4353 2586
rect 4295 2398 4353 2410
rect 4413 2586 4471 2598
rect 4413 2410 4425 2586
rect 4459 2410 4471 2586
rect 4413 2398 4471 2410
rect 4531 2586 4589 2598
rect 4531 2410 4543 2586
rect 4577 2410 4589 2586
rect 4531 2398 4589 2410
rect 4649 2586 4707 2598
rect 4649 2410 4661 2586
rect 4695 2410 4707 2586
rect 4649 2398 4707 2410
rect 4779 2410 4791 2786
rect 4825 2410 4837 2786
rect 4779 2398 4837 2410
rect 4897 2786 4955 2798
rect 4897 2410 4909 2786
rect 4943 2410 4955 2786
rect 4897 2398 4955 2410
rect 5015 2786 5073 2798
rect 5015 2410 5027 2786
rect 5061 2410 5073 2786
rect 5015 2398 5073 2410
rect 5133 2786 5191 2798
rect 5133 2410 5145 2786
rect 5179 2410 5191 2786
rect 5133 2398 5191 2410
rect 5251 2786 5309 2798
rect 5251 2410 5263 2786
rect 5297 2410 5309 2786
rect 5251 2398 5309 2410
rect 5369 2786 5427 2798
rect 5369 2410 5381 2786
rect 5415 2410 5427 2786
rect 5369 2398 5427 2410
rect 5487 2786 5545 2798
rect 5487 2410 5499 2786
rect 5533 2410 5545 2786
rect 13980 3007 14038 3019
rect 14098 3195 14156 3207
rect 14098 3019 14110 3195
rect 14144 3019 14156 3195
rect 14098 3007 14156 3019
rect 14216 3195 14274 3207
rect 14216 3019 14228 3195
rect 14262 3019 14274 3195
rect 14216 3007 14274 3019
rect 14334 3195 14392 3207
rect 14334 3019 14346 3195
rect 14380 3019 14392 3195
rect 14334 3007 14392 3019
rect 14452 3195 14510 3207
rect 14452 3019 14464 3195
rect 14498 3019 14510 3195
rect 14452 3007 14510 3019
rect 14570 3195 14628 3207
rect 14570 3019 14582 3195
rect 14616 3019 14628 3195
rect 14570 3007 14628 3019
rect 14688 3195 14746 3207
rect 14688 3019 14700 3195
rect 14734 3019 14746 3195
rect 14688 3007 14746 3019
rect 14806 3195 14864 3207
rect 14806 3019 14818 3195
rect 14852 3019 14864 3195
rect 14806 3007 14864 3019
rect 14924 3195 14982 3207
rect 14924 3019 14936 3195
rect 14970 3019 14982 3195
rect 14924 3007 14982 3019
rect 15042 3195 15100 3207
rect 15042 3019 15054 3195
rect 15088 3019 15100 3195
rect 20538 3199 20596 3211
rect 15042 3007 15100 3019
rect 20538 3023 20550 3199
rect 20584 3023 20596 3199
rect 20538 3011 20596 3023
rect 20656 3199 20714 3211
rect 20656 3023 20668 3199
rect 20702 3023 20714 3199
rect 20656 3011 20714 3023
rect 20774 3199 20832 3211
rect 20774 3023 20786 3199
rect 20820 3023 20832 3199
rect 20774 3011 20832 3023
rect 20892 3199 20950 3211
rect 20892 3023 20904 3199
rect 20938 3023 20950 3199
rect 20892 3011 20950 3023
rect 21010 3199 21068 3211
rect 21010 3023 21022 3199
rect 21056 3023 21068 3199
rect 21010 3011 21068 3023
rect 21128 3199 21186 3211
rect 21128 3023 21140 3199
rect 21174 3023 21186 3199
rect 21128 3011 21186 3023
rect 21246 3199 21304 3211
rect 21246 3023 21258 3199
rect 21292 3023 21304 3199
rect 21246 3011 21304 3023
rect 21364 3199 21422 3211
rect 21364 3023 21376 3199
rect 21410 3023 21422 3199
rect 21364 3011 21422 3023
rect 21482 3199 21540 3211
rect 21482 3023 21494 3199
rect 21528 3023 21540 3199
rect 21482 3011 21540 3023
rect 21600 3199 21658 3211
rect 21600 3023 21612 3199
rect 21646 3023 21658 3199
rect 21600 3011 21658 3023
rect 9394 2783 9452 2795
rect 5487 2398 5545 2410
rect 5616 2586 5674 2598
rect 5616 2410 5628 2586
rect 5662 2410 5674 2586
rect 5616 2398 5674 2410
rect 5734 2586 5792 2598
rect 5734 2410 5746 2586
rect 5780 2410 5792 2586
rect 5734 2398 5792 2410
rect 5852 2586 5910 2598
rect 5852 2410 5864 2586
rect 5898 2410 5910 2586
rect 5852 2398 5910 2410
rect 5970 2586 6028 2598
rect 5970 2410 5982 2586
rect 6016 2410 6028 2586
rect 5970 2398 6028 2410
rect 928 1599 986 1611
rect 928 1423 940 1599
rect 974 1423 986 1599
rect 928 1411 986 1423
rect 1046 1599 1104 1611
rect 1046 1423 1058 1599
rect 1092 1423 1104 1599
rect 1046 1411 1104 1423
rect 1164 1599 1222 1611
rect 1164 1423 1176 1599
rect 1210 1423 1222 1599
rect 1164 1411 1222 1423
rect 1282 1599 1340 1611
rect 1282 1423 1294 1599
rect 1328 1423 1340 1599
rect 1282 1411 1340 1423
rect 1400 1599 1458 1611
rect 1400 1423 1412 1599
rect 1446 1423 1458 1599
rect 1400 1411 1458 1423
rect 1518 1599 1576 1611
rect 1518 1423 1530 1599
rect 1564 1423 1576 1599
rect 1518 1411 1576 1423
rect 1636 1599 1694 1611
rect 1636 1423 1648 1599
rect 1682 1423 1694 1599
rect 1636 1411 1694 1423
rect 1754 1599 1812 1611
rect 1754 1423 1766 1599
rect 1800 1423 1812 1599
rect 1754 1411 1812 1423
rect 1872 1599 1930 1611
rect 1872 1423 1884 1599
rect 1918 1423 1930 1599
rect 1872 1411 1930 1423
rect 1990 1599 2048 1611
rect 1990 1423 2002 1599
rect 2036 1423 2048 1599
rect 1990 1411 2048 1423
rect 2824 2093 2882 2105
rect 2824 1717 2836 2093
rect 2870 1717 2882 2093
rect 2824 1705 2882 1717
rect 2942 2093 3000 2105
rect 2942 1717 2954 2093
rect 2988 1717 3000 2093
rect 2942 1705 3000 1717
rect 3060 2093 3118 2105
rect 3060 1717 3072 2093
rect 3106 1717 3118 2093
rect 3060 1705 3118 1717
rect 3178 2093 3236 2105
rect 3178 1717 3190 2093
rect 3224 1717 3236 2093
rect 3178 1705 3236 1717
rect 3296 2093 3354 2105
rect 3296 1717 3308 2093
rect 3342 1717 3354 2093
rect 3296 1705 3354 1717
rect 3414 2093 3472 2105
rect 3414 1717 3426 2093
rect 3460 1717 3472 2093
rect 3414 1705 3472 1717
rect 3532 2093 3590 2105
rect 3532 1717 3544 2093
rect 3578 1717 3590 2093
rect 3532 1705 3590 1717
rect 8910 2583 8968 2595
rect 8910 2407 8922 2583
rect 8956 2407 8968 2583
rect 8910 2395 8968 2407
rect 9028 2583 9086 2595
rect 9028 2407 9040 2583
rect 9074 2407 9086 2583
rect 9028 2395 9086 2407
rect 9146 2583 9204 2595
rect 9146 2407 9158 2583
rect 9192 2407 9204 2583
rect 9146 2395 9204 2407
rect 9264 2583 9322 2595
rect 9264 2407 9276 2583
rect 9310 2407 9322 2583
rect 9264 2395 9322 2407
rect 9394 2407 9406 2783
rect 9440 2407 9452 2783
rect 9394 2395 9452 2407
rect 9512 2783 9570 2795
rect 9512 2407 9524 2783
rect 9558 2407 9570 2783
rect 9512 2395 9570 2407
rect 9630 2783 9688 2795
rect 9630 2407 9642 2783
rect 9676 2407 9688 2783
rect 9630 2395 9688 2407
rect 9748 2783 9806 2795
rect 9748 2407 9760 2783
rect 9794 2407 9806 2783
rect 9748 2395 9806 2407
rect 9866 2783 9924 2795
rect 9866 2407 9878 2783
rect 9912 2407 9924 2783
rect 9866 2395 9924 2407
rect 9984 2783 10042 2795
rect 9984 2407 9996 2783
rect 10030 2407 10042 2783
rect 9984 2395 10042 2407
rect 10102 2783 10160 2795
rect 10102 2407 10114 2783
rect 10148 2407 10160 2783
rect 11292 2783 11350 2795
rect 10102 2395 10160 2407
rect 10231 2583 10289 2595
rect 10231 2407 10243 2583
rect 10277 2407 10289 2583
rect 10231 2395 10289 2407
rect 10349 2583 10407 2595
rect 10349 2407 10361 2583
rect 10395 2407 10407 2583
rect 10349 2395 10407 2407
rect 10467 2583 10525 2595
rect 10467 2407 10479 2583
rect 10513 2407 10525 2583
rect 10467 2395 10525 2407
rect 10585 2583 10643 2595
rect 10585 2407 10597 2583
rect 10631 2407 10643 2583
rect 10585 2395 10643 2407
rect 10808 2583 10866 2595
rect 10808 2407 10820 2583
rect 10854 2407 10866 2583
rect 10808 2395 10866 2407
rect 10926 2583 10984 2595
rect 10926 2407 10938 2583
rect 10972 2407 10984 2583
rect 10926 2395 10984 2407
rect 11044 2583 11102 2595
rect 11044 2407 11056 2583
rect 11090 2407 11102 2583
rect 11044 2395 11102 2407
rect 11162 2583 11220 2595
rect 11162 2407 11174 2583
rect 11208 2407 11220 2583
rect 11162 2395 11220 2407
rect 11292 2407 11304 2783
rect 11338 2407 11350 2783
rect 11292 2395 11350 2407
rect 11410 2783 11468 2795
rect 11410 2407 11422 2783
rect 11456 2407 11468 2783
rect 11410 2395 11468 2407
rect 11528 2783 11586 2795
rect 11528 2407 11540 2783
rect 11574 2407 11586 2783
rect 11528 2395 11586 2407
rect 11646 2783 11704 2795
rect 11646 2407 11658 2783
rect 11692 2407 11704 2783
rect 11646 2395 11704 2407
rect 11764 2783 11822 2795
rect 11764 2407 11776 2783
rect 11810 2407 11822 2783
rect 11764 2395 11822 2407
rect 11882 2783 11940 2795
rect 11882 2407 11894 2783
rect 11928 2407 11940 2783
rect 11882 2395 11940 2407
rect 12000 2783 12058 2795
rect 12000 2407 12012 2783
rect 12046 2407 12058 2783
rect 15928 2778 15986 2790
rect 12000 2395 12058 2407
rect 12129 2583 12187 2595
rect 12129 2407 12141 2583
rect 12175 2407 12187 2583
rect 12129 2395 12187 2407
rect 12247 2583 12305 2595
rect 12247 2407 12259 2583
rect 12293 2407 12305 2583
rect 12247 2395 12305 2407
rect 12365 2583 12423 2595
rect 12365 2407 12377 2583
rect 12411 2407 12423 2583
rect 12365 2395 12423 2407
rect 12483 2583 12541 2595
rect 12483 2407 12495 2583
rect 12529 2407 12541 2583
rect 12483 2395 12541 2407
rect 4722 2093 4780 2105
rect 4722 1717 4734 2093
rect 4768 1717 4780 2093
rect 4722 1705 4780 1717
rect 4840 2093 4898 2105
rect 4840 1717 4852 2093
rect 4886 1717 4898 2093
rect 4840 1705 4898 1717
rect 4958 2093 5016 2105
rect 4958 1717 4970 2093
rect 5004 1717 5016 2093
rect 4958 1705 5016 1717
rect 5076 2093 5134 2105
rect 5076 1717 5088 2093
rect 5122 1717 5134 2093
rect 5076 1705 5134 1717
rect 5194 2093 5252 2105
rect 5194 1717 5206 2093
rect 5240 1717 5252 2093
rect 5194 1705 5252 1717
rect 5312 2093 5370 2105
rect 5312 1717 5324 2093
rect 5358 1717 5370 2093
rect 5312 1705 5370 1717
rect 5430 2093 5488 2105
rect 5430 1717 5442 2093
rect 5476 1717 5488 2093
rect 5430 1705 5488 1717
rect 7441 1596 7499 1608
rect 7441 1420 7453 1596
rect 7487 1420 7499 1596
rect 7441 1408 7499 1420
rect 7559 1596 7617 1608
rect 7559 1420 7571 1596
rect 7605 1420 7617 1596
rect 7559 1408 7617 1420
rect 7677 1596 7735 1608
rect 7677 1420 7689 1596
rect 7723 1420 7735 1596
rect 7677 1408 7735 1420
rect 7795 1596 7853 1608
rect 7795 1420 7807 1596
rect 7841 1420 7853 1596
rect 7795 1408 7853 1420
rect 7913 1596 7971 1608
rect 7913 1420 7925 1596
rect 7959 1420 7971 1596
rect 7913 1408 7971 1420
rect 8031 1596 8089 1608
rect 8031 1420 8043 1596
rect 8077 1420 8089 1596
rect 8031 1408 8089 1420
rect 8149 1596 8207 1608
rect 8149 1420 8161 1596
rect 8195 1420 8207 1596
rect 8149 1408 8207 1420
rect 8267 1596 8325 1608
rect 8267 1420 8279 1596
rect 8313 1420 8325 1596
rect 8267 1408 8325 1420
rect 8385 1596 8443 1608
rect 8385 1420 8397 1596
rect 8431 1420 8443 1596
rect 8385 1408 8443 1420
rect 8503 1596 8561 1608
rect 8503 1420 8515 1596
rect 8549 1420 8561 1596
rect 8503 1408 8561 1420
rect 9337 2090 9395 2102
rect 9337 1714 9349 2090
rect 9383 1714 9395 2090
rect 9337 1702 9395 1714
rect 9455 2090 9513 2102
rect 9455 1714 9467 2090
rect 9501 1714 9513 2090
rect 9455 1702 9513 1714
rect 9573 2090 9631 2102
rect 9573 1714 9585 2090
rect 9619 1714 9631 2090
rect 9573 1702 9631 1714
rect 9691 2090 9749 2102
rect 9691 1714 9703 2090
rect 9737 1714 9749 2090
rect 9691 1702 9749 1714
rect 9809 2090 9867 2102
rect 9809 1714 9821 2090
rect 9855 1714 9867 2090
rect 9809 1702 9867 1714
rect 9927 2090 9985 2102
rect 9927 1714 9939 2090
rect 9973 1714 9985 2090
rect 9927 1702 9985 1714
rect 10045 2090 10103 2102
rect 10045 1714 10057 2090
rect 10091 1714 10103 2090
rect 10045 1702 10103 1714
rect 15444 2578 15502 2590
rect 15444 2402 15456 2578
rect 15490 2402 15502 2578
rect 15444 2390 15502 2402
rect 15562 2578 15620 2590
rect 15562 2402 15574 2578
rect 15608 2402 15620 2578
rect 15562 2390 15620 2402
rect 15680 2578 15738 2590
rect 15680 2402 15692 2578
rect 15726 2402 15738 2578
rect 15680 2390 15738 2402
rect 15798 2578 15856 2590
rect 15798 2402 15810 2578
rect 15844 2402 15856 2578
rect 15798 2390 15856 2402
rect 15928 2402 15940 2778
rect 15974 2402 15986 2778
rect 15928 2390 15986 2402
rect 16046 2778 16104 2790
rect 16046 2402 16058 2778
rect 16092 2402 16104 2778
rect 16046 2390 16104 2402
rect 16164 2778 16222 2790
rect 16164 2402 16176 2778
rect 16210 2402 16222 2778
rect 16164 2390 16222 2402
rect 16282 2778 16340 2790
rect 16282 2402 16294 2778
rect 16328 2402 16340 2778
rect 16282 2390 16340 2402
rect 16400 2778 16458 2790
rect 16400 2402 16412 2778
rect 16446 2402 16458 2778
rect 16400 2390 16458 2402
rect 16518 2778 16576 2790
rect 16518 2402 16530 2778
rect 16564 2402 16576 2778
rect 16518 2390 16576 2402
rect 16636 2778 16694 2790
rect 16636 2402 16648 2778
rect 16682 2402 16694 2778
rect 17826 2778 17884 2790
rect 16636 2390 16694 2402
rect 16765 2578 16823 2590
rect 16765 2402 16777 2578
rect 16811 2402 16823 2578
rect 16765 2390 16823 2402
rect 16883 2578 16941 2590
rect 16883 2402 16895 2578
rect 16929 2402 16941 2578
rect 16883 2390 16941 2402
rect 17001 2578 17059 2590
rect 17001 2402 17013 2578
rect 17047 2402 17059 2578
rect 17001 2390 17059 2402
rect 17119 2578 17177 2590
rect 17119 2402 17131 2578
rect 17165 2402 17177 2578
rect 17119 2390 17177 2402
rect 17342 2578 17400 2590
rect 17342 2402 17354 2578
rect 17388 2402 17400 2578
rect 17342 2390 17400 2402
rect 17460 2578 17518 2590
rect 17460 2402 17472 2578
rect 17506 2402 17518 2578
rect 17460 2390 17518 2402
rect 17578 2578 17636 2590
rect 17578 2402 17590 2578
rect 17624 2402 17636 2578
rect 17578 2390 17636 2402
rect 17696 2578 17754 2590
rect 17696 2402 17708 2578
rect 17742 2402 17754 2578
rect 17696 2390 17754 2402
rect 17826 2402 17838 2778
rect 17872 2402 17884 2778
rect 17826 2390 17884 2402
rect 17944 2778 18002 2790
rect 17944 2402 17956 2778
rect 17990 2402 18002 2778
rect 17944 2390 18002 2402
rect 18062 2778 18120 2790
rect 18062 2402 18074 2778
rect 18108 2402 18120 2778
rect 18062 2390 18120 2402
rect 18180 2778 18238 2790
rect 18180 2402 18192 2778
rect 18226 2402 18238 2778
rect 18180 2390 18238 2402
rect 18298 2778 18356 2790
rect 18298 2402 18310 2778
rect 18344 2402 18356 2778
rect 18298 2390 18356 2402
rect 18416 2778 18474 2790
rect 18416 2402 18428 2778
rect 18462 2402 18474 2778
rect 18416 2390 18474 2402
rect 18534 2778 18592 2790
rect 18534 2402 18546 2778
rect 18580 2402 18592 2778
rect 22486 2782 22544 2794
rect 18534 2390 18592 2402
rect 18663 2578 18721 2590
rect 18663 2402 18675 2578
rect 18709 2402 18721 2578
rect 18663 2390 18721 2402
rect 18781 2578 18839 2590
rect 18781 2402 18793 2578
rect 18827 2402 18839 2578
rect 18781 2390 18839 2402
rect 18899 2578 18957 2590
rect 18899 2402 18911 2578
rect 18945 2402 18957 2578
rect 18899 2390 18957 2402
rect 19017 2578 19075 2590
rect 19017 2402 19029 2578
rect 19063 2402 19075 2578
rect 19017 2390 19075 2402
rect 11235 2090 11293 2102
rect 11235 1714 11247 2090
rect 11281 1714 11293 2090
rect 11235 1702 11293 1714
rect 11353 2090 11411 2102
rect 11353 1714 11365 2090
rect 11399 1714 11411 2090
rect 11353 1702 11411 1714
rect 11471 2090 11529 2102
rect 11471 1714 11483 2090
rect 11517 1714 11529 2090
rect 11471 1702 11529 1714
rect 11589 2090 11647 2102
rect 11589 1714 11601 2090
rect 11635 1714 11647 2090
rect 11589 1702 11647 1714
rect 11707 2090 11765 2102
rect 11707 1714 11719 2090
rect 11753 1714 11765 2090
rect 11707 1702 11765 1714
rect 11825 2090 11883 2102
rect 11825 1714 11837 2090
rect 11871 1714 11883 2090
rect 11825 1702 11883 1714
rect 11943 2090 12001 2102
rect 11943 1714 11955 2090
rect 11989 1714 12001 2090
rect 11943 1702 12001 1714
rect 13975 1591 14033 1603
rect 13975 1415 13987 1591
rect 14021 1415 14033 1591
rect 13975 1403 14033 1415
rect 14093 1591 14151 1603
rect 14093 1415 14105 1591
rect 14139 1415 14151 1591
rect 14093 1403 14151 1415
rect 14211 1591 14269 1603
rect 14211 1415 14223 1591
rect 14257 1415 14269 1591
rect 14211 1403 14269 1415
rect 14329 1591 14387 1603
rect 14329 1415 14341 1591
rect 14375 1415 14387 1591
rect 14329 1403 14387 1415
rect 14447 1591 14505 1603
rect 14447 1415 14459 1591
rect 14493 1415 14505 1591
rect 14447 1403 14505 1415
rect 14565 1591 14623 1603
rect 14565 1415 14577 1591
rect 14611 1415 14623 1591
rect 14565 1403 14623 1415
rect 14683 1591 14741 1603
rect 14683 1415 14695 1591
rect 14729 1415 14741 1591
rect 14683 1403 14741 1415
rect 14801 1591 14859 1603
rect 14801 1415 14813 1591
rect 14847 1415 14859 1591
rect 14801 1403 14859 1415
rect 14919 1591 14977 1603
rect 14919 1415 14931 1591
rect 14965 1415 14977 1591
rect 14919 1403 14977 1415
rect 15037 1591 15095 1603
rect 15037 1415 15049 1591
rect 15083 1415 15095 1591
rect 15037 1403 15095 1415
rect 15871 2085 15929 2097
rect 15871 1709 15883 2085
rect 15917 1709 15929 2085
rect 15871 1697 15929 1709
rect 15989 2085 16047 2097
rect 15989 1709 16001 2085
rect 16035 1709 16047 2085
rect 15989 1697 16047 1709
rect 16107 2085 16165 2097
rect 16107 1709 16119 2085
rect 16153 1709 16165 2085
rect 16107 1697 16165 1709
rect 16225 2085 16283 2097
rect 16225 1709 16237 2085
rect 16271 1709 16283 2085
rect 16225 1697 16283 1709
rect 16343 2085 16401 2097
rect 16343 1709 16355 2085
rect 16389 1709 16401 2085
rect 16343 1697 16401 1709
rect 16461 2085 16519 2097
rect 16461 1709 16473 2085
rect 16507 1709 16519 2085
rect 16461 1697 16519 1709
rect 16579 2085 16637 2097
rect 16579 1709 16591 2085
rect 16625 1709 16637 2085
rect 16579 1697 16637 1709
rect 22002 2582 22060 2594
rect 22002 2406 22014 2582
rect 22048 2406 22060 2582
rect 22002 2394 22060 2406
rect 22120 2582 22178 2594
rect 22120 2406 22132 2582
rect 22166 2406 22178 2582
rect 22120 2394 22178 2406
rect 22238 2582 22296 2594
rect 22238 2406 22250 2582
rect 22284 2406 22296 2582
rect 22238 2394 22296 2406
rect 22356 2582 22414 2594
rect 22356 2406 22368 2582
rect 22402 2406 22414 2582
rect 22356 2394 22414 2406
rect 22486 2406 22498 2782
rect 22532 2406 22544 2782
rect 22486 2394 22544 2406
rect 22604 2782 22662 2794
rect 22604 2406 22616 2782
rect 22650 2406 22662 2782
rect 22604 2394 22662 2406
rect 22722 2782 22780 2794
rect 22722 2406 22734 2782
rect 22768 2406 22780 2782
rect 22722 2394 22780 2406
rect 22840 2782 22898 2794
rect 22840 2406 22852 2782
rect 22886 2406 22898 2782
rect 22840 2394 22898 2406
rect 22958 2782 23016 2794
rect 22958 2406 22970 2782
rect 23004 2406 23016 2782
rect 22958 2394 23016 2406
rect 23076 2782 23134 2794
rect 23076 2406 23088 2782
rect 23122 2406 23134 2782
rect 23076 2394 23134 2406
rect 23194 2782 23252 2794
rect 23194 2406 23206 2782
rect 23240 2406 23252 2782
rect 24384 2782 24442 2794
rect 23194 2394 23252 2406
rect 23323 2582 23381 2594
rect 23323 2406 23335 2582
rect 23369 2406 23381 2582
rect 23323 2394 23381 2406
rect 23441 2582 23499 2594
rect 23441 2406 23453 2582
rect 23487 2406 23499 2582
rect 23441 2394 23499 2406
rect 23559 2582 23617 2594
rect 23559 2406 23571 2582
rect 23605 2406 23617 2582
rect 23559 2394 23617 2406
rect 23677 2582 23735 2594
rect 23677 2406 23689 2582
rect 23723 2406 23735 2582
rect 23677 2394 23735 2406
rect 23900 2582 23958 2594
rect 23900 2406 23912 2582
rect 23946 2406 23958 2582
rect 23900 2394 23958 2406
rect 24018 2582 24076 2594
rect 24018 2406 24030 2582
rect 24064 2406 24076 2582
rect 24018 2394 24076 2406
rect 24136 2582 24194 2594
rect 24136 2406 24148 2582
rect 24182 2406 24194 2582
rect 24136 2394 24194 2406
rect 24254 2582 24312 2594
rect 24254 2406 24266 2582
rect 24300 2406 24312 2582
rect 24254 2394 24312 2406
rect 24384 2406 24396 2782
rect 24430 2406 24442 2782
rect 24384 2394 24442 2406
rect 24502 2782 24560 2794
rect 24502 2406 24514 2782
rect 24548 2406 24560 2782
rect 24502 2394 24560 2406
rect 24620 2782 24678 2794
rect 24620 2406 24632 2782
rect 24666 2406 24678 2782
rect 24620 2394 24678 2406
rect 24738 2782 24796 2794
rect 24738 2406 24750 2782
rect 24784 2406 24796 2782
rect 24738 2394 24796 2406
rect 24856 2782 24914 2794
rect 24856 2406 24868 2782
rect 24902 2406 24914 2782
rect 24856 2394 24914 2406
rect 24974 2782 25032 2794
rect 24974 2406 24986 2782
rect 25020 2406 25032 2782
rect 24974 2394 25032 2406
rect 25092 2782 25150 2794
rect 25092 2406 25104 2782
rect 25138 2406 25150 2782
rect 25092 2394 25150 2406
rect 25221 2582 25279 2594
rect 25221 2406 25233 2582
rect 25267 2406 25279 2582
rect 25221 2394 25279 2406
rect 25339 2582 25397 2594
rect 25339 2406 25351 2582
rect 25385 2406 25397 2582
rect 25339 2394 25397 2406
rect 25457 2582 25515 2594
rect 25457 2406 25469 2582
rect 25503 2406 25515 2582
rect 25457 2394 25515 2406
rect 25575 2582 25633 2594
rect 25575 2406 25587 2582
rect 25621 2406 25633 2582
rect 25575 2394 25633 2406
rect 17769 2085 17827 2097
rect 17769 1709 17781 2085
rect 17815 1709 17827 2085
rect 17769 1697 17827 1709
rect 17887 2085 17945 2097
rect 17887 1709 17899 2085
rect 17933 1709 17945 2085
rect 17887 1697 17945 1709
rect 18005 2085 18063 2097
rect 18005 1709 18017 2085
rect 18051 1709 18063 2085
rect 18005 1697 18063 1709
rect 18123 2085 18181 2097
rect 18123 1709 18135 2085
rect 18169 1709 18181 2085
rect 18123 1697 18181 1709
rect 18241 2085 18299 2097
rect 18241 1709 18253 2085
rect 18287 1709 18299 2085
rect 18241 1697 18299 1709
rect 18359 2085 18417 2097
rect 18359 1709 18371 2085
rect 18405 1709 18417 2085
rect 18359 1697 18417 1709
rect 18477 2085 18535 2097
rect 18477 1709 18489 2085
rect 18523 1709 18535 2085
rect 18477 1697 18535 1709
rect 20533 1595 20591 1607
rect 20533 1419 20545 1595
rect 20579 1419 20591 1595
rect 20533 1407 20591 1419
rect 20651 1595 20709 1607
rect 20651 1419 20663 1595
rect 20697 1419 20709 1595
rect 20651 1407 20709 1419
rect 20769 1595 20827 1607
rect 20769 1419 20781 1595
rect 20815 1419 20827 1595
rect 20769 1407 20827 1419
rect 20887 1595 20945 1607
rect 20887 1419 20899 1595
rect 20933 1419 20945 1595
rect 20887 1407 20945 1419
rect 21005 1595 21063 1607
rect 21005 1419 21017 1595
rect 21051 1419 21063 1595
rect 21005 1407 21063 1419
rect 21123 1595 21181 1607
rect 21123 1419 21135 1595
rect 21169 1419 21181 1595
rect 21123 1407 21181 1419
rect 21241 1595 21299 1607
rect 21241 1419 21253 1595
rect 21287 1419 21299 1595
rect 21241 1407 21299 1419
rect 21359 1595 21417 1607
rect 21359 1419 21371 1595
rect 21405 1419 21417 1595
rect 21359 1407 21417 1419
rect 21477 1595 21535 1607
rect 21477 1419 21489 1595
rect 21523 1419 21535 1595
rect 21477 1407 21535 1419
rect 21595 1595 21653 1607
rect 21595 1419 21607 1595
rect 21641 1419 21653 1595
rect 21595 1407 21653 1419
rect 22429 2089 22487 2101
rect 22429 1713 22441 2089
rect 22475 1713 22487 2089
rect 22429 1701 22487 1713
rect 22547 2089 22605 2101
rect 22547 1713 22559 2089
rect 22593 1713 22605 2089
rect 22547 1701 22605 1713
rect 22665 2089 22723 2101
rect 22665 1713 22677 2089
rect 22711 1713 22723 2089
rect 22665 1701 22723 1713
rect 22783 2089 22841 2101
rect 22783 1713 22795 2089
rect 22829 1713 22841 2089
rect 22783 1701 22841 1713
rect 22901 2089 22959 2101
rect 22901 1713 22913 2089
rect 22947 1713 22959 2089
rect 22901 1701 22959 1713
rect 23019 2089 23077 2101
rect 23019 1713 23031 2089
rect 23065 1713 23077 2089
rect 23019 1701 23077 1713
rect 23137 2089 23195 2101
rect 23137 1713 23149 2089
rect 23183 1713 23195 2089
rect 23137 1701 23195 1713
rect 24327 2089 24385 2101
rect 24327 1713 24339 2089
rect 24373 1713 24385 2089
rect 24327 1701 24385 1713
rect 24445 2089 24503 2101
rect 24445 1713 24457 2089
rect 24491 1713 24503 2089
rect 24445 1701 24503 1713
rect 24563 2089 24621 2101
rect 24563 1713 24575 2089
rect 24609 1713 24621 2089
rect 24563 1701 24621 1713
rect 24681 2089 24739 2101
rect 24681 1713 24693 2089
rect 24727 1713 24739 2089
rect 24681 1701 24739 1713
rect 24799 2089 24857 2101
rect 24799 1713 24811 2089
rect 24845 1713 24857 2089
rect 24799 1701 24857 1713
rect 24917 2089 24975 2101
rect 24917 1713 24929 2089
rect 24963 1713 24975 2089
rect 24917 1701 24975 1713
rect 25035 2089 25093 2101
rect 25035 1713 25047 2089
rect 25081 1713 25093 2089
rect 25035 1701 25093 1713
rect 930 -679 988 -667
rect 930 -1055 942 -679
rect 976 -1055 988 -679
rect 930 -1067 988 -1055
rect 1048 -679 1106 -667
rect 1048 -1055 1060 -679
rect 1094 -1055 1106 -679
rect 1048 -1067 1106 -1055
rect 1166 -679 1224 -667
rect 1166 -1055 1178 -679
rect 1212 -1055 1224 -679
rect 1166 -1067 1224 -1055
rect 1284 -679 1342 -667
rect 1284 -1055 1296 -679
rect 1330 -1055 1342 -679
rect 1284 -1067 1342 -1055
rect 1402 -679 1460 -667
rect 1402 -1055 1414 -679
rect 1448 -1055 1460 -679
rect 1402 -1067 1460 -1055
rect 1520 -679 1578 -667
rect 1520 -1055 1532 -679
rect 1566 -1055 1578 -679
rect 1520 -1067 1578 -1055
rect 1638 -679 1696 -667
rect 1638 -1055 1650 -679
rect 1684 -1055 1696 -679
rect 1638 -1067 1696 -1055
rect 2072 -683 2130 -671
rect 2072 -1059 2084 -683
rect 2118 -1059 2130 -683
rect 2072 -1071 2130 -1059
rect 2190 -683 2248 -671
rect 2190 -1059 2202 -683
rect 2236 -1059 2248 -683
rect 2190 -1071 2248 -1059
rect 2308 -683 2366 -671
rect 2308 -1059 2320 -683
rect 2354 -1059 2366 -683
rect 2308 -1071 2366 -1059
rect 2426 -683 2484 -671
rect 2426 -1059 2438 -683
rect 2472 -1059 2484 -683
rect 2426 -1071 2484 -1059
rect 2544 -683 2602 -671
rect 2544 -1059 2556 -683
rect 2590 -1059 2602 -683
rect 2544 -1071 2602 -1059
rect 2662 -683 2720 -671
rect 2662 -1059 2674 -683
rect 2708 -1059 2720 -683
rect 2662 -1071 2720 -1059
rect 2780 -683 2838 -671
rect 2780 -1059 2792 -683
rect 2826 -1059 2838 -683
rect 7488 -683 7546 -671
rect 4043 -755 4101 -743
rect 4043 -931 4055 -755
rect 4089 -931 4101 -755
rect 4043 -943 4101 -931
rect 4161 -755 4219 -743
rect 4161 -931 4173 -755
rect 4207 -931 4219 -755
rect 4161 -943 4219 -931
rect 4279 -755 4337 -743
rect 4279 -931 4291 -755
rect 4325 -931 4337 -755
rect 4279 -943 4337 -931
rect 4397 -755 4455 -743
rect 4397 -931 4409 -755
rect 4443 -931 4455 -755
rect 4397 -943 4455 -931
rect 4515 -755 4573 -743
rect 4515 -931 4527 -755
rect 4561 -931 4573 -755
rect 4515 -943 4573 -931
rect 4633 -755 4691 -743
rect 4633 -931 4645 -755
rect 4679 -931 4691 -755
rect 4633 -943 4691 -931
rect 4751 -755 4809 -743
rect 4751 -931 4763 -755
rect 4797 -931 4809 -755
rect 4751 -943 4809 -931
rect 4869 -755 4927 -743
rect 4869 -931 4881 -755
rect 4915 -931 4927 -755
rect 4869 -943 4927 -931
rect 4987 -755 5045 -743
rect 4987 -931 4999 -755
rect 5033 -931 5045 -755
rect 4987 -943 5045 -931
rect 5105 -755 5163 -743
rect 5105 -931 5117 -755
rect 5151 -931 5163 -755
rect 5105 -943 5163 -931
rect 2780 -1071 2838 -1059
rect 7488 -1059 7500 -683
rect 7534 -1059 7546 -683
rect 7488 -1071 7546 -1059
rect 7606 -683 7664 -671
rect 7606 -1059 7618 -683
rect 7652 -1059 7664 -683
rect 7606 -1071 7664 -1059
rect 7724 -683 7782 -671
rect 7724 -1059 7736 -683
rect 7770 -1059 7782 -683
rect 7724 -1071 7782 -1059
rect 7842 -683 7900 -671
rect 7842 -1059 7854 -683
rect 7888 -1059 7900 -683
rect 7842 -1071 7900 -1059
rect 7960 -683 8018 -671
rect 7960 -1059 7972 -683
rect 8006 -1059 8018 -683
rect 7960 -1071 8018 -1059
rect 8078 -683 8136 -671
rect 8078 -1059 8090 -683
rect 8124 -1059 8136 -683
rect 8078 -1071 8136 -1059
rect 8196 -683 8254 -671
rect 8196 -1059 8208 -683
rect 8242 -1059 8254 -683
rect 8196 -1071 8254 -1059
rect 8630 -687 8688 -675
rect 8630 -1063 8642 -687
rect 8676 -1063 8688 -687
rect 855 -1462 913 -1450
rect 855 -1638 867 -1462
rect 901 -1638 913 -1462
rect 855 -1650 913 -1638
rect 973 -1462 1031 -1450
rect 973 -1638 985 -1462
rect 1019 -1638 1031 -1462
rect 973 -1650 1031 -1638
rect 1091 -1462 1149 -1450
rect 1091 -1638 1103 -1462
rect 1137 -1638 1149 -1462
rect 1091 -1650 1149 -1638
rect 1209 -1462 1267 -1450
rect 1209 -1638 1221 -1462
rect 1255 -1638 1267 -1462
rect 1209 -1650 1267 -1638
rect 1997 -1466 2055 -1454
rect 1997 -1642 2009 -1466
rect 2043 -1642 2055 -1466
rect 1997 -1654 2055 -1642
rect 2115 -1466 2173 -1454
rect 2115 -1642 2127 -1466
rect 2161 -1642 2173 -1466
rect 2115 -1654 2173 -1642
rect 2233 -1466 2291 -1454
rect 2233 -1642 2245 -1466
rect 2279 -1642 2291 -1466
rect 2233 -1654 2291 -1642
rect 2351 -1466 2409 -1454
rect 2351 -1642 2363 -1466
rect 2397 -1642 2409 -1466
rect 2351 -1654 2409 -1642
rect 8630 -1075 8688 -1063
rect 8748 -687 8806 -675
rect 8748 -1063 8760 -687
rect 8794 -1063 8806 -687
rect 8748 -1075 8806 -1063
rect 8866 -687 8924 -675
rect 8866 -1063 8878 -687
rect 8912 -1063 8924 -687
rect 8866 -1075 8924 -1063
rect 8984 -687 9042 -675
rect 8984 -1063 8996 -687
rect 9030 -1063 9042 -687
rect 8984 -1075 9042 -1063
rect 9102 -687 9160 -675
rect 9102 -1063 9114 -687
rect 9148 -1063 9160 -687
rect 9102 -1075 9160 -1063
rect 9220 -687 9278 -675
rect 9220 -1063 9232 -687
rect 9266 -1063 9278 -687
rect 9220 -1075 9278 -1063
rect 9338 -687 9396 -675
rect 14022 -678 14080 -666
rect 9338 -1063 9350 -687
rect 9384 -1063 9396 -687
rect 10601 -759 10659 -747
rect 10601 -935 10613 -759
rect 10647 -935 10659 -759
rect 10601 -947 10659 -935
rect 10719 -759 10777 -747
rect 10719 -935 10731 -759
rect 10765 -935 10777 -759
rect 10719 -947 10777 -935
rect 10837 -759 10895 -747
rect 10837 -935 10849 -759
rect 10883 -935 10895 -759
rect 10837 -947 10895 -935
rect 10955 -759 11013 -747
rect 10955 -935 10967 -759
rect 11001 -935 11013 -759
rect 10955 -947 11013 -935
rect 11073 -759 11131 -747
rect 11073 -935 11085 -759
rect 11119 -935 11131 -759
rect 11073 -947 11131 -935
rect 11191 -759 11249 -747
rect 11191 -935 11203 -759
rect 11237 -935 11249 -759
rect 11191 -947 11249 -935
rect 11309 -759 11367 -747
rect 11309 -935 11321 -759
rect 11355 -935 11367 -759
rect 11309 -947 11367 -935
rect 11427 -759 11485 -747
rect 11427 -935 11439 -759
rect 11473 -935 11485 -759
rect 11427 -947 11485 -935
rect 11545 -759 11603 -747
rect 11545 -935 11557 -759
rect 11591 -935 11603 -759
rect 11545 -947 11603 -935
rect 11663 -759 11721 -747
rect 11663 -935 11675 -759
rect 11709 -935 11721 -759
rect 11663 -947 11721 -935
rect 9338 -1075 9396 -1063
rect 14022 -1054 14034 -678
rect 14068 -1054 14080 -678
rect 14022 -1066 14080 -1054
rect 14140 -678 14198 -666
rect 14140 -1054 14152 -678
rect 14186 -1054 14198 -678
rect 14140 -1066 14198 -1054
rect 14258 -678 14316 -666
rect 14258 -1054 14270 -678
rect 14304 -1054 14316 -678
rect 14258 -1066 14316 -1054
rect 14376 -678 14434 -666
rect 14376 -1054 14388 -678
rect 14422 -1054 14434 -678
rect 14376 -1066 14434 -1054
rect 14494 -678 14552 -666
rect 14494 -1054 14506 -678
rect 14540 -1054 14552 -678
rect 14494 -1066 14552 -1054
rect 14612 -678 14670 -666
rect 14612 -1054 14624 -678
rect 14658 -1054 14670 -678
rect 14612 -1066 14670 -1054
rect 14730 -678 14788 -666
rect 14730 -1054 14742 -678
rect 14776 -1054 14788 -678
rect 14730 -1066 14788 -1054
rect 15164 -682 15222 -670
rect 15164 -1058 15176 -682
rect 15210 -1058 15222 -682
rect 7413 -1466 7471 -1454
rect 7413 -1642 7425 -1466
rect 7459 -1642 7471 -1466
rect 7413 -1654 7471 -1642
rect 7531 -1466 7589 -1454
rect 7531 -1642 7543 -1466
rect 7577 -1642 7589 -1466
rect 7531 -1654 7589 -1642
rect 7649 -1466 7707 -1454
rect 7649 -1642 7661 -1466
rect 7695 -1642 7707 -1466
rect 7649 -1654 7707 -1642
rect 7767 -1466 7825 -1454
rect 7767 -1642 7779 -1466
rect 7813 -1642 7825 -1466
rect 7767 -1654 7825 -1642
rect 8555 -1470 8613 -1458
rect 8555 -1646 8567 -1470
rect 8601 -1646 8613 -1470
rect 8555 -1658 8613 -1646
rect 8673 -1470 8731 -1458
rect 8673 -1646 8685 -1470
rect 8719 -1646 8731 -1470
rect 8673 -1658 8731 -1646
rect 8791 -1470 8849 -1458
rect 8791 -1646 8803 -1470
rect 8837 -1646 8849 -1470
rect 8791 -1658 8849 -1646
rect 8909 -1470 8967 -1458
rect 8909 -1646 8921 -1470
rect 8955 -1646 8967 -1470
rect 8909 -1658 8967 -1646
rect 15164 -1070 15222 -1058
rect 15282 -682 15340 -670
rect 15282 -1058 15294 -682
rect 15328 -1058 15340 -682
rect 15282 -1070 15340 -1058
rect 15400 -682 15458 -670
rect 15400 -1058 15412 -682
rect 15446 -1058 15458 -682
rect 15400 -1070 15458 -1058
rect 15518 -682 15576 -670
rect 15518 -1058 15530 -682
rect 15564 -1058 15576 -682
rect 15518 -1070 15576 -1058
rect 15636 -682 15694 -670
rect 15636 -1058 15648 -682
rect 15682 -1058 15694 -682
rect 15636 -1070 15694 -1058
rect 15754 -682 15812 -670
rect 15754 -1058 15766 -682
rect 15800 -1058 15812 -682
rect 15754 -1070 15812 -1058
rect 15872 -682 15930 -670
rect 15872 -1058 15884 -682
rect 15918 -1058 15930 -682
rect 20535 -675 20593 -663
rect 17135 -754 17193 -742
rect 17135 -930 17147 -754
rect 17181 -930 17193 -754
rect 17135 -942 17193 -930
rect 17253 -754 17311 -742
rect 17253 -930 17265 -754
rect 17299 -930 17311 -754
rect 17253 -942 17311 -930
rect 17371 -754 17429 -742
rect 17371 -930 17383 -754
rect 17417 -930 17429 -754
rect 17371 -942 17429 -930
rect 17489 -754 17547 -742
rect 17489 -930 17501 -754
rect 17535 -930 17547 -754
rect 17489 -942 17547 -930
rect 17607 -754 17665 -742
rect 17607 -930 17619 -754
rect 17653 -930 17665 -754
rect 17607 -942 17665 -930
rect 17725 -754 17783 -742
rect 17725 -930 17737 -754
rect 17771 -930 17783 -754
rect 17725 -942 17783 -930
rect 17843 -754 17901 -742
rect 17843 -930 17855 -754
rect 17889 -930 17901 -754
rect 17843 -942 17901 -930
rect 17961 -754 18019 -742
rect 17961 -930 17973 -754
rect 18007 -930 18019 -754
rect 17961 -942 18019 -930
rect 18079 -754 18137 -742
rect 18079 -930 18091 -754
rect 18125 -930 18137 -754
rect 18079 -942 18137 -930
rect 18197 -754 18255 -742
rect 18197 -930 18209 -754
rect 18243 -930 18255 -754
rect 18197 -942 18255 -930
rect 15872 -1070 15930 -1058
rect 20535 -1051 20547 -675
rect 20581 -1051 20593 -675
rect 20535 -1063 20593 -1051
rect 20653 -675 20711 -663
rect 20653 -1051 20665 -675
rect 20699 -1051 20711 -675
rect 20653 -1063 20711 -1051
rect 20771 -675 20829 -663
rect 20771 -1051 20783 -675
rect 20817 -1051 20829 -675
rect 20771 -1063 20829 -1051
rect 20889 -675 20947 -663
rect 20889 -1051 20901 -675
rect 20935 -1051 20947 -675
rect 20889 -1063 20947 -1051
rect 21007 -675 21065 -663
rect 21007 -1051 21019 -675
rect 21053 -1051 21065 -675
rect 21007 -1063 21065 -1051
rect 21125 -675 21183 -663
rect 21125 -1051 21137 -675
rect 21171 -1051 21183 -675
rect 21125 -1063 21183 -1051
rect 21243 -675 21301 -663
rect 21243 -1051 21255 -675
rect 21289 -1051 21301 -675
rect 21243 -1063 21301 -1051
rect 21677 -679 21735 -667
rect 21677 -1055 21689 -679
rect 21723 -1055 21735 -679
rect 13947 -1461 14005 -1449
rect 13947 -1637 13959 -1461
rect 13993 -1637 14005 -1461
rect 13947 -1649 14005 -1637
rect 14065 -1461 14123 -1449
rect 14065 -1637 14077 -1461
rect 14111 -1637 14123 -1461
rect 14065 -1649 14123 -1637
rect 14183 -1461 14241 -1449
rect 14183 -1637 14195 -1461
rect 14229 -1637 14241 -1461
rect 14183 -1649 14241 -1637
rect 14301 -1461 14359 -1449
rect 14301 -1637 14313 -1461
rect 14347 -1637 14359 -1461
rect 14301 -1649 14359 -1637
rect 15089 -1465 15147 -1453
rect 15089 -1641 15101 -1465
rect 15135 -1641 15147 -1465
rect 15089 -1653 15147 -1641
rect 15207 -1465 15265 -1453
rect 15207 -1641 15219 -1465
rect 15253 -1641 15265 -1465
rect 15207 -1653 15265 -1641
rect 15325 -1465 15383 -1453
rect 15325 -1641 15337 -1465
rect 15371 -1641 15383 -1465
rect 15325 -1653 15383 -1641
rect 15443 -1465 15501 -1453
rect 15443 -1641 15455 -1465
rect 15489 -1641 15501 -1465
rect 15443 -1653 15501 -1641
rect 21677 -1067 21735 -1055
rect 21795 -679 21853 -667
rect 21795 -1055 21807 -679
rect 21841 -1055 21853 -679
rect 21795 -1067 21853 -1055
rect 21913 -679 21971 -667
rect 21913 -1055 21925 -679
rect 21959 -1055 21971 -679
rect 21913 -1067 21971 -1055
rect 22031 -679 22089 -667
rect 22031 -1055 22043 -679
rect 22077 -1055 22089 -679
rect 22031 -1067 22089 -1055
rect 22149 -679 22207 -667
rect 22149 -1055 22161 -679
rect 22195 -1055 22207 -679
rect 22149 -1067 22207 -1055
rect 22267 -679 22325 -667
rect 22267 -1055 22279 -679
rect 22313 -1055 22325 -679
rect 22267 -1067 22325 -1055
rect 22385 -679 22443 -667
rect 22385 -1055 22397 -679
rect 22431 -1055 22443 -679
rect 23648 -751 23706 -739
rect 23648 -927 23660 -751
rect 23694 -927 23706 -751
rect 23648 -939 23706 -927
rect 23766 -751 23824 -739
rect 23766 -927 23778 -751
rect 23812 -927 23824 -751
rect 23766 -939 23824 -927
rect 23884 -751 23942 -739
rect 23884 -927 23896 -751
rect 23930 -927 23942 -751
rect 23884 -939 23942 -927
rect 24002 -751 24060 -739
rect 24002 -927 24014 -751
rect 24048 -927 24060 -751
rect 24002 -939 24060 -927
rect 24120 -751 24178 -739
rect 24120 -927 24132 -751
rect 24166 -927 24178 -751
rect 24120 -939 24178 -927
rect 24238 -751 24296 -739
rect 24238 -927 24250 -751
rect 24284 -927 24296 -751
rect 24238 -939 24296 -927
rect 24356 -751 24414 -739
rect 24356 -927 24368 -751
rect 24402 -927 24414 -751
rect 24356 -939 24414 -927
rect 24474 -751 24532 -739
rect 24474 -927 24486 -751
rect 24520 -927 24532 -751
rect 24474 -939 24532 -927
rect 24592 -751 24650 -739
rect 24592 -927 24604 -751
rect 24638 -927 24650 -751
rect 24592 -939 24650 -927
rect 24710 -751 24768 -739
rect 24710 -927 24722 -751
rect 24756 -927 24768 -751
rect 24710 -939 24768 -927
rect 22385 -1067 22443 -1055
rect 20460 -1458 20518 -1446
rect 20460 -1634 20472 -1458
rect 20506 -1634 20518 -1458
rect 20460 -1646 20518 -1634
rect 20578 -1458 20636 -1446
rect 20578 -1634 20590 -1458
rect 20624 -1634 20636 -1458
rect 20578 -1646 20636 -1634
rect 20696 -1458 20754 -1446
rect 20696 -1634 20708 -1458
rect 20742 -1634 20754 -1458
rect 20696 -1646 20754 -1634
rect 20814 -1458 20872 -1446
rect 20814 -1634 20826 -1458
rect 20860 -1634 20872 -1458
rect 20814 -1646 20872 -1634
rect 21602 -1462 21660 -1450
rect 21602 -1638 21614 -1462
rect 21648 -1638 21660 -1462
rect 21602 -1650 21660 -1638
rect 21720 -1462 21778 -1450
rect 21720 -1638 21732 -1462
rect 21766 -1638 21778 -1462
rect 21720 -1650 21778 -1638
rect 21838 -1462 21896 -1450
rect 21838 -1638 21850 -1462
rect 21884 -1638 21896 -1462
rect 21838 -1650 21896 -1638
rect 21956 -1462 22014 -1450
rect 21956 -1638 21968 -1462
rect 22002 -1638 22014 -1462
rect 21956 -1650 22014 -1638
rect 4029 -2405 4087 -2393
rect 4029 -2581 4041 -2405
rect 4075 -2581 4087 -2405
rect 4029 -2593 4087 -2581
rect 4147 -2405 4205 -2393
rect 4147 -2581 4159 -2405
rect 4193 -2581 4205 -2405
rect 4147 -2593 4205 -2581
rect 4265 -2405 4323 -2393
rect 4265 -2581 4277 -2405
rect 4311 -2581 4323 -2405
rect 4265 -2593 4323 -2581
rect 4383 -2405 4441 -2393
rect 4383 -2581 4395 -2405
rect 4429 -2581 4441 -2405
rect 4383 -2593 4441 -2581
rect 4501 -2405 4559 -2393
rect 4501 -2581 4513 -2405
rect 4547 -2581 4559 -2405
rect 4501 -2593 4559 -2581
rect 4619 -2405 4677 -2393
rect 4619 -2581 4631 -2405
rect 4665 -2581 4677 -2405
rect 4619 -2593 4677 -2581
rect 4737 -2405 4795 -2393
rect 4737 -2581 4749 -2405
rect 4783 -2581 4795 -2405
rect 4737 -2593 4795 -2581
rect 4855 -2405 4913 -2393
rect 4855 -2581 4867 -2405
rect 4901 -2581 4913 -2405
rect 4855 -2593 4913 -2581
rect 4973 -2405 5031 -2393
rect 4973 -2581 4985 -2405
rect 5019 -2581 5031 -2405
rect 4973 -2593 5031 -2581
rect 5091 -2405 5149 -2393
rect 5091 -2581 5103 -2405
rect 5137 -2581 5149 -2405
rect 10587 -2409 10645 -2397
rect 5091 -2593 5149 -2581
rect 10587 -2585 10599 -2409
rect 10633 -2585 10645 -2409
rect 10587 -2597 10645 -2585
rect 10705 -2409 10763 -2397
rect 10705 -2585 10717 -2409
rect 10751 -2585 10763 -2409
rect 10705 -2597 10763 -2585
rect 10823 -2409 10881 -2397
rect 10823 -2585 10835 -2409
rect 10869 -2585 10881 -2409
rect 10823 -2597 10881 -2585
rect 10941 -2409 10999 -2397
rect 10941 -2585 10953 -2409
rect 10987 -2585 10999 -2409
rect 10941 -2597 10999 -2585
rect 11059 -2409 11117 -2397
rect 11059 -2585 11071 -2409
rect 11105 -2585 11117 -2409
rect 11059 -2597 11117 -2585
rect 11177 -2409 11235 -2397
rect 11177 -2585 11189 -2409
rect 11223 -2585 11235 -2409
rect 11177 -2597 11235 -2585
rect 11295 -2409 11353 -2397
rect 11295 -2585 11307 -2409
rect 11341 -2585 11353 -2409
rect 11295 -2597 11353 -2585
rect 11413 -2409 11471 -2397
rect 11413 -2585 11425 -2409
rect 11459 -2585 11471 -2409
rect 11413 -2597 11471 -2585
rect 11531 -2409 11589 -2397
rect 11531 -2585 11543 -2409
rect 11577 -2585 11589 -2409
rect 11531 -2597 11589 -2585
rect 11649 -2409 11707 -2397
rect 11649 -2585 11661 -2409
rect 11695 -2585 11707 -2409
rect 17121 -2404 17179 -2392
rect 11649 -2597 11707 -2585
rect 17121 -2580 17133 -2404
rect 17167 -2580 17179 -2404
rect 17121 -2592 17179 -2580
rect 17239 -2404 17297 -2392
rect 17239 -2580 17251 -2404
rect 17285 -2580 17297 -2404
rect 17239 -2592 17297 -2580
rect 17357 -2404 17415 -2392
rect 17357 -2580 17369 -2404
rect 17403 -2580 17415 -2404
rect 17357 -2592 17415 -2580
rect 17475 -2404 17533 -2392
rect 17475 -2580 17487 -2404
rect 17521 -2580 17533 -2404
rect 17475 -2592 17533 -2580
rect 17593 -2404 17651 -2392
rect 17593 -2580 17605 -2404
rect 17639 -2580 17651 -2404
rect 17593 -2592 17651 -2580
rect 17711 -2404 17769 -2392
rect 17711 -2580 17723 -2404
rect 17757 -2580 17769 -2404
rect 17711 -2592 17769 -2580
rect 17829 -2404 17887 -2392
rect 17829 -2580 17841 -2404
rect 17875 -2580 17887 -2404
rect 17829 -2592 17887 -2580
rect 17947 -2404 18005 -2392
rect 17947 -2580 17959 -2404
rect 17993 -2580 18005 -2404
rect 17947 -2592 18005 -2580
rect 18065 -2404 18123 -2392
rect 18065 -2580 18077 -2404
rect 18111 -2580 18123 -2404
rect 18065 -2592 18123 -2580
rect 18183 -2404 18241 -2392
rect 18183 -2580 18195 -2404
rect 18229 -2580 18241 -2404
rect 23634 -2401 23692 -2389
rect 18183 -2592 18241 -2580
rect 23634 -2577 23646 -2401
rect 23680 -2577 23692 -2401
rect 23634 -2589 23692 -2577
rect 23752 -2401 23810 -2389
rect 23752 -2577 23764 -2401
rect 23798 -2577 23810 -2401
rect 23752 -2589 23810 -2577
rect 23870 -2401 23928 -2389
rect 23870 -2577 23882 -2401
rect 23916 -2577 23928 -2401
rect 23870 -2589 23928 -2577
rect 23988 -2401 24046 -2389
rect 23988 -2577 24000 -2401
rect 24034 -2577 24046 -2401
rect 23988 -2589 24046 -2577
rect 24106 -2401 24164 -2389
rect 24106 -2577 24118 -2401
rect 24152 -2577 24164 -2401
rect 24106 -2589 24164 -2577
rect 24224 -2401 24282 -2389
rect 24224 -2577 24236 -2401
rect 24270 -2577 24282 -2401
rect 24224 -2589 24282 -2577
rect 24342 -2401 24400 -2389
rect 24342 -2577 24354 -2401
rect 24388 -2577 24400 -2401
rect 24342 -2589 24400 -2577
rect 24460 -2401 24518 -2389
rect 24460 -2577 24472 -2401
rect 24506 -2577 24518 -2401
rect 24460 -2589 24518 -2577
rect 24578 -2401 24636 -2389
rect 24578 -2577 24590 -2401
rect 24624 -2577 24636 -2401
rect 24578 -2589 24636 -2577
rect 24696 -2401 24754 -2389
rect 24696 -2577 24708 -2401
rect 24742 -2577 24754 -2401
rect 24696 -2589 24754 -2577
rect 537 -2822 595 -2810
rect 54 -3022 112 -3010
rect 54 -3198 66 -3022
rect 100 -3198 112 -3022
rect 54 -3210 112 -3198
rect 172 -3022 230 -3010
rect 172 -3198 184 -3022
rect 218 -3198 230 -3022
rect 172 -3210 230 -3198
rect 290 -3022 348 -3010
rect 290 -3198 302 -3022
rect 336 -3198 348 -3022
rect 290 -3210 348 -3198
rect 408 -3022 466 -3010
rect 408 -3198 420 -3022
rect 454 -3198 466 -3022
rect 408 -3210 466 -3198
rect 537 -3198 549 -2822
rect 583 -3198 595 -2822
rect 537 -3210 595 -3198
rect 655 -2822 713 -2810
rect 655 -3198 667 -2822
rect 701 -3198 713 -2822
rect 655 -3210 713 -3198
rect 773 -2822 831 -2810
rect 773 -3198 785 -2822
rect 819 -3198 831 -2822
rect 773 -3210 831 -3198
rect 891 -2822 949 -2810
rect 891 -3198 903 -2822
rect 937 -3198 949 -2822
rect 891 -3210 949 -3198
rect 1009 -2822 1067 -2810
rect 1009 -3198 1021 -2822
rect 1055 -3198 1067 -2822
rect 1009 -3210 1067 -3198
rect 1127 -2822 1185 -2810
rect 1127 -3198 1139 -2822
rect 1173 -3198 1185 -2822
rect 1127 -3210 1185 -3198
rect 1245 -2822 1303 -2810
rect 1245 -3198 1257 -2822
rect 1291 -3198 1303 -2822
rect 2435 -2822 2493 -2810
rect 1245 -3210 1303 -3198
rect 1375 -3022 1433 -3010
rect 1375 -3198 1387 -3022
rect 1421 -3198 1433 -3022
rect 1375 -3210 1433 -3198
rect 1493 -3022 1551 -3010
rect 1493 -3198 1505 -3022
rect 1539 -3198 1551 -3022
rect 1493 -3210 1551 -3198
rect 1611 -3022 1669 -3010
rect 1611 -3198 1623 -3022
rect 1657 -3198 1669 -3022
rect 1611 -3210 1669 -3198
rect 1729 -3022 1787 -3010
rect 1729 -3198 1741 -3022
rect 1775 -3198 1787 -3022
rect 1729 -3210 1787 -3198
rect 1952 -3022 2010 -3010
rect 1952 -3198 1964 -3022
rect 1998 -3198 2010 -3022
rect 1952 -3210 2010 -3198
rect 2070 -3022 2128 -3010
rect 2070 -3198 2082 -3022
rect 2116 -3198 2128 -3022
rect 2070 -3210 2128 -3198
rect 2188 -3022 2246 -3010
rect 2188 -3198 2200 -3022
rect 2234 -3198 2246 -3022
rect 2188 -3210 2246 -3198
rect 2306 -3022 2364 -3010
rect 2306 -3198 2318 -3022
rect 2352 -3198 2364 -3022
rect 2306 -3210 2364 -3198
rect 2435 -3198 2447 -2822
rect 2481 -3198 2493 -2822
rect 2435 -3210 2493 -3198
rect 2553 -2822 2611 -2810
rect 2553 -3198 2565 -2822
rect 2599 -3198 2611 -2822
rect 2553 -3210 2611 -3198
rect 2671 -2822 2729 -2810
rect 2671 -3198 2683 -2822
rect 2717 -3198 2729 -2822
rect 2671 -3210 2729 -3198
rect 2789 -2822 2847 -2810
rect 2789 -3198 2801 -2822
rect 2835 -3198 2847 -2822
rect 2789 -3210 2847 -3198
rect 2907 -2822 2965 -2810
rect 2907 -3198 2919 -2822
rect 2953 -3198 2965 -2822
rect 2907 -3210 2965 -3198
rect 3025 -2822 3083 -2810
rect 3025 -3198 3037 -2822
rect 3071 -3198 3083 -2822
rect 3025 -3210 3083 -3198
rect 3143 -2822 3201 -2810
rect 3143 -3198 3155 -2822
rect 3189 -3198 3201 -2822
rect 7095 -2826 7153 -2814
rect 3143 -3210 3201 -3198
rect 3273 -3022 3331 -3010
rect 3273 -3198 3285 -3022
rect 3319 -3198 3331 -3022
rect 3273 -3210 3331 -3198
rect 3391 -3022 3449 -3010
rect 3391 -3198 3403 -3022
rect 3437 -3198 3449 -3022
rect 3391 -3210 3449 -3198
rect 3509 -3022 3567 -3010
rect 3509 -3198 3521 -3022
rect 3555 -3198 3567 -3022
rect 3509 -3210 3567 -3198
rect 3627 -3022 3685 -3010
rect 3627 -3198 3639 -3022
rect 3673 -3198 3685 -3022
rect 3627 -3210 3685 -3198
rect 594 -3515 652 -3503
rect 594 -3891 606 -3515
rect 640 -3891 652 -3515
rect 594 -3903 652 -3891
rect 712 -3515 770 -3503
rect 712 -3891 724 -3515
rect 758 -3891 770 -3515
rect 712 -3903 770 -3891
rect 830 -3515 888 -3503
rect 830 -3891 842 -3515
rect 876 -3891 888 -3515
rect 830 -3903 888 -3891
rect 948 -3515 1006 -3503
rect 948 -3891 960 -3515
rect 994 -3891 1006 -3515
rect 948 -3903 1006 -3891
rect 1066 -3515 1124 -3503
rect 1066 -3891 1078 -3515
rect 1112 -3891 1124 -3515
rect 1066 -3903 1124 -3891
rect 1184 -3515 1242 -3503
rect 1184 -3891 1196 -3515
rect 1230 -3891 1242 -3515
rect 1184 -3903 1242 -3891
rect 1302 -3515 1360 -3503
rect 1302 -3891 1314 -3515
rect 1348 -3891 1360 -3515
rect 1302 -3903 1360 -3891
rect 6612 -3026 6670 -3014
rect 6612 -3202 6624 -3026
rect 6658 -3202 6670 -3026
rect 6612 -3214 6670 -3202
rect 6730 -3026 6788 -3014
rect 6730 -3202 6742 -3026
rect 6776 -3202 6788 -3026
rect 6730 -3214 6788 -3202
rect 6848 -3026 6906 -3014
rect 6848 -3202 6860 -3026
rect 6894 -3202 6906 -3026
rect 6848 -3214 6906 -3202
rect 6966 -3026 7024 -3014
rect 6966 -3202 6978 -3026
rect 7012 -3202 7024 -3026
rect 6966 -3214 7024 -3202
rect 7095 -3202 7107 -2826
rect 7141 -3202 7153 -2826
rect 7095 -3214 7153 -3202
rect 7213 -2826 7271 -2814
rect 7213 -3202 7225 -2826
rect 7259 -3202 7271 -2826
rect 7213 -3214 7271 -3202
rect 7331 -2826 7389 -2814
rect 7331 -3202 7343 -2826
rect 7377 -3202 7389 -2826
rect 7331 -3214 7389 -3202
rect 7449 -2826 7507 -2814
rect 7449 -3202 7461 -2826
rect 7495 -3202 7507 -2826
rect 7449 -3214 7507 -3202
rect 7567 -2826 7625 -2814
rect 7567 -3202 7579 -2826
rect 7613 -3202 7625 -2826
rect 7567 -3214 7625 -3202
rect 7685 -2826 7743 -2814
rect 7685 -3202 7697 -2826
rect 7731 -3202 7743 -2826
rect 7685 -3214 7743 -3202
rect 7803 -2826 7861 -2814
rect 7803 -3202 7815 -2826
rect 7849 -3202 7861 -2826
rect 8993 -2826 9051 -2814
rect 7803 -3214 7861 -3202
rect 7933 -3026 7991 -3014
rect 7933 -3202 7945 -3026
rect 7979 -3202 7991 -3026
rect 7933 -3214 7991 -3202
rect 8051 -3026 8109 -3014
rect 8051 -3202 8063 -3026
rect 8097 -3202 8109 -3026
rect 8051 -3214 8109 -3202
rect 8169 -3026 8227 -3014
rect 8169 -3202 8181 -3026
rect 8215 -3202 8227 -3026
rect 8169 -3214 8227 -3202
rect 8287 -3026 8345 -3014
rect 8287 -3202 8299 -3026
rect 8333 -3202 8345 -3026
rect 8287 -3214 8345 -3202
rect 8510 -3026 8568 -3014
rect 8510 -3202 8522 -3026
rect 8556 -3202 8568 -3026
rect 8510 -3214 8568 -3202
rect 8628 -3026 8686 -3014
rect 8628 -3202 8640 -3026
rect 8674 -3202 8686 -3026
rect 8628 -3214 8686 -3202
rect 8746 -3026 8804 -3014
rect 8746 -3202 8758 -3026
rect 8792 -3202 8804 -3026
rect 8746 -3214 8804 -3202
rect 8864 -3026 8922 -3014
rect 8864 -3202 8876 -3026
rect 8910 -3202 8922 -3026
rect 8864 -3214 8922 -3202
rect 8993 -3202 9005 -2826
rect 9039 -3202 9051 -2826
rect 8993 -3214 9051 -3202
rect 9111 -2826 9169 -2814
rect 9111 -3202 9123 -2826
rect 9157 -3202 9169 -2826
rect 9111 -3214 9169 -3202
rect 9229 -2826 9287 -2814
rect 9229 -3202 9241 -2826
rect 9275 -3202 9287 -2826
rect 9229 -3214 9287 -3202
rect 9347 -2826 9405 -2814
rect 9347 -3202 9359 -2826
rect 9393 -3202 9405 -2826
rect 9347 -3214 9405 -3202
rect 9465 -2826 9523 -2814
rect 9465 -3202 9477 -2826
rect 9511 -3202 9523 -2826
rect 9465 -3214 9523 -3202
rect 9583 -2826 9641 -2814
rect 9583 -3202 9595 -2826
rect 9629 -3202 9641 -2826
rect 9583 -3214 9641 -3202
rect 9701 -2826 9759 -2814
rect 9701 -3202 9713 -2826
rect 9747 -3202 9759 -2826
rect 13629 -2821 13687 -2809
rect 9701 -3214 9759 -3202
rect 9831 -3026 9889 -3014
rect 9831 -3202 9843 -3026
rect 9877 -3202 9889 -3026
rect 9831 -3214 9889 -3202
rect 9949 -3026 10007 -3014
rect 9949 -3202 9961 -3026
rect 9995 -3202 10007 -3026
rect 9949 -3214 10007 -3202
rect 10067 -3026 10125 -3014
rect 10067 -3202 10079 -3026
rect 10113 -3202 10125 -3026
rect 10067 -3214 10125 -3202
rect 10185 -3026 10243 -3014
rect 10185 -3202 10197 -3026
rect 10231 -3202 10243 -3026
rect 10185 -3214 10243 -3202
rect 2492 -3515 2550 -3503
rect 2492 -3891 2504 -3515
rect 2538 -3891 2550 -3515
rect 2492 -3903 2550 -3891
rect 2610 -3515 2668 -3503
rect 2610 -3891 2622 -3515
rect 2656 -3891 2668 -3515
rect 2610 -3903 2668 -3891
rect 2728 -3515 2786 -3503
rect 2728 -3891 2740 -3515
rect 2774 -3891 2786 -3515
rect 2728 -3903 2786 -3891
rect 2846 -3515 2904 -3503
rect 2846 -3891 2858 -3515
rect 2892 -3891 2904 -3515
rect 2846 -3903 2904 -3891
rect 2964 -3515 3022 -3503
rect 2964 -3891 2976 -3515
rect 3010 -3891 3022 -3515
rect 2964 -3903 3022 -3891
rect 3082 -3515 3140 -3503
rect 3082 -3891 3094 -3515
rect 3128 -3891 3140 -3515
rect 3082 -3903 3140 -3891
rect 3200 -3515 3258 -3503
rect 3200 -3891 3212 -3515
rect 3246 -3891 3258 -3515
rect 3200 -3903 3258 -3891
rect 4034 -4009 4092 -3997
rect 4034 -4185 4046 -4009
rect 4080 -4185 4092 -4009
rect 4034 -4197 4092 -4185
rect 4152 -4009 4210 -3997
rect 4152 -4185 4164 -4009
rect 4198 -4185 4210 -4009
rect 4152 -4197 4210 -4185
rect 4270 -4009 4328 -3997
rect 4270 -4185 4282 -4009
rect 4316 -4185 4328 -4009
rect 4270 -4197 4328 -4185
rect 4388 -4009 4446 -3997
rect 4388 -4185 4400 -4009
rect 4434 -4185 4446 -4009
rect 4388 -4197 4446 -4185
rect 4506 -4009 4564 -3997
rect 4506 -4185 4518 -4009
rect 4552 -4185 4564 -4009
rect 4506 -4197 4564 -4185
rect 4624 -4009 4682 -3997
rect 4624 -4185 4636 -4009
rect 4670 -4185 4682 -4009
rect 4624 -4197 4682 -4185
rect 4742 -4009 4800 -3997
rect 4742 -4185 4754 -4009
rect 4788 -4185 4800 -4009
rect 4742 -4197 4800 -4185
rect 4860 -4009 4918 -3997
rect 4860 -4185 4872 -4009
rect 4906 -4185 4918 -4009
rect 4860 -4197 4918 -4185
rect 4978 -4009 5036 -3997
rect 4978 -4185 4990 -4009
rect 5024 -4185 5036 -4009
rect 4978 -4197 5036 -4185
rect 5096 -4009 5154 -3997
rect 5096 -4185 5108 -4009
rect 5142 -4185 5154 -4009
rect 5096 -4197 5154 -4185
rect 7152 -3519 7210 -3507
rect 7152 -3895 7164 -3519
rect 7198 -3895 7210 -3519
rect 7152 -3907 7210 -3895
rect 7270 -3519 7328 -3507
rect 7270 -3895 7282 -3519
rect 7316 -3895 7328 -3519
rect 7270 -3907 7328 -3895
rect 7388 -3519 7446 -3507
rect 7388 -3895 7400 -3519
rect 7434 -3895 7446 -3519
rect 7388 -3907 7446 -3895
rect 7506 -3519 7564 -3507
rect 7506 -3895 7518 -3519
rect 7552 -3895 7564 -3519
rect 7506 -3907 7564 -3895
rect 7624 -3519 7682 -3507
rect 7624 -3895 7636 -3519
rect 7670 -3895 7682 -3519
rect 7624 -3907 7682 -3895
rect 7742 -3519 7800 -3507
rect 7742 -3895 7754 -3519
rect 7788 -3895 7800 -3519
rect 7742 -3907 7800 -3895
rect 7860 -3519 7918 -3507
rect 7860 -3895 7872 -3519
rect 7906 -3895 7918 -3519
rect 7860 -3907 7918 -3895
rect 13146 -3021 13204 -3009
rect 13146 -3197 13158 -3021
rect 13192 -3197 13204 -3021
rect 13146 -3209 13204 -3197
rect 13264 -3021 13322 -3009
rect 13264 -3197 13276 -3021
rect 13310 -3197 13322 -3021
rect 13264 -3209 13322 -3197
rect 13382 -3021 13440 -3009
rect 13382 -3197 13394 -3021
rect 13428 -3197 13440 -3021
rect 13382 -3209 13440 -3197
rect 13500 -3021 13558 -3009
rect 13500 -3197 13512 -3021
rect 13546 -3197 13558 -3021
rect 13500 -3209 13558 -3197
rect 13629 -3197 13641 -2821
rect 13675 -3197 13687 -2821
rect 13629 -3209 13687 -3197
rect 13747 -2821 13805 -2809
rect 13747 -3197 13759 -2821
rect 13793 -3197 13805 -2821
rect 13747 -3209 13805 -3197
rect 13865 -2821 13923 -2809
rect 13865 -3197 13877 -2821
rect 13911 -3197 13923 -2821
rect 13865 -3209 13923 -3197
rect 13983 -2821 14041 -2809
rect 13983 -3197 13995 -2821
rect 14029 -3197 14041 -2821
rect 13983 -3209 14041 -3197
rect 14101 -2821 14159 -2809
rect 14101 -3197 14113 -2821
rect 14147 -3197 14159 -2821
rect 14101 -3209 14159 -3197
rect 14219 -2821 14277 -2809
rect 14219 -3197 14231 -2821
rect 14265 -3197 14277 -2821
rect 14219 -3209 14277 -3197
rect 14337 -2821 14395 -2809
rect 14337 -3197 14349 -2821
rect 14383 -3197 14395 -2821
rect 15527 -2821 15585 -2809
rect 14337 -3209 14395 -3197
rect 14467 -3021 14525 -3009
rect 14467 -3197 14479 -3021
rect 14513 -3197 14525 -3021
rect 14467 -3209 14525 -3197
rect 14585 -3021 14643 -3009
rect 14585 -3197 14597 -3021
rect 14631 -3197 14643 -3021
rect 14585 -3209 14643 -3197
rect 14703 -3021 14761 -3009
rect 14703 -3197 14715 -3021
rect 14749 -3197 14761 -3021
rect 14703 -3209 14761 -3197
rect 14821 -3021 14879 -3009
rect 14821 -3197 14833 -3021
rect 14867 -3197 14879 -3021
rect 14821 -3209 14879 -3197
rect 15044 -3021 15102 -3009
rect 15044 -3197 15056 -3021
rect 15090 -3197 15102 -3021
rect 15044 -3209 15102 -3197
rect 15162 -3021 15220 -3009
rect 15162 -3197 15174 -3021
rect 15208 -3197 15220 -3021
rect 15162 -3209 15220 -3197
rect 15280 -3021 15338 -3009
rect 15280 -3197 15292 -3021
rect 15326 -3197 15338 -3021
rect 15280 -3209 15338 -3197
rect 15398 -3021 15456 -3009
rect 15398 -3197 15410 -3021
rect 15444 -3197 15456 -3021
rect 15398 -3209 15456 -3197
rect 15527 -3197 15539 -2821
rect 15573 -3197 15585 -2821
rect 15527 -3209 15585 -3197
rect 15645 -2821 15703 -2809
rect 15645 -3197 15657 -2821
rect 15691 -3197 15703 -2821
rect 15645 -3209 15703 -3197
rect 15763 -2821 15821 -2809
rect 15763 -3197 15775 -2821
rect 15809 -3197 15821 -2821
rect 15763 -3209 15821 -3197
rect 15881 -2821 15939 -2809
rect 15881 -3197 15893 -2821
rect 15927 -3197 15939 -2821
rect 15881 -3209 15939 -3197
rect 15999 -2821 16057 -2809
rect 15999 -3197 16011 -2821
rect 16045 -3197 16057 -2821
rect 15999 -3209 16057 -3197
rect 16117 -2821 16175 -2809
rect 16117 -3197 16129 -2821
rect 16163 -3197 16175 -2821
rect 16117 -3209 16175 -3197
rect 16235 -2821 16293 -2809
rect 16235 -3197 16247 -2821
rect 16281 -3197 16293 -2821
rect 20142 -2818 20200 -2806
rect 16235 -3209 16293 -3197
rect 16365 -3021 16423 -3009
rect 16365 -3197 16377 -3021
rect 16411 -3197 16423 -3021
rect 16365 -3209 16423 -3197
rect 16483 -3021 16541 -3009
rect 16483 -3197 16495 -3021
rect 16529 -3197 16541 -3021
rect 16483 -3209 16541 -3197
rect 16601 -3021 16659 -3009
rect 16601 -3197 16613 -3021
rect 16647 -3197 16659 -3021
rect 16601 -3209 16659 -3197
rect 16719 -3021 16777 -3009
rect 16719 -3197 16731 -3021
rect 16765 -3197 16777 -3021
rect 16719 -3209 16777 -3197
rect 9050 -3519 9108 -3507
rect 9050 -3895 9062 -3519
rect 9096 -3895 9108 -3519
rect 9050 -3907 9108 -3895
rect 9168 -3519 9226 -3507
rect 9168 -3895 9180 -3519
rect 9214 -3895 9226 -3519
rect 9168 -3907 9226 -3895
rect 9286 -3519 9344 -3507
rect 9286 -3895 9298 -3519
rect 9332 -3895 9344 -3519
rect 9286 -3907 9344 -3895
rect 9404 -3519 9462 -3507
rect 9404 -3895 9416 -3519
rect 9450 -3895 9462 -3519
rect 9404 -3907 9462 -3895
rect 9522 -3519 9580 -3507
rect 9522 -3895 9534 -3519
rect 9568 -3895 9580 -3519
rect 9522 -3907 9580 -3895
rect 9640 -3519 9698 -3507
rect 9640 -3895 9652 -3519
rect 9686 -3895 9698 -3519
rect 9640 -3907 9698 -3895
rect 9758 -3519 9816 -3507
rect 9758 -3895 9770 -3519
rect 9804 -3895 9816 -3519
rect 9758 -3907 9816 -3895
rect 10592 -4013 10650 -4001
rect 10592 -4189 10604 -4013
rect 10638 -4189 10650 -4013
rect 10592 -4201 10650 -4189
rect 10710 -4013 10768 -4001
rect 10710 -4189 10722 -4013
rect 10756 -4189 10768 -4013
rect 10710 -4201 10768 -4189
rect 10828 -4013 10886 -4001
rect 10828 -4189 10840 -4013
rect 10874 -4189 10886 -4013
rect 10828 -4201 10886 -4189
rect 10946 -4013 11004 -4001
rect 10946 -4189 10958 -4013
rect 10992 -4189 11004 -4013
rect 10946 -4201 11004 -4189
rect 11064 -4013 11122 -4001
rect 11064 -4189 11076 -4013
rect 11110 -4189 11122 -4013
rect 11064 -4201 11122 -4189
rect 11182 -4013 11240 -4001
rect 11182 -4189 11194 -4013
rect 11228 -4189 11240 -4013
rect 11182 -4201 11240 -4189
rect 11300 -4013 11358 -4001
rect 11300 -4189 11312 -4013
rect 11346 -4189 11358 -4013
rect 11300 -4201 11358 -4189
rect 11418 -4013 11476 -4001
rect 11418 -4189 11430 -4013
rect 11464 -4189 11476 -4013
rect 11418 -4201 11476 -4189
rect 11536 -4013 11594 -4001
rect 11536 -4189 11548 -4013
rect 11582 -4189 11594 -4013
rect 11536 -4201 11594 -4189
rect 11654 -4013 11712 -4001
rect 11654 -4189 11666 -4013
rect 11700 -4189 11712 -4013
rect 11654 -4201 11712 -4189
rect 13686 -3514 13744 -3502
rect 13686 -3890 13698 -3514
rect 13732 -3890 13744 -3514
rect 13686 -3902 13744 -3890
rect 13804 -3514 13862 -3502
rect 13804 -3890 13816 -3514
rect 13850 -3890 13862 -3514
rect 13804 -3902 13862 -3890
rect 13922 -3514 13980 -3502
rect 13922 -3890 13934 -3514
rect 13968 -3890 13980 -3514
rect 13922 -3902 13980 -3890
rect 14040 -3514 14098 -3502
rect 14040 -3890 14052 -3514
rect 14086 -3890 14098 -3514
rect 14040 -3902 14098 -3890
rect 14158 -3514 14216 -3502
rect 14158 -3890 14170 -3514
rect 14204 -3890 14216 -3514
rect 14158 -3902 14216 -3890
rect 14276 -3514 14334 -3502
rect 14276 -3890 14288 -3514
rect 14322 -3890 14334 -3514
rect 14276 -3902 14334 -3890
rect 14394 -3514 14452 -3502
rect 14394 -3890 14406 -3514
rect 14440 -3890 14452 -3514
rect 14394 -3902 14452 -3890
rect 19659 -3018 19717 -3006
rect 19659 -3194 19671 -3018
rect 19705 -3194 19717 -3018
rect 19659 -3206 19717 -3194
rect 19777 -3018 19835 -3006
rect 19777 -3194 19789 -3018
rect 19823 -3194 19835 -3018
rect 19777 -3206 19835 -3194
rect 19895 -3018 19953 -3006
rect 19895 -3194 19907 -3018
rect 19941 -3194 19953 -3018
rect 19895 -3206 19953 -3194
rect 20013 -3018 20071 -3006
rect 20013 -3194 20025 -3018
rect 20059 -3194 20071 -3018
rect 20013 -3206 20071 -3194
rect 20142 -3194 20154 -2818
rect 20188 -3194 20200 -2818
rect 20142 -3206 20200 -3194
rect 20260 -2818 20318 -2806
rect 20260 -3194 20272 -2818
rect 20306 -3194 20318 -2818
rect 20260 -3206 20318 -3194
rect 20378 -2818 20436 -2806
rect 20378 -3194 20390 -2818
rect 20424 -3194 20436 -2818
rect 20378 -3206 20436 -3194
rect 20496 -2818 20554 -2806
rect 20496 -3194 20508 -2818
rect 20542 -3194 20554 -2818
rect 20496 -3206 20554 -3194
rect 20614 -2818 20672 -2806
rect 20614 -3194 20626 -2818
rect 20660 -3194 20672 -2818
rect 20614 -3206 20672 -3194
rect 20732 -2818 20790 -2806
rect 20732 -3194 20744 -2818
rect 20778 -3194 20790 -2818
rect 20732 -3206 20790 -3194
rect 20850 -2818 20908 -2806
rect 20850 -3194 20862 -2818
rect 20896 -3194 20908 -2818
rect 22040 -2818 22098 -2806
rect 20850 -3206 20908 -3194
rect 20980 -3018 21038 -3006
rect 20980 -3194 20992 -3018
rect 21026 -3194 21038 -3018
rect 20980 -3206 21038 -3194
rect 21098 -3018 21156 -3006
rect 21098 -3194 21110 -3018
rect 21144 -3194 21156 -3018
rect 21098 -3206 21156 -3194
rect 21216 -3018 21274 -3006
rect 21216 -3194 21228 -3018
rect 21262 -3194 21274 -3018
rect 21216 -3206 21274 -3194
rect 21334 -3018 21392 -3006
rect 21334 -3194 21346 -3018
rect 21380 -3194 21392 -3018
rect 21334 -3206 21392 -3194
rect 21557 -3018 21615 -3006
rect 21557 -3194 21569 -3018
rect 21603 -3194 21615 -3018
rect 21557 -3206 21615 -3194
rect 21675 -3018 21733 -3006
rect 21675 -3194 21687 -3018
rect 21721 -3194 21733 -3018
rect 21675 -3206 21733 -3194
rect 21793 -3018 21851 -3006
rect 21793 -3194 21805 -3018
rect 21839 -3194 21851 -3018
rect 21793 -3206 21851 -3194
rect 21911 -3018 21969 -3006
rect 21911 -3194 21923 -3018
rect 21957 -3194 21969 -3018
rect 21911 -3206 21969 -3194
rect 22040 -3194 22052 -2818
rect 22086 -3194 22098 -2818
rect 22040 -3206 22098 -3194
rect 22158 -2818 22216 -2806
rect 22158 -3194 22170 -2818
rect 22204 -3194 22216 -2818
rect 22158 -3206 22216 -3194
rect 22276 -2818 22334 -2806
rect 22276 -3194 22288 -2818
rect 22322 -3194 22334 -2818
rect 22276 -3206 22334 -3194
rect 22394 -2818 22452 -2806
rect 22394 -3194 22406 -2818
rect 22440 -3194 22452 -2818
rect 22394 -3206 22452 -3194
rect 22512 -2818 22570 -2806
rect 22512 -3194 22524 -2818
rect 22558 -3194 22570 -2818
rect 22512 -3206 22570 -3194
rect 22630 -2818 22688 -2806
rect 22630 -3194 22642 -2818
rect 22676 -3194 22688 -2818
rect 22630 -3206 22688 -3194
rect 22748 -2818 22806 -2806
rect 22748 -3194 22760 -2818
rect 22794 -3194 22806 -2818
rect 22748 -3206 22806 -3194
rect 22878 -3018 22936 -3006
rect 22878 -3194 22890 -3018
rect 22924 -3194 22936 -3018
rect 22878 -3206 22936 -3194
rect 22996 -3018 23054 -3006
rect 22996 -3194 23008 -3018
rect 23042 -3194 23054 -3018
rect 22996 -3206 23054 -3194
rect 23114 -3018 23172 -3006
rect 23114 -3194 23126 -3018
rect 23160 -3194 23172 -3018
rect 23114 -3206 23172 -3194
rect 23232 -3018 23290 -3006
rect 23232 -3194 23244 -3018
rect 23278 -3194 23290 -3018
rect 23232 -3206 23290 -3194
rect 15584 -3514 15642 -3502
rect 15584 -3890 15596 -3514
rect 15630 -3890 15642 -3514
rect 15584 -3902 15642 -3890
rect 15702 -3514 15760 -3502
rect 15702 -3890 15714 -3514
rect 15748 -3890 15760 -3514
rect 15702 -3902 15760 -3890
rect 15820 -3514 15878 -3502
rect 15820 -3890 15832 -3514
rect 15866 -3890 15878 -3514
rect 15820 -3902 15878 -3890
rect 15938 -3514 15996 -3502
rect 15938 -3890 15950 -3514
rect 15984 -3890 15996 -3514
rect 15938 -3902 15996 -3890
rect 16056 -3514 16114 -3502
rect 16056 -3890 16068 -3514
rect 16102 -3890 16114 -3514
rect 16056 -3902 16114 -3890
rect 16174 -3514 16232 -3502
rect 16174 -3890 16186 -3514
rect 16220 -3890 16232 -3514
rect 16174 -3902 16232 -3890
rect 16292 -3514 16350 -3502
rect 16292 -3890 16304 -3514
rect 16338 -3890 16350 -3514
rect 16292 -3902 16350 -3890
rect 17126 -4008 17184 -3996
rect 17126 -4184 17138 -4008
rect 17172 -4184 17184 -4008
rect 17126 -4196 17184 -4184
rect 17244 -4008 17302 -3996
rect 17244 -4184 17256 -4008
rect 17290 -4184 17302 -4008
rect 17244 -4196 17302 -4184
rect 17362 -4008 17420 -3996
rect 17362 -4184 17374 -4008
rect 17408 -4184 17420 -4008
rect 17362 -4196 17420 -4184
rect 17480 -4008 17538 -3996
rect 17480 -4184 17492 -4008
rect 17526 -4184 17538 -4008
rect 17480 -4196 17538 -4184
rect 17598 -4008 17656 -3996
rect 17598 -4184 17610 -4008
rect 17644 -4184 17656 -4008
rect 17598 -4196 17656 -4184
rect 17716 -4008 17774 -3996
rect 17716 -4184 17728 -4008
rect 17762 -4184 17774 -4008
rect 17716 -4196 17774 -4184
rect 17834 -4008 17892 -3996
rect 17834 -4184 17846 -4008
rect 17880 -4184 17892 -4008
rect 17834 -4196 17892 -4184
rect 17952 -4008 18010 -3996
rect 17952 -4184 17964 -4008
rect 17998 -4184 18010 -4008
rect 17952 -4196 18010 -4184
rect 18070 -4008 18128 -3996
rect 18070 -4184 18082 -4008
rect 18116 -4184 18128 -4008
rect 18070 -4196 18128 -4184
rect 18188 -4008 18246 -3996
rect 18188 -4184 18200 -4008
rect 18234 -4184 18246 -4008
rect 18188 -4196 18246 -4184
rect 20199 -3511 20257 -3499
rect 20199 -3887 20211 -3511
rect 20245 -3887 20257 -3511
rect 20199 -3899 20257 -3887
rect 20317 -3511 20375 -3499
rect 20317 -3887 20329 -3511
rect 20363 -3887 20375 -3511
rect 20317 -3899 20375 -3887
rect 20435 -3511 20493 -3499
rect 20435 -3887 20447 -3511
rect 20481 -3887 20493 -3511
rect 20435 -3899 20493 -3887
rect 20553 -3511 20611 -3499
rect 20553 -3887 20565 -3511
rect 20599 -3887 20611 -3511
rect 20553 -3899 20611 -3887
rect 20671 -3511 20729 -3499
rect 20671 -3887 20683 -3511
rect 20717 -3887 20729 -3511
rect 20671 -3899 20729 -3887
rect 20789 -3511 20847 -3499
rect 20789 -3887 20801 -3511
rect 20835 -3887 20847 -3511
rect 20789 -3899 20847 -3887
rect 20907 -3511 20965 -3499
rect 20907 -3887 20919 -3511
rect 20953 -3887 20965 -3511
rect 20907 -3899 20965 -3887
rect 22097 -3511 22155 -3499
rect 22097 -3887 22109 -3511
rect 22143 -3887 22155 -3511
rect 22097 -3899 22155 -3887
rect 22215 -3511 22273 -3499
rect 22215 -3887 22227 -3511
rect 22261 -3887 22273 -3511
rect 22215 -3899 22273 -3887
rect 22333 -3511 22391 -3499
rect 22333 -3887 22345 -3511
rect 22379 -3887 22391 -3511
rect 22333 -3899 22391 -3887
rect 22451 -3511 22509 -3499
rect 22451 -3887 22463 -3511
rect 22497 -3887 22509 -3511
rect 22451 -3899 22509 -3887
rect 22569 -3511 22627 -3499
rect 22569 -3887 22581 -3511
rect 22615 -3887 22627 -3511
rect 22569 -3899 22627 -3887
rect 22687 -3511 22745 -3499
rect 22687 -3887 22699 -3511
rect 22733 -3887 22745 -3511
rect 22687 -3899 22745 -3887
rect 22805 -3511 22863 -3499
rect 22805 -3887 22817 -3511
rect 22851 -3887 22863 -3511
rect 22805 -3899 22863 -3887
rect 23639 -4005 23697 -3993
rect 23639 -4181 23651 -4005
rect 23685 -4181 23697 -4005
rect 23639 -4193 23697 -4181
rect 23757 -4005 23815 -3993
rect 23757 -4181 23769 -4005
rect 23803 -4181 23815 -4005
rect 23757 -4193 23815 -4181
rect 23875 -4005 23933 -3993
rect 23875 -4181 23887 -4005
rect 23921 -4181 23933 -4005
rect 23875 -4193 23933 -4181
rect 23993 -4005 24051 -3993
rect 23993 -4181 24005 -4005
rect 24039 -4181 24051 -4005
rect 23993 -4193 24051 -4181
rect 24111 -4005 24169 -3993
rect 24111 -4181 24123 -4005
rect 24157 -4181 24169 -4005
rect 24111 -4193 24169 -4181
rect 24229 -4005 24287 -3993
rect 24229 -4181 24241 -4005
rect 24275 -4181 24287 -4005
rect 24229 -4193 24287 -4181
rect 24347 -4005 24405 -3993
rect 24347 -4181 24359 -4005
rect 24393 -4181 24405 -4005
rect 24347 -4193 24405 -4181
rect 24465 -4005 24523 -3993
rect 24465 -4181 24477 -4005
rect 24511 -4181 24523 -4005
rect 24465 -4193 24523 -4181
rect 24583 -4005 24641 -3993
rect 24583 -4181 24595 -4005
rect 24629 -4181 24641 -4005
rect 24583 -4193 24641 -4181
rect 24701 -4005 24759 -3993
rect 24701 -4181 24713 -4005
rect 24747 -4181 24759 -4005
rect 24701 -4193 24759 -4181
<< ndiffc >>
rect 1168 4040 1202 4416
rect 1286 4040 1320 4416
rect 1404 4040 1438 4416
rect 1521 4240 1555 4416
rect 1639 4240 1673 4416
rect 3166 3966 3200 4142
rect 3284 3966 3318 4142
rect 3402 3966 3436 4142
rect 3520 3966 3554 4142
rect 4308 3970 4342 4146
rect 4426 3970 4460 4146
rect 4544 3970 4578 4146
rect 4662 3970 4696 4146
rect 7681 4037 7715 4413
rect 7799 4037 7833 4413
rect 7917 4037 7951 4413
rect 8034 4237 8068 4413
rect 8152 4237 8186 4413
rect 9679 3963 9713 4139
rect 9797 3963 9831 4139
rect 9915 3963 9949 4139
rect 10033 3963 10067 4139
rect 10821 3967 10855 4143
rect 10939 3967 10973 4143
rect 11057 3967 11091 4143
rect 11175 3967 11209 4143
rect 14215 4032 14249 4408
rect 14333 4032 14367 4408
rect 14451 4032 14485 4408
rect 14568 4232 14602 4408
rect 14686 4232 14720 4408
rect 16213 3958 16247 4134
rect 16331 3958 16365 4134
rect 16449 3958 16483 4134
rect 16567 3958 16601 4134
rect 17355 3962 17389 4138
rect 17473 3962 17507 4138
rect 17591 3962 17625 4138
rect 17709 3962 17743 4138
rect 20773 4036 20807 4412
rect 20891 4036 20925 4412
rect 21009 4036 21043 4412
rect 21126 4236 21160 4412
rect 21244 4236 21278 4412
rect 22771 3962 22805 4138
rect 22889 3962 22923 4138
rect 23007 3962 23041 4138
rect 23125 3962 23159 4138
rect 23913 3966 23947 4142
rect 24031 3966 24065 4142
rect 24149 3966 24183 4142
rect 24267 3966 24301 4142
rect 1182 2390 1216 2766
rect 1300 2390 1334 2766
rect 1418 2390 1452 2766
rect 1535 2590 1569 2766
rect 1653 2590 1687 2766
rect 7695 2387 7729 2763
rect 7813 2387 7847 2763
rect 7931 2387 7965 2763
rect 8048 2587 8082 2763
rect 8166 2587 8200 2763
rect 2534 1185 2568 1361
rect 1177 786 1211 1162
rect 1295 786 1329 1162
rect 1413 786 1447 1162
rect 1530 986 1564 1162
rect 2652 1185 2686 1361
rect 1648 986 1682 1162
rect 2954 985 2988 1361
rect 3072 985 3106 1361
rect 3190 985 3224 1361
rect 3308 985 3342 1361
rect 3426 985 3460 1361
rect 3832 1185 3866 1361
rect 3950 1185 3984 1361
rect 4432 1185 4466 1361
rect 4550 1185 4584 1361
rect 4852 985 4886 1361
rect 4970 985 5004 1361
rect 5088 985 5122 1361
rect 5206 985 5240 1361
rect 5324 985 5358 1361
rect 5730 1185 5764 1361
rect 5848 1185 5882 1361
rect 14229 2382 14263 2758
rect 14347 2382 14381 2758
rect 14465 2382 14499 2758
rect 14582 2582 14616 2758
rect 14700 2582 14734 2758
rect 9047 1182 9081 1358
rect 7690 783 7724 1159
rect 7808 783 7842 1159
rect 7926 783 7960 1159
rect 8043 983 8077 1159
rect 9165 1182 9199 1358
rect 8161 983 8195 1159
rect 9467 982 9501 1358
rect 9585 982 9619 1358
rect 9703 982 9737 1358
rect 9821 982 9855 1358
rect 9939 982 9973 1358
rect 10345 1182 10379 1358
rect 10463 1182 10497 1358
rect 10945 1182 10979 1358
rect 11063 1182 11097 1358
rect 11365 982 11399 1358
rect 11483 982 11517 1358
rect 11601 982 11635 1358
rect 11719 982 11753 1358
rect 11837 982 11871 1358
rect 12243 1182 12277 1358
rect 12361 1182 12395 1358
rect 20787 2386 20821 2762
rect 20905 2386 20939 2762
rect 21023 2386 21057 2762
rect 21140 2586 21174 2762
rect 21258 2586 21292 2762
rect 15581 1177 15615 1353
rect 14224 778 14258 1154
rect 14342 778 14376 1154
rect 14460 778 14494 1154
rect 14577 978 14611 1154
rect 15699 1177 15733 1353
rect 14695 978 14729 1154
rect 16001 977 16035 1353
rect 16119 977 16153 1353
rect 16237 977 16271 1353
rect 16355 977 16389 1353
rect 16473 977 16507 1353
rect 16879 1177 16913 1353
rect 16997 1177 17031 1353
rect 17479 1177 17513 1353
rect 17597 1177 17631 1353
rect 17899 977 17933 1353
rect 18017 977 18051 1353
rect 18135 977 18169 1353
rect 18253 977 18287 1353
rect 18371 977 18405 1353
rect 18777 1177 18811 1353
rect 18895 1177 18929 1353
rect 22139 1181 22173 1357
rect 20782 782 20816 1158
rect 20900 782 20934 1158
rect 21018 782 21052 1158
rect 21135 982 21169 1158
rect 22257 1181 22291 1357
rect 21253 982 21287 1158
rect 22559 981 22593 1357
rect 22677 981 22711 1357
rect 22795 981 22829 1357
rect 22913 981 22947 1357
rect 23031 981 23065 1357
rect 23437 1181 23471 1357
rect 23555 1181 23589 1357
rect 24037 1181 24071 1357
rect 24155 1181 24189 1357
rect 24457 981 24491 1357
rect 24575 981 24609 1357
rect 24693 981 24727 1357
rect 24811 981 24845 1357
rect 24929 981 24963 1357
rect 25335 1181 25369 1357
rect 25453 1181 25487 1357
rect 1386 -1638 1420 -1462
rect 1504 -1638 1538 -1462
rect 1622 -1638 1656 -1462
rect 4409 -1368 4443 -1192
rect 4527 -1368 4561 -1192
rect 1740 -1638 1774 -1462
rect 2528 -1642 2562 -1466
rect 2646 -1642 2680 -1466
rect 2764 -1642 2798 -1466
rect 2882 -1642 2916 -1466
rect 4644 -1568 4678 -1192
rect 4762 -1568 4796 -1192
rect 4880 -1568 4914 -1192
rect 7944 -1642 7978 -1466
rect 8062 -1642 8096 -1466
rect 8180 -1642 8214 -1466
rect 10967 -1372 11001 -1196
rect 11085 -1372 11119 -1196
rect 8298 -1642 8332 -1466
rect 9086 -1646 9120 -1470
rect 9204 -1646 9238 -1470
rect 9322 -1646 9356 -1470
rect 9440 -1646 9474 -1470
rect 11202 -1572 11236 -1196
rect 11320 -1572 11354 -1196
rect 11438 -1572 11472 -1196
rect 14478 -1637 14512 -1461
rect 14596 -1637 14630 -1461
rect 14714 -1637 14748 -1461
rect 17501 -1367 17535 -1191
rect 17619 -1367 17653 -1191
rect 14832 -1637 14866 -1461
rect 15620 -1641 15654 -1465
rect 15738 -1641 15772 -1465
rect 15856 -1641 15890 -1465
rect 15974 -1641 16008 -1465
rect 17736 -1567 17770 -1191
rect 17854 -1567 17888 -1191
rect 17972 -1567 18006 -1191
rect 20991 -1634 21025 -1458
rect 21109 -1634 21143 -1458
rect 21227 -1634 21261 -1458
rect 24014 -1364 24048 -1188
rect 24132 -1364 24166 -1188
rect 21345 -1634 21379 -1458
rect 22133 -1638 22167 -1462
rect 22251 -1638 22285 -1462
rect 22369 -1638 22403 -1462
rect 22487 -1638 22521 -1462
rect 24249 -1564 24283 -1188
rect 24367 -1564 24401 -1188
rect 24485 -1564 24519 -1188
rect 4395 -3018 4429 -2842
rect 4513 -3018 4547 -2842
rect 4630 -3218 4664 -2842
rect 4748 -3218 4782 -2842
rect 4866 -3218 4900 -2842
rect 10953 -3022 10987 -2846
rect 11071 -3022 11105 -2846
rect 200 -4423 234 -4247
rect 318 -4423 352 -4247
rect 724 -4623 758 -4247
rect 842 -4623 876 -4247
rect 960 -4623 994 -4247
rect 1078 -4623 1112 -4247
rect 1196 -4623 1230 -4247
rect 1498 -4423 1532 -4247
rect 1616 -4423 1650 -4247
rect 2098 -4423 2132 -4247
rect 2216 -4423 2250 -4247
rect 2622 -4623 2656 -4247
rect 2740 -4623 2774 -4247
rect 2858 -4623 2892 -4247
rect 2976 -4623 3010 -4247
rect 3094 -4623 3128 -4247
rect 3396 -4423 3430 -4247
rect 3514 -4423 3548 -4247
rect 11188 -3222 11222 -2846
rect 11306 -3222 11340 -2846
rect 11424 -3222 11458 -2846
rect 17487 -3017 17521 -2841
rect 17605 -3017 17639 -2841
rect 6758 -4427 6792 -4251
rect 4400 -4622 4434 -4446
rect 4518 -4622 4552 -4446
rect 4635 -4822 4669 -4446
rect 4753 -4822 4787 -4446
rect 6876 -4427 6910 -4251
rect 4871 -4822 4905 -4446
rect 7282 -4627 7316 -4251
rect 7400 -4627 7434 -4251
rect 7518 -4627 7552 -4251
rect 7636 -4627 7670 -4251
rect 7754 -4627 7788 -4251
rect 8056 -4427 8090 -4251
rect 8174 -4427 8208 -4251
rect 8656 -4427 8690 -4251
rect 8774 -4427 8808 -4251
rect 9180 -4627 9214 -4251
rect 9298 -4627 9332 -4251
rect 9416 -4627 9450 -4251
rect 9534 -4627 9568 -4251
rect 9652 -4627 9686 -4251
rect 9954 -4427 9988 -4251
rect 10072 -4427 10106 -4251
rect 17722 -3217 17756 -2841
rect 17840 -3217 17874 -2841
rect 17958 -3217 17992 -2841
rect 24000 -3014 24034 -2838
rect 24118 -3014 24152 -2838
rect 13292 -4422 13326 -4246
rect 13410 -4422 13444 -4246
rect 10958 -4626 10992 -4450
rect 11076 -4626 11110 -4450
rect 11193 -4826 11227 -4450
rect 11311 -4826 11345 -4450
rect 11429 -4826 11463 -4450
rect 13816 -4622 13850 -4246
rect 13934 -4622 13968 -4246
rect 14052 -4622 14086 -4246
rect 14170 -4622 14204 -4246
rect 14288 -4622 14322 -4246
rect 14590 -4422 14624 -4246
rect 14708 -4422 14742 -4246
rect 15190 -4422 15224 -4246
rect 15308 -4422 15342 -4246
rect 15714 -4622 15748 -4246
rect 15832 -4622 15866 -4246
rect 15950 -4622 15984 -4246
rect 16068 -4622 16102 -4246
rect 16186 -4622 16220 -4246
rect 16488 -4422 16522 -4246
rect 16606 -4422 16640 -4246
rect 24235 -3214 24269 -2838
rect 24353 -3214 24387 -2838
rect 24471 -3214 24505 -2838
rect 19805 -4419 19839 -4243
rect 19923 -4419 19957 -4243
rect 17492 -4621 17526 -4445
rect 17610 -4621 17644 -4445
rect 17727 -4821 17761 -4445
rect 17845 -4821 17879 -4445
rect 17963 -4821 17997 -4445
rect 20329 -4619 20363 -4243
rect 20447 -4619 20481 -4243
rect 20565 -4619 20599 -4243
rect 20683 -4619 20717 -4243
rect 20801 -4619 20835 -4243
rect 21103 -4419 21137 -4243
rect 21221 -4419 21255 -4243
rect 21703 -4419 21737 -4243
rect 21821 -4419 21855 -4243
rect 22227 -4619 22261 -4243
rect 22345 -4619 22379 -4243
rect 22463 -4619 22497 -4243
rect 22581 -4619 22615 -4243
rect 22699 -4619 22733 -4243
rect 23001 -4419 23035 -4243
rect 23119 -4419 23153 -4243
rect 24005 -4618 24039 -4442
rect 24123 -4618 24157 -4442
rect 24240 -4818 24274 -4442
rect 24358 -4818 24392 -4442
rect 24476 -4818 24510 -4442
<< pdiffc >>
rect 931 4677 965 4853
rect 1049 4677 1083 4853
rect 1167 4677 1201 4853
rect 1285 4677 1319 4853
rect 1403 4677 1437 4853
rect 1521 4677 1555 4853
rect 1639 4677 1673 4853
rect 1757 4677 1791 4853
rect 1875 4677 1909 4853
rect 1993 4677 2027 4853
rect 3256 4549 3290 4925
rect 3374 4549 3408 4925
rect 3492 4549 3526 4925
rect 3610 4549 3644 4925
rect 3728 4549 3762 4925
rect 3846 4549 3880 4925
rect 3964 4549 3998 4925
rect 4398 4553 4432 4929
rect 4516 4553 4550 4929
rect 4634 4553 4668 4929
rect 4752 4553 4786 4929
rect 4870 4553 4904 4929
rect 4988 4553 5022 4929
rect 5106 4553 5140 4929
rect 7444 4674 7478 4850
rect 7562 4674 7596 4850
rect 7680 4674 7714 4850
rect 7798 4674 7832 4850
rect 7916 4674 7950 4850
rect 8034 4674 8068 4850
rect 8152 4674 8186 4850
rect 8270 4674 8304 4850
rect 8388 4674 8422 4850
rect 8506 4674 8540 4850
rect 9769 4546 9803 4922
rect 9887 4546 9921 4922
rect 10005 4546 10039 4922
rect 10123 4546 10157 4922
rect 10241 4546 10275 4922
rect 10359 4546 10393 4922
rect 10477 4546 10511 4922
rect 10911 4550 10945 4926
rect 11029 4550 11063 4926
rect 11147 4550 11181 4926
rect 11265 4550 11299 4926
rect 11383 4550 11417 4926
rect 11501 4550 11535 4926
rect 11619 4550 11653 4926
rect 13978 4669 14012 4845
rect 14096 4669 14130 4845
rect 14214 4669 14248 4845
rect 14332 4669 14366 4845
rect 14450 4669 14484 4845
rect 14568 4669 14602 4845
rect 14686 4669 14720 4845
rect 14804 4669 14838 4845
rect 14922 4669 14956 4845
rect 15040 4669 15074 4845
rect 3685 3966 3719 4142
rect 3803 3966 3837 4142
rect 3921 3966 3955 4142
rect 4039 3966 4073 4142
rect 4827 3970 4861 4146
rect 4945 3970 4979 4146
rect 5063 3970 5097 4146
rect 5181 3970 5215 4146
rect 16303 4541 16337 4917
rect 16421 4541 16455 4917
rect 16539 4541 16573 4917
rect 16657 4541 16691 4917
rect 16775 4541 16809 4917
rect 16893 4541 16927 4917
rect 17011 4541 17045 4917
rect 17445 4545 17479 4921
rect 17563 4545 17597 4921
rect 17681 4545 17715 4921
rect 17799 4545 17833 4921
rect 17917 4545 17951 4921
rect 18035 4545 18069 4921
rect 18153 4545 18187 4921
rect 20536 4673 20570 4849
rect 20654 4673 20688 4849
rect 20772 4673 20806 4849
rect 20890 4673 20924 4849
rect 21008 4673 21042 4849
rect 21126 4673 21160 4849
rect 21244 4673 21278 4849
rect 21362 4673 21396 4849
rect 21480 4673 21514 4849
rect 21598 4673 21632 4849
rect 10198 3963 10232 4139
rect 10316 3963 10350 4139
rect 10434 3963 10468 4139
rect 10552 3963 10586 4139
rect 11340 3967 11374 4143
rect 11458 3967 11492 4143
rect 11576 3967 11610 4143
rect 11694 3967 11728 4143
rect 22861 4545 22895 4921
rect 22979 4545 23013 4921
rect 23097 4545 23131 4921
rect 23215 4545 23249 4921
rect 23333 4545 23367 4921
rect 23451 4545 23485 4921
rect 23569 4545 23603 4921
rect 24003 4549 24037 4925
rect 24121 4549 24155 4925
rect 24239 4549 24273 4925
rect 24357 4549 24391 4925
rect 24475 4549 24509 4925
rect 24593 4549 24627 4925
rect 24711 4549 24745 4925
rect 16732 3958 16766 4134
rect 16850 3958 16884 4134
rect 16968 3958 17002 4134
rect 17086 3958 17120 4134
rect 17874 3962 17908 4138
rect 17992 3962 18026 4138
rect 18110 3962 18144 4138
rect 18228 3962 18262 4138
rect 23290 3962 23324 4138
rect 23408 3962 23442 4138
rect 23526 3962 23560 4138
rect 23644 3962 23678 4138
rect 24432 3966 24466 4142
rect 24550 3966 24584 4142
rect 24668 3966 24702 4142
rect 24786 3966 24820 4142
rect 945 3027 979 3203
rect 1063 3027 1097 3203
rect 1181 3027 1215 3203
rect 1299 3027 1333 3203
rect 1417 3027 1451 3203
rect 1535 3027 1569 3203
rect 1653 3027 1687 3203
rect 1771 3027 1805 3203
rect 1889 3027 1923 3203
rect 2007 3027 2041 3203
rect 7458 3024 7492 3200
rect 7576 3024 7610 3200
rect 7694 3024 7728 3200
rect 7812 3024 7846 3200
rect 7930 3024 7964 3200
rect 8048 3024 8082 3200
rect 8166 3024 8200 3200
rect 8284 3024 8318 3200
rect 8402 3024 8436 3200
rect 8520 3024 8554 3200
rect 13992 3019 14026 3195
rect 2409 2410 2443 2586
rect 2527 2410 2561 2586
rect 2645 2410 2679 2586
rect 2763 2410 2797 2586
rect 2893 2410 2927 2786
rect 3011 2410 3045 2786
rect 3129 2410 3163 2786
rect 3247 2410 3281 2786
rect 3365 2410 3399 2786
rect 3483 2410 3517 2786
rect 3601 2410 3635 2786
rect 3730 2410 3764 2586
rect 3848 2410 3882 2586
rect 3966 2410 4000 2586
rect 4084 2410 4118 2586
rect 4307 2410 4341 2586
rect 4425 2410 4459 2586
rect 4543 2410 4577 2586
rect 4661 2410 4695 2586
rect 4791 2410 4825 2786
rect 4909 2410 4943 2786
rect 5027 2410 5061 2786
rect 5145 2410 5179 2786
rect 5263 2410 5297 2786
rect 5381 2410 5415 2786
rect 5499 2410 5533 2786
rect 14110 3019 14144 3195
rect 14228 3019 14262 3195
rect 14346 3019 14380 3195
rect 14464 3019 14498 3195
rect 14582 3019 14616 3195
rect 14700 3019 14734 3195
rect 14818 3019 14852 3195
rect 14936 3019 14970 3195
rect 15054 3019 15088 3195
rect 20550 3023 20584 3199
rect 20668 3023 20702 3199
rect 20786 3023 20820 3199
rect 20904 3023 20938 3199
rect 21022 3023 21056 3199
rect 21140 3023 21174 3199
rect 21258 3023 21292 3199
rect 21376 3023 21410 3199
rect 21494 3023 21528 3199
rect 21612 3023 21646 3199
rect 5628 2410 5662 2586
rect 5746 2410 5780 2586
rect 5864 2410 5898 2586
rect 5982 2410 6016 2586
rect 940 1423 974 1599
rect 1058 1423 1092 1599
rect 1176 1423 1210 1599
rect 1294 1423 1328 1599
rect 1412 1423 1446 1599
rect 1530 1423 1564 1599
rect 1648 1423 1682 1599
rect 1766 1423 1800 1599
rect 1884 1423 1918 1599
rect 2002 1423 2036 1599
rect 2836 1717 2870 2093
rect 2954 1717 2988 2093
rect 3072 1717 3106 2093
rect 3190 1717 3224 2093
rect 3308 1717 3342 2093
rect 3426 1717 3460 2093
rect 3544 1717 3578 2093
rect 8922 2407 8956 2583
rect 9040 2407 9074 2583
rect 9158 2407 9192 2583
rect 9276 2407 9310 2583
rect 9406 2407 9440 2783
rect 9524 2407 9558 2783
rect 9642 2407 9676 2783
rect 9760 2407 9794 2783
rect 9878 2407 9912 2783
rect 9996 2407 10030 2783
rect 10114 2407 10148 2783
rect 10243 2407 10277 2583
rect 10361 2407 10395 2583
rect 10479 2407 10513 2583
rect 10597 2407 10631 2583
rect 10820 2407 10854 2583
rect 10938 2407 10972 2583
rect 11056 2407 11090 2583
rect 11174 2407 11208 2583
rect 11304 2407 11338 2783
rect 11422 2407 11456 2783
rect 11540 2407 11574 2783
rect 11658 2407 11692 2783
rect 11776 2407 11810 2783
rect 11894 2407 11928 2783
rect 12012 2407 12046 2783
rect 12141 2407 12175 2583
rect 12259 2407 12293 2583
rect 12377 2407 12411 2583
rect 12495 2407 12529 2583
rect 4734 1717 4768 2093
rect 4852 1717 4886 2093
rect 4970 1717 5004 2093
rect 5088 1717 5122 2093
rect 5206 1717 5240 2093
rect 5324 1717 5358 2093
rect 5442 1717 5476 2093
rect 7453 1420 7487 1596
rect 7571 1420 7605 1596
rect 7689 1420 7723 1596
rect 7807 1420 7841 1596
rect 7925 1420 7959 1596
rect 8043 1420 8077 1596
rect 8161 1420 8195 1596
rect 8279 1420 8313 1596
rect 8397 1420 8431 1596
rect 8515 1420 8549 1596
rect 9349 1714 9383 2090
rect 9467 1714 9501 2090
rect 9585 1714 9619 2090
rect 9703 1714 9737 2090
rect 9821 1714 9855 2090
rect 9939 1714 9973 2090
rect 10057 1714 10091 2090
rect 15456 2402 15490 2578
rect 15574 2402 15608 2578
rect 15692 2402 15726 2578
rect 15810 2402 15844 2578
rect 15940 2402 15974 2778
rect 16058 2402 16092 2778
rect 16176 2402 16210 2778
rect 16294 2402 16328 2778
rect 16412 2402 16446 2778
rect 16530 2402 16564 2778
rect 16648 2402 16682 2778
rect 16777 2402 16811 2578
rect 16895 2402 16929 2578
rect 17013 2402 17047 2578
rect 17131 2402 17165 2578
rect 17354 2402 17388 2578
rect 17472 2402 17506 2578
rect 17590 2402 17624 2578
rect 17708 2402 17742 2578
rect 17838 2402 17872 2778
rect 17956 2402 17990 2778
rect 18074 2402 18108 2778
rect 18192 2402 18226 2778
rect 18310 2402 18344 2778
rect 18428 2402 18462 2778
rect 18546 2402 18580 2778
rect 18675 2402 18709 2578
rect 18793 2402 18827 2578
rect 18911 2402 18945 2578
rect 19029 2402 19063 2578
rect 11247 1714 11281 2090
rect 11365 1714 11399 2090
rect 11483 1714 11517 2090
rect 11601 1714 11635 2090
rect 11719 1714 11753 2090
rect 11837 1714 11871 2090
rect 11955 1714 11989 2090
rect 13987 1415 14021 1591
rect 14105 1415 14139 1591
rect 14223 1415 14257 1591
rect 14341 1415 14375 1591
rect 14459 1415 14493 1591
rect 14577 1415 14611 1591
rect 14695 1415 14729 1591
rect 14813 1415 14847 1591
rect 14931 1415 14965 1591
rect 15049 1415 15083 1591
rect 15883 1709 15917 2085
rect 16001 1709 16035 2085
rect 16119 1709 16153 2085
rect 16237 1709 16271 2085
rect 16355 1709 16389 2085
rect 16473 1709 16507 2085
rect 16591 1709 16625 2085
rect 22014 2406 22048 2582
rect 22132 2406 22166 2582
rect 22250 2406 22284 2582
rect 22368 2406 22402 2582
rect 22498 2406 22532 2782
rect 22616 2406 22650 2782
rect 22734 2406 22768 2782
rect 22852 2406 22886 2782
rect 22970 2406 23004 2782
rect 23088 2406 23122 2782
rect 23206 2406 23240 2782
rect 23335 2406 23369 2582
rect 23453 2406 23487 2582
rect 23571 2406 23605 2582
rect 23689 2406 23723 2582
rect 23912 2406 23946 2582
rect 24030 2406 24064 2582
rect 24148 2406 24182 2582
rect 24266 2406 24300 2582
rect 24396 2406 24430 2782
rect 24514 2406 24548 2782
rect 24632 2406 24666 2782
rect 24750 2406 24784 2782
rect 24868 2406 24902 2782
rect 24986 2406 25020 2782
rect 25104 2406 25138 2782
rect 25233 2406 25267 2582
rect 25351 2406 25385 2582
rect 25469 2406 25503 2582
rect 25587 2406 25621 2582
rect 17781 1709 17815 2085
rect 17899 1709 17933 2085
rect 18017 1709 18051 2085
rect 18135 1709 18169 2085
rect 18253 1709 18287 2085
rect 18371 1709 18405 2085
rect 18489 1709 18523 2085
rect 20545 1419 20579 1595
rect 20663 1419 20697 1595
rect 20781 1419 20815 1595
rect 20899 1419 20933 1595
rect 21017 1419 21051 1595
rect 21135 1419 21169 1595
rect 21253 1419 21287 1595
rect 21371 1419 21405 1595
rect 21489 1419 21523 1595
rect 21607 1419 21641 1595
rect 22441 1713 22475 2089
rect 22559 1713 22593 2089
rect 22677 1713 22711 2089
rect 22795 1713 22829 2089
rect 22913 1713 22947 2089
rect 23031 1713 23065 2089
rect 23149 1713 23183 2089
rect 24339 1713 24373 2089
rect 24457 1713 24491 2089
rect 24575 1713 24609 2089
rect 24693 1713 24727 2089
rect 24811 1713 24845 2089
rect 24929 1713 24963 2089
rect 25047 1713 25081 2089
rect 942 -1055 976 -679
rect 1060 -1055 1094 -679
rect 1178 -1055 1212 -679
rect 1296 -1055 1330 -679
rect 1414 -1055 1448 -679
rect 1532 -1055 1566 -679
rect 1650 -1055 1684 -679
rect 2084 -1059 2118 -683
rect 2202 -1059 2236 -683
rect 2320 -1059 2354 -683
rect 2438 -1059 2472 -683
rect 2556 -1059 2590 -683
rect 2674 -1059 2708 -683
rect 2792 -1059 2826 -683
rect 4055 -931 4089 -755
rect 4173 -931 4207 -755
rect 4291 -931 4325 -755
rect 4409 -931 4443 -755
rect 4527 -931 4561 -755
rect 4645 -931 4679 -755
rect 4763 -931 4797 -755
rect 4881 -931 4915 -755
rect 4999 -931 5033 -755
rect 5117 -931 5151 -755
rect 7500 -1059 7534 -683
rect 7618 -1059 7652 -683
rect 7736 -1059 7770 -683
rect 7854 -1059 7888 -683
rect 7972 -1059 8006 -683
rect 8090 -1059 8124 -683
rect 8208 -1059 8242 -683
rect 8642 -1063 8676 -687
rect 867 -1638 901 -1462
rect 985 -1638 1019 -1462
rect 1103 -1638 1137 -1462
rect 1221 -1638 1255 -1462
rect 2009 -1642 2043 -1466
rect 2127 -1642 2161 -1466
rect 2245 -1642 2279 -1466
rect 2363 -1642 2397 -1466
rect 8760 -1063 8794 -687
rect 8878 -1063 8912 -687
rect 8996 -1063 9030 -687
rect 9114 -1063 9148 -687
rect 9232 -1063 9266 -687
rect 9350 -1063 9384 -687
rect 10613 -935 10647 -759
rect 10731 -935 10765 -759
rect 10849 -935 10883 -759
rect 10967 -935 11001 -759
rect 11085 -935 11119 -759
rect 11203 -935 11237 -759
rect 11321 -935 11355 -759
rect 11439 -935 11473 -759
rect 11557 -935 11591 -759
rect 11675 -935 11709 -759
rect 14034 -1054 14068 -678
rect 14152 -1054 14186 -678
rect 14270 -1054 14304 -678
rect 14388 -1054 14422 -678
rect 14506 -1054 14540 -678
rect 14624 -1054 14658 -678
rect 14742 -1054 14776 -678
rect 15176 -1058 15210 -682
rect 7425 -1642 7459 -1466
rect 7543 -1642 7577 -1466
rect 7661 -1642 7695 -1466
rect 7779 -1642 7813 -1466
rect 8567 -1646 8601 -1470
rect 8685 -1646 8719 -1470
rect 8803 -1646 8837 -1470
rect 8921 -1646 8955 -1470
rect 15294 -1058 15328 -682
rect 15412 -1058 15446 -682
rect 15530 -1058 15564 -682
rect 15648 -1058 15682 -682
rect 15766 -1058 15800 -682
rect 15884 -1058 15918 -682
rect 17147 -930 17181 -754
rect 17265 -930 17299 -754
rect 17383 -930 17417 -754
rect 17501 -930 17535 -754
rect 17619 -930 17653 -754
rect 17737 -930 17771 -754
rect 17855 -930 17889 -754
rect 17973 -930 18007 -754
rect 18091 -930 18125 -754
rect 18209 -930 18243 -754
rect 20547 -1051 20581 -675
rect 20665 -1051 20699 -675
rect 20783 -1051 20817 -675
rect 20901 -1051 20935 -675
rect 21019 -1051 21053 -675
rect 21137 -1051 21171 -675
rect 21255 -1051 21289 -675
rect 21689 -1055 21723 -679
rect 13959 -1637 13993 -1461
rect 14077 -1637 14111 -1461
rect 14195 -1637 14229 -1461
rect 14313 -1637 14347 -1461
rect 15101 -1641 15135 -1465
rect 15219 -1641 15253 -1465
rect 15337 -1641 15371 -1465
rect 15455 -1641 15489 -1465
rect 21807 -1055 21841 -679
rect 21925 -1055 21959 -679
rect 22043 -1055 22077 -679
rect 22161 -1055 22195 -679
rect 22279 -1055 22313 -679
rect 22397 -1055 22431 -679
rect 23660 -927 23694 -751
rect 23778 -927 23812 -751
rect 23896 -927 23930 -751
rect 24014 -927 24048 -751
rect 24132 -927 24166 -751
rect 24250 -927 24284 -751
rect 24368 -927 24402 -751
rect 24486 -927 24520 -751
rect 24604 -927 24638 -751
rect 24722 -927 24756 -751
rect 20472 -1634 20506 -1458
rect 20590 -1634 20624 -1458
rect 20708 -1634 20742 -1458
rect 20826 -1634 20860 -1458
rect 21614 -1638 21648 -1462
rect 21732 -1638 21766 -1462
rect 21850 -1638 21884 -1462
rect 21968 -1638 22002 -1462
rect 4041 -2581 4075 -2405
rect 4159 -2581 4193 -2405
rect 4277 -2581 4311 -2405
rect 4395 -2581 4429 -2405
rect 4513 -2581 4547 -2405
rect 4631 -2581 4665 -2405
rect 4749 -2581 4783 -2405
rect 4867 -2581 4901 -2405
rect 4985 -2581 5019 -2405
rect 5103 -2581 5137 -2405
rect 10599 -2585 10633 -2409
rect 10717 -2585 10751 -2409
rect 10835 -2585 10869 -2409
rect 10953 -2585 10987 -2409
rect 11071 -2585 11105 -2409
rect 11189 -2585 11223 -2409
rect 11307 -2585 11341 -2409
rect 11425 -2585 11459 -2409
rect 11543 -2585 11577 -2409
rect 11661 -2585 11695 -2409
rect 17133 -2580 17167 -2404
rect 17251 -2580 17285 -2404
rect 17369 -2580 17403 -2404
rect 17487 -2580 17521 -2404
rect 17605 -2580 17639 -2404
rect 17723 -2580 17757 -2404
rect 17841 -2580 17875 -2404
rect 17959 -2580 17993 -2404
rect 18077 -2580 18111 -2404
rect 18195 -2580 18229 -2404
rect 23646 -2577 23680 -2401
rect 23764 -2577 23798 -2401
rect 23882 -2577 23916 -2401
rect 24000 -2577 24034 -2401
rect 24118 -2577 24152 -2401
rect 24236 -2577 24270 -2401
rect 24354 -2577 24388 -2401
rect 24472 -2577 24506 -2401
rect 24590 -2577 24624 -2401
rect 24708 -2577 24742 -2401
rect 66 -3198 100 -3022
rect 184 -3198 218 -3022
rect 302 -3198 336 -3022
rect 420 -3198 454 -3022
rect 549 -3198 583 -2822
rect 667 -3198 701 -2822
rect 785 -3198 819 -2822
rect 903 -3198 937 -2822
rect 1021 -3198 1055 -2822
rect 1139 -3198 1173 -2822
rect 1257 -3198 1291 -2822
rect 1387 -3198 1421 -3022
rect 1505 -3198 1539 -3022
rect 1623 -3198 1657 -3022
rect 1741 -3198 1775 -3022
rect 1964 -3198 1998 -3022
rect 2082 -3198 2116 -3022
rect 2200 -3198 2234 -3022
rect 2318 -3198 2352 -3022
rect 2447 -3198 2481 -2822
rect 2565 -3198 2599 -2822
rect 2683 -3198 2717 -2822
rect 2801 -3198 2835 -2822
rect 2919 -3198 2953 -2822
rect 3037 -3198 3071 -2822
rect 3155 -3198 3189 -2822
rect 3285 -3198 3319 -3022
rect 3403 -3198 3437 -3022
rect 3521 -3198 3555 -3022
rect 3639 -3198 3673 -3022
rect 606 -3891 640 -3515
rect 724 -3891 758 -3515
rect 842 -3891 876 -3515
rect 960 -3891 994 -3515
rect 1078 -3891 1112 -3515
rect 1196 -3891 1230 -3515
rect 1314 -3891 1348 -3515
rect 6624 -3202 6658 -3026
rect 6742 -3202 6776 -3026
rect 6860 -3202 6894 -3026
rect 6978 -3202 7012 -3026
rect 7107 -3202 7141 -2826
rect 7225 -3202 7259 -2826
rect 7343 -3202 7377 -2826
rect 7461 -3202 7495 -2826
rect 7579 -3202 7613 -2826
rect 7697 -3202 7731 -2826
rect 7815 -3202 7849 -2826
rect 7945 -3202 7979 -3026
rect 8063 -3202 8097 -3026
rect 8181 -3202 8215 -3026
rect 8299 -3202 8333 -3026
rect 8522 -3202 8556 -3026
rect 8640 -3202 8674 -3026
rect 8758 -3202 8792 -3026
rect 8876 -3202 8910 -3026
rect 9005 -3202 9039 -2826
rect 9123 -3202 9157 -2826
rect 9241 -3202 9275 -2826
rect 9359 -3202 9393 -2826
rect 9477 -3202 9511 -2826
rect 9595 -3202 9629 -2826
rect 9713 -3202 9747 -2826
rect 9843 -3202 9877 -3026
rect 9961 -3202 9995 -3026
rect 10079 -3202 10113 -3026
rect 10197 -3202 10231 -3026
rect 2504 -3891 2538 -3515
rect 2622 -3891 2656 -3515
rect 2740 -3891 2774 -3515
rect 2858 -3891 2892 -3515
rect 2976 -3891 3010 -3515
rect 3094 -3891 3128 -3515
rect 3212 -3891 3246 -3515
rect 4046 -4185 4080 -4009
rect 4164 -4185 4198 -4009
rect 4282 -4185 4316 -4009
rect 4400 -4185 4434 -4009
rect 4518 -4185 4552 -4009
rect 4636 -4185 4670 -4009
rect 4754 -4185 4788 -4009
rect 4872 -4185 4906 -4009
rect 4990 -4185 5024 -4009
rect 5108 -4185 5142 -4009
rect 7164 -3895 7198 -3519
rect 7282 -3895 7316 -3519
rect 7400 -3895 7434 -3519
rect 7518 -3895 7552 -3519
rect 7636 -3895 7670 -3519
rect 7754 -3895 7788 -3519
rect 7872 -3895 7906 -3519
rect 13158 -3197 13192 -3021
rect 13276 -3197 13310 -3021
rect 13394 -3197 13428 -3021
rect 13512 -3197 13546 -3021
rect 13641 -3197 13675 -2821
rect 13759 -3197 13793 -2821
rect 13877 -3197 13911 -2821
rect 13995 -3197 14029 -2821
rect 14113 -3197 14147 -2821
rect 14231 -3197 14265 -2821
rect 14349 -3197 14383 -2821
rect 14479 -3197 14513 -3021
rect 14597 -3197 14631 -3021
rect 14715 -3197 14749 -3021
rect 14833 -3197 14867 -3021
rect 15056 -3197 15090 -3021
rect 15174 -3197 15208 -3021
rect 15292 -3197 15326 -3021
rect 15410 -3197 15444 -3021
rect 15539 -3197 15573 -2821
rect 15657 -3197 15691 -2821
rect 15775 -3197 15809 -2821
rect 15893 -3197 15927 -2821
rect 16011 -3197 16045 -2821
rect 16129 -3197 16163 -2821
rect 16247 -3197 16281 -2821
rect 16377 -3197 16411 -3021
rect 16495 -3197 16529 -3021
rect 16613 -3197 16647 -3021
rect 16731 -3197 16765 -3021
rect 9062 -3895 9096 -3519
rect 9180 -3895 9214 -3519
rect 9298 -3895 9332 -3519
rect 9416 -3895 9450 -3519
rect 9534 -3895 9568 -3519
rect 9652 -3895 9686 -3519
rect 9770 -3895 9804 -3519
rect 10604 -4189 10638 -4013
rect 10722 -4189 10756 -4013
rect 10840 -4189 10874 -4013
rect 10958 -4189 10992 -4013
rect 11076 -4189 11110 -4013
rect 11194 -4189 11228 -4013
rect 11312 -4189 11346 -4013
rect 11430 -4189 11464 -4013
rect 11548 -4189 11582 -4013
rect 11666 -4189 11700 -4013
rect 13698 -3890 13732 -3514
rect 13816 -3890 13850 -3514
rect 13934 -3890 13968 -3514
rect 14052 -3890 14086 -3514
rect 14170 -3890 14204 -3514
rect 14288 -3890 14322 -3514
rect 14406 -3890 14440 -3514
rect 19671 -3194 19705 -3018
rect 19789 -3194 19823 -3018
rect 19907 -3194 19941 -3018
rect 20025 -3194 20059 -3018
rect 20154 -3194 20188 -2818
rect 20272 -3194 20306 -2818
rect 20390 -3194 20424 -2818
rect 20508 -3194 20542 -2818
rect 20626 -3194 20660 -2818
rect 20744 -3194 20778 -2818
rect 20862 -3194 20896 -2818
rect 20992 -3194 21026 -3018
rect 21110 -3194 21144 -3018
rect 21228 -3194 21262 -3018
rect 21346 -3194 21380 -3018
rect 21569 -3194 21603 -3018
rect 21687 -3194 21721 -3018
rect 21805 -3194 21839 -3018
rect 21923 -3194 21957 -3018
rect 22052 -3194 22086 -2818
rect 22170 -3194 22204 -2818
rect 22288 -3194 22322 -2818
rect 22406 -3194 22440 -2818
rect 22524 -3194 22558 -2818
rect 22642 -3194 22676 -2818
rect 22760 -3194 22794 -2818
rect 22890 -3194 22924 -3018
rect 23008 -3194 23042 -3018
rect 23126 -3194 23160 -3018
rect 23244 -3194 23278 -3018
rect 15596 -3890 15630 -3514
rect 15714 -3890 15748 -3514
rect 15832 -3890 15866 -3514
rect 15950 -3890 15984 -3514
rect 16068 -3890 16102 -3514
rect 16186 -3890 16220 -3514
rect 16304 -3890 16338 -3514
rect 17138 -4184 17172 -4008
rect 17256 -4184 17290 -4008
rect 17374 -4184 17408 -4008
rect 17492 -4184 17526 -4008
rect 17610 -4184 17644 -4008
rect 17728 -4184 17762 -4008
rect 17846 -4184 17880 -4008
rect 17964 -4184 17998 -4008
rect 18082 -4184 18116 -4008
rect 18200 -4184 18234 -4008
rect 20211 -3887 20245 -3511
rect 20329 -3887 20363 -3511
rect 20447 -3887 20481 -3511
rect 20565 -3887 20599 -3511
rect 20683 -3887 20717 -3511
rect 20801 -3887 20835 -3511
rect 20919 -3887 20953 -3511
rect 22109 -3887 22143 -3511
rect 22227 -3887 22261 -3511
rect 22345 -3887 22379 -3511
rect 22463 -3887 22497 -3511
rect 22581 -3887 22615 -3511
rect 22699 -3887 22733 -3511
rect 22817 -3887 22851 -3511
rect 23651 -4181 23685 -4005
rect 23769 -4181 23803 -4005
rect 23887 -4181 23921 -4005
rect 24005 -4181 24039 -4005
rect 24123 -4181 24157 -4005
rect 24241 -4181 24275 -4005
rect 24359 -4181 24393 -4005
rect 24477 -4181 24511 -4005
rect 24595 -4181 24629 -4005
rect 24713 -4181 24747 -4005
<< psubdiff >>
rect 1692 4090 1926 4124
rect 1692 4000 1738 4090
rect 1901 4000 1926 4090
rect 1692 3969 1926 4000
rect 8205 4087 8439 4121
rect 8205 3997 8251 4087
rect 8414 3997 8439 4087
rect 8205 3966 8439 3997
rect 14739 4082 14973 4116
rect 14739 3992 14785 4082
rect 14948 3992 14973 4082
rect 14739 3961 14973 3992
rect 21297 4086 21531 4120
rect 21297 3996 21343 4086
rect 21506 3996 21531 4086
rect 21297 3965 21531 3996
rect 3189 3719 3344 3765
rect 3189 3556 3220 3719
rect 3310 3556 3344 3719
rect 3189 3531 3344 3556
rect 4331 3717 4486 3763
rect 4331 3554 4362 3717
rect 4452 3554 4486 3717
rect 9702 3716 9857 3762
rect 4331 3529 4486 3554
rect 9702 3553 9733 3716
rect 9823 3553 9857 3716
rect 9702 3528 9857 3553
rect 10844 3714 10999 3760
rect 10844 3551 10875 3714
rect 10965 3551 10999 3714
rect 16236 3711 16391 3757
rect 10844 3526 10999 3551
rect 16236 3548 16267 3711
rect 16357 3548 16391 3711
rect 16236 3523 16391 3548
rect 17378 3709 17533 3755
rect 17378 3546 17409 3709
rect 17499 3546 17533 3709
rect 22794 3715 22949 3761
rect 17378 3521 17533 3546
rect 22794 3552 22825 3715
rect 22915 3552 22949 3715
rect 22794 3527 22949 3552
rect 23936 3713 24091 3759
rect 23936 3550 23967 3713
rect 24057 3550 24091 3713
rect 23936 3525 24091 3550
rect 1706 2440 1940 2474
rect 1706 2350 1752 2440
rect 1915 2350 1940 2440
rect 1706 2319 1940 2350
rect 8219 2437 8453 2471
rect 8219 2347 8265 2437
rect 8428 2347 8453 2437
rect 8219 2316 8453 2347
rect 14753 2432 14987 2466
rect 14753 2342 14799 2432
rect 14962 2342 14987 2432
rect 14753 2311 14987 2342
rect 1701 836 1935 870
rect 1701 746 1747 836
rect 1910 746 1935 836
rect 21311 2436 21545 2470
rect 21311 2346 21357 2436
rect 21520 2346 21545 2436
rect 21311 2315 21545 2346
rect 8214 833 8448 867
rect 1701 715 1935 746
rect 3133 676 3288 722
rect 8214 743 8260 833
rect 8423 743 8448 833
rect 14748 828 14982 862
rect 8214 712 8448 743
rect 3133 513 3164 676
rect 3254 513 3288 676
rect 3133 488 3288 513
rect 9646 673 9801 719
rect 14748 738 14794 828
rect 14957 738 14982 828
rect 21306 832 21540 866
rect 14748 707 14982 738
rect 9646 510 9677 673
rect 9767 510 9801 673
rect 9646 485 9801 510
rect 16180 668 16335 714
rect 21306 742 21352 832
rect 21515 742 21540 832
rect 21306 711 21540 742
rect 16180 505 16211 668
rect 16301 505 16335 668
rect 16180 480 16335 505
rect 22738 672 22893 718
rect 22738 509 22769 672
rect 22859 509 22893 672
rect 22738 484 22893 509
rect 4156 -1518 4390 -1484
rect 4156 -1608 4181 -1518
rect 4344 -1608 4390 -1518
rect 4156 -1639 4390 -1608
rect 10714 -1522 10948 -1488
rect 10714 -1612 10739 -1522
rect 10902 -1612 10948 -1522
rect 10714 -1643 10948 -1612
rect 17248 -1517 17482 -1483
rect 17248 -1607 17273 -1517
rect 17436 -1607 17482 -1517
rect 17248 -1638 17482 -1607
rect 23761 -1514 23995 -1480
rect 23761 -1604 23786 -1514
rect 23949 -1604 23995 -1514
rect 23761 -1635 23995 -1604
rect 1596 -1891 1751 -1845
rect 1596 -2054 1630 -1891
rect 1720 -2054 1751 -1891
rect 1596 -2079 1751 -2054
rect 2738 -1889 2893 -1843
rect 2738 -2052 2772 -1889
rect 2862 -2052 2893 -1889
rect 8154 -1895 8309 -1849
rect 2738 -2077 2893 -2052
rect 8154 -2058 8188 -1895
rect 8278 -2058 8309 -1895
rect 8154 -2083 8309 -2058
rect 9296 -1893 9451 -1847
rect 9296 -2056 9330 -1893
rect 9420 -2056 9451 -1893
rect 14688 -1890 14843 -1844
rect 9296 -2081 9451 -2056
rect 14688 -2053 14722 -1890
rect 14812 -2053 14843 -1890
rect 14688 -2078 14843 -2053
rect 15830 -1888 15985 -1842
rect 15830 -2051 15864 -1888
rect 15954 -2051 15985 -1888
rect 21201 -1887 21356 -1841
rect 15830 -2076 15985 -2051
rect 21201 -2050 21235 -1887
rect 21325 -2050 21356 -1887
rect 21201 -2075 21356 -2050
rect 22343 -1885 22498 -1839
rect 22343 -2048 22377 -1885
rect 22467 -2048 22498 -1885
rect 22343 -2073 22498 -2048
rect 4142 -3168 4376 -3134
rect 4142 -3258 4167 -3168
rect 4330 -3258 4376 -3168
rect 10700 -3172 10934 -3138
rect 4142 -3289 4376 -3258
rect 10700 -3262 10725 -3172
rect 10888 -3262 10934 -3172
rect 17234 -3167 17468 -3133
rect 10700 -3293 10934 -3262
rect 4147 -4772 4381 -4738
rect 4147 -4862 4172 -4772
rect 4335 -4862 4381 -4772
rect 17234 -3257 17259 -3167
rect 17422 -3257 17468 -3167
rect 23747 -3164 23981 -3130
rect 17234 -3288 17468 -3257
rect 10705 -4776 10939 -4742
rect 2794 -4932 2949 -4886
rect 4147 -4893 4381 -4862
rect 10705 -4866 10730 -4776
rect 10893 -4866 10939 -4776
rect 23747 -3254 23772 -3164
rect 23935 -3254 23981 -3164
rect 23747 -3285 23981 -3254
rect 17239 -4771 17473 -4737
rect 2794 -5095 2828 -4932
rect 2918 -5095 2949 -4932
rect 2794 -5120 2949 -5095
rect 9352 -4936 9507 -4890
rect 10705 -4897 10939 -4866
rect 17239 -4861 17264 -4771
rect 17427 -4861 17473 -4771
rect 23752 -4768 23986 -4734
rect 9352 -5099 9386 -4936
rect 9476 -5099 9507 -4936
rect 9352 -5124 9507 -5099
rect 15886 -4931 16041 -4885
rect 17239 -4892 17473 -4861
rect 23752 -4858 23777 -4768
rect 23940 -4858 23986 -4768
rect 15886 -5094 15920 -4931
rect 16010 -5094 16041 -4931
rect 15886 -5119 16041 -5094
rect 22399 -4928 22554 -4882
rect 23752 -4889 23986 -4858
rect 22399 -5091 22433 -4928
rect 22523 -5091 22554 -4928
rect 22399 -5116 22554 -5091
<< nsubdiff >>
rect 3844 5321 3997 5361
rect 1362 5267 1515 5307
rect 1362 5118 1405 5267
rect 1472 5118 1515 5267
rect 1362 5049 1515 5118
rect 3844 5172 3887 5321
rect 3954 5172 3997 5321
rect 3844 5103 3997 5172
rect 4991 5321 5144 5361
rect 4991 5172 5034 5321
rect 5101 5172 5144 5321
rect 10357 5318 10510 5358
rect 4991 5103 5144 5172
rect 7875 5264 8028 5304
rect 7875 5115 7918 5264
rect 7985 5115 8028 5264
rect 7875 5046 8028 5115
rect 10357 5169 10400 5318
rect 10467 5169 10510 5318
rect 10357 5100 10510 5169
rect 11504 5318 11657 5358
rect 11504 5169 11547 5318
rect 11614 5169 11657 5318
rect 16891 5313 17044 5353
rect 11504 5100 11657 5169
rect 14409 5259 14562 5299
rect 14409 5110 14452 5259
rect 14519 5110 14562 5259
rect 14409 5041 14562 5110
rect 16891 5164 16934 5313
rect 17001 5164 17044 5313
rect 16891 5095 17044 5164
rect 18038 5313 18191 5353
rect 18038 5164 18081 5313
rect 18148 5164 18191 5313
rect 23449 5317 23602 5357
rect 18038 5095 18191 5164
rect 20967 5263 21120 5303
rect 20967 5114 21010 5263
rect 21077 5114 21120 5263
rect 20967 5045 21120 5114
rect 23449 5168 23492 5317
rect 23559 5168 23602 5317
rect 23449 5099 23602 5168
rect 24596 5317 24749 5357
rect 24596 5168 24639 5317
rect 24706 5168 24749 5317
rect 24596 5099 24749 5168
rect 1376 3617 1529 3657
rect 1376 3468 1419 3617
rect 1486 3468 1529 3617
rect 7889 3614 8042 3654
rect 1376 3399 1529 3468
rect 7889 3465 7932 3614
rect 7999 3465 8042 3614
rect 14423 3609 14576 3649
rect 7889 3396 8042 3465
rect 14423 3460 14466 3609
rect 14533 3460 14576 3609
rect 20981 3613 21134 3653
rect 14423 3391 14576 3460
rect 20981 3464 21024 3613
rect 21091 3464 21134 3613
rect 20981 3395 21134 3464
rect 5087 3274 5240 3314
rect 5087 3125 5130 3274
rect 5197 3125 5240 3274
rect 11600 3271 11753 3311
rect 5087 3056 5240 3125
rect 11600 3122 11643 3271
rect 11710 3122 11753 3271
rect 18134 3266 18287 3306
rect 24692 3270 24845 3310
rect 11600 3053 11753 3122
rect 18134 3117 18177 3266
rect 18244 3117 18287 3266
rect 18134 3048 18287 3117
rect 24692 3121 24735 3270
rect 24802 3121 24845 3270
rect 24692 3052 24845 3121
rect 1371 2013 1524 2053
rect 1371 1864 1414 2013
rect 1481 1864 1524 2013
rect 1371 1795 1524 1864
rect 7884 2010 8037 2050
rect 7884 1861 7927 2010
rect 7994 1861 8037 2010
rect 7884 1792 8037 1861
rect 14418 2005 14571 2045
rect 14418 1856 14461 2005
rect 14528 1856 14571 2005
rect 14418 1787 14571 1856
rect 20976 2009 21129 2049
rect 20976 1860 21019 2009
rect 21086 1860 21129 2009
rect 20976 1791 21129 1860
rect 938 -287 1091 -247
rect 938 -436 981 -287
rect 1048 -436 1091 -287
rect 938 -505 1091 -436
rect 2085 -287 2238 -247
rect 2085 -436 2128 -287
rect 2195 -436 2238 -287
rect 7496 -291 7649 -251
rect 2085 -505 2238 -436
rect 4567 -341 4720 -301
rect 4567 -490 4610 -341
rect 4677 -490 4720 -341
rect 4567 -559 4720 -490
rect 7496 -440 7539 -291
rect 7606 -440 7649 -291
rect 7496 -509 7649 -440
rect 8643 -291 8796 -251
rect 8643 -440 8686 -291
rect 8753 -440 8796 -291
rect 14030 -286 14183 -246
rect 8643 -509 8796 -440
rect 11125 -345 11278 -305
rect 11125 -494 11168 -345
rect 11235 -494 11278 -345
rect 11125 -563 11278 -494
rect 14030 -435 14073 -286
rect 14140 -435 14183 -286
rect 14030 -504 14183 -435
rect 15177 -286 15330 -246
rect 15177 -435 15220 -286
rect 15287 -435 15330 -286
rect 20543 -283 20696 -243
rect 15177 -504 15330 -435
rect 17659 -340 17812 -300
rect 17659 -489 17702 -340
rect 17769 -489 17812 -340
rect 17659 -558 17812 -489
rect 20543 -432 20586 -283
rect 20653 -432 20696 -283
rect 20543 -501 20696 -432
rect 21690 -283 21843 -243
rect 21690 -432 21733 -283
rect 21800 -432 21843 -283
rect 21690 -501 21843 -432
rect 24172 -337 24325 -297
rect 24172 -486 24215 -337
rect 24282 -486 24325 -337
rect 24172 -555 24325 -486
rect 4553 -1991 4706 -1951
rect 4553 -2140 4596 -1991
rect 4663 -2140 4706 -1991
rect 11111 -1995 11264 -1955
rect 4553 -2209 4706 -2140
rect 11111 -2144 11154 -1995
rect 11221 -2144 11264 -1995
rect 17645 -1990 17798 -1950
rect 11111 -2213 11264 -2144
rect 17645 -2139 17688 -1990
rect 17755 -2139 17798 -1990
rect 24158 -1987 24311 -1947
rect 17645 -2208 17798 -2139
rect 24158 -2136 24201 -1987
rect 24268 -2136 24311 -1987
rect 24158 -2205 24311 -2136
rect 842 -2334 995 -2294
rect 842 -2483 885 -2334
rect 952 -2483 995 -2334
rect 7400 -2338 7553 -2298
rect 842 -2552 995 -2483
rect 7400 -2487 7443 -2338
rect 7510 -2487 7553 -2338
rect 13934 -2333 14087 -2293
rect 7400 -2556 7553 -2487
rect 13934 -2482 13977 -2333
rect 14044 -2482 14087 -2333
rect 20447 -2330 20600 -2290
rect 13934 -2551 14087 -2482
rect 20447 -2479 20490 -2330
rect 20557 -2479 20600 -2330
rect 20447 -2548 20600 -2479
rect 4558 -3595 4711 -3555
rect 4558 -3744 4601 -3595
rect 4668 -3744 4711 -3595
rect 4558 -3813 4711 -3744
rect 11116 -3599 11269 -3559
rect 11116 -3748 11159 -3599
rect 11226 -3748 11269 -3599
rect 11116 -3817 11269 -3748
rect 17650 -3594 17803 -3554
rect 17650 -3743 17693 -3594
rect 17760 -3743 17803 -3594
rect 17650 -3812 17803 -3743
rect 24163 -3591 24316 -3551
rect 24163 -3740 24206 -3591
rect 24273 -3740 24316 -3591
rect 24163 -3809 24316 -3740
<< psubdiffcont >>
rect 1738 4000 1901 4090
rect 8251 3997 8414 4087
rect 14785 3992 14948 4082
rect 21343 3996 21506 4086
rect 3220 3556 3310 3719
rect 4362 3554 4452 3717
rect 9733 3553 9823 3716
rect 10875 3551 10965 3714
rect 16267 3548 16357 3711
rect 17409 3546 17499 3709
rect 22825 3552 22915 3715
rect 23967 3550 24057 3713
rect 1752 2350 1915 2440
rect 8265 2347 8428 2437
rect 14799 2342 14962 2432
rect 1747 746 1910 836
rect 21357 2346 21520 2436
rect 8260 743 8423 833
rect 3164 513 3254 676
rect 14794 738 14957 828
rect 9677 510 9767 673
rect 21352 742 21515 832
rect 16211 505 16301 668
rect 22769 509 22859 672
rect 4181 -1608 4344 -1518
rect 10739 -1612 10902 -1522
rect 17273 -1607 17436 -1517
rect 23786 -1604 23949 -1514
rect 1630 -2054 1720 -1891
rect 2772 -2052 2862 -1889
rect 8188 -2058 8278 -1895
rect 9330 -2056 9420 -1893
rect 14722 -2053 14812 -1890
rect 15864 -2051 15954 -1888
rect 21235 -2050 21325 -1887
rect 22377 -2048 22467 -1885
rect 4167 -3258 4330 -3168
rect 10725 -3262 10888 -3172
rect 4172 -4862 4335 -4772
rect 17259 -3257 17422 -3167
rect 10730 -4866 10893 -4776
rect 23772 -3254 23935 -3164
rect 2828 -5095 2918 -4932
rect 17264 -4861 17427 -4771
rect 9386 -5099 9476 -4936
rect 23777 -4858 23940 -4768
rect 15920 -5094 16010 -4931
rect 22433 -5091 22523 -4928
<< nsubdiffcont >>
rect 1405 5118 1472 5267
rect 3887 5172 3954 5321
rect 5034 5172 5101 5321
rect 7918 5115 7985 5264
rect 10400 5169 10467 5318
rect 11547 5169 11614 5318
rect 14452 5110 14519 5259
rect 16934 5164 17001 5313
rect 18081 5164 18148 5313
rect 21010 5114 21077 5263
rect 23492 5168 23559 5317
rect 24639 5168 24706 5317
rect 1419 3468 1486 3617
rect 7932 3465 7999 3614
rect 14466 3460 14533 3609
rect 21024 3464 21091 3613
rect 5130 3125 5197 3274
rect 11643 3122 11710 3271
rect 18177 3117 18244 3266
rect 24735 3121 24802 3270
rect 1414 1864 1481 2013
rect 7927 1861 7994 2010
rect 14461 1856 14528 2005
rect 21019 1860 21086 2009
rect 981 -436 1048 -287
rect 2128 -436 2195 -287
rect 4610 -490 4677 -341
rect 7539 -440 7606 -291
rect 8686 -440 8753 -291
rect 11168 -494 11235 -345
rect 14073 -435 14140 -286
rect 15220 -435 15287 -286
rect 17702 -489 17769 -340
rect 20586 -432 20653 -283
rect 21733 -432 21800 -283
rect 24215 -486 24282 -337
rect 4596 -2140 4663 -1991
rect 11154 -2144 11221 -1995
rect 17688 -2139 17755 -1990
rect 24201 -2136 24268 -1987
rect 885 -2483 952 -2334
rect 7443 -2487 7510 -2338
rect 13977 -2482 14044 -2333
rect 20490 -2479 20557 -2330
rect 4601 -3744 4668 -3595
rect 11159 -3748 11226 -3599
rect 17693 -3743 17760 -3594
rect 24206 -3740 24273 -3591
<< poly >>
rect 3125 5101 3191 5117
rect 4255 5107 4321 5123
rect 3125 5067 3141 5101
rect 3175 5094 3191 5101
rect 3175 5067 3700 5094
rect 3125 5051 3700 5067
rect 4255 5073 4271 5107
rect 4305 5098 4321 5107
rect 4305 5073 4842 5098
rect 4255 5055 4842 5073
rect 3656 4999 3700 5051
rect 4798 5003 4842 5055
rect 9638 5098 9704 5114
rect 10768 5104 10834 5120
rect 9638 5064 9654 5098
rect 9688 5091 9704 5098
rect 9688 5064 10213 5091
rect 9638 5048 10213 5064
rect 10768 5070 10784 5104
rect 10818 5095 10834 5104
rect 10818 5070 11355 5095
rect 10768 5052 11355 5070
rect 3125 4983 3598 4999
rect 3125 4949 3141 4983
rect 3175 4958 3598 4983
rect 3175 4957 3362 4958
rect 3175 4949 3191 4957
rect 3125 4933 3191 4949
rect 3302 4937 3362 4957
rect 3420 4937 3480 4958
rect 3538 4937 3598 4958
rect 3656 4958 3952 4999
rect 3656 4937 3716 4958
rect 3774 4937 3834 4958
rect 3892 4937 3952 4958
rect 4255 4987 4740 5003
rect 4255 4953 4271 4987
rect 4305 4962 4740 4987
rect 4305 4961 4504 4962
rect 4305 4953 4321 4961
rect 4255 4937 4321 4953
rect 4444 4941 4504 4961
rect 4562 4941 4622 4962
rect 4680 4941 4740 4962
rect 4798 4962 5094 5003
rect 10169 4996 10213 5048
rect 11311 5000 11355 5052
rect 16172 5093 16238 5109
rect 17302 5099 17368 5115
rect 16172 5059 16188 5093
rect 16222 5086 16238 5093
rect 16222 5059 16747 5086
rect 16172 5043 16747 5059
rect 17302 5065 17318 5099
rect 17352 5090 17368 5099
rect 17352 5065 17889 5090
rect 17302 5047 17889 5065
rect 4798 4941 4858 4962
rect 4916 4941 4976 4962
rect 5034 4941 5094 4962
rect 9638 4980 10111 4996
rect 9638 4946 9654 4980
rect 9688 4955 10111 4980
rect 9688 4954 9875 4955
rect 9688 4946 9704 4954
rect 977 4886 1273 4922
rect 977 4865 1037 4886
rect 1095 4865 1155 4886
rect 1213 4865 1273 4886
rect 1331 4885 1627 4921
rect 1331 4865 1391 4885
rect 1449 4865 1509 4885
rect 1567 4865 1627 4885
rect 1685 4885 1981 4921
rect 1685 4865 1745 4885
rect 1803 4865 1863 4885
rect 1921 4865 1981 4885
rect 977 4639 1037 4665
rect 1095 4639 1155 4665
rect 1213 4639 1273 4665
rect 1331 4645 1391 4665
rect 1331 4639 1392 4645
rect 1449 4639 1509 4665
rect 1567 4639 1627 4665
rect 1214 4454 1272 4639
rect 1214 4428 1274 4454
rect 1332 4428 1392 4639
rect 1685 4633 1745 4665
rect 1803 4639 1863 4665
rect 1921 4639 1981 4665
rect 1682 4617 1748 4633
rect 1682 4583 1698 4617
rect 1732 4583 1748 4617
rect 1682 4567 1748 4583
rect 9638 4930 9704 4946
rect 9815 4934 9875 4954
rect 9933 4934 9993 4955
rect 10051 4934 10111 4955
rect 10169 4955 10465 4996
rect 10169 4934 10229 4955
rect 10287 4934 10347 4955
rect 10405 4934 10465 4955
rect 10768 4984 11253 5000
rect 10768 4950 10784 4984
rect 10818 4959 11253 4984
rect 10818 4958 11017 4959
rect 10818 4950 10834 4958
rect 10768 4934 10834 4950
rect 10957 4938 11017 4958
rect 11075 4938 11135 4959
rect 11193 4938 11253 4959
rect 11311 4959 11607 5000
rect 16703 4991 16747 5043
rect 17845 4995 17889 5047
rect 22730 5097 22796 5113
rect 23860 5103 23926 5119
rect 22730 5063 22746 5097
rect 22780 5090 22796 5097
rect 22780 5063 23305 5090
rect 22730 5047 23305 5063
rect 23860 5069 23876 5103
rect 23910 5094 23926 5103
rect 23910 5069 24447 5094
rect 23860 5051 24447 5069
rect 23261 4995 23305 5047
rect 24403 4999 24447 5051
rect 11311 4938 11371 4959
rect 11429 4938 11489 4959
rect 11547 4938 11607 4959
rect 16172 4975 16645 4991
rect 16172 4941 16188 4975
rect 16222 4950 16645 4975
rect 16222 4949 16409 4950
rect 16222 4941 16238 4949
rect 7490 4883 7786 4919
rect 7490 4862 7550 4883
rect 7608 4862 7668 4883
rect 7726 4862 7786 4883
rect 7844 4882 8140 4918
rect 7844 4862 7904 4882
rect 7962 4862 8022 4882
rect 8080 4862 8140 4882
rect 8198 4882 8494 4918
rect 8198 4862 8258 4882
rect 8316 4862 8376 4882
rect 8434 4862 8494 4882
rect 7490 4636 7550 4662
rect 7608 4636 7668 4662
rect 7726 4636 7786 4662
rect 7844 4642 7904 4662
rect 7844 4636 7905 4642
rect 7962 4636 8022 4662
rect 8080 4636 8140 4662
rect 3302 4520 3362 4537
rect 1564 4500 1630 4516
rect 1564 4466 1580 4500
rect 1614 4466 1630 4500
rect 1564 4450 1630 4466
rect 1567 4428 1627 4450
rect 3302 4431 3363 4520
rect 3420 4511 3480 4537
rect 3538 4511 3598 4537
rect 3212 4378 3363 4431
rect 1567 4202 1627 4228
rect 3212 4154 3272 4378
rect 3656 4336 3716 4537
rect 3774 4511 3834 4537
rect 3892 4511 3952 4537
rect 4444 4524 4504 4541
rect 4444 4435 4505 4524
rect 4562 4515 4622 4541
rect 4680 4515 4740 4541
rect 3330 4285 3716 4336
rect 4354 4382 4505 4435
rect 3330 4154 3390 4285
rect 3445 4227 3511 4243
rect 3445 4193 3461 4227
rect 3495 4193 3511 4227
rect 3445 4177 3511 4193
rect 3448 4154 3508 4177
rect 3731 4154 3791 4180
rect 3849 4154 3909 4180
rect 3967 4154 4027 4180
rect 4354 4158 4414 4382
rect 4798 4340 4858 4541
rect 4916 4515 4976 4541
rect 5034 4515 5094 4541
rect 7727 4451 7785 4636
rect 7727 4425 7787 4451
rect 7845 4425 7905 4636
rect 8198 4630 8258 4662
rect 8316 4636 8376 4662
rect 8434 4636 8494 4662
rect 8195 4614 8261 4630
rect 8195 4580 8211 4614
rect 8245 4580 8261 4614
rect 8195 4564 8261 4580
rect 16172 4925 16238 4941
rect 16349 4929 16409 4949
rect 16467 4929 16527 4950
rect 16585 4929 16645 4950
rect 16703 4950 16999 4991
rect 16703 4929 16763 4950
rect 16821 4929 16881 4950
rect 16939 4929 16999 4950
rect 17302 4979 17787 4995
rect 17302 4945 17318 4979
rect 17352 4954 17787 4979
rect 17352 4953 17551 4954
rect 17352 4945 17368 4953
rect 17302 4929 17368 4945
rect 17491 4933 17551 4953
rect 17609 4933 17669 4954
rect 17727 4933 17787 4954
rect 17845 4954 18141 4995
rect 17845 4933 17905 4954
rect 17963 4933 18023 4954
rect 18081 4933 18141 4954
rect 22730 4979 23203 4995
rect 22730 4945 22746 4979
rect 22780 4954 23203 4979
rect 22780 4953 22967 4954
rect 22780 4945 22796 4953
rect 14024 4878 14320 4914
rect 14024 4857 14084 4878
rect 14142 4857 14202 4878
rect 14260 4857 14320 4878
rect 14378 4877 14674 4913
rect 14378 4857 14438 4877
rect 14496 4857 14556 4877
rect 14614 4857 14674 4877
rect 14732 4877 15028 4913
rect 14732 4857 14792 4877
rect 14850 4857 14910 4877
rect 14968 4857 15028 4877
rect 14024 4631 14084 4657
rect 14142 4631 14202 4657
rect 14260 4631 14320 4657
rect 14378 4637 14438 4657
rect 14378 4631 14439 4637
rect 14496 4631 14556 4657
rect 14614 4631 14674 4657
rect 9815 4517 9875 4534
rect 8077 4497 8143 4513
rect 8077 4463 8093 4497
rect 8127 4463 8143 4497
rect 8077 4447 8143 4463
rect 8080 4425 8140 4447
rect 9815 4428 9876 4517
rect 9933 4508 9993 4534
rect 10051 4508 10111 4534
rect 4472 4289 4858 4340
rect 4472 4158 4532 4289
rect 4587 4231 4653 4247
rect 4587 4197 4603 4231
rect 4637 4197 4653 4231
rect 4587 4181 4653 4197
rect 4590 4158 4650 4181
rect 4873 4158 4933 4184
rect 4991 4158 5051 4184
rect 5109 4158 5169 4184
rect 1214 4006 1274 4028
rect 1332 4006 1392 4028
rect 1211 3990 1277 4006
rect 1211 3956 1227 3990
rect 1261 3956 1277 3990
rect 1211 3940 1277 3956
rect 1329 3990 1395 4006
rect 1329 3956 1345 3990
rect 1379 3956 1395 3990
rect 1329 3940 1395 3956
rect 9725 4375 9876 4428
rect 8080 4199 8140 4225
rect 9725 4151 9785 4375
rect 10169 4333 10229 4534
rect 10287 4508 10347 4534
rect 10405 4508 10465 4534
rect 10957 4521 11017 4538
rect 10957 4432 11018 4521
rect 11075 4512 11135 4538
rect 11193 4512 11253 4538
rect 9843 4282 10229 4333
rect 10867 4379 11018 4432
rect 9843 4151 9903 4282
rect 9958 4224 10024 4240
rect 9958 4190 9974 4224
rect 10008 4190 10024 4224
rect 9958 4174 10024 4190
rect 9961 4151 10021 4174
rect 10244 4151 10304 4177
rect 10362 4151 10422 4177
rect 10480 4151 10540 4177
rect 10867 4155 10927 4379
rect 11311 4337 11371 4538
rect 11429 4512 11489 4538
rect 11547 4512 11607 4538
rect 14261 4446 14319 4631
rect 14261 4420 14321 4446
rect 14379 4420 14439 4631
rect 14732 4625 14792 4657
rect 14850 4631 14910 4657
rect 14968 4631 15028 4657
rect 14729 4609 14795 4625
rect 14729 4575 14745 4609
rect 14779 4575 14795 4609
rect 14729 4559 14795 4575
rect 22730 4929 22796 4945
rect 22907 4933 22967 4953
rect 23025 4933 23085 4954
rect 23143 4933 23203 4954
rect 23261 4954 23557 4995
rect 23261 4933 23321 4954
rect 23379 4933 23439 4954
rect 23497 4933 23557 4954
rect 23860 4983 24345 4999
rect 23860 4949 23876 4983
rect 23910 4958 24345 4983
rect 23910 4957 24109 4958
rect 23910 4949 23926 4957
rect 23860 4933 23926 4949
rect 24049 4937 24109 4957
rect 24167 4937 24227 4958
rect 24285 4937 24345 4958
rect 24403 4958 24699 4999
rect 24403 4937 24463 4958
rect 24521 4937 24581 4958
rect 24639 4937 24699 4958
rect 20582 4882 20878 4918
rect 20582 4861 20642 4882
rect 20700 4861 20760 4882
rect 20818 4861 20878 4882
rect 20936 4881 21232 4917
rect 20936 4861 20996 4881
rect 21054 4861 21114 4881
rect 21172 4861 21232 4881
rect 21290 4881 21586 4917
rect 21290 4861 21350 4881
rect 21408 4861 21468 4881
rect 21526 4861 21586 4881
rect 20582 4635 20642 4661
rect 20700 4635 20760 4661
rect 20818 4635 20878 4661
rect 20936 4641 20996 4661
rect 20936 4635 20997 4641
rect 21054 4635 21114 4661
rect 21172 4635 21232 4661
rect 16349 4512 16409 4529
rect 14611 4492 14677 4508
rect 14611 4458 14627 4492
rect 14661 4458 14677 4492
rect 14611 4442 14677 4458
rect 14614 4420 14674 4442
rect 16349 4423 16410 4512
rect 16467 4503 16527 4529
rect 16585 4503 16645 4529
rect 10985 4286 11371 4337
rect 10985 4155 11045 4286
rect 11100 4228 11166 4244
rect 11100 4194 11116 4228
rect 11150 4194 11166 4228
rect 11100 4178 11166 4194
rect 11103 4155 11163 4178
rect 11386 4155 11446 4181
rect 11504 4155 11564 4181
rect 11622 4155 11682 4181
rect 7727 4003 7787 4025
rect 7845 4003 7905 4025
rect 7724 3987 7790 4003
rect 3212 3928 3272 3954
rect 3330 3928 3390 3954
rect 3448 3922 3508 3954
rect 3731 3922 3791 3954
rect 3849 3922 3909 3954
rect 3967 3922 4027 3954
rect 4354 3932 4414 3958
rect 4472 3932 4532 3958
rect 3448 3881 4027 3922
rect 4590 3926 4650 3958
rect 4873 3926 4933 3958
rect 4991 3926 5051 3958
rect 5109 3926 5169 3958
rect 7724 3953 7740 3987
rect 7774 3953 7790 3987
rect 7724 3937 7790 3953
rect 7842 3987 7908 4003
rect 7842 3953 7858 3987
rect 7892 3953 7908 3987
rect 7842 3937 7908 3953
rect 16259 4370 16410 4423
rect 14614 4194 14674 4220
rect 16259 4146 16319 4370
rect 16703 4328 16763 4529
rect 16821 4503 16881 4529
rect 16939 4503 16999 4529
rect 17491 4516 17551 4533
rect 17491 4427 17552 4516
rect 17609 4507 17669 4533
rect 17727 4507 17787 4533
rect 16377 4277 16763 4328
rect 17401 4374 17552 4427
rect 16377 4146 16437 4277
rect 16492 4219 16558 4235
rect 16492 4185 16508 4219
rect 16542 4185 16558 4219
rect 16492 4169 16558 4185
rect 16495 4146 16555 4169
rect 16778 4146 16838 4172
rect 16896 4146 16956 4172
rect 17014 4146 17074 4172
rect 17401 4150 17461 4374
rect 17845 4332 17905 4533
rect 17963 4507 18023 4533
rect 18081 4507 18141 4533
rect 20819 4450 20877 4635
rect 20819 4424 20879 4450
rect 20937 4424 20997 4635
rect 21290 4629 21350 4661
rect 21408 4635 21468 4661
rect 21526 4635 21586 4661
rect 21287 4613 21353 4629
rect 21287 4579 21303 4613
rect 21337 4579 21353 4613
rect 21287 4563 21353 4579
rect 22907 4516 22967 4533
rect 21169 4496 21235 4512
rect 21169 4462 21185 4496
rect 21219 4462 21235 4496
rect 21169 4446 21235 4462
rect 21172 4424 21232 4446
rect 22907 4427 22968 4516
rect 23025 4507 23085 4533
rect 23143 4507 23203 4533
rect 17519 4281 17905 4332
rect 17519 4150 17579 4281
rect 17634 4223 17700 4239
rect 17634 4189 17650 4223
rect 17684 4189 17700 4223
rect 17634 4173 17700 4189
rect 17637 4150 17697 4173
rect 17920 4150 17980 4176
rect 18038 4150 18098 4176
rect 18156 4150 18216 4176
rect 14261 3998 14321 4020
rect 14379 3998 14439 4020
rect 14258 3982 14324 3998
rect 4590 3885 5169 3926
rect 9725 3925 9785 3951
rect 9843 3925 9903 3951
rect 9961 3919 10021 3951
rect 10244 3919 10304 3951
rect 10362 3919 10422 3951
rect 10480 3919 10540 3951
rect 10867 3929 10927 3955
rect 10985 3929 11045 3955
rect 9961 3878 10540 3919
rect 11103 3923 11163 3955
rect 11386 3923 11446 3955
rect 11504 3923 11564 3955
rect 11622 3923 11682 3955
rect 14258 3948 14274 3982
rect 14308 3948 14324 3982
rect 14258 3932 14324 3948
rect 14376 3982 14442 3998
rect 14376 3948 14392 3982
rect 14426 3948 14442 3982
rect 14376 3932 14442 3948
rect 22817 4374 22968 4427
rect 21172 4198 21232 4224
rect 22817 4150 22877 4374
rect 23261 4332 23321 4533
rect 23379 4507 23439 4533
rect 23497 4507 23557 4533
rect 24049 4520 24109 4537
rect 24049 4431 24110 4520
rect 24167 4511 24227 4537
rect 24285 4511 24345 4537
rect 22935 4281 23321 4332
rect 23959 4378 24110 4431
rect 22935 4150 22995 4281
rect 23050 4223 23116 4239
rect 23050 4189 23066 4223
rect 23100 4189 23116 4223
rect 23050 4173 23116 4189
rect 23053 4150 23113 4173
rect 23336 4150 23396 4176
rect 23454 4150 23514 4176
rect 23572 4150 23632 4176
rect 23959 4154 24019 4378
rect 24403 4336 24463 4537
rect 24521 4511 24581 4537
rect 24639 4511 24699 4537
rect 24077 4285 24463 4336
rect 24077 4154 24137 4285
rect 24192 4227 24258 4243
rect 24192 4193 24208 4227
rect 24242 4193 24258 4227
rect 24192 4177 24258 4193
rect 24195 4154 24255 4177
rect 24478 4154 24538 4180
rect 24596 4154 24656 4180
rect 24714 4154 24774 4180
rect 20819 4002 20879 4024
rect 20937 4002 20997 4024
rect 20816 3986 20882 4002
rect 20816 3952 20832 3986
rect 20866 3952 20882 3986
rect 11103 3882 11682 3923
rect 16259 3920 16319 3946
rect 16377 3920 16437 3946
rect 16495 3914 16555 3946
rect 16778 3914 16838 3946
rect 16896 3914 16956 3946
rect 17014 3914 17074 3946
rect 17401 3924 17461 3950
rect 17519 3924 17579 3950
rect 16495 3873 17074 3914
rect 17637 3918 17697 3950
rect 17920 3918 17980 3950
rect 18038 3918 18098 3950
rect 18156 3918 18216 3950
rect 20816 3936 20882 3952
rect 20934 3986 21000 4002
rect 20934 3952 20950 3986
rect 20984 3952 21000 3986
rect 20934 3936 21000 3952
rect 22817 3924 22877 3950
rect 22935 3924 22995 3950
rect 17637 3877 18216 3918
rect 23053 3918 23113 3950
rect 23336 3918 23396 3950
rect 23454 3918 23514 3950
rect 23572 3918 23632 3950
rect 23959 3928 24019 3954
rect 24077 3928 24137 3954
rect 23053 3877 23632 3918
rect 24195 3922 24255 3954
rect 24478 3922 24538 3954
rect 24596 3922 24656 3954
rect 24714 3922 24774 3954
rect 24195 3881 24774 3922
rect 991 3236 1287 3272
rect 991 3215 1051 3236
rect 1109 3215 1169 3236
rect 1227 3215 1287 3236
rect 1345 3235 1641 3271
rect 1345 3215 1405 3235
rect 1463 3215 1523 3235
rect 1581 3215 1641 3235
rect 1699 3235 1995 3271
rect 1699 3215 1759 3235
rect 1817 3215 1877 3235
rect 1935 3215 1995 3235
rect 7504 3233 7800 3269
rect 7504 3212 7564 3233
rect 7622 3212 7682 3233
rect 7740 3212 7800 3233
rect 7858 3232 8154 3268
rect 7858 3212 7918 3232
rect 7976 3212 8036 3232
rect 8094 3212 8154 3232
rect 8212 3232 8508 3268
rect 8212 3212 8272 3232
rect 8330 3212 8390 3232
rect 8448 3212 8508 3232
rect 991 2989 1051 3015
rect 1109 2989 1169 3015
rect 1227 2989 1287 3015
rect 1345 2995 1405 3015
rect 1345 2989 1406 2995
rect 1463 2989 1523 3015
rect 1581 2989 1641 3015
rect 1228 2804 1286 2989
rect 1228 2778 1288 2804
rect 1346 2778 1406 2989
rect 1699 2983 1759 3015
rect 1817 2989 1877 3015
rect 1935 2989 1995 3015
rect 14038 3228 14334 3264
rect 14038 3207 14098 3228
rect 14156 3207 14216 3228
rect 14274 3207 14334 3228
rect 14392 3227 14688 3263
rect 14392 3207 14452 3227
rect 14510 3207 14570 3227
rect 14628 3207 14688 3227
rect 14746 3227 15042 3263
rect 14746 3207 14806 3227
rect 14864 3207 14924 3227
rect 14982 3207 15042 3227
rect 7504 2986 7564 3012
rect 7622 2986 7682 3012
rect 7740 2986 7800 3012
rect 7858 2992 7918 3012
rect 7858 2986 7919 2992
rect 7976 2986 8036 3012
rect 8094 2986 8154 3012
rect 1696 2967 1762 2983
rect 1696 2933 1712 2967
rect 1746 2933 1762 2967
rect 1696 2917 1762 2933
rect 1578 2850 1644 2866
rect 1578 2816 1594 2850
rect 1628 2816 1644 2850
rect 1578 2800 1644 2816
rect 2939 2813 3235 2864
rect 1581 2778 1641 2800
rect 2939 2798 2999 2813
rect 3057 2798 3117 2813
rect 3175 2798 3235 2813
rect 3293 2798 3353 2824
rect 3411 2798 3471 2824
rect 3529 2798 3589 2824
rect 4837 2813 5133 2864
rect 4837 2798 4897 2813
rect 4955 2798 5015 2813
rect 5073 2798 5133 2813
rect 5191 2798 5251 2824
rect 5309 2798 5369 2824
rect 5427 2798 5487 2824
rect 7741 2801 7799 2986
rect 2455 2598 2515 2624
rect 2573 2598 2633 2624
rect 2691 2598 2751 2624
rect 1581 2552 1641 2578
rect 1228 2356 1288 2378
rect 1346 2362 1406 2378
rect 1225 2340 1291 2356
rect 1225 2306 1241 2340
rect 1275 2306 1291 2340
rect 1225 2290 1291 2306
rect 1340 2340 1414 2362
rect 1340 2306 1359 2340
rect 1393 2306 1414 2340
rect 3776 2615 4072 2666
rect 3776 2598 3836 2615
rect 3894 2598 3954 2615
rect 4012 2598 4072 2615
rect 4353 2598 4413 2624
rect 4471 2598 4531 2624
rect 4589 2598 4649 2624
rect 7741 2775 7801 2801
rect 7859 2775 7919 2986
rect 8212 2980 8272 3012
rect 8330 2986 8390 3012
rect 8448 2986 8508 3012
rect 20596 3232 20892 3268
rect 20596 3211 20656 3232
rect 20714 3211 20774 3232
rect 20832 3211 20892 3232
rect 20950 3231 21246 3267
rect 20950 3211 21010 3231
rect 21068 3211 21128 3231
rect 21186 3211 21246 3231
rect 21304 3231 21600 3267
rect 21304 3211 21364 3231
rect 21422 3211 21482 3231
rect 21540 3211 21600 3231
rect 14038 2981 14098 3007
rect 14156 2981 14216 3007
rect 14274 2981 14334 3007
rect 14392 2987 14452 3007
rect 14392 2981 14453 2987
rect 14510 2981 14570 3007
rect 14628 2981 14688 3007
rect 8209 2964 8275 2980
rect 8209 2930 8225 2964
rect 8259 2930 8275 2964
rect 8209 2914 8275 2930
rect 8091 2847 8157 2863
rect 8091 2813 8107 2847
rect 8141 2813 8157 2847
rect 8091 2797 8157 2813
rect 9452 2810 9748 2861
rect 8094 2775 8154 2797
rect 9452 2795 9512 2810
rect 9570 2795 9630 2810
rect 9688 2795 9748 2810
rect 9806 2795 9866 2821
rect 9924 2795 9984 2821
rect 10042 2795 10102 2821
rect 11350 2810 11646 2861
rect 11350 2795 11410 2810
rect 11468 2795 11528 2810
rect 11586 2795 11646 2810
rect 11704 2795 11764 2821
rect 11822 2795 11882 2821
rect 11940 2795 12000 2821
rect 14275 2796 14333 2981
rect 5674 2615 5970 2666
rect 5674 2598 5734 2615
rect 5792 2598 5852 2615
rect 5910 2598 5970 2615
rect 2455 2381 2515 2398
rect 2573 2381 2633 2398
rect 2691 2381 2751 2398
rect 2939 2381 2999 2398
rect 2455 2330 2999 2381
rect 3057 2372 3117 2398
rect 3175 2372 3235 2398
rect 3293 2379 3353 2398
rect 3411 2379 3471 2398
rect 3529 2379 3589 2398
rect 3776 2379 3836 2398
rect 3894 2379 3954 2398
rect 1340 2249 1414 2306
rect 2580 2249 2640 2330
rect 3293 2328 3836 2379
rect 3878 2372 3954 2379
rect 4012 2372 4072 2398
rect 4353 2381 4413 2398
rect 4471 2381 4531 2398
rect 4589 2381 4649 2398
rect 4837 2381 4897 2398
rect 3878 2328 3953 2372
rect 4353 2330 4897 2381
rect 4955 2372 5015 2398
rect 5073 2372 5133 2398
rect 5191 2379 5251 2398
rect 5309 2379 5369 2398
rect 5427 2379 5487 2398
rect 5674 2379 5734 2398
rect 5792 2379 5852 2398
rect 1340 2224 2640 2249
rect 1339 2176 2640 2224
rect 3878 2208 3938 2328
rect 986 1632 1282 1668
rect 986 1611 1046 1632
rect 1104 1611 1164 1632
rect 1222 1611 1282 1632
rect 1340 1631 1636 1667
rect 1340 1611 1400 1631
rect 1458 1611 1518 1631
rect 1576 1611 1636 1631
rect 1694 1631 1990 1667
rect 1694 1611 1754 1631
rect 1812 1611 1872 1631
rect 1930 1611 1990 1631
rect 2580 1478 2640 2176
rect 2882 2128 3178 2188
rect 2882 2105 2942 2128
rect 3000 2105 3060 2128
rect 3118 2105 3178 2128
rect 3236 2129 3532 2189
rect 3877 2188 3938 2208
rect 3236 2105 3296 2129
rect 3354 2105 3414 2129
rect 3472 2105 3532 2129
rect 3858 2172 3938 2188
rect 3858 2138 3873 2172
rect 3907 2138 3938 2172
rect 3858 2122 3938 2138
rect 3877 2099 3938 2122
rect 3878 1953 3938 2099
rect 3877 1780 3938 1953
rect 2882 1679 2942 1705
rect 2850 1538 2917 1545
rect 3000 1538 3060 1705
rect 3118 1679 3178 1705
rect 3236 1679 3296 1705
rect 2850 1529 3060 1538
rect 2850 1495 2866 1529
rect 2900 1495 3060 1529
rect 2850 1479 3060 1495
rect 2580 1462 2731 1478
rect 2580 1428 2681 1462
rect 2715 1428 2731 1462
rect 2580 1412 2731 1428
rect 986 1385 1046 1411
rect 1104 1385 1164 1411
rect 1222 1385 1282 1411
rect 1340 1391 1400 1411
rect 1340 1385 1401 1391
rect 1458 1385 1518 1411
rect 1576 1385 1636 1411
rect 1223 1200 1281 1385
rect 1223 1174 1283 1200
rect 1341 1174 1401 1385
rect 1694 1379 1754 1411
rect 1812 1385 1872 1411
rect 1930 1385 1990 1411
rect 1691 1363 1757 1379
rect 2580 1373 2640 1412
rect 3000 1373 3060 1479
rect 3354 1538 3414 1705
rect 3472 1679 3532 1705
rect 3497 1538 3564 1545
rect 3354 1529 3564 1538
rect 3354 1495 3514 1529
rect 3548 1495 3564 1529
rect 3354 1479 3564 1495
rect 3116 1445 3182 1461
rect 3116 1411 3132 1445
rect 3166 1411 3182 1445
rect 3116 1395 3182 1411
rect 3234 1446 3300 1461
rect 3234 1412 3250 1446
rect 3284 1412 3300 1446
rect 3234 1396 3300 1412
rect 3118 1373 3178 1395
rect 3236 1373 3296 1396
rect 3354 1373 3414 1479
rect 3878 1477 3938 1780
rect 3788 1461 3938 1477
rect 3788 1427 3804 1461
rect 3838 1427 3938 1461
rect 3788 1411 3938 1427
rect 3878 1373 3938 1411
rect 4478 1672 4538 2330
rect 5191 2328 5734 2379
rect 5776 2372 5852 2379
rect 5910 2372 5970 2398
rect 8968 2595 9028 2621
rect 9086 2595 9146 2621
rect 9204 2595 9264 2621
rect 8094 2549 8154 2575
rect 5776 2328 5851 2372
rect 7741 2353 7801 2375
rect 7859 2359 7919 2375
rect 7738 2337 7804 2353
rect 4780 2128 5076 2188
rect 4780 2105 4840 2128
rect 4898 2105 4958 2128
rect 5016 2105 5076 2128
rect 5134 2129 5430 2189
rect 5134 2105 5194 2129
rect 5252 2105 5312 2129
rect 5370 2105 5430 2129
rect 5776 2175 5836 2328
rect 7738 2303 7754 2337
rect 7788 2303 7804 2337
rect 7738 2287 7804 2303
rect 7853 2337 7927 2359
rect 7853 2303 7872 2337
rect 7906 2303 7927 2337
rect 10289 2612 10585 2663
rect 10289 2595 10349 2612
rect 10407 2595 10467 2612
rect 10525 2595 10585 2612
rect 10866 2595 10926 2621
rect 10984 2595 11044 2621
rect 11102 2595 11162 2621
rect 14275 2770 14335 2796
rect 14393 2770 14453 2981
rect 14746 2975 14806 3007
rect 14864 2981 14924 3007
rect 14982 2981 15042 3007
rect 20596 2985 20656 3011
rect 20714 2985 20774 3011
rect 20832 2985 20892 3011
rect 20950 2991 21010 3011
rect 20950 2985 21011 2991
rect 21068 2985 21128 3011
rect 21186 2985 21246 3011
rect 14743 2959 14809 2975
rect 14743 2925 14759 2959
rect 14793 2925 14809 2959
rect 14743 2909 14809 2925
rect 14625 2842 14691 2858
rect 14625 2808 14641 2842
rect 14675 2808 14691 2842
rect 14625 2792 14691 2808
rect 15986 2805 16282 2856
rect 14628 2770 14688 2792
rect 15986 2790 16046 2805
rect 16104 2790 16164 2805
rect 16222 2790 16282 2805
rect 16340 2790 16400 2816
rect 16458 2790 16518 2816
rect 16576 2790 16636 2816
rect 17884 2805 18180 2856
rect 17884 2790 17944 2805
rect 18002 2790 18062 2805
rect 18120 2790 18180 2805
rect 18238 2790 18298 2816
rect 18356 2790 18416 2816
rect 18474 2790 18534 2816
rect 20833 2800 20891 2985
rect 12187 2612 12483 2663
rect 12187 2595 12247 2612
rect 12305 2595 12365 2612
rect 12423 2595 12483 2612
rect 8968 2378 9028 2395
rect 9086 2378 9146 2395
rect 9204 2378 9264 2395
rect 9452 2378 9512 2395
rect 8968 2327 9512 2378
rect 9570 2369 9630 2395
rect 9688 2369 9748 2395
rect 9806 2376 9866 2395
rect 9924 2376 9984 2395
rect 10042 2376 10102 2395
rect 10289 2376 10349 2395
rect 10407 2376 10467 2395
rect 7853 2246 7927 2303
rect 9093 2246 9153 2327
rect 9806 2325 10349 2376
rect 10391 2369 10467 2376
rect 10525 2369 10585 2395
rect 10866 2378 10926 2395
rect 10984 2378 11044 2395
rect 11102 2378 11162 2395
rect 11350 2378 11410 2395
rect 10391 2325 10466 2369
rect 10866 2327 11410 2378
rect 11468 2369 11528 2395
rect 11586 2369 11646 2395
rect 11704 2376 11764 2395
rect 11822 2376 11882 2395
rect 11940 2376 12000 2395
rect 12187 2376 12247 2395
rect 12305 2376 12365 2395
rect 7853 2221 9153 2246
rect 5776 2151 6030 2175
rect 7852 2173 9153 2221
rect 10391 2205 10451 2325
rect 5776 2117 5980 2151
rect 6014 2117 6030 2151
rect 5776 2101 6030 2117
rect 4780 1679 4840 1705
rect 4478 1656 4545 1672
rect 4478 1622 4494 1656
rect 4528 1622 4545 1656
rect 4478 1606 4545 1622
rect 4478 1478 4538 1606
rect 4748 1538 4815 1545
rect 4898 1538 4958 1705
rect 5016 1679 5076 1705
rect 5134 1679 5194 1705
rect 4748 1529 4958 1538
rect 4748 1495 4764 1529
rect 4798 1495 4958 1529
rect 4748 1479 4958 1495
rect 4478 1462 4629 1478
rect 4478 1428 4579 1462
rect 4613 1428 4629 1462
rect 4478 1412 4629 1428
rect 4478 1373 4538 1412
rect 4898 1373 4958 1479
rect 5252 1538 5312 1705
rect 5370 1679 5430 1705
rect 5393 1539 5460 1546
rect 5387 1538 5460 1539
rect 5252 1530 5460 1538
rect 5252 1496 5410 1530
rect 5444 1496 5460 1530
rect 5252 1480 5460 1496
rect 5252 1479 5449 1480
rect 5014 1445 5080 1461
rect 5014 1411 5030 1445
rect 5064 1411 5080 1445
rect 5014 1395 5080 1411
rect 5132 1446 5198 1461
rect 5132 1412 5148 1446
rect 5182 1412 5198 1446
rect 5132 1396 5198 1412
rect 5016 1373 5076 1395
rect 5134 1373 5194 1396
rect 5252 1373 5312 1479
rect 5776 1477 5836 2101
rect 7499 1629 7795 1665
rect 7499 1608 7559 1629
rect 7617 1608 7677 1629
rect 7735 1608 7795 1629
rect 7853 1628 8149 1664
rect 7853 1608 7913 1628
rect 7971 1608 8031 1628
rect 8089 1608 8149 1628
rect 8207 1628 8503 1664
rect 8207 1608 8267 1628
rect 8325 1608 8385 1628
rect 8443 1608 8503 1628
rect 5686 1461 5836 1477
rect 5686 1427 5702 1461
rect 5736 1427 5836 1461
rect 5686 1411 5836 1427
rect 5776 1373 5836 1411
rect 9093 1475 9153 2173
rect 9395 2125 9691 2185
rect 9395 2102 9455 2125
rect 9513 2102 9573 2125
rect 9631 2102 9691 2125
rect 9749 2126 10045 2186
rect 10390 2185 10451 2205
rect 9749 2102 9809 2126
rect 9867 2102 9927 2126
rect 9985 2102 10045 2126
rect 10371 2169 10451 2185
rect 10371 2135 10386 2169
rect 10420 2135 10451 2169
rect 10371 2119 10451 2135
rect 10390 2096 10451 2119
rect 10391 1950 10451 2096
rect 10390 1777 10451 1950
rect 9395 1676 9455 1702
rect 9363 1535 9430 1542
rect 9513 1535 9573 1702
rect 9631 1676 9691 1702
rect 9749 1676 9809 1702
rect 9363 1526 9573 1535
rect 9363 1492 9379 1526
rect 9413 1492 9573 1526
rect 9363 1476 9573 1492
rect 9093 1459 9244 1475
rect 9093 1425 9194 1459
rect 9228 1425 9244 1459
rect 9093 1409 9244 1425
rect 7499 1382 7559 1408
rect 7617 1382 7677 1408
rect 7735 1382 7795 1408
rect 7853 1388 7913 1408
rect 7853 1382 7914 1388
rect 7971 1382 8031 1408
rect 8089 1382 8149 1408
rect 1691 1329 1707 1363
rect 1741 1329 1757 1363
rect 1691 1313 1757 1329
rect 1573 1246 1639 1262
rect 1573 1212 1589 1246
rect 1623 1212 1639 1246
rect 1573 1196 1639 1212
rect 1576 1174 1636 1196
rect 2580 1147 2640 1173
rect 1576 948 1636 974
rect 3878 1147 3938 1173
rect 4478 1147 4538 1173
rect 7736 1197 7794 1382
rect 5776 1147 5836 1173
rect 7736 1171 7796 1197
rect 7854 1171 7914 1382
rect 8207 1376 8267 1408
rect 8325 1382 8385 1408
rect 8443 1382 8503 1408
rect 8204 1360 8270 1376
rect 9093 1370 9153 1409
rect 9513 1370 9573 1476
rect 9867 1535 9927 1702
rect 9985 1676 10045 1702
rect 10010 1535 10077 1542
rect 9867 1526 10077 1535
rect 9867 1492 10027 1526
rect 10061 1492 10077 1526
rect 9867 1476 10077 1492
rect 9629 1442 9695 1458
rect 9629 1408 9645 1442
rect 9679 1408 9695 1442
rect 9629 1392 9695 1408
rect 9747 1443 9813 1458
rect 9747 1409 9763 1443
rect 9797 1409 9813 1443
rect 9747 1393 9813 1409
rect 9631 1370 9691 1392
rect 9749 1370 9809 1393
rect 9867 1370 9927 1476
rect 10391 1474 10451 1777
rect 10301 1458 10451 1474
rect 10301 1424 10317 1458
rect 10351 1424 10451 1458
rect 10301 1408 10451 1424
rect 10391 1370 10451 1408
rect 10991 1669 11051 2327
rect 11704 2325 12247 2376
rect 12289 2369 12365 2376
rect 12423 2369 12483 2395
rect 15502 2590 15562 2616
rect 15620 2590 15680 2616
rect 15738 2590 15798 2616
rect 14628 2544 14688 2570
rect 12289 2325 12364 2369
rect 14275 2348 14335 2370
rect 14393 2354 14453 2370
rect 14272 2332 14338 2348
rect 11293 2125 11589 2185
rect 11293 2102 11353 2125
rect 11411 2102 11471 2125
rect 11529 2102 11589 2125
rect 11647 2126 11943 2186
rect 11647 2102 11707 2126
rect 11765 2102 11825 2126
rect 11883 2102 11943 2126
rect 12289 2172 12349 2325
rect 14272 2298 14288 2332
rect 14322 2298 14338 2332
rect 14272 2282 14338 2298
rect 14387 2332 14461 2354
rect 14387 2298 14406 2332
rect 14440 2298 14461 2332
rect 16823 2607 17119 2658
rect 16823 2590 16883 2607
rect 16941 2590 17001 2607
rect 17059 2590 17119 2607
rect 17400 2590 17460 2616
rect 17518 2590 17578 2616
rect 17636 2590 17696 2616
rect 20833 2774 20893 2800
rect 20951 2774 21011 2985
rect 21304 2979 21364 3011
rect 21422 2985 21482 3011
rect 21540 2985 21600 3011
rect 21301 2963 21367 2979
rect 21301 2929 21317 2963
rect 21351 2929 21367 2963
rect 21301 2913 21367 2929
rect 21183 2846 21249 2862
rect 21183 2812 21199 2846
rect 21233 2812 21249 2846
rect 21183 2796 21249 2812
rect 22544 2809 22840 2860
rect 21186 2774 21246 2796
rect 22544 2794 22604 2809
rect 22662 2794 22722 2809
rect 22780 2794 22840 2809
rect 22898 2794 22958 2820
rect 23016 2794 23076 2820
rect 23134 2794 23194 2820
rect 24442 2809 24738 2860
rect 24442 2794 24502 2809
rect 24560 2794 24620 2809
rect 24678 2794 24738 2809
rect 24796 2794 24856 2820
rect 24914 2794 24974 2820
rect 25032 2794 25092 2820
rect 18721 2607 19017 2658
rect 18721 2590 18781 2607
rect 18839 2590 18899 2607
rect 18957 2590 19017 2607
rect 15502 2373 15562 2390
rect 15620 2373 15680 2390
rect 15738 2373 15798 2390
rect 15986 2373 16046 2390
rect 15502 2322 16046 2373
rect 16104 2364 16164 2390
rect 16222 2364 16282 2390
rect 16340 2371 16400 2390
rect 16458 2371 16518 2390
rect 16576 2371 16636 2390
rect 16823 2371 16883 2390
rect 16941 2371 17001 2390
rect 14387 2241 14461 2298
rect 15627 2241 15687 2322
rect 16340 2320 16883 2371
rect 16925 2364 17001 2371
rect 17059 2364 17119 2390
rect 17400 2373 17460 2390
rect 17518 2373 17578 2390
rect 17636 2373 17696 2390
rect 17884 2373 17944 2390
rect 16925 2320 17000 2364
rect 17400 2322 17944 2373
rect 18002 2364 18062 2390
rect 18120 2364 18180 2390
rect 18238 2371 18298 2390
rect 18356 2371 18416 2390
rect 18474 2371 18534 2390
rect 18721 2371 18781 2390
rect 18839 2371 18899 2390
rect 14387 2216 15687 2241
rect 12289 2148 12543 2172
rect 14386 2168 15687 2216
rect 16925 2200 16985 2320
rect 12289 2114 12493 2148
rect 12527 2114 12543 2148
rect 12289 2098 12543 2114
rect 11293 1676 11353 1702
rect 10991 1653 11058 1669
rect 10991 1619 11007 1653
rect 11041 1619 11058 1653
rect 10991 1603 11058 1619
rect 10991 1475 11051 1603
rect 11261 1535 11328 1542
rect 11411 1535 11471 1702
rect 11529 1676 11589 1702
rect 11647 1676 11707 1702
rect 11261 1526 11471 1535
rect 11261 1492 11277 1526
rect 11311 1492 11471 1526
rect 11261 1476 11471 1492
rect 10991 1459 11142 1475
rect 10991 1425 11092 1459
rect 11126 1425 11142 1459
rect 10991 1409 11142 1425
rect 10991 1370 11051 1409
rect 11411 1370 11471 1476
rect 11765 1535 11825 1702
rect 11883 1676 11943 1702
rect 11906 1536 11973 1543
rect 11900 1535 11973 1536
rect 11765 1527 11973 1535
rect 11765 1493 11923 1527
rect 11957 1493 11973 1527
rect 11765 1477 11973 1493
rect 11765 1476 11962 1477
rect 11527 1442 11593 1458
rect 11527 1408 11543 1442
rect 11577 1408 11593 1442
rect 11527 1392 11593 1408
rect 11645 1443 11711 1458
rect 11645 1409 11661 1443
rect 11695 1409 11711 1443
rect 11645 1393 11711 1409
rect 11529 1370 11589 1392
rect 11647 1370 11707 1393
rect 11765 1370 11825 1476
rect 12289 1474 12349 2098
rect 14033 1624 14329 1660
rect 14033 1603 14093 1624
rect 14151 1603 14211 1624
rect 14269 1603 14329 1624
rect 14387 1623 14683 1659
rect 14387 1603 14447 1623
rect 14505 1603 14565 1623
rect 14623 1603 14683 1623
rect 14741 1623 15037 1659
rect 14741 1603 14801 1623
rect 14859 1603 14919 1623
rect 14977 1603 15037 1623
rect 12199 1458 12349 1474
rect 12199 1424 12215 1458
rect 12249 1424 12349 1458
rect 12199 1408 12349 1424
rect 12289 1370 12349 1408
rect 15627 1470 15687 2168
rect 15929 2120 16225 2180
rect 15929 2097 15989 2120
rect 16047 2097 16107 2120
rect 16165 2097 16225 2120
rect 16283 2121 16579 2181
rect 16924 2180 16985 2200
rect 16283 2097 16343 2121
rect 16401 2097 16461 2121
rect 16519 2097 16579 2121
rect 16905 2164 16985 2180
rect 16905 2130 16920 2164
rect 16954 2130 16985 2164
rect 16905 2114 16985 2130
rect 16924 2091 16985 2114
rect 16925 1945 16985 2091
rect 16924 1772 16985 1945
rect 15929 1671 15989 1697
rect 15897 1530 15964 1537
rect 16047 1530 16107 1697
rect 16165 1671 16225 1697
rect 16283 1671 16343 1697
rect 15897 1521 16107 1530
rect 15897 1487 15913 1521
rect 15947 1487 16107 1521
rect 15897 1471 16107 1487
rect 15627 1454 15778 1470
rect 15627 1420 15728 1454
rect 15762 1420 15778 1454
rect 15627 1404 15778 1420
rect 14033 1377 14093 1403
rect 14151 1377 14211 1403
rect 14269 1377 14329 1403
rect 14387 1383 14447 1403
rect 14387 1377 14448 1383
rect 14505 1377 14565 1403
rect 14623 1377 14683 1403
rect 8204 1326 8220 1360
rect 8254 1326 8270 1360
rect 8204 1310 8270 1326
rect 8086 1243 8152 1259
rect 8086 1209 8102 1243
rect 8136 1209 8152 1243
rect 8086 1193 8152 1209
rect 8089 1171 8149 1193
rect 3000 947 3060 973
rect 3118 947 3178 973
rect 3236 947 3296 973
rect 3354 947 3414 973
rect 4898 947 4958 973
rect 5016 947 5076 973
rect 5134 947 5194 973
rect 5252 947 5312 973
rect 1223 752 1283 774
rect 1341 752 1401 774
rect 1220 736 1286 752
rect 1220 702 1236 736
rect 1270 702 1286 736
rect 1220 686 1286 702
rect 1338 736 1404 752
rect 1338 702 1354 736
rect 1388 702 1404 736
rect 9093 1144 9153 1170
rect 8089 945 8149 971
rect 10391 1144 10451 1170
rect 10991 1144 11051 1170
rect 14270 1192 14328 1377
rect 12289 1144 12349 1170
rect 14270 1166 14330 1192
rect 14388 1166 14448 1377
rect 14741 1371 14801 1403
rect 14859 1377 14919 1403
rect 14977 1377 15037 1403
rect 14738 1355 14804 1371
rect 15627 1365 15687 1404
rect 16047 1365 16107 1471
rect 16401 1530 16461 1697
rect 16519 1671 16579 1697
rect 16544 1530 16611 1537
rect 16401 1521 16611 1530
rect 16401 1487 16561 1521
rect 16595 1487 16611 1521
rect 16401 1471 16611 1487
rect 16163 1437 16229 1453
rect 16163 1403 16179 1437
rect 16213 1403 16229 1437
rect 16163 1387 16229 1403
rect 16281 1438 16347 1453
rect 16281 1404 16297 1438
rect 16331 1404 16347 1438
rect 16281 1388 16347 1404
rect 16165 1365 16225 1387
rect 16283 1365 16343 1388
rect 16401 1365 16461 1471
rect 16925 1469 16985 1772
rect 16835 1453 16985 1469
rect 16835 1419 16851 1453
rect 16885 1419 16985 1453
rect 16835 1403 16985 1419
rect 16925 1365 16985 1403
rect 17525 1664 17585 2322
rect 18238 2320 18781 2371
rect 18823 2364 18899 2371
rect 18957 2364 19017 2390
rect 22060 2594 22120 2620
rect 22178 2594 22238 2620
rect 22296 2594 22356 2620
rect 21186 2548 21246 2574
rect 18823 2320 18898 2364
rect 20833 2352 20893 2374
rect 20951 2358 21011 2374
rect 20830 2336 20896 2352
rect 17827 2120 18123 2180
rect 17827 2097 17887 2120
rect 17945 2097 18005 2120
rect 18063 2097 18123 2120
rect 18181 2121 18477 2181
rect 18181 2097 18241 2121
rect 18299 2097 18359 2121
rect 18417 2097 18477 2121
rect 18823 2167 18883 2320
rect 20830 2302 20846 2336
rect 20880 2302 20896 2336
rect 20830 2286 20896 2302
rect 20945 2336 21019 2358
rect 20945 2302 20964 2336
rect 20998 2302 21019 2336
rect 23381 2611 23677 2662
rect 23381 2594 23441 2611
rect 23499 2594 23559 2611
rect 23617 2594 23677 2611
rect 23958 2594 24018 2620
rect 24076 2594 24136 2620
rect 24194 2594 24254 2620
rect 25279 2611 25575 2662
rect 25279 2594 25339 2611
rect 25397 2594 25457 2611
rect 25515 2594 25575 2611
rect 22060 2377 22120 2394
rect 22178 2377 22238 2394
rect 22296 2377 22356 2394
rect 22544 2377 22604 2394
rect 22060 2326 22604 2377
rect 22662 2368 22722 2394
rect 22780 2368 22840 2394
rect 22898 2375 22958 2394
rect 23016 2375 23076 2394
rect 23134 2375 23194 2394
rect 23381 2375 23441 2394
rect 23499 2375 23559 2394
rect 20945 2245 21019 2302
rect 22185 2245 22245 2326
rect 22898 2324 23441 2375
rect 23483 2368 23559 2375
rect 23617 2368 23677 2394
rect 23958 2377 24018 2394
rect 24076 2377 24136 2394
rect 24194 2377 24254 2394
rect 24442 2377 24502 2394
rect 23483 2324 23558 2368
rect 23958 2326 24502 2377
rect 24560 2368 24620 2394
rect 24678 2368 24738 2394
rect 24796 2375 24856 2394
rect 24914 2375 24974 2394
rect 25032 2375 25092 2394
rect 25279 2375 25339 2394
rect 25397 2375 25457 2394
rect 20945 2220 22245 2245
rect 20944 2172 22245 2220
rect 23483 2204 23543 2324
rect 18823 2143 19077 2167
rect 18823 2109 19027 2143
rect 19061 2109 19077 2143
rect 18823 2093 19077 2109
rect 17827 1671 17887 1697
rect 17525 1648 17592 1664
rect 17525 1614 17541 1648
rect 17575 1614 17592 1648
rect 17525 1598 17592 1614
rect 17525 1470 17585 1598
rect 17795 1530 17862 1537
rect 17945 1530 18005 1697
rect 18063 1671 18123 1697
rect 18181 1671 18241 1697
rect 17795 1521 18005 1530
rect 17795 1487 17811 1521
rect 17845 1487 18005 1521
rect 17795 1471 18005 1487
rect 17525 1454 17676 1470
rect 17525 1420 17626 1454
rect 17660 1420 17676 1454
rect 17525 1404 17676 1420
rect 17525 1365 17585 1404
rect 17945 1365 18005 1471
rect 18299 1530 18359 1697
rect 18417 1671 18477 1697
rect 18440 1531 18507 1538
rect 18434 1530 18507 1531
rect 18299 1522 18507 1530
rect 18299 1488 18457 1522
rect 18491 1488 18507 1522
rect 18299 1472 18507 1488
rect 18299 1471 18496 1472
rect 18061 1437 18127 1453
rect 18061 1403 18077 1437
rect 18111 1403 18127 1437
rect 18061 1387 18127 1403
rect 18179 1438 18245 1453
rect 18179 1404 18195 1438
rect 18229 1404 18245 1438
rect 18179 1388 18245 1404
rect 18063 1365 18123 1387
rect 18181 1365 18241 1388
rect 18299 1365 18359 1471
rect 18823 1469 18883 2093
rect 20591 1628 20887 1664
rect 20591 1607 20651 1628
rect 20709 1607 20769 1628
rect 20827 1607 20887 1628
rect 20945 1627 21241 1663
rect 20945 1607 21005 1627
rect 21063 1607 21123 1627
rect 21181 1607 21241 1627
rect 21299 1627 21595 1663
rect 21299 1607 21359 1627
rect 21417 1607 21477 1627
rect 21535 1607 21595 1627
rect 18733 1453 18883 1469
rect 18733 1419 18749 1453
rect 18783 1419 18883 1453
rect 18733 1403 18883 1419
rect 22185 1474 22245 2172
rect 22487 2124 22783 2184
rect 22487 2101 22547 2124
rect 22605 2101 22665 2124
rect 22723 2101 22783 2124
rect 22841 2125 23137 2185
rect 23482 2184 23543 2204
rect 22841 2101 22901 2125
rect 22959 2101 23019 2125
rect 23077 2101 23137 2125
rect 23463 2168 23543 2184
rect 23463 2134 23478 2168
rect 23512 2134 23543 2168
rect 23463 2118 23543 2134
rect 23482 2095 23543 2118
rect 23483 1949 23543 2095
rect 23482 1776 23543 1949
rect 22487 1675 22547 1701
rect 22455 1534 22522 1541
rect 22605 1534 22665 1701
rect 22723 1675 22783 1701
rect 22841 1675 22901 1701
rect 22455 1525 22665 1534
rect 22455 1491 22471 1525
rect 22505 1491 22665 1525
rect 22455 1475 22665 1491
rect 22185 1458 22336 1474
rect 22185 1424 22286 1458
rect 22320 1424 22336 1458
rect 22185 1408 22336 1424
rect 18823 1365 18883 1403
rect 20591 1381 20651 1407
rect 20709 1381 20769 1407
rect 20827 1381 20887 1407
rect 20945 1387 21005 1407
rect 20945 1381 21006 1387
rect 21063 1381 21123 1407
rect 21181 1381 21241 1407
rect 14738 1321 14754 1355
rect 14788 1321 14804 1355
rect 14738 1305 14804 1321
rect 14620 1238 14686 1254
rect 14620 1204 14636 1238
rect 14670 1204 14686 1238
rect 14620 1188 14686 1204
rect 14623 1166 14683 1188
rect 9513 944 9573 970
rect 9631 944 9691 970
rect 9749 944 9809 970
rect 9867 944 9927 970
rect 11411 944 11471 970
rect 11529 944 11589 970
rect 11647 944 11707 970
rect 11765 944 11825 970
rect 7736 749 7796 771
rect 7854 749 7914 771
rect 7733 733 7799 749
rect 1338 686 1404 702
rect 7733 699 7749 733
rect 7783 699 7799 733
rect 7733 683 7799 699
rect 7851 733 7917 749
rect 7851 699 7867 733
rect 7901 699 7917 733
rect 15627 1139 15687 1165
rect 14623 940 14683 966
rect 16925 1139 16985 1165
rect 17525 1139 17585 1165
rect 20828 1196 20886 1381
rect 20828 1170 20888 1196
rect 20946 1170 21006 1381
rect 21299 1375 21359 1407
rect 21417 1381 21477 1407
rect 21535 1381 21595 1407
rect 21296 1359 21362 1375
rect 22185 1369 22245 1408
rect 22605 1369 22665 1475
rect 22959 1534 23019 1701
rect 23077 1675 23137 1701
rect 23102 1534 23169 1541
rect 22959 1525 23169 1534
rect 22959 1491 23119 1525
rect 23153 1491 23169 1525
rect 22959 1475 23169 1491
rect 22721 1441 22787 1457
rect 22721 1407 22737 1441
rect 22771 1407 22787 1441
rect 22721 1391 22787 1407
rect 22839 1442 22905 1457
rect 22839 1408 22855 1442
rect 22889 1408 22905 1442
rect 22839 1392 22905 1408
rect 22723 1369 22783 1391
rect 22841 1369 22901 1392
rect 22959 1369 23019 1475
rect 23483 1473 23543 1776
rect 23393 1457 23543 1473
rect 23393 1423 23409 1457
rect 23443 1423 23543 1457
rect 23393 1407 23543 1423
rect 23483 1369 23543 1407
rect 24083 1668 24143 2326
rect 24796 2324 25339 2375
rect 25381 2368 25457 2375
rect 25515 2368 25575 2394
rect 25381 2324 25456 2368
rect 24385 2124 24681 2184
rect 24385 2101 24445 2124
rect 24503 2101 24563 2124
rect 24621 2101 24681 2124
rect 24739 2125 25035 2185
rect 24739 2101 24799 2125
rect 24857 2101 24917 2125
rect 24975 2101 25035 2125
rect 25381 2171 25441 2324
rect 25381 2147 25635 2171
rect 25381 2113 25585 2147
rect 25619 2113 25635 2147
rect 25381 2097 25635 2113
rect 24385 1675 24445 1701
rect 24083 1652 24150 1668
rect 24083 1618 24099 1652
rect 24133 1618 24150 1652
rect 24083 1602 24150 1618
rect 24083 1474 24143 1602
rect 24353 1534 24420 1541
rect 24503 1534 24563 1701
rect 24621 1675 24681 1701
rect 24739 1675 24799 1701
rect 24353 1525 24563 1534
rect 24353 1491 24369 1525
rect 24403 1491 24563 1525
rect 24353 1475 24563 1491
rect 24083 1458 24234 1474
rect 24083 1424 24184 1458
rect 24218 1424 24234 1458
rect 24083 1408 24234 1424
rect 24083 1369 24143 1408
rect 24503 1369 24563 1475
rect 24857 1534 24917 1701
rect 24975 1675 25035 1701
rect 24998 1535 25065 1542
rect 24992 1534 25065 1535
rect 24857 1526 25065 1534
rect 24857 1492 25015 1526
rect 25049 1492 25065 1526
rect 24857 1476 25065 1492
rect 24857 1475 25054 1476
rect 24619 1441 24685 1457
rect 24619 1407 24635 1441
rect 24669 1407 24685 1441
rect 24619 1391 24685 1407
rect 24737 1442 24803 1457
rect 24737 1408 24753 1442
rect 24787 1408 24803 1442
rect 24737 1392 24803 1408
rect 24621 1369 24681 1391
rect 24739 1369 24799 1392
rect 24857 1369 24917 1475
rect 25381 1473 25441 2097
rect 25291 1457 25441 1473
rect 25291 1423 25307 1457
rect 25341 1423 25441 1457
rect 25291 1407 25441 1423
rect 25381 1369 25441 1407
rect 21296 1325 21312 1359
rect 21346 1325 21362 1359
rect 21296 1309 21362 1325
rect 21178 1242 21244 1258
rect 21178 1208 21194 1242
rect 21228 1208 21244 1242
rect 21178 1192 21244 1208
rect 21181 1170 21241 1192
rect 18823 1139 18883 1165
rect 16047 939 16107 965
rect 16165 939 16225 965
rect 16283 939 16343 965
rect 16401 939 16461 965
rect 17945 939 18005 965
rect 18063 939 18123 965
rect 18181 939 18241 965
rect 18299 939 18359 965
rect 14270 744 14330 766
rect 14388 744 14448 766
rect 14267 728 14333 744
rect 7851 683 7917 699
rect 14267 694 14283 728
rect 14317 694 14333 728
rect 14267 678 14333 694
rect 14385 728 14451 744
rect 14385 694 14401 728
rect 14435 694 14451 728
rect 22185 1143 22245 1169
rect 21181 944 21241 970
rect 23483 1143 23543 1169
rect 24083 1143 24143 1169
rect 25381 1143 25441 1169
rect 22605 943 22665 969
rect 22723 943 22783 969
rect 22841 943 22901 969
rect 22959 943 23019 969
rect 24503 943 24563 969
rect 24621 943 24681 969
rect 24739 943 24799 969
rect 24857 943 24917 969
rect 20828 748 20888 770
rect 20946 748 21006 770
rect 20825 732 20891 748
rect 14385 678 14451 694
rect 20825 698 20841 732
rect 20875 698 20891 732
rect 20825 682 20891 698
rect 20943 732 21009 748
rect 20943 698 20959 732
rect 20993 698 21009 732
rect 20943 682 21009 698
rect 1761 -501 1827 -485
rect 1761 -510 1777 -501
rect 1240 -535 1777 -510
rect 1811 -535 1827 -501
rect 2891 -507 2957 -491
rect 2891 -514 2907 -507
rect 1240 -553 1827 -535
rect 2382 -541 2907 -514
rect 2941 -541 2957 -507
rect 1240 -605 1284 -553
rect 2382 -557 2957 -541
rect 988 -646 1284 -605
rect 988 -667 1048 -646
rect 1106 -667 1166 -646
rect 1224 -667 1284 -646
rect 1342 -621 1827 -605
rect 2382 -609 2426 -557
rect 8319 -505 8385 -489
rect 8319 -514 8335 -505
rect 7798 -539 8335 -514
rect 8369 -539 8385 -505
rect 9449 -511 9515 -495
rect 9449 -518 9465 -511
rect 7798 -557 8385 -539
rect 8940 -545 9465 -518
rect 9499 -545 9515 -511
rect 7798 -609 7842 -557
rect 8940 -561 9515 -545
rect 1342 -646 1777 -621
rect 1342 -667 1402 -646
rect 1460 -667 1520 -646
rect 1578 -647 1777 -646
rect 1578 -667 1638 -647
rect 1761 -655 1777 -647
rect 1811 -655 1827 -621
rect 1761 -671 1827 -655
rect 2130 -650 2426 -609
rect 2130 -671 2190 -650
rect 2248 -671 2308 -650
rect 2366 -671 2426 -650
rect 2484 -625 2957 -609
rect 2484 -650 2907 -625
rect 2484 -671 2544 -650
rect 2602 -671 2662 -650
rect 2720 -651 2907 -650
rect 2720 -671 2780 -651
rect 2891 -659 2907 -651
rect 2941 -659 2957 -625
rect 988 -1093 1048 -1067
rect 1106 -1093 1166 -1067
rect 1224 -1268 1284 -1067
rect 1342 -1093 1402 -1067
rect 1460 -1093 1520 -1067
rect 1578 -1084 1638 -1067
rect 2891 -675 2957 -659
rect 7546 -650 7842 -609
rect 7546 -671 7606 -650
rect 7664 -671 7724 -650
rect 7782 -671 7842 -650
rect 7900 -625 8385 -609
rect 8940 -613 8984 -561
rect 14853 -500 14919 -484
rect 14853 -509 14869 -500
rect 14332 -534 14869 -509
rect 14903 -534 14919 -500
rect 15983 -506 16049 -490
rect 15983 -513 15999 -506
rect 14332 -552 14919 -534
rect 15474 -540 15999 -513
rect 16033 -540 16049 -506
rect 14332 -604 14376 -552
rect 15474 -556 16049 -540
rect 7900 -650 8335 -625
rect 7900 -671 7960 -650
rect 8018 -671 8078 -650
rect 8136 -651 8335 -650
rect 8136 -671 8196 -651
rect 8319 -659 8335 -651
rect 8369 -659 8385 -625
rect 4101 -723 4397 -687
rect 4101 -743 4161 -723
rect 4219 -743 4279 -723
rect 4337 -743 4397 -723
rect 4455 -723 4751 -687
rect 4455 -743 4515 -723
rect 4573 -743 4633 -723
rect 4691 -743 4751 -723
rect 4809 -722 5105 -686
rect 4809 -743 4869 -722
rect 4927 -743 4987 -722
rect 5045 -743 5105 -722
rect 4101 -969 4161 -943
rect 4219 -969 4279 -943
rect 4337 -975 4397 -943
rect 4455 -969 4515 -943
rect 4573 -969 4633 -943
rect 4691 -963 4751 -943
rect 4690 -969 4751 -963
rect 4809 -969 4869 -943
rect 4927 -969 4987 -943
rect 5045 -969 5105 -943
rect 4334 -991 4400 -975
rect 4334 -1025 4350 -991
rect 4384 -1025 4400 -991
rect 4334 -1041 4400 -1025
rect 1577 -1173 1638 -1084
rect 2130 -1097 2190 -1071
rect 2248 -1097 2308 -1071
rect 1577 -1226 1728 -1173
rect 1224 -1319 1610 -1268
rect 1429 -1377 1495 -1361
rect 1429 -1411 1445 -1377
rect 1479 -1411 1495 -1377
rect 913 -1450 973 -1424
rect 1031 -1450 1091 -1424
rect 1149 -1450 1209 -1424
rect 1429 -1427 1495 -1411
rect 1432 -1450 1492 -1427
rect 1550 -1450 1610 -1319
rect 1668 -1450 1728 -1226
rect 2366 -1272 2426 -1071
rect 2484 -1097 2544 -1071
rect 2602 -1097 2662 -1071
rect 2720 -1088 2780 -1071
rect 2719 -1177 2780 -1088
rect 4452 -1108 4518 -1092
rect 4452 -1142 4468 -1108
rect 4502 -1142 4518 -1108
rect 4452 -1158 4518 -1142
rect 2719 -1230 2870 -1177
rect 4455 -1180 4515 -1158
rect 4690 -1180 4750 -969
rect 4810 -1154 4868 -969
rect 8319 -675 8385 -659
rect 8688 -654 8984 -613
rect 8688 -675 8748 -654
rect 8806 -675 8866 -654
rect 8924 -675 8984 -654
rect 9042 -629 9515 -613
rect 9042 -654 9465 -629
rect 9042 -675 9102 -654
rect 9160 -675 9220 -654
rect 9278 -655 9465 -654
rect 9278 -675 9338 -655
rect 9449 -663 9465 -655
rect 9499 -663 9515 -629
rect 7546 -1097 7606 -1071
rect 7664 -1097 7724 -1071
rect 4808 -1180 4868 -1154
rect 2366 -1323 2752 -1272
rect 2571 -1381 2637 -1365
rect 2571 -1415 2587 -1381
rect 2621 -1415 2637 -1381
rect 2055 -1454 2115 -1428
rect 2173 -1454 2233 -1428
rect 2291 -1454 2351 -1428
rect 2571 -1431 2637 -1415
rect 2574 -1454 2634 -1431
rect 2692 -1454 2752 -1323
rect 2810 -1454 2870 -1230
rect 4455 -1406 4515 -1380
rect 913 -1682 973 -1650
rect 1031 -1682 1091 -1650
rect 1149 -1682 1209 -1650
rect 1432 -1682 1492 -1650
rect 1550 -1676 1610 -1650
rect 1668 -1676 1728 -1650
rect 7782 -1272 7842 -1071
rect 7900 -1097 7960 -1071
rect 8018 -1097 8078 -1071
rect 8136 -1088 8196 -1071
rect 9449 -679 9515 -663
rect 14080 -645 14376 -604
rect 14080 -666 14140 -645
rect 14198 -666 14258 -645
rect 14316 -666 14376 -645
rect 14434 -620 14919 -604
rect 15474 -608 15518 -556
rect 21366 -497 21432 -481
rect 21366 -506 21382 -497
rect 20845 -531 21382 -506
rect 21416 -531 21432 -497
rect 22496 -503 22562 -487
rect 22496 -510 22512 -503
rect 20845 -549 21432 -531
rect 21987 -537 22512 -510
rect 22546 -537 22562 -503
rect 20845 -601 20889 -549
rect 21987 -553 22562 -537
rect 14434 -645 14869 -620
rect 14434 -666 14494 -645
rect 14552 -666 14612 -645
rect 14670 -646 14869 -645
rect 14670 -666 14730 -646
rect 14853 -654 14869 -646
rect 14903 -654 14919 -620
rect 10659 -727 10955 -691
rect 10659 -747 10719 -727
rect 10777 -747 10837 -727
rect 10895 -747 10955 -727
rect 11013 -727 11309 -691
rect 11013 -747 11073 -727
rect 11131 -747 11191 -727
rect 11249 -747 11309 -727
rect 11367 -726 11663 -690
rect 11367 -747 11427 -726
rect 11485 -747 11545 -726
rect 11603 -747 11663 -726
rect 10659 -973 10719 -947
rect 10777 -973 10837 -947
rect 10895 -979 10955 -947
rect 11013 -973 11073 -947
rect 11131 -973 11191 -947
rect 11249 -967 11309 -947
rect 11248 -973 11309 -967
rect 11367 -973 11427 -947
rect 11485 -973 11545 -947
rect 11603 -973 11663 -947
rect 10892 -995 10958 -979
rect 10892 -1029 10908 -995
rect 10942 -1029 10958 -995
rect 10892 -1045 10958 -1029
rect 8135 -1177 8196 -1088
rect 8688 -1101 8748 -1075
rect 8806 -1101 8866 -1075
rect 8135 -1230 8286 -1177
rect 7782 -1323 8168 -1272
rect 7987 -1381 8053 -1365
rect 7987 -1415 8003 -1381
rect 8037 -1415 8053 -1381
rect 7471 -1454 7531 -1428
rect 7589 -1454 7649 -1428
rect 7707 -1454 7767 -1428
rect 7987 -1431 8053 -1415
rect 7990 -1454 8050 -1431
rect 8108 -1454 8168 -1323
rect 8226 -1454 8286 -1230
rect 8924 -1276 8984 -1075
rect 9042 -1101 9102 -1075
rect 9160 -1101 9220 -1075
rect 9278 -1092 9338 -1075
rect 9277 -1181 9338 -1092
rect 11010 -1112 11076 -1096
rect 11010 -1146 11026 -1112
rect 11060 -1146 11076 -1112
rect 11010 -1162 11076 -1146
rect 9277 -1234 9428 -1181
rect 11013 -1184 11073 -1162
rect 11248 -1184 11308 -973
rect 11368 -1158 11426 -973
rect 14853 -670 14919 -654
rect 15222 -649 15518 -608
rect 15222 -670 15282 -649
rect 15340 -670 15400 -649
rect 15458 -670 15518 -649
rect 15576 -624 16049 -608
rect 15576 -649 15999 -624
rect 15576 -670 15636 -649
rect 15694 -670 15754 -649
rect 15812 -650 15999 -649
rect 15812 -670 15872 -650
rect 15983 -658 15999 -650
rect 16033 -658 16049 -624
rect 14080 -1092 14140 -1066
rect 14198 -1092 14258 -1066
rect 11366 -1184 11426 -1158
rect 8924 -1327 9310 -1276
rect 9129 -1385 9195 -1369
rect 9129 -1419 9145 -1385
rect 9179 -1419 9195 -1385
rect 4690 -1602 4750 -1580
rect 4808 -1602 4868 -1580
rect 4687 -1618 4753 -1602
rect 4687 -1652 4703 -1618
rect 4737 -1652 4753 -1618
rect 913 -1723 1492 -1682
rect 2055 -1686 2115 -1654
rect 2173 -1686 2233 -1654
rect 2291 -1686 2351 -1654
rect 2574 -1686 2634 -1654
rect 2692 -1680 2752 -1654
rect 2810 -1680 2870 -1654
rect 4687 -1668 4753 -1652
rect 4805 -1618 4871 -1602
rect 4805 -1652 4821 -1618
rect 4855 -1652 4871 -1618
rect 4805 -1668 4871 -1652
rect 8613 -1458 8673 -1432
rect 8731 -1458 8791 -1432
rect 8849 -1458 8909 -1432
rect 9129 -1435 9195 -1419
rect 9132 -1458 9192 -1435
rect 9250 -1458 9310 -1327
rect 9368 -1458 9428 -1234
rect 11013 -1410 11073 -1384
rect 2055 -1727 2634 -1686
rect 7471 -1686 7531 -1654
rect 7589 -1686 7649 -1654
rect 7707 -1686 7767 -1654
rect 7990 -1686 8050 -1654
rect 8108 -1680 8168 -1654
rect 8226 -1680 8286 -1654
rect 14316 -1267 14376 -1066
rect 14434 -1092 14494 -1066
rect 14552 -1092 14612 -1066
rect 14670 -1083 14730 -1066
rect 15983 -674 16049 -658
rect 20593 -642 20889 -601
rect 20593 -663 20653 -642
rect 20711 -663 20771 -642
rect 20829 -663 20889 -642
rect 20947 -617 21432 -601
rect 21987 -605 22031 -553
rect 20947 -642 21382 -617
rect 20947 -663 21007 -642
rect 21065 -663 21125 -642
rect 21183 -643 21382 -642
rect 21183 -663 21243 -643
rect 21366 -651 21382 -643
rect 21416 -651 21432 -617
rect 17193 -722 17489 -686
rect 17193 -742 17253 -722
rect 17311 -742 17371 -722
rect 17429 -742 17489 -722
rect 17547 -722 17843 -686
rect 17547 -742 17607 -722
rect 17665 -742 17725 -722
rect 17783 -742 17843 -722
rect 17901 -721 18197 -685
rect 17901 -742 17961 -721
rect 18019 -742 18079 -721
rect 18137 -742 18197 -721
rect 17193 -968 17253 -942
rect 17311 -968 17371 -942
rect 17429 -974 17489 -942
rect 17547 -968 17607 -942
rect 17665 -968 17725 -942
rect 17783 -962 17843 -942
rect 17782 -968 17843 -962
rect 17901 -968 17961 -942
rect 18019 -968 18079 -942
rect 18137 -968 18197 -942
rect 17426 -990 17492 -974
rect 17426 -1024 17442 -990
rect 17476 -1024 17492 -990
rect 17426 -1040 17492 -1024
rect 14669 -1172 14730 -1083
rect 15222 -1096 15282 -1070
rect 15340 -1096 15400 -1070
rect 14669 -1225 14820 -1172
rect 14316 -1318 14702 -1267
rect 14521 -1376 14587 -1360
rect 14521 -1410 14537 -1376
rect 14571 -1410 14587 -1376
rect 14005 -1449 14065 -1423
rect 14123 -1449 14183 -1423
rect 14241 -1449 14301 -1423
rect 14521 -1426 14587 -1410
rect 14524 -1449 14584 -1426
rect 14642 -1449 14702 -1318
rect 14760 -1449 14820 -1225
rect 15458 -1271 15518 -1070
rect 15576 -1096 15636 -1070
rect 15694 -1096 15754 -1070
rect 15812 -1087 15872 -1070
rect 15811 -1176 15872 -1087
rect 17544 -1107 17610 -1091
rect 17544 -1141 17560 -1107
rect 17594 -1141 17610 -1107
rect 17544 -1157 17610 -1141
rect 15811 -1229 15962 -1176
rect 17547 -1179 17607 -1157
rect 17782 -1179 17842 -968
rect 17902 -1153 17960 -968
rect 21366 -667 21432 -651
rect 21735 -646 22031 -605
rect 21735 -667 21795 -646
rect 21853 -667 21913 -646
rect 21971 -667 22031 -646
rect 22089 -621 22562 -605
rect 22089 -646 22512 -621
rect 22089 -667 22149 -646
rect 22207 -667 22267 -646
rect 22325 -647 22512 -646
rect 22325 -667 22385 -647
rect 22496 -655 22512 -647
rect 22546 -655 22562 -621
rect 20593 -1089 20653 -1063
rect 20711 -1089 20771 -1063
rect 17900 -1179 17960 -1153
rect 15458 -1322 15844 -1271
rect 15663 -1380 15729 -1364
rect 15663 -1414 15679 -1380
rect 15713 -1414 15729 -1380
rect 11248 -1606 11308 -1584
rect 11366 -1606 11426 -1584
rect 11245 -1622 11311 -1606
rect 11245 -1656 11261 -1622
rect 11295 -1656 11311 -1622
rect 7471 -1727 8050 -1686
rect 8613 -1690 8673 -1658
rect 8731 -1690 8791 -1658
rect 8849 -1690 8909 -1658
rect 9132 -1690 9192 -1658
rect 9250 -1684 9310 -1658
rect 9368 -1684 9428 -1658
rect 11245 -1672 11311 -1656
rect 11363 -1622 11429 -1606
rect 11363 -1656 11379 -1622
rect 11413 -1656 11429 -1622
rect 15147 -1453 15207 -1427
rect 15265 -1453 15325 -1427
rect 15383 -1453 15443 -1427
rect 15663 -1430 15729 -1414
rect 15666 -1453 15726 -1430
rect 15784 -1453 15844 -1322
rect 15902 -1453 15962 -1229
rect 17547 -1405 17607 -1379
rect 11363 -1672 11429 -1656
rect 14005 -1681 14065 -1649
rect 14123 -1681 14183 -1649
rect 14241 -1681 14301 -1649
rect 14524 -1681 14584 -1649
rect 14642 -1675 14702 -1649
rect 14760 -1675 14820 -1649
rect 20829 -1264 20889 -1063
rect 20947 -1089 21007 -1063
rect 21065 -1089 21125 -1063
rect 21183 -1080 21243 -1063
rect 22496 -671 22562 -655
rect 23706 -719 24002 -683
rect 23706 -739 23766 -719
rect 23824 -739 23884 -719
rect 23942 -739 24002 -719
rect 24060 -719 24356 -683
rect 24060 -739 24120 -719
rect 24178 -739 24238 -719
rect 24296 -739 24356 -719
rect 24414 -718 24710 -682
rect 24414 -739 24474 -718
rect 24532 -739 24592 -718
rect 24650 -739 24710 -718
rect 23706 -965 23766 -939
rect 23824 -965 23884 -939
rect 23942 -971 24002 -939
rect 24060 -965 24120 -939
rect 24178 -965 24238 -939
rect 24296 -959 24356 -939
rect 24295 -965 24356 -959
rect 24414 -965 24474 -939
rect 24532 -965 24592 -939
rect 24650 -965 24710 -939
rect 23939 -987 24005 -971
rect 23939 -1021 23955 -987
rect 23989 -1021 24005 -987
rect 23939 -1037 24005 -1021
rect 21182 -1169 21243 -1080
rect 21735 -1093 21795 -1067
rect 21853 -1093 21913 -1067
rect 21182 -1222 21333 -1169
rect 20829 -1315 21215 -1264
rect 21034 -1373 21100 -1357
rect 21034 -1407 21050 -1373
rect 21084 -1407 21100 -1373
rect 20518 -1446 20578 -1420
rect 20636 -1446 20696 -1420
rect 20754 -1446 20814 -1420
rect 21034 -1423 21100 -1407
rect 21037 -1446 21097 -1423
rect 21155 -1446 21215 -1315
rect 21273 -1446 21333 -1222
rect 21971 -1268 22031 -1067
rect 22089 -1093 22149 -1067
rect 22207 -1093 22267 -1067
rect 22325 -1084 22385 -1067
rect 22324 -1173 22385 -1084
rect 24057 -1104 24123 -1088
rect 24057 -1138 24073 -1104
rect 24107 -1138 24123 -1104
rect 24057 -1154 24123 -1138
rect 22324 -1226 22475 -1173
rect 24060 -1176 24120 -1154
rect 24295 -1176 24355 -965
rect 24415 -1150 24473 -965
rect 24413 -1176 24473 -1150
rect 21971 -1319 22357 -1268
rect 22176 -1377 22242 -1361
rect 22176 -1411 22192 -1377
rect 22226 -1411 22242 -1377
rect 17782 -1601 17842 -1579
rect 17900 -1601 17960 -1579
rect 17779 -1617 17845 -1601
rect 17779 -1651 17795 -1617
rect 17829 -1651 17845 -1617
rect 8613 -1731 9192 -1690
rect 14005 -1722 14584 -1681
rect 15147 -1685 15207 -1653
rect 15265 -1685 15325 -1653
rect 15383 -1685 15443 -1653
rect 15666 -1685 15726 -1653
rect 15784 -1679 15844 -1653
rect 15902 -1679 15962 -1653
rect 17779 -1667 17845 -1651
rect 17897 -1617 17963 -1601
rect 17897 -1651 17913 -1617
rect 17947 -1651 17963 -1617
rect 21660 -1450 21720 -1424
rect 21778 -1450 21838 -1424
rect 21896 -1450 21956 -1424
rect 22176 -1427 22242 -1411
rect 22179 -1450 22239 -1427
rect 22297 -1450 22357 -1319
rect 22415 -1450 22475 -1226
rect 24060 -1402 24120 -1376
rect 17897 -1667 17963 -1651
rect 20518 -1678 20578 -1646
rect 20636 -1678 20696 -1646
rect 20754 -1678 20814 -1646
rect 21037 -1678 21097 -1646
rect 21155 -1672 21215 -1646
rect 21273 -1672 21333 -1646
rect 24295 -1598 24355 -1576
rect 24413 -1598 24473 -1576
rect 24292 -1614 24358 -1598
rect 24292 -1648 24308 -1614
rect 24342 -1648 24358 -1614
rect 15147 -1726 15726 -1685
rect 20518 -1719 21097 -1678
rect 21660 -1682 21720 -1650
rect 21778 -1682 21838 -1650
rect 21896 -1682 21956 -1650
rect 22179 -1682 22239 -1650
rect 22297 -1676 22357 -1650
rect 22415 -1676 22475 -1650
rect 24292 -1664 24358 -1648
rect 24410 -1614 24476 -1598
rect 24410 -1648 24426 -1614
rect 24460 -1648 24476 -1614
rect 24410 -1664 24476 -1648
rect 21660 -1723 22239 -1682
rect 4087 -2373 4383 -2337
rect 4087 -2393 4147 -2373
rect 4205 -2393 4265 -2373
rect 4323 -2393 4383 -2373
rect 4441 -2373 4737 -2337
rect 4441 -2393 4501 -2373
rect 4559 -2393 4619 -2373
rect 4677 -2393 4737 -2373
rect 4795 -2372 5091 -2336
rect 4795 -2393 4855 -2372
rect 4913 -2393 4973 -2372
rect 5031 -2393 5091 -2372
rect 10645 -2377 10941 -2341
rect 10645 -2397 10705 -2377
rect 10763 -2397 10823 -2377
rect 10881 -2397 10941 -2377
rect 10999 -2377 11295 -2341
rect 10999 -2397 11059 -2377
rect 11117 -2397 11177 -2377
rect 11235 -2397 11295 -2377
rect 11353 -2376 11649 -2340
rect 11353 -2397 11413 -2376
rect 11471 -2397 11531 -2376
rect 11589 -2397 11649 -2376
rect 4087 -2619 4147 -2593
rect 4205 -2619 4265 -2593
rect 4323 -2625 4383 -2593
rect 4441 -2619 4501 -2593
rect 4559 -2619 4619 -2593
rect 4677 -2613 4737 -2593
rect 4676 -2619 4737 -2613
rect 4795 -2619 4855 -2593
rect 4913 -2619 4973 -2593
rect 5031 -2619 5091 -2593
rect 17179 -2372 17475 -2336
rect 17179 -2392 17239 -2372
rect 17297 -2392 17357 -2372
rect 17415 -2392 17475 -2372
rect 17533 -2372 17829 -2336
rect 17533 -2392 17593 -2372
rect 17651 -2392 17711 -2372
rect 17769 -2392 17829 -2372
rect 17887 -2371 18183 -2335
rect 17887 -2392 17947 -2371
rect 18005 -2392 18065 -2371
rect 18123 -2392 18183 -2371
rect 23692 -2369 23988 -2333
rect 23692 -2389 23752 -2369
rect 23810 -2389 23870 -2369
rect 23928 -2389 23988 -2369
rect 24046 -2369 24342 -2333
rect 24046 -2389 24106 -2369
rect 24164 -2389 24224 -2369
rect 24282 -2389 24342 -2369
rect 24400 -2368 24696 -2332
rect 24400 -2389 24460 -2368
rect 24518 -2389 24578 -2368
rect 24636 -2389 24696 -2368
rect 4320 -2641 4386 -2625
rect 4320 -2675 4336 -2641
rect 4370 -2675 4386 -2641
rect 4320 -2691 4386 -2675
rect 595 -2810 655 -2784
rect 713 -2810 773 -2784
rect 831 -2810 891 -2784
rect 949 -2795 1245 -2744
rect 949 -2810 1009 -2795
rect 1067 -2810 1127 -2795
rect 1185 -2810 1245 -2795
rect 2493 -2810 2553 -2784
rect 2611 -2810 2671 -2784
rect 2729 -2810 2789 -2784
rect 2847 -2795 3143 -2744
rect 2847 -2810 2907 -2795
rect 2965 -2810 3025 -2795
rect 3083 -2810 3143 -2795
rect 4438 -2758 4504 -2742
rect 4438 -2792 4454 -2758
rect 4488 -2792 4504 -2758
rect 4438 -2808 4504 -2792
rect 112 -2993 408 -2942
rect 112 -3010 172 -2993
rect 230 -3010 290 -2993
rect 348 -3010 408 -2993
rect 1433 -3010 1493 -2984
rect 1551 -3010 1611 -2984
rect 1669 -3010 1729 -2984
rect 2010 -2993 2306 -2942
rect 2010 -3010 2070 -2993
rect 2128 -3010 2188 -2993
rect 2246 -3010 2306 -2993
rect 4441 -2830 4501 -2808
rect 4676 -2830 4736 -2619
rect 4796 -2804 4854 -2619
rect 10645 -2623 10705 -2597
rect 10763 -2623 10823 -2597
rect 10881 -2629 10941 -2597
rect 10999 -2623 11059 -2597
rect 11117 -2623 11177 -2597
rect 11235 -2617 11295 -2597
rect 11234 -2623 11295 -2617
rect 11353 -2623 11413 -2597
rect 11471 -2623 11531 -2597
rect 11589 -2623 11649 -2597
rect 17179 -2618 17239 -2592
rect 17297 -2618 17357 -2592
rect 10878 -2645 10944 -2629
rect 10878 -2679 10894 -2645
rect 10928 -2679 10944 -2645
rect 10878 -2695 10944 -2679
rect 4794 -2830 4854 -2804
rect 7153 -2814 7213 -2788
rect 7271 -2814 7331 -2788
rect 7389 -2814 7449 -2788
rect 7507 -2799 7803 -2748
rect 7507 -2814 7567 -2799
rect 7625 -2814 7685 -2799
rect 7743 -2814 7803 -2799
rect 9051 -2814 9111 -2788
rect 9169 -2814 9229 -2788
rect 9287 -2814 9347 -2788
rect 9405 -2799 9701 -2748
rect 9405 -2814 9465 -2799
rect 9523 -2814 9583 -2799
rect 9641 -2814 9701 -2799
rect 10996 -2762 11062 -2746
rect 10996 -2796 11012 -2762
rect 11046 -2796 11062 -2762
rect 10996 -2812 11062 -2796
rect 3331 -3010 3391 -2984
rect 3449 -3010 3509 -2984
rect 3567 -3010 3627 -2984
rect 4441 -3056 4501 -3030
rect 112 -3236 172 -3210
rect 230 -3229 290 -3210
rect 348 -3229 408 -3210
rect 595 -3229 655 -3210
rect 713 -3229 773 -3210
rect 831 -3229 891 -3210
rect 230 -3236 306 -3229
rect 231 -3280 306 -3236
rect 348 -3280 891 -3229
rect 949 -3236 1009 -3210
rect 1067 -3236 1127 -3210
rect 1185 -3227 1245 -3210
rect 1433 -3227 1493 -3210
rect 1551 -3227 1611 -3210
rect 1669 -3227 1729 -3210
rect 1185 -3278 1729 -3227
rect 2010 -3236 2070 -3210
rect 2128 -3229 2188 -3210
rect 2246 -3229 2306 -3210
rect 2493 -3229 2553 -3210
rect 2611 -3229 2671 -3210
rect 2729 -3229 2789 -3210
rect 2128 -3236 2204 -3229
rect 246 -3433 306 -3280
rect 52 -3457 306 -3433
rect 52 -3491 68 -3457
rect 102 -3491 306 -3457
rect 52 -3507 306 -3491
rect 652 -3479 948 -3419
rect 652 -3503 712 -3479
rect 770 -3503 830 -3479
rect 888 -3503 948 -3479
rect 1006 -3480 1302 -3420
rect 1006 -3503 1066 -3480
rect 1124 -3503 1184 -3480
rect 1242 -3503 1302 -3480
rect 246 -4131 306 -3507
rect 652 -3929 712 -3903
rect 622 -4069 689 -4062
rect 622 -4070 695 -4069
rect 770 -4070 830 -3903
rect 888 -3929 948 -3903
rect 1006 -3929 1066 -3903
rect 622 -4078 830 -4070
rect 622 -4112 638 -4078
rect 672 -4112 830 -4078
rect 622 -4128 830 -4112
rect 633 -4129 830 -4128
rect 246 -4147 396 -4131
rect 246 -4181 346 -4147
rect 380 -4181 396 -4147
rect 246 -4197 396 -4181
rect 246 -4235 306 -4197
rect 770 -4235 830 -4129
rect 1124 -4070 1184 -3903
rect 1242 -3929 1302 -3903
rect 1544 -3936 1604 -3278
rect 2129 -3280 2204 -3236
rect 2246 -3280 2789 -3229
rect 2847 -3236 2907 -3210
rect 2965 -3236 3025 -3210
rect 3083 -3227 3143 -3210
rect 3331 -3227 3391 -3210
rect 3449 -3227 3509 -3210
rect 3567 -3227 3627 -3210
rect 3083 -3278 3627 -3227
rect 6670 -2997 6966 -2946
rect 6670 -3014 6730 -2997
rect 6788 -3014 6848 -2997
rect 6906 -3014 6966 -2997
rect 7991 -3014 8051 -2988
rect 8109 -3014 8169 -2988
rect 8227 -3014 8287 -2988
rect 8568 -2997 8864 -2946
rect 8568 -3014 8628 -2997
rect 8686 -3014 8746 -2997
rect 8804 -3014 8864 -2997
rect 10999 -2834 11059 -2812
rect 11234 -2834 11294 -2623
rect 11354 -2808 11412 -2623
rect 17415 -2624 17475 -2592
rect 17533 -2618 17593 -2592
rect 17651 -2618 17711 -2592
rect 17769 -2612 17829 -2592
rect 17768 -2618 17829 -2612
rect 17887 -2618 17947 -2592
rect 18005 -2618 18065 -2592
rect 18123 -2618 18183 -2592
rect 23692 -2615 23752 -2589
rect 23810 -2615 23870 -2589
rect 17412 -2640 17478 -2624
rect 17412 -2674 17428 -2640
rect 17462 -2674 17478 -2640
rect 17412 -2690 17478 -2674
rect 11352 -2834 11412 -2808
rect 13687 -2809 13747 -2783
rect 13805 -2809 13865 -2783
rect 13923 -2809 13983 -2783
rect 14041 -2794 14337 -2743
rect 14041 -2809 14101 -2794
rect 14159 -2809 14219 -2794
rect 14277 -2809 14337 -2794
rect 15585 -2809 15645 -2783
rect 15703 -2809 15763 -2783
rect 15821 -2809 15881 -2783
rect 15939 -2794 16235 -2743
rect 15939 -2809 15999 -2794
rect 16057 -2809 16117 -2794
rect 16175 -2809 16235 -2794
rect 17530 -2757 17596 -2741
rect 17530 -2791 17546 -2757
rect 17580 -2791 17596 -2757
rect 17530 -2807 17596 -2791
rect 9889 -3014 9949 -2988
rect 10007 -3014 10067 -2988
rect 10125 -3014 10185 -2988
rect 10999 -3060 11059 -3034
rect 4676 -3246 4736 -3230
rect 1537 -3952 1604 -3936
rect 1537 -3986 1554 -3952
rect 1588 -3986 1604 -3952
rect 1537 -4002 1604 -3986
rect 1267 -4070 1334 -4063
rect 1124 -4079 1334 -4070
rect 1124 -4113 1284 -4079
rect 1318 -4113 1334 -4079
rect 1124 -4129 1334 -4113
rect 884 -4162 950 -4147
rect 884 -4196 900 -4162
rect 934 -4196 950 -4162
rect 884 -4212 950 -4196
rect 1002 -4163 1068 -4147
rect 1002 -4197 1018 -4163
rect 1052 -4197 1068 -4163
rect 888 -4235 948 -4212
rect 1002 -4213 1068 -4197
rect 1006 -4235 1066 -4213
rect 1124 -4235 1184 -4129
rect 1544 -4130 1604 -4002
rect 1453 -4146 1604 -4130
rect 1453 -4180 1469 -4146
rect 1503 -4180 1604 -4146
rect 1453 -4196 1604 -4180
rect 1544 -4235 1604 -4196
rect 2144 -3400 2204 -3280
rect 3442 -3359 3502 -3278
rect 4668 -3268 4742 -3246
rect 4794 -3252 4854 -3230
rect 6670 -3240 6730 -3214
rect 6788 -3233 6848 -3214
rect 6906 -3233 6966 -3214
rect 7153 -3233 7213 -3214
rect 7271 -3233 7331 -3214
rect 7389 -3233 7449 -3214
rect 6788 -3240 6864 -3233
rect 4668 -3302 4689 -3268
rect 4723 -3302 4742 -3268
rect 4668 -3359 4742 -3302
rect 4791 -3268 4857 -3252
rect 4791 -3302 4807 -3268
rect 4841 -3302 4857 -3268
rect 6789 -3284 6864 -3240
rect 6906 -3284 7449 -3233
rect 7507 -3240 7567 -3214
rect 7625 -3240 7685 -3214
rect 7743 -3231 7803 -3214
rect 7991 -3231 8051 -3214
rect 8109 -3231 8169 -3214
rect 8227 -3231 8287 -3214
rect 7743 -3282 8287 -3231
rect 8568 -3240 8628 -3214
rect 8686 -3233 8746 -3214
rect 8804 -3233 8864 -3214
rect 9051 -3233 9111 -3214
rect 9169 -3233 9229 -3214
rect 9287 -3233 9347 -3214
rect 8686 -3240 8762 -3233
rect 4791 -3318 4857 -3302
rect 3442 -3384 4742 -3359
rect 2144 -3420 2205 -3400
rect 2144 -3436 2224 -3420
rect 2144 -3470 2175 -3436
rect 2209 -3470 2224 -3436
rect 2144 -3486 2224 -3470
rect 2550 -3479 2846 -3419
rect 2144 -3509 2205 -3486
rect 2550 -3503 2610 -3479
rect 2668 -3503 2728 -3479
rect 2786 -3503 2846 -3479
rect 2904 -3480 3200 -3420
rect 2904 -3503 2964 -3480
rect 3022 -3503 3082 -3480
rect 3140 -3503 3200 -3480
rect 3442 -3432 4743 -3384
rect 2144 -3655 2204 -3509
rect 2144 -3828 2205 -3655
rect 2144 -4131 2204 -3828
rect 2550 -3929 2610 -3903
rect 2518 -4070 2585 -4063
rect 2668 -4070 2728 -3903
rect 2786 -3929 2846 -3903
rect 2904 -3929 2964 -3903
rect 2518 -4079 2728 -4070
rect 2518 -4113 2534 -4079
rect 2568 -4113 2728 -4079
rect 2518 -4129 2728 -4113
rect 2144 -4147 2294 -4131
rect 2144 -4181 2244 -4147
rect 2278 -4181 2294 -4147
rect 2144 -4197 2294 -4181
rect 2144 -4235 2204 -4197
rect 2668 -4235 2728 -4129
rect 3022 -4070 3082 -3903
rect 3140 -3929 3200 -3903
rect 3165 -4070 3232 -4063
rect 3022 -4079 3232 -4070
rect 3022 -4113 3182 -4079
rect 3216 -4113 3232 -4079
rect 3022 -4129 3232 -4113
rect 2782 -4162 2848 -4147
rect 2782 -4196 2798 -4162
rect 2832 -4196 2848 -4162
rect 2782 -4212 2848 -4196
rect 2900 -4163 2966 -4147
rect 2900 -4197 2916 -4163
rect 2950 -4197 2966 -4163
rect 2786 -4235 2846 -4212
rect 2900 -4213 2966 -4197
rect 2904 -4235 2964 -4213
rect 3022 -4235 3082 -4129
rect 3442 -4130 3502 -3432
rect 6804 -3437 6864 -3284
rect 6610 -3461 6864 -3437
rect 6610 -3495 6626 -3461
rect 6660 -3495 6864 -3461
rect 6610 -3511 6864 -3495
rect 7210 -3483 7506 -3423
rect 7210 -3507 7270 -3483
rect 7328 -3507 7388 -3483
rect 7446 -3507 7506 -3483
rect 7564 -3484 7860 -3424
rect 7564 -3507 7624 -3484
rect 7682 -3507 7742 -3484
rect 7800 -3507 7860 -3484
rect 4092 -3977 4388 -3941
rect 4092 -3997 4152 -3977
rect 4210 -3997 4270 -3977
rect 4328 -3997 4388 -3977
rect 4446 -3977 4742 -3941
rect 4446 -3997 4506 -3977
rect 4564 -3997 4624 -3977
rect 4682 -3997 4742 -3977
rect 4800 -3976 5096 -3940
rect 4800 -3997 4860 -3976
rect 4918 -3997 4978 -3976
rect 5036 -3997 5096 -3976
rect 3351 -4146 3502 -4130
rect 3351 -4180 3367 -4146
rect 3401 -4180 3502 -4146
rect 3351 -4196 3502 -4180
rect 3442 -4235 3502 -4196
rect 6804 -4135 6864 -3511
rect 7210 -3933 7270 -3907
rect 7180 -4073 7247 -4066
rect 7180 -4074 7253 -4073
rect 7328 -4074 7388 -3907
rect 7446 -3933 7506 -3907
rect 7564 -3933 7624 -3907
rect 7180 -4082 7388 -4074
rect 7180 -4116 7196 -4082
rect 7230 -4116 7388 -4082
rect 7180 -4132 7388 -4116
rect 7191 -4133 7388 -4132
rect 6804 -4151 6954 -4135
rect 6804 -4185 6904 -4151
rect 6938 -4185 6954 -4151
rect 4092 -4223 4152 -4197
rect 4210 -4223 4270 -4197
rect 4328 -4229 4388 -4197
rect 4446 -4223 4506 -4197
rect 4564 -4223 4624 -4197
rect 4682 -4217 4742 -4197
rect 4681 -4223 4742 -4217
rect 4800 -4223 4860 -4197
rect 4918 -4223 4978 -4197
rect 5036 -4223 5096 -4197
rect 6804 -4201 6954 -4185
rect 246 -4461 306 -4435
rect 1544 -4461 1604 -4435
rect 2144 -4461 2204 -4435
rect 4325 -4245 4391 -4229
rect 4325 -4279 4341 -4245
rect 4375 -4279 4391 -4245
rect 4325 -4295 4391 -4279
rect 4443 -4362 4509 -4346
rect 4443 -4396 4459 -4362
rect 4493 -4396 4509 -4362
rect 4443 -4412 4509 -4396
rect 4446 -4434 4506 -4412
rect 4681 -4434 4741 -4223
rect 4801 -4408 4859 -4223
rect 6804 -4239 6864 -4201
rect 7328 -4239 7388 -4133
rect 7682 -4074 7742 -3907
rect 7800 -3933 7860 -3907
rect 8102 -3940 8162 -3282
rect 8687 -3284 8762 -3240
rect 8804 -3284 9347 -3233
rect 9405 -3240 9465 -3214
rect 9523 -3240 9583 -3214
rect 9641 -3231 9701 -3214
rect 9889 -3231 9949 -3214
rect 10007 -3231 10067 -3214
rect 10125 -3231 10185 -3214
rect 9641 -3282 10185 -3231
rect 13204 -2992 13500 -2941
rect 13204 -3009 13264 -2992
rect 13322 -3009 13382 -2992
rect 13440 -3009 13500 -2992
rect 14525 -3009 14585 -2983
rect 14643 -3009 14703 -2983
rect 14761 -3009 14821 -2983
rect 15102 -2992 15398 -2941
rect 15102 -3009 15162 -2992
rect 15220 -3009 15280 -2992
rect 15338 -3009 15398 -2992
rect 17533 -2829 17593 -2807
rect 17768 -2829 17828 -2618
rect 17888 -2803 17946 -2618
rect 23928 -2621 23988 -2589
rect 24046 -2615 24106 -2589
rect 24164 -2615 24224 -2589
rect 24282 -2609 24342 -2589
rect 24281 -2615 24342 -2609
rect 24400 -2615 24460 -2589
rect 24518 -2615 24578 -2589
rect 24636 -2615 24696 -2589
rect 23925 -2637 23991 -2621
rect 23925 -2671 23941 -2637
rect 23975 -2671 23991 -2637
rect 23925 -2687 23991 -2671
rect 17886 -2829 17946 -2803
rect 20200 -2806 20260 -2780
rect 20318 -2806 20378 -2780
rect 20436 -2806 20496 -2780
rect 20554 -2791 20850 -2740
rect 20554 -2806 20614 -2791
rect 20672 -2806 20732 -2791
rect 20790 -2806 20850 -2791
rect 22098 -2806 22158 -2780
rect 22216 -2806 22276 -2780
rect 22334 -2806 22394 -2780
rect 22452 -2791 22748 -2740
rect 22452 -2806 22512 -2791
rect 22570 -2806 22630 -2791
rect 22688 -2806 22748 -2791
rect 24043 -2754 24109 -2738
rect 24043 -2788 24059 -2754
rect 24093 -2788 24109 -2754
rect 24043 -2804 24109 -2788
rect 16423 -3009 16483 -2983
rect 16541 -3009 16601 -2983
rect 16659 -3009 16719 -2983
rect 17533 -3055 17593 -3029
rect 11234 -3250 11294 -3234
rect 8095 -3956 8162 -3940
rect 8095 -3990 8112 -3956
rect 8146 -3990 8162 -3956
rect 8095 -4006 8162 -3990
rect 7825 -4074 7892 -4067
rect 7682 -4083 7892 -4074
rect 7682 -4117 7842 -4083
rect 7876 -4117 7892 -4083
rect 7682 -4133 7892 -4117
rect 7442 -4166 7508 -4151
rect 7442 -4200 7458 -4166
rect 7492 -4200 7508 -4166
rect 7442 -4216 7508 -4200
rect 7560 -4167 7626 -4151
rect 7560 -4201 7576 -4167
rect 7610 -4201 7626 -4167
rect 7446 -4239 7506 -4216
rect 7560 -4217 7626 -4201
rect 7564 -4239 7624 -4217
rect 7682 -4239 7742 -4133
rect 8102 -4134 8162 -4006
rect 8011 -4150 8162 -4134
rect 8011 -4184 8027 -4150
rect 8061 -4184 8162 -4150
rect 8011 -4200 8162 -4184
rect 8102 -4239 8162 -4200
rect 8702 -3404 8762 -3284
rect 10000 -3363 10060 -3282
rect 11226 -3272 11300 -3250
rect 11352 -3256 11412 -3234
rect 13204 -3235 13264 -3209
rect 13322 -3228 13382 -3209
rect 13440 -3228 13500 -3209
rect 13687 -3228 13747 -3209
rect 13805 -3228 13865 -3209
rect 13923 -3228 13983 -3209
rect 13322 -3235 13398 -3228
rect 11226 -3306 11247 -3272
rect 11281 -3306 11300 -3272
rect 11226 -3363 11300 -3306
rect 11349 -3272 11415 -3256
rect 11349 -3306 11365 -3272
rect 11399 -3306 11415 -3272
rect 13323 -3279 13398 -3235
rect 13440 -3279 13983 -3228
rect 14041 -3235 14101 -3209
rect 14159 -3235 14219 -3209
rect 14277 -3226 14337 -3209
rect 14525 -3226 14585 -3209
rect 14643 -3226 14703 -3209
rect 14761 -3226 14821 -3209
rect 14277 -3277 14821 -3226
rect 15102 -3235 15162 -3209
rect 15220 -3228 15280 -3209
rect 15338 -3228 15398 -3209
rect 15585 -3228 15645 -3209
rect 15703 -3228 15763 -3209
rect 15821 -3228 15881 -3209
rect 15220 -3235 15296 -3228
rect 11349 -3322 11415 -3306
rect 10000 -3388 11300 -3363
rect 8702 -3424 8763 -3404
rect 8702 -3440 8782 -3424
rect 8702 -3474 8733 -3440
rect 8767 -3474 8782 -3440
rect 8702 -3490 8782 -3474
rect 9108 -3483 9404 -3423
rect 8702 -3513 8763 -3490
rect 9108 -3507 9168 -3483
rect 9226 -3507 9286 -3483
rect 9344 -3507 9404 -3483
rect 9462 -3484 9758 -3424
rect 9462 -3507 9522 -3484
rect 9580 -3507 9640 -3484
rect 9698 -3507 9758 -3484
rect 10000 -3436 11301 -3388
rect 13338 -3432 13398 -3279
rect 8702 -3659 8762 -3513
rect 8702 -3832 8763 -3659
rect 8702 -4135 8762 -3832
rect 9108 -3933 9168 -3907
rect 9076 -4074 9143 -4067
rect 9226 -4074 9286 -3907
rect 9344 -3933 9404 -3907
rect 9462 -3933 9522 -3907
rect 9076 -4083 9286 -4074
rect 9076 -4117 9092 -4083
rect 9126 -4117 9286 -4083
rect 9076 -4133 9286 -4117
rect 8702 -4151 8852 -4135
rect 8702 -4185 8802 -4151
rect 8836 -4185 8852 -4151
rect 8702 -4201 8852 -4185
rect 8702 -4239 8762 -4201
rect 9226 -4239 9286 -4133
rect 9580 -4074 9640 -3907
rect 9698 -3933 9758 -3907
rect 9723 -4074 9790 -4067
rect 9580 -4083 9790 -4074
rect 9580 -4117 9740 -4083
rect 9774 -4117 9790 -4083
rect 9580 -4133 9790 -4117
rect 9340 -4166 9406 -4151
rect 9340 -4200 9356 -4166
rect 9390 -4200 9406 -4166
rect 9340 -4216 9406 -4200
rect 9458 -4167 9524 -4151
rect 9458 -4201 9474 -4167
rect 9508 -4201 9524 -4167
rect 9344 -4239 9404 -4216
rect 9458 -4217 9524 -4201
rect 9462 -4239 9522 -4217
rect 9580 -4239 9640 -4133
rect 10000 -4134 10060 -3436
rect 13144 -3456 13398 -3432
rect 13144 -3490 13160 -3456
rect 13194 -3490 13398 -3456
rect 13144 -3506 13398 -3490
rect 13744 -3478 14040 -3418
rect 13744 -3502 13804 -3478
rect 13862 -3502 13922 -3478
rect 13980 -3502 14040 -3478
rect 14098 -3479 14394 -3419
rect 14098 -3502 14158 -3479
rect 14216 -3502 14276 -3479
rect 14334 -3502 14394 -3479
rect 10650 -3981 10946 -3945
rect 10650 -4001 10710 -3981
rect 10768 -4001 10828 -3981
rect 10886 -4001 10946 -3981
rect 11004 -3981 11300 -3945
rect 11004 -4001 11064 -3981
rect 11122 -4001 11182 -3981
rect 11240 -4001 11300 -3981
rect 11358 -3980 11654 -3944
rect 11358 -4001 11418 -3980
rect 11476 -4001 11536 -3980
rect 11594 -4001 11654 -3980
rect 9909 -4150 10060 -4134
rect 9909 -4184 9925 -4150
rect 9959 -4184 10060 -4150
rect 9909 -4200 10060 -4184
rect 10000 -4239 10060 -4200
rect 13338 -4130 13398 -3506
rect 13744 -3928 13804 -3902
rect 13714 -4068 13781 -4061
rect 13714 -4069 13787 -4068
rect 13862 -4069 13922 -3902
rect 13980 -3928 14040 -3902
rect 14098 -3928 14158 -3902
rect 13714 -4077 13922 -4069
rect 13714 -4111 13730 -4077
rect 13764 -4111 13922 -4077
rect 13714 -4127 13922 -4111
rect 13725 -4128 13922 -4127
rect 13338 -4146 13488 -4130
rect 13338 -4180 13438 -4146
rect 13472 -4180 13488 -4146
rect 13338 -4196 13488 -4180
rect 10650 -4227 10710 -4201
rect 10768 -4227 10828 -4201
rect 10886 -4233 10946 -4201
rect 11004 -4227 11064 -4201
rect 11122 -4227 11182 -4201
rect 11240 -4221 11300 -4201
rect 11239 -4227 11300 -4221
rect 11358 -4227 11418 -4201
rect 11476 -4227 11536 -4201
rect 11594 -4227 11654 -4201
rect 4799 -4434 4859 -4408
rect 3442 -4461 3502 -4435
rect 770 -4661 830 -4635
rect 888 -4661 948 -4635
rect 1006 -4661 1066 -4635
rect 1124 -4661 1184 -4635
rect 2668 -4661 2728 -4635
rect 2786 -4661 2846 -4635
rect 2904 -4661 2964 -4635
rect 3022 -4661 3082 -4635
rect 4446 -4660 4506 -4634
rect 6804 -4465 6864 -4439
rect 8102 -4465 8162 -4439
rect 8702 -4465 8762 -4439
rect 10883 -4249 10949 -4233
rect 10883 -4283 10899 -4249
rect 10933 -4283 10949 -4249
rect 10883 -4299 10949 -4283
rect 11001 -4366 11067 -4350
rect 11001 -4400 11017 -4366
rect 11051 -4400 11067 -4366
rect 11001 -4416 11067 -4400
rect 11004 -4438 11064 -4416
rect 11239 -4438 11299 -4227
rect 11359 -4412 11417 -4227
rect 13338 -4234 13398 -4196
rect 13862 -4234 13922 -4128
rect 14216 -4069 14276 -3902
rect 14334 -3928 14394 -3902
rect 14636 -3935 14696 -3277
rect 15221 -3279 15296 -3235
rect 15338 -3279 15881 -3228
rect 15939 -3235 15999 -3209
rect 16057 -3235 16117 -3209
rect 16175 -3226 16235 -3209
rect 16423 -3226 16483 -3209
rect 16541 -3226 16601 -3209
rect 16659 -3226 16719 -3209
rect 16175 -3277 16719 -3226
rect 19717 -2989 20013 -2938
rect 19717 -3006 19777 -2989
rect 19835 -3006 19895 -2989
rect 19953 -3006 20013 -2989
rect 21038 -3006 21098 -2980
rect 21156 -3006 21216 -2980
rect 21274 -3006 21334 -2980
rect 21615 -2989 21911 -2938
rect 21615 -3006 21675 -2989
rect 21733 -3006 21793 -2989
rect 21851 -3006 21911 -2989
rect 24046 -2826 24106 -2804
rect 24281 -2826 24341 -2615
rect 24401 -2800 24459 -2615
rect 24399 -2826 24459 -2800
rect 22936 -3006 22996 -2980
rect 23054 -3006 23114 -2980
rect 23172 -3006 23232 -2980
rect 24046 -3052 24106 -3026
rect 17768 -3245 17828 -3229
rect 14629 -3951 14696 -3935
rect 14629 -3985 14646 -3951
rect 14680 -3985 14696 -3951
rect 14629 -4001 14696 -3985
rect 14359 -4069 14426 -4062
rect 14216 -4078 14426 -4069
rect 14216 -4112 14376 -4078
rect 14410 -4112 14426 -4078
rect 14216 -4128 14426 -4112
rect 13976 -4161 14042 -4146
rect 13976 -4195 13992 -4161
rect 14026 -4195 14042 -4161
rect 13976 -4211 14042 -4195
rect 14094 -4162 14160 -4146
rect 14094 -4196 14110 -4162
rect 14144 -4196 14160 -4162
rect 13980 -4234 14040 -4211
rect 14094 -4212 14160 -4196
rect 14098 -4234 14158 -4212
rect 14216 -4234 14276 -4128
rect 14636 -4129 14696 -4001
rect 14545 -4145 14696 -4129
rect 14545 -4179 14561 -4145
rect 14595 -4179 14696 -4145
rect 14545 -4195 14696 -4179
rect 14636 -4234 14696 -4195
rect 15236 -3399 15296 -3279
rect 16534 -3358 16594 -3277
rect 17760 -3267 17834 -3245
rect 17886 -3251 17946 -3229
rect 19717 -3232 19777 -3206
rect 19835 -3225 19895 -3206
rect 19953 -3225 20013 -3206
rect 20200 -3225 20260 -3206
rect 20318 -3225 20378 -3206
rect 20436 -3225 20496 -3206
rect 19835 -3232 19911 -3225
rect 17760 -3301 17781 -3267
rect 17815 -3301 17834 -3267
rect 17760 -3358 17834 -3301
rect 17883 -3267 17949 -3251
rect 17883 -3301 17899 -3267
rect 17933 -3301 17949 -3267
rect 19836 -3276 19911 -3232
rect 19953 -3276 20496 -3225
rect 20554 -3232 20614 -3206
rect 20672 -3232 20732 -3206
rect 20790 -3223 20850 -3206
rect 21038 -3223 21098 -3206
rect 21156 -3223 21216 -3206
rect 21274 -3223 21334 -3206
rect 20790 -3274 21334 -3223
rect 21615 -3232 21675 -3206
rect 21733 -3225 21793 -3206
rect 21851 -3225 21911 -3206
rect 22098 -3225 22158 -3206
rect 22216 -3225 22276 -3206
rect 22334 -3225 22394 -3206
rect 21733 -3232 21809 -3225
rect 17883 -3317 17949 -3301
rect 16534 -3383 17834 -3358
rect 15236 -3419 15297 -3399
rect 15236 -3435 15316 -3419
rect 15236 -3469 15267 -3435
rect 15301 -3469 15316 -3435
rect 15236 -3485 15316 -3469
rect 15642 -3478 15938 -3418
rect 15236 -3508 15297 -3485
rect 15642 -3502 15702 -3478
rect 15760 -3502 15820 -3478
rect 15878 -3502 15938 -3478
rect 15996 -3479 16292 -3419
rect 15996 -3502 16056 -3479
rect 16114 -3502 16174 -3479
rect 16232 -3502 16292 -3479
rect 16534 -3431 17835 -3383
rect 19851 -3429 19911 -3276
rect 15236 -3654 15296 -3508
rect 15236 -3827 15297 -3654
rect 15236 -4130 15296 -3827
rect 15642 -3928 15702 -3902
rect 15610 -4069 15677 -4062
rect 15760 -4069 15820 -3902
rect 15878 -3928 15938 -3902
rect 15996 -3928 16056 -3902
rect 15610 -4078 15820 -4069
rect 15610 -4112 15626 -4078
rect 15660 -4112 15820 -4078
rect 15610 -4128 15820 -4112
rect 15236 -4146 15386 -4130
rect 15236 -4180 15336 -4146
rect 15370 -4180 15386 -4146
rect 15236 -4196 15386 -4180
rect 15236 -4234 15296 -4196
rect 15760 -4234 15820 -4128
rect 16114 -4069 16174 -3902
rect 16232 -3928 16292 -3902
rect 16257 -4069 16324 -4062
rect 16114 -4078 16324 -4069
rect 16114 -4112 16274 -4078
rect 16308 -4112 16324 -4078
rect 16114 -4128 16324 -4112
rect 15874 -4161 15940 -4146
rect 15874 -4195 15890 -4161
rect 15924 -4195 15940 -4161
rect 15874 -4211 15940 -4195
rect 15992 -4162 16058 -4146
rect 15992 -4196 16008 -4162
rect 16042 -4196 16058 -4162
rect 15878 -4234 15938 -4211
rect 15992 -4212 16058 -4196
rect 15996 -4234 16056 -4212
rect 16114 -4234 16174 -4128
rect 16534 -4129 16594 -3431
rect 19657 -3453 19911 -3429
rect 19657 -3487 19673 -3453
rect 19707 -3487 19911 -3453
rect 19657 -3503 19911 -3487
rect 20257 -3475 20553 -3415
rect 20257 -3499 20317 -3475
rect 20375 -3499 20435 -3475
rect 20493 -3499 20553 -3475
rect 20611 -3476 20907 -3416
rect 20611 -3499 20671 -3476
rect 20729 -3499 20789 -3476
rect 20847 -3499 20907 -3476
rect 17184 -3976 17480 -3940
rect 17184 -3996 17244 -3976
rect 17302 -3996 17362 -3976
rect 17420 -3996 17480 -3976
rect 17538 -3976 17834 -3940
rect 17538 -3996 17598 -3976
rect 17656 -3996 17716 -3976
rect 17774 -3996 17834 -3976
rect 17892 -3975 18188 -3939
rect 17892 -3996 17952 -3975
rect 18010 -3996 18070 -3975
rect 18128 -3996 18188 -3975
rect 16443 -4145 16594 -4129
rect 16443 -4179 16459 -4145
rect 16493 -4179 16594 -4145
rect 16443 -4195 16594 -4179
rect 16534 -4234 16594 -4195
rect 19851 -4127 19911 -3503
rect 20257 -3925 20317 -3899
rect 20227 -4065 20294 -4058
rect 20227 -4066 20300 -4065
rect 20375 -4066 20435 -3899
rect 20493 -3925 20553 -3899
rect 20611 -3925 20671 -3899
rect 20227 -4074 20435 -4066
rect 20227 -4108 20243 -4074
rect 20277 -4108 20435 -4074
rect 20227 -4124 20435 -4108
rect 20238 -4125 20435 -4124
rect 19851 -4143 20001 -4127
rect 19851 -4177 19951 -4143
rect 19985 -4177 20001 -4143
rect 19851 -4193 20001 -4177
rect 17184 -4222 17244 -4196
rect 17302 -4222 17362 -4196
rect 17420 -4228 17480 -4196
rect 17538 -4222 17598 -4196
rect 17656 -4222 17716 -4196
rect 17774 -4216 17834 -4196
rect 17773 -4222 17834 -4216
rect 17892 -4222 17952 -4196
rect 18010 -4222 18070 -4196
rect 18128 -4222 18188 -4196
rect 11357 -4438 11417 -4412
rect 10000 -4465 10060 -4439
rect 7328 -4665 7388 -4639
rect 7446 -4665 7506 -4639
rect 7564 -4665 7624 -4639
rect 7682 -4665 7742 -4639
rect 9226 -4665 9286 -4639
rect 9344 -4665 9404 -4639
rect 9462 -4665 9522 -4639
rect 9580 -4665 9640 -4639
rect 11004 -4664 11064 -4638
rect 4681 -4856 4741 -4834
rect 4799 -4856 4859 -4834
rect 4678 -4872 4744 -4856
rect 4678 -4906 4694 -4872
rect 4728 -4906 4744 -4872
rect 4678 -4922 4744 -4906
rect 4796 -4872 4862 -4856
rect 4796 -4906 4812 -4872
rect 4846 -4906 4862 -4872
rect 13338 -4460 13398 -4434
rect 14636 -4460 14696 -4434
rect 15236 -4460 15296 -4434
rect 17417 -4244 17483 -4228
rect 17417 -4278 17433 -4244
rect 17467 -4278 17483 -4244
rect 17417 -4294 17483 -4278
rect 17535 -4361 17601 -4345
rect 17535 -4395 17551 -4361
rect 17585 -4395 17601 -4361
rect 17535 -4411 17601 -4395
rect 17538 -4433 17598 -4411
rect 17773 -4433 17833 -4222
rect 17893 -4407 17951 -4222
rect 19851 -4231 19911 -4193
rect 20375 -4231 20435 -4125
rect 20729 -4066 20789 -3899
rect 20847 -3925 20907 -3899
rect 21149 -3932 21209 -3274
rect 21734 -3276 21809 -3232
rect 21851 -3276 22394 -3225
rect 22452 -3232 22512 -3206
rect 22570 -3232 22630 -3206
rect 22688 -3223 22748 -3206
rect 22936 -3223 22996 -3206
rect 23054 -3223 23114 -3206
rect 23172 -3223 23232 -3206
rect 22688 -3274 23232 -3223
rect 24281 -3242 24341 -3226
rect 21142 -3948 21209 -3932
rect 21142 -3982 21159 -3948
rect 21193 -3982 21209 -3948
rect 21142 -3998 21209 -3982
rect 20872 -4066 20939 -4059
rect 20729 -4075 20939 -4066
rect 20729 -4109 20889 -4075
rect 20923 -4109 20939 -4075
rect 20729 -4125 20939 -4109
rect 20489 -4158 20555 -4143
rect 20489 -4192 20505 -4158
rect 20539 -4192 20555 -4158
rect 20489 -4208 20555 -4192
rect 20607 -4159 20673 -4143
rect 20607 -4193 20623 -4159
rect 20657 -4193 20673 -4159
rect 20493 -4231 20553 -4208
rect 20607 -4209 20673 -4193
rect 20611 -4231 20671 -4209
rect 20729 -4231 20789 -4125
rect 21149 -4126 21209 -3998
rect 21058 -4142 21209 -4126
rect 21058 -4176 21074 -4142
rect 21108 -4176 21209 -4142
rect 21058 -4192 21209 -4176
rect 21149 -4231 21209 -4192
rect 21749 -3396 21809 -3276
rect 23047 -3355 23107 -3274
rect 24273 -3264 24347 -3242
rect 24399 -3248 24459 -3226
rect 24273 -3298 24294 -3264
rect 24328 -3298 24347 -3264
rect 24273 -3355 24347 -3298
rect 24396 -3264 24462 -3248
rect 24396 -3298 24412 -3264
rect 24446 -3298 24462 -3264
rect 24396 -3314 24462 -3298
rect 23047 -3380 24347 -3355
rect 21749 -3416 21810 -3396
rect 21749 -3432 21829 -3416
rect 21749 -3466 21780 -3432
rect 21814 -3466 21829 -3432
rect 21749 -3482 21829 -3466
rect 22155 -3475 22451 -3415
rect 21749 -3505 21810 -3482
rect 22155 -3499 22215 -3475
rect 22273 -3499 22333 -3475
rect 22391 -3499 22451 -3475
rect 22509 -3476 22805 -3416
rect 22509 -3499 22569 -3476
rect 22627 -3499 22687 -3476
rect 22745 -3499 22805 -3476
rect 23047 -3428 24348 -3380
rect 21749 -3651 21809 -3505
rect 21749 -3824 21810 -3651
rect 21749 -4127 21809 -3824
rect 22155 -3925 22215 -3899
rect 22123 -4066 22190 -4059
rect 22273 -4066 22333 -3899
rect 22391 -3925 22451 -3899
rect 22509 -3925 22569 -3899
rect 22123 -4075 22333 -4066
rect 22123 -4109 22139 -4075
rect 22173 -4109 22333 -4075
rect 22123 -4125 22333 -4109
rect 21749 -4143 21899 -4127
rect 21749 -4177 21849 -4143
rect 21883 -4177 21899 -4143
rect 21749 -4193 21899 -4177
rect 21749 -4231 21809 -4193
rect 22273 -4231 22333 -4125
rect 22627 -4066 22687 -3899
rect 22745 -3925 22805 -3899
rect 22770 -4066 22837 -4059
rect 22627 -4075 22837 -4066
rect 22627 -4109 22787 -4075
rect 22821 -4109 22837 -4075
rect 22627 -4125 22837 -4109
rect 22387 -4158 22453 -4143
rect 22387 -4192 22403 -4158
rect 22437 -4192 22453 -4158
rect 22387 -4208 22453 -4192
rect 22505 -4159 22571 -4143
rect 22505 -4193 22521 -4159
rect 22555 -4193 22571 -4159
rect 22391 -4231 22451 -4208
rect 22505 -4209 22571 -4193
rect 22509 -4231 22569 -4209
rect 22627 -4231 22687 -4125
rect 23047 -4126 23107 -3428
rect 23697 -3973 23993 -3937
rect 23697 -3993 23757 -3973
rect 23815 -3993 23875 -3973
rect 23933 -3993 23993 -3973
rect 24051 -3973 24347 -3937
rect 24051 -3993 24111 -3973
rect 24169 -3993 24229 -3973
rect 24287 -3993 24347 -3973
rect 24405 -3972 24701 -3936
rect 24405 -3993 24465 -3972
rect 24523 -3993 24583 -3972
rect 24641 -3993 24701 -3972
rect 22956 -4142 23107 -4126
rect 22956 -4176 22972 -4142
rect 23006 -4176 23107 -4142
rect 22956 -4192 23107 -4176
rect 23047 -4231 23107 -4192
rect 23697 -4219 23757 -4193
rect 23815 -4219 23875 -4193
rect 23933 -4225 23993 -4193
rect 24051 -4219 24111 -4193
rect 24169 -4219 24229 -4193
rect 24287 -4213 24347 -4193
rect 24286 -4219 24347 -4213
rect 24405 -4219 24465 -4193
rect 24523 -4219 24583 -4193
rect 24641 -4219 24701 -4193
rect 17891 -4433 17951 -4407
rect 16534 -4460 16594 -4434
rect 13862 -4660 13922 -4634
rect 13980 -4660 14040 -4634
rect 14098 -4660 14158 -4634
rect 14216 -4660 14276 -4634
rect 15760 -4660 15820 -4634
rect 15878 -4660 15938 -4634
rect 15996 -4660 16056 -4634
rect 16114 -4660 16174 -4634
rect 17538 -4659 17598 -4633
rect 11239 -4860 11299 -4838
rect 11357 -4860 11417 -4838
rect 4796 -4922 4862 -4906
rect 11236 -4876 11302 -4860
rect 11236 -4910 11252 -4876
rect 11286 -4910 11302 -4876
rect 11236 -4926 11302 -4910
rect 11354 -4876 11420 -4860
rect 11354 -4910 11370 -4876
rect 11404 -4910 11420 -4876
rect 19851 -4457 19911 -4431
rect 21149 -4457 21209 -4431
rect 21749 -4457 21809 -4431
rect 23930 -4241 23996 -4225
rect 23930 -4275 23946 -4241
rect 23980 -4275 23996 -4241
rect 23930 -4291 23996 -4275
rect 24048 -4358 24114 -4342
rect 24048 -4392 24064 -4358
rect 24098 -4392 24114 -4358
rect 24048 -4408 24114 -4392
rect 24051 -4430 24111 -4408
rect 24286 -4430 24346 -4219
rect 24406 -4404 24464 -4219
rect 24404 -4430 24464 -4404
rect 23047 -4457 23107 -4431
rect 20375 -4657 20435 -4631
rect 20493 -4657 20553 -4631
rect 20611 -4657 20671 -4631
rect 20729 -4657 20789 -4631
rect 22273 -4657 22333 -4631
rect 22391 -4657 22451 -4631
rect 22509 -4657 22569 -4631
rect 22627 -4657 22687 -4631
rect 24051 -4656 24111 -4630
rect 17773 -4855 17833 -4833
rect 17891 -4855 17951 -4833
rect 11354 -4926 11420 -4910
rect 17770 -4871 17836 -4855
rect 17770 -4905 17786 -4871
rect 17820 -4905 17836 -4871
rect 17770 -4921 17836 -4905
rect 17888 -4871 17954 -4855
rect 17888 -4905 17904 -4871
rect 17938 -4905 17954 -4871
rect 24286 -4852 24346 -4830
rect 24404 -4852 24464 -4830
rect 17888 -4921 17954 -4905
rect 24283 -4868 24349 -4852
rect 24283 -4902 24299 -4868
rect 24333 -4902 24349 -4868
rect 24283 -4918 24349 -4902
rect 24401 -4868 24467 -4852
rect 24401 -4902 24417 -4868
rect 24451 -4902 24467 -4868
rect 24401 -4918 24467 -4902
<< polycont >>
rect 3141 5067 3175 5101
rect 4271 5073 4305 5107
rect 9654 5064 9688 5098
rect 10784 5070 10818 5104
rect 3141 4949 3175 4983
rect 4271 4953 4305 4987
rect 16188 5059 16222 5093
rect 17318 5065 17352 5099
rect 9654 4946 9688 4980
rect 1698 4583 1732 4617
rect 10784 4950 10818 4984
rect 22746 5063 22780 5097
rect 23876 5069 23910 5103
rect 16188 4941 16222 4975
rect 1580 4466 1614 4500
rect 3461 4193 3495 4227
rect 8211 4580 8245 4614
rect 17318 4945 17352 4979
rect 22746 4945 22780 4979
rect 8093 4463 8127 4497
rect 4603 4197 4637 4231
rect 1227 3956 1261 3990
rect 1345 3956 1379 3990
rect 9974 4190 10008 4224
rect 14745 4575 14779 4609
rect 23876 4949 23910 4983
rect 14627 4458 14661 4492
rect 11116 4194 11150 4228
rect 7740 3953 7774 3987
rect 7858 3953 7892 3987
rect 16508 4185 16542 4219
rect 21303 4579 21337 4613
rect 21185 4462 21219 4496
rect 17650 4189 17684 4223
rect 14274 3948 14308 3982
rect 14392 3948 14426 3982
rect 23066 4189 23100 4223
rect 24208 4193 24242 4227
rect 20832 3952 20866 3986
rect 20950 3952 20984 3986
rect 1712 2933 1746 2967
rect 1594 2816 1628 2850
rect 1241 2306 1275 2340
rect 1359 2306 1393 2340
rect 8225 2930 8259 2964
rect 8107 2813 8141 2847
rect 3873 2138 3907 2172
rect 2866 1495 2900 1529
rect 2681 1428 2715 1462
rect 3514 1495 3548 1529
rect 3132 1411 3166 1445
rect 3250 1412 3284 1446
rect 3804 1427 3838 1461
rect 7754 2303 7788 2337
rect 7872 2303 7906 2337
rect 14759 2925 14793 2959
rect 14641 2808 14675 2842
rect 5980 2117 6014 2151
rect 4494 1622 4528 1656
rect 4764 1495 4798 1529
rect 4579 1428 4613 1462
rect 5410 1496 5444 1530
rect 5030 1411 5064 1445
rect 5148 1412 5182 1446
rect 5702 1427 5736 1461
rect 10386 2135 10420 2169
rect 9379 1492 9413 1526
rect 9194 1425 9228 1459
rect 1707 1329 1741 1363
rect 1589 1212 1623 1246
rect 10027 1492 10061 1526
rect 9645 1408 9679 1442
rect 9763 1409 9797 1443
rect 10317 1424 10351 1458
rect 14288 2298 14322 2332
rect 14406 2298 14440 2332
rect 21317 2929 21351 2963
rect 21199 2812 21233 2846
rect 12493 2114 12527 2148
rect 11007 1619 11041 1653
rect 11277 1492 11311 1526
rect 11092 1425 11126 1459
rect 11923 1493 11957 1527
rect 11543 1408 11577 1442
rect 11661 1409 11695 1443
rect 12215 1424 12249 1458
rect 16920 2130 16954 2164
rect 15913 1487 15947 1521
rect 15728 1420 15762 1454
rect 8220 1326 8254 1360
rect 8102 1209 8136 1243
rect 1236 702 1270 736
rect 1354 702 1388 736
rect 16561 1487 16595 1521
rect 16179 1403 16213 1437
rect 16297 1404 16331 1438
rect 16851 1419 16885 1453
rect 20846 2302 20880 2336
rect 20964 2302 20998 2336
rect 19027 2109 19061 2143
rect 17541 1614 17575 1648
rect 17811 1487 17845 1521
rect 17626 1420 17660 1454
rect 18457 1488 18491 1522
rect 18077 1403 18111 1437
rect 18195 1404 18229 1438
rect 18749 1419 18783 1453
rect 23478 2134 23512 2168
rect 22471 1491 22505 1525
rect 22286 1424 22320 1458
rect 14754 1321 14788 1355
rect 14636 1204 14670 1238
rect 7749 699 7783 733
rect 7867 699 7901 733
rect 23119 1491 23153 1525
rect 22737 1407 22771 1441
rect 22855 1408 22889 1442
rect 23409 1423 23443 1457
rect 25585 2113 25619 2147
rect 24099 1618 24133 1652
rect 24369 1491 24403 1525
rect 24184 1424 24218 1458
rect 25015 1492 25049 1526
rect 24635 1407 24669 1441
rect 24753 1408 24787 1442
rect 25307 1423 25341 1457
rect 21312 1325 21346 1359
rect 21194 1208 21228 1242
rect 14283 694 14317 728
rect 14401 694 14435 728
rect 20841 698 20875 732
rect 20959 698 20993 732
rect 1777 -535 1811 -501
rect 2907 -541 2941 -507
rect 8335 -539 8369 -505
rect 9465 -545 9499 -511
rect 1777 -655 1811 -621
rect 2907 -659 2941 -625
rect 14869 -534 14903 -500
rect 15999 -540 16033 -506
rect 8335 -659 8369 -625
rect 4350 -1025 4384 -991
rect 1445 -1411 1479 -1377
rect 4468 -1142 4502 -1108
rect 9465 -663 9499 -629
rect 2587 -1415 2621 -1381
rect 21382 -531 21416 -497
rect 22512 -537 22546 -503
rect 14869 -654 14903 -620
rect 10908 -1029 10942 -995
rect 8003 -1415 8037 -1381
rect 11026 -1146 11060 -1112
rect 15999 -658 16033 -624
rect 9145 -1419 9179 -1385
rect 4703 -1652 4737 -1618
rect 4821 -1652 4855 -1618
rect 21382 -651 21416 -617
rect 17442 -1024 17476 -990
rect 14537 -1410 14571 -1376
rect 17560 -1141 17594 -1107
rect 22512 -655 22546 -621
rect 15679 -1414 15713 -1380
rect 11261 -1656 11295 -1622
rect 11379 -1656 11413 -1622
rect 23955 -1021 23989 -987
rect 21050 -1407 21084 -1373
rect 24073 -1138 24107 -1104
rect 22192 -1411 22226 -1377
rect 17795 -1651 17829 -1617
rect 17913 -1651 17947 -1617
rect 24308 -1648 24342 -1614
rect 24426 -1648 24460 -1614
rect 4336 -2675 4370 -2641
rect 4454 -2792 4488 -2758
rect 10894 -2679 10928 -2645
rect 11012 -2796 11046 -2762
rect 68 -3491 102 -3457
rect 638 -4112 672 -4078
rect 346 -4181 380 -4147
rect 17428 -2674 17462 -2640
rect 17546 -2791 17580 -2757
rect 1554 -3986 1588 -3952
rect 1284 -4113 1318 -4079
rect 900 -4196 934 -4162
rect 1018 -4197 1052 -4163
rect 1469 -4180 1503 -4146
rect 4689 -3302 4723 -3268
rect 4807 -3302 4841 -3268
rect 2175 -3470 2209 -3436
rect 2534 -4113 2568 -4079
rect 2244 -4181 2278 -4147
rect 3182 -4113 3216 -4079
rect 2798 -4196 2832 -4162
rect 2916 -4197 2950 -4163
rect 6626 -3495 6660 -3461
rect 3367 -4180 3401 -4146
rect 7196 -4116 7230 -4082
rect 6904 -4185 6938 -4151
rect 4341 -4279 4375 -4245
rect 4459 -4396 4493 -4362
rect 23941 -2671 23975 -2637
rect 24059 -2788 24093 -2754
rect 8112 -3990 8146 -3956
rect 7842 -4117 7876 -4083
rect 7458 -4200 7492 -4166
rect 7576 -4201 7610 -4167
rect 8027 -4184 8061 -4150
rect 11247 -3306 11281 -3272
rect 11365 -3306 11399 -3272
rect 8733 -3474 8767 -3440
rect 9092 -4117 9126 -4083
rect 8802 -4185 8836 -4151
rect 9740 -4117 9774 -4083
rect 9356 -4200 9390 -4166
rect 9474 -4201 9508 -4167
rect 13160 -3490 13194 -3456
rect 9925 -4184 9959 -4150
rect 13730 -4111 13764 -4077
rect 13438 -4180 13472 -4146
rect 10899 -4283 10933 -4249
rect 11017 -4400 11051 -4366
rect 14646 -3985 14680 -3951
rect 14376 -4112 14410 -4078
rect 13992 -4195 14026 -4161
rect 14110 -4196 14144 -4162
rect 14561 -4179 14595 -4145
rect 17781 -3301 17815 -3267
rect 17899 -3301 17933 -3267
rect 15267 -3469 15301 -3435
rect 15626 -4112 15660 -4078
rect 15336 -4180 15370 -4146
rect 16274 -4112 16308 -4078
rect 15890 -4195 15924 -4161
rect 16008 -4196 16042 -4162
rect 19673 -3487 19707 -3453
rect 16459 -4179 16493 -4145
rect 20243 -4108 20277 -4074
rect 19951 -4177 19985 -4143
rect 4694 -4906 4728 -4872
rect 4812 -4906 4846 -4872
rect 17433 -4278 17467 -4244
rect 17551 -4395 17585 -4361
rect 21159 -3982 21193 -3948
rect 20889 -4109 20923 -4075
rect 20505 -4192 20539 -4158
rect 20623 -4193 20657 -4159
rect 21074 -4176 21108 -4142
rect 24294 -3298 24328 -3264
rect 24412 -3298 24446 -3264
rect 21780 -3466 21814 -3432
rect 22139 -4109 22173 -4075
rect 21849 -4177 21883 -4143
rect 22787 -4109 22821 -4075
rect 22403 -4192 22437 -4158
rect 22521 -4193 22555 -4159
rect 22972 -4176 23006 -4142
rect 11252 -4910 11286 -4876
rect 11370 -4910 11404 -4876
rect 23946 -4275 23980 -4241
rect 24064 -4392 24098 -4358
rect 17786 -4905 17820 -4871
rect 17904 -4905 17938 -4871
rect 24299 -4902 24333 -4868
rect 24417 -4902 24451 -4868
<< locali >>
rect 1326 5267 1549 5343
rect 1326 5118 1405 5267
rect 1472 5118 1549 5267
rect 1326 5012 1549 5118
rect 3808 5321 4031 5397
rect 3808 5172 3887 5321
rect 3954 5172 4031 5321
rect 3141 5101 3175 5117
rect 3141 5051 3175 5067
rect 3808 5066 4031 5172
rect 4955 5321 5178 5397
rect 4955 5172 5034 5321
rect 5101 5172 5178 5321
rect 4271 5107 4305 5123
rect 4271 5057 4305 5073
rect 4955 5066 5178 5172
rect 7839 5264 8062 5340
rect 7839 5115 7918 5264
rect 7985 5115 8062 5264
rect 7839 5009 8062 5115
rect 10321 5318 10544 5394
rect 10321 5169 10400 5318
rect 10467 5169 10544 5318
rect 9654 5098 9688 5114
rect 9654 5048 9688 5064
rect 10321 5063 10544 5169
rect 11468 5318 11691 5394
rect 11468 5169 11547 5318
rect 11614 5169 11691 5318
rect 10784 5104 10818 5120
rect 10784 5054 10818 5070
rect 11468 5063 11691 5169
rect 14373 5259 14596 5335
rect 14373 5110 14452 5259
rect 14519 5110 14596 5259
rect 14373 5004 14596 5110
rect 16855 5313 17078 5389
rect 16855 5164 16934 5313
rect 17001 5164 17078 5313
rect 16188 5093 16222 5109
rect 16188 5043 16222 5059
rect 16855 5058 17078 5164
rect 18002 5313 18225 5389
rect 18002 5164 18081 5313
rect 18148 5164 18225 5313
rect 17318 5099 17352 5115
rect 17318 5049 17352 5065
rect 18002 5058 18225 5164
rect 20931 5263 21154 5339
rect 20931 5114 21010 5263
rect 21077 5114 21154 5263
rect 20931 5008 21154 5114
rect 23413 5317 23636 5393
rect 23413 5168 23492 5317
rect 23559 5168 23636 5317
rect 22746 5097 22780 5113
rect 22746 5047 22780 5063
rect 23413 5062 23636 5168
rect 24560 5317 24783 5393
rect 24560 5168 24639 5317
rect 24706 5168 24783 5317
rect 23876 5103 23910 5119
rect 23876 5053 23910 5069
rect 24560 5062 24783 5168
rect 3141 4983 3175 4999
rect 1757 4903 2027 4937
rect 3141 4933 3175 4949
rect 4271 4987 4305 5003
rect 931 4853 965 4869
rect 931 4661 965 4677
rect 1049 4853 1083 4869
rect 1049 4661 1083 4677
rect 1167 4853 1201 4869
rect 1167 4661 1201 4677
rect 1285 4853 1319 4869
rect 1285 4661 1319 4677
rect 1403 4853 1437 4869
rect 1403 4661 1437 4677
rect 1521 4853 1555 4869
rect 1521 4661 1555 4677
rect 1639 4853 1673 4869
rect 1639 4661 1673 4677
rect 1757 4853 1791 4903
rect 1757 4661 1791 4677
rect 1875 4853 1909 4869
rect 1875 4661 1909 4677
rect 1993 4853 2027 4903
rect 1993 4661 2027 4677
rect 3256 4925 3290 4941
rect 1682 4583 1698 4617
rect 1732 4583 1748 4617
rect 3256 4533 3290 4549
rect 3374 4925 3408 4941
rect 3374 4533 3408 4549
rect 3492 4925 3526 4941
rect 3492 4533 3526 4549
rect 3610 4925 3644 4941
rect 3610 4533 3644 4549
rect 3728 4925 3762 4941
rect 3728 4533 3762 4549
rect 3846 4925 3880 4941
rect 3846 4533 3880 4549
rect 3964 4925 3998 4941
rect 4271 4937 4305 4953
rect 9654 4980 9688 4996
rect 3964 4533 3998 4549
rect 4398 4929 4432 4945
rect 4398 4537 4432 4553
rect 4516 4929 4550 4945
rect 4516 4537 4550 4553
rect 4634 4929 4668 4945
rect 4634 4537 4668 4553
rect 4752 4929 4786 4945
rect 4752 4537 4786 4553
rect 4870 4929 4904 4945
rect 4870 4537 4904 4553
rect 4988 4929 5022 4945
rect 4988 4537 5022 4553
rect 5106 4929 5140 4945
rect 8270 4900 8540 4934
rect 9654 4930 9688 4946
rect 10784 4984 10818 5000
rect 7444 4850 7478 4866
rect 7444 4658 7478 4674
rect 7562 4850 7596 4866
rect 7562 4658 7596 4674
rect 7680 4850 7714 4866
rect 7680 4658 7714 4674
rect 7798 4850 7832 4866
rect 7798 4658 7832 4674
rect 7916 4850 7950 4866
rect 7916 4658 7950 4674
rect 8034 4850 8068 4866
rect 8034 4658 8068 4674
rect 8152 4850 8186 4866
rect 8152 4658 8186 4674
rect 8270 4850 8304 4900
rect 8270 4658 8304 4674
rect 8388 4850 8422 4866
rect 8388 4658 8422 4674
rect 8506 4850 8540 4900
rect 8506 4658 8540 4674
rect 9769 4922 9803 4938
rect 8195 4580 8211 4614
rect 8245 4580 8261 4614
rect 5106 4537 5140 4553
rect 9769 4530 9803 4546
rect 9887 4922 9921 4938
rect 9887 4530 9921 4546
rect 10005 4922 10039 4938
rect 10005 4530 10039 4546
rect 10123 4922 10157 4938
rect 10123 4530 10157 4546
rect 10241 4922 10275 4938
rect 10241 4530 10275 4546
rect 10359 4922 10393 4938
rect 10359 4530 10393 4546
rect 10477 4922 10511 4938
rect 10784 4934 10818 4950
rect 16188 4975 16222 4991
rect 10477 4530 10511 4546
rect 10911 4926 10945 4942
rect 10911 4534 10945 4550
rect 11029 4926 11063 4942
rect 11029 4534 11063 4550
rect 11147 4926 11181 4942
rect 11147 4534 11181 4550
rect 11265 4926 11299 4942
rect 11265 4534 11299 4550
rect 11383 4926 11417 4942
rect 11383 4534 11417 4550
rect 11501 4926 11535 4942
rect 11501 4534 11535 4550
rect 11619 4926 11653 4942
rect 14804 4895 15074 4929
rect 16188 4925 16222 4941
rect 17318 4979 17352 4995
rect 13978 4845 14012 4861
rect 13978 4653 14012 4669
rect 14096 4845 14130 4861
rect 14096 4653 14130 4669
rect 14214 4845 14248 4861
rect 14214 4653 14248 4669
rect 14332 4845 14366 4861
rect 14332 4653 14366 4669
rect 14450 4845 14484 4861
rect 14450 4653 14484 4669
rect 14568 4845 14602 4861
rect 14568 4653 14602 4669
rect 14686 4845 14720 4861
rect 14686 4653 14720 4669
rect 14804 4845 14838 4895
rect 14804 4653 14838 4669
rect 14922 4845 14956 4861
rect 14922 4653 14956 4669
rect 15040 4845 15074 4895
rect 15040 4653 15074 4669
rect 16303 4917 16337 4933
rect 14729 4575 14745 4609
rect 14779 4575 14795 4609
rect 11619 4534 11653 4550
rect 16303 4525 16337 4541
rect 16421 4917 16455 4933
rect 16421 4525 16455 4541
rect 16539 4917 16573 4933
rect 16539 4525 16573 4541
rect 16657 4917 16691 4933
rect 16657 4525 16691 4541
rect 16775 4917 16809 4933
rect 16775 4525 16809 4541
rect 16893 4917 16927 4933
rect 16893 4525 16927 4541
rect 17011 4917 17045 4933
rect 17318 4929 17352 4945
rect 22746 4979 22780 4995
rect 17011 4525 17045 4541
rect 17445 4921 17479 4937
rect 17445 4529 17479 4545
rect 17563 4921 17597 4937
rect 17563 4529 17597 4545
rect 17681 4921 17715 4937
rect 17681 4529 17715 4545
rect 17799 4921 17833 4937
rect 17799 4529 17833 4545
rect 17917 4921 17951 4937
rect 17917 4529 17951 4545
rect 18035 4921 18069 4937
rect 18035 4529 18069 4545
rect 18153 4921 18187 4937
rect 21362 4899 21632 4933
rect 22746 4929 22780 4945
rect 23876 4983 23910 4999
rect 20536 4849 20570 4865
rect 20536 4657 20570 4673
rect 20654 4849 20688 4865
rect 20654 4657 20688 4673
rect 20772 4849 20806 4865
rect 20772 4657 20806 4673
rect 20890 4849 20924 4865
rect 20890 4657 20924 4673
rect 21008 4849 21042 4865
rect 21008 4657 21042 4673
rect 21126 4849 21160 4865
rect 21126 4657 21160 4673
rect 21244 4849 21278 4865
rect 21244 4657 21278 4673
rect 21362 4849 21396 4899
rect 21362 4657 21396 4673
rect 21480 4849 21514 4865
rect 21480 4657 21514 4673
rect 21598 4849 21632 4899
rect 21598 4657 21632 4673
rect 22861 4921 22895 4937
rect 21287 4579 21303 4613
rect 21337 4579 21353 4613
rect 18153 4529 18187 4545
rect 22861 4529 22895 4545
rect 22979 4921 23013 4937
rect 22979 4529 23013 4545
rect 23097 4921 23131 4937
rect 23097 4529 23131 4545
rect 23215 4921 23249 4937
rect 23215 4529 23249 4545
rect 23333 4921 23367 4937
rect 23333 4529 23367 4545
rect 23451 4921 23485 4937
rect 23451 4529 23485 4545
rect 23569 4921 23603 4937
rect 23876 4933 23910 4949
rect 23569 4529 23603 4545
rect 24003 4925 24037 4941
rect 24003 4533 24037 4549
rect 24121 4925 24155 4941
rect 24121 4533 24155 4549
rect 24239 4925 24273 4941
rect 24239 4533 24273 4549
rect 24357 4925 24391 4941
rect 24357 4533 24391 4549
rect 24475 4925 24509 4941
rect 24475 4533 24509 4549
rect 24593 4925 24627 4941
rect 24593 4533 24627 4549
rect 24711 4925 24745 4941
rect 24711 4533 24745 4549
rect 1564 4466 1580 4500
rect 1614 4466 1630 4500
rect 8077 4463 8093 4497
rect 8127 4463 8143 4497
rect 14611 4458 14627 4492
rect 14661 4458 14677 4492
rect 21169 4462 21185 4496
rect 21219 4462 21235 4496
rect 1168 4416 1202 4432
rect 1168 4024 1202 4040
rect 1286 4416 1320 4432
rect 1286 4024 1320 4040
rect 1404 4416 1438 4432
rect 1521 4416 1555 4432
rect 1521 4224 1555 4240
rect 1639 4416 1673 4432
rect 1639 4224 1673 4240
rect 7681 4413 7715 4429
rect 3445 4193 3461 4227
rect 3495 4193 3511 4227
rect 4587 4197 4603 4231
rect 4637 4197 4653 4231
rect 3166 4142 3200 4158
rect 1404 4024 1438 4040
rect 1691 4090 1940 4133
rect 1691 4000 1738 4090
rect 1901 4000 1940 4090
rect 1211 3956 1227 3990
rect 1261 3956 1277 3990
rect 1329 3956 1345 3990
rect 1379 3956 1395 3990
rect 1691 3961 1940 4000
rect 3166 3950 3200 3966
rect 3284 4142 3318 4158
rect 3284 3950 3318 3966
rect 3402 4142 3436 4158
rect 3402 3950 3436 3966
rect 3520 4142 3554 4158
rect 3520 3950 3554 3966
rect 3685 4142 3719 4158
rect 3685 3950 3719 3966
rect 3803 4142 3837 4158
rect 3803 3950 3837 3966
rect 3921 4142 3955 4158
rect 3921 3950 3955 3966
rect 4039 4142 4073 4158
rect 4039 3950 4073 3966
rect 4308 4146 4342 4162
rect 4308 3954 4342 3970
rect 4426 4146 4460 4162
rect 4426 3954 4460 3970
rect 4544 4146 4578 4162
rect 4544 3954 4578 3970
rect 4662 4146 4696 4162
rect 4662 3954 4696 3970
rect 4827 4146 4861 4162
rect 4827 3954 4861 3970
rect 4945 4146 4979 4162
rect 4945 3954 4979 3970
rect 5063 4146 5097 4162
rect 5063 3954 5097 3970
rect 5181 4146 5215 4162
rect 7681 4021 7715 4037
rect 7799 4413 7833 4429
rect 7799 4021 7833 4037
rect 7917 4413 7951 4429
rect 8034 4413 8068 4429
rect 8034 4221 8068 4237
rect 8152 4413 8186 4429
rect 8152 4221 8186 4237
rect 14215 4408 14249 4424
rect 9958 4190 9974 4224
rect 10008 4190 10024 4224
rect 11100 4194 11116 4228
rect 11150 4194 11166 4228
rect 9679 4139 9713 4155
rect 7917 4021 7951 4037
rect 8204 4087 8453 4130
rect 8204 3997 8251 4087
rect 8414 3997 8453 4087
rect 5181 3954 5215 3970
rect 7724 3953 7740 3987
rect 7774 3953 7790 3987
rect 7842 3953 7858 3987
rect 7892 3953 7908 3987
rect 8204 3958 8453 3997
rect 9679 3947 9713 3963
rect 9797 4139 9831 4155
rect 9797 3947 9831 3963
rect 9915 4139 9949 4155
rect 9915 3947 9949 3963
rect 10033 4139 10067 4155
rect 10033 3947 10067 3963
rect 10198 4139 10232 4155
rect 10198 3947 10232 3963
rect 10316 4139 10350 4155
rect 10316 3947 10350 3963
rect 10434 4139 10468 4155
rect 10434 3947 10468 3963
rect 10552 4139 10586 4155
rect 10552 3947 10586 3963
rect 10821 4143 10855 4159
rect 10821 3951 10855 3967
rect 10939 4143 10973 4159
rect 10939 3951 10973 3967
rect 11057 4143 11091 4159
rect 11057 3951 11091 3967
rect 11175 4143 11209 4159
rect 11175 3951 11209 3967
rect 11340 4143 11374 4159
rect 11340 3951 11374 3967
rect 11458 4143 11492 4159
rect 11458 3951 11492 3967
rect 11576 4143 11610 4159
rect 11576 3951 11610 3967
rect 11694 4143 11728 4159
rect 14215 4016 14249 4032
rect 14333 4408 14367 4424
rect 14333 4016 14367 4032
rect 14451 4408 14485 4424
rect 14568 4408 14602 4424
rect 14568 4216 14602 4232
rect 14686 4408 14720 4424
rect 14686 4216 14720 4232
rect 20773 4412 20807 4428
rect 16492 4185 16508 4219
rect 16542 4185 16558 4219
rect 17634 4189 17650 4223
rect 17684 4189 17700 4223
rect 16213 4134 16247 4150
rect 14451 4016 14485 4032
rect 14738 4082 14987 4125
rect 14738 3992 14785 4082
rect 14948 3992 14987 4082
rect 11694 3951 11728 3967
rect 14258 3948 14274 3982
rect 14308 3948 14324 3982
rect 14376 3948 14392 3982
rect 14426 3948 14442 3982
rect 14738 3953 14987 3992
rect 16213 3942 16247 3958
rect 16331 4134 16365 4150
rect 16331 3942 16365 3958
rect 16449 4134 16483 4150
rect 16449 3942 16483 3958
rect 16567 4134 16601 4150
rect 16567 3942 16601 3958
rect 16732 4134 16766 4150
rect 16732 3942 16766 3958
rect 16850 4134 16884 4150
rect 16850 3942 16884 3958
rect 16968 4134 17002 4150
rect 16968 3942 17002 3958
rect 17086 4134 17120 4150
rect 17086 3942 17120 3958
rect 17355 4138 17389 4154
rect 17355 3946 17389 3962
rect 17473 4138 17507 4154
rect 17473 3946 17507 3962
rect 17591 4138 17625 4154
rect 17591 3946 17625 3962
rect 17709 4138 17743 4154
rect 17709 3946 17743 3962
rect 17874 4138 17908 4154
rect 17874 3946 17908 3962
rect 17992 4138 18026 4154
rect 17992 3946 18026 3962
rect 18110 4138 18144 4154
rect 18110 3946 18144 3962
rect 18228 4138 18262 4154
rect 20773 4020 20807 4036
rect 20891 4412 20925 4428
rect 20891 4020 20925 4036
rect 21009 4412 21043 4428
rect 21126 4412 21160 4428
rect 21126 4220 21160 4236
rect 21244 4412 21278 4428
rect 21244 4220 21278 4236
rect 23050 4189 23066 4223
rect 23100 4189 23116 4223
rect 24192 4193 24208 4227
rect 24242 4193 24258 4227
rect 22771 4138 22805 4154
rect 21009 4020 21043 4036
rect 21296 4086 21545 4129
rect 21296 3996 21343 4086
rect 21506 3996 21545 4086
rect 18228 3946 18262 3962
rect 20816 3952 20832 3986
rect 20866 3952 20882 3986
rect 20934 3952 20950 3986
rect 20984 3952 21000 3986
rect 21296 3957 21545 3996
rect 22771 3946 22805 3962
rect 22889 4138 22923 4154
rect 22889 3946 22923 3962
rect 23007 4138 23041 4154
rect 23007 3946 23041 3962
rect 23125 4138 23159 4154
rect 23125 3946 23159 3962
rect 23290 4138 23324 4154
rect 23290 3946 23324 3962
rect 23408 4138 23442 4154
rect 23408 3946 23442 3962
rect 23526 4138 23560 4154
rect 23526 3946 23560 3962
rect 23644 4138 23678 4154
rect 23644 3946 23678 3962
rect 23913 4142 23947 4158
rect 23913 3950 23947 3966
rect 24031 4142 24065 4158
rect 24031 3950 24065 3966
rect 24149 4142 24183 4158
rect 24149 3950 24183 3966
rect 24267 4142 24301 4158
rect 24267 3950 24301 3966
rect 24432 4142 24466 4158
rect 24432 3950 24466 3966
rect 24550 4142 24584 4158
rect 24550 3950 24584 3966
rect 24668 4142 24702 4158
rect 24668 3950 24702 3966
rect 24786 4142 24820 4158
rect 24786 3950 24820 3966
rect 3181 3719 3353 3766
rect 1340 3617 1563 3693
rect 1340 3468 1419 3617
rect 1486 3468 1563 3617
rect 3181 3556 3220 3719
rect 3310 3556 3353 3719
rect 3181 3517 3353 3556
rect 4323 3717 4495 3764
rect 4323 3554 4362 3717
rect 4452 3554 4495 3717
rect 9694 3716 9866 3763
rect 4323 3515 4495 3554
rect 7853 3614 8076 3690
rect 1340 3362 1563 3468
rect 7853 3465 7932 3614
rect 7999 3465 8076 3614
rect 9694 3553 9733 3716
rect 9823 3553 9866 3716
rect 9694 3514 9866 3553
rect 10836 3714 11008 3761
rect 10836 3551 10875 3714
rect 10965 3551 11008 3714
rect 16228 3711 16400 3758
rect 10836 3512 11008 3551
rect 14387 3609 14610 3685
rect 7853 3359 8076 3465
rect 14387 3460 14466 3609
rect 14533 3460 14610 3609
rect 16228 3548 16267 3711
rect 16357 3548 16400 3711
rect 16228 3509 16400 3548
rect 17370 3709 17542 3756
rect 17370 3546 17409 3709
rect 17499 3546 17542 3709
rect 22786 3715 22958 3762
rect 17370 3507 17542 3546
rect 20945 3613 21168 3689
rect 14387 3354 14610 3460
rect 20945 3464 21024 3613
rect 21091 3464 21168 3613
rect 22786 3552 22825 3715
rect 22915 3552 22958 3715
rect 22786 3513 22958 3552
rect 23928 3713 24100 3760
rect 23928 3550 23967 3713
rect 24057 3550 24100 3713
rect 23928 3511 24100 3550
rect 20945 3358 21168 3464
rect 1771 3253 2041 3287
rect 945 3203 979 3219
rect 945 3011 979 3027
rect 1063 3203 1097 3219
rect 1063 3011 1097 3027
rect 1181 3203 1215 3219
rect 1181 3011 1215 3027
rect 1299 3203 1333 3219
rect 1299 3011 1333 3027
rect 1417 3203 1451 3219
rect 1417 3011 1451 3027
rect 1535 3203 1569 3219
rect 1535 3011 1569 3027
rect 1653 3203 1687 3219
rect 1653 3011 1687 3027
rect 1771 3203 1805 3253
rect 1771 3011 1805 3027
rect 1889 3203 1923 3219
rect 1889 3011 1923 3027
rect 2007 3203 2041 3253
rect 2007 3011 2041 3027
rect 5051 3274 5276 3350
rect 5051 3125 5130 3274
rect 5197 3125 5276 3274
rect 8284 3250 8554 3284
rect 5051 3019 5276 3125
rect 7458 3200 7492 3216
rect 7458 3008 7492 3024
rect 7576 3200 7610 3216
rect 7576 3008 7610 3024
rect 7694 3200 7728 3216
rect 7694 3008 7728 3024
rect 7812 3200 7846 3216
rect 7812 3008 7846 3024
rect 7930 3200 7964 3216
rect 7930 3008 7964 3024
rect 8048 3200 8082 3216
rect 8048 3008 8082 3024
rect 8166 3200 8200 3216
rect 8166 3008 8200 3024
rect 8284 3200 8318 3250
rect 8284 3008 8318 3024
rect 8402 3200 8436 3216
rect 8402 3008 8436 3024
rect 8520 3200 8554 3250
rect 8520 3008 8554 3024
rect 11564 3271 11789 3347
rect 11564 3122 11643 3271
rect 11710 3122 11789 3271
rect 14818 3245 15088 3279
rect 11564 3016 11789 3122
rect 13992 3195 14026 3211
rect 13992 3003 14026 3019
rect 14110 3195 14144 3211
rect 14110 3003 14144 3019
rect 14228 3195 14262 3211
rect 14228 3003 14262 3019
rect 14346 3195 14380 3211
rect 14346 3003 14380 3019
rect 14464 3195 14498 3211
rect 14464 3003 14498 3019
rect 14582 3195 14616 3211
rect 14582 3003 14616 3019
rect 14700 3195 14734 3211
rect 14700 3003 14734 3019
rect 14818 3195 14852 3245
rect 14818 3003 14852 3019
rect 14936 3195 14970 3211
rect 14936 3003 14970 3019
rect 15054 3195 15088 3245
rect 15054 3003 15088 3019
rect 18098 3266 18323 3342
rect 18098 3117 18177 3266
rect 18244 3117 18323 3266
rect 21376 3249 21646 3283
rect 18098 3011 18323 3117
rect 20550 3199 20584 3215
rect 20550 3007 20584 3023
rect 20668 3199 20702 3215
rect 20668 3007 20702 3023
rect 20786 3199 20820 3215
rect 20786 3007 20820 3023
rect 20904 3199 20938 3215
rect 20904 3007 20938 3023
rect 21022 3199 21056 3215
rect 21022 3007 21056 3023
rect 21140 3199 21174 3215
rect 21140 3007 21174 3023
rect 21258 3199 21292 3215
rect 21258 3007 21292 3023
rect 21376 3199 21410 3249
rect 21376 3007 21410 3023
rect 21494 3199 21528 3215
rect 21494 3007 21528 3023
rect 21612 3199 21646 3249
rect 21612 3007 21646 3023
rect 24656 3270 24881 3346
rect 24656 3121 24735 3270
rect 24802 3121 24881 3270
rect 24656 3015 24881 3121
rect 1696 2933 1712 2967
rect 1746 2933 1762 2967
rect 8209 2930 8225 2964
rect 8259 2930 8275 2964
rect 14743 2925 14759 2959
rect 14793 2925 14809 2959
rect 21301 2929 21317 2963
rect 21351 2929 21367 2963
rect 1578 2816 1594 2850
rect 1628 2816 1644 2850
rect 3247 2839 3517 2874
rect 2893 2786 2927 2802
rect 1182 2766 1216 2782
rect 1182 2374 1216 2390
rect 1300 2766 1334 2782
rect 1300 2374 1334 2390
rect 1418 2766 1452 2782
rect 1535 2766 1569 2782
rect 1535 2574 1569 2590
rect 1653 2766 1687 2782
rect 1653 2574 1687 2590
rect 2409 2640 2679 2675
rect 2409 2586 2443 2640
rect 1418 2374 1452 2390
rect 1705 2440 1954 2483
rect 1705 2350 1752 2440
rect 1915 2350 1954 2440
rect 2409 2394 2443 2410
rect 2527 2586 2561 2602
rect 2527 2394 2561 2410
rect 2645 2586 2679 2640
rect 2645 2394 2679 2410
rect 2763 2586 2797 2602
rect 2763 2394 2797 2410
rect 2893 2394 2927 2410
rect 3011 2786 3045 2802
rect 3011 2394 3045 2410
rect 3129 2786 3163 2802
rect 3129 2394 3163 2410
rect 3247 2786 3281 2839
rect 3247 2394 3281 2410
rect 3365 2786 3399 2802
rect 3365 2394 3399 2410
rect 3483 2786 3517 2839
rect 5145 2839 5415 2874
rect 3483 2394 3517 2410
rect 3601 2786 3635 2802
rect 4791 2786 4825 2802
rect 4307 2640 4577 2675
rect 3601 2394 3635 2410
rect 3730 2586 3764 2602
rect 3730 2394 3764 2410
rect 3848 2586 3882 2602
rect 3848 2394 3882 2410
rect 3966 2586 4000 2602
rect 3966 2394 4000 2410
rect 4084 2586 4118 2602
rect 4084 2394 4118 2410
rect 4307 2586 4341 2640
rect 4307 2394 4341 2410
rect 4425 2586 4459 2602
rect 4425 2394 4459 2410
rect 4543 2586 4577 2640
rect 4543 2394 4577 2410
rect 4661 2586 4695 2602
rect 4661 2394 4695 2410
rect 4791 2394 4825 2410
rect 4909 2786 4943 2802
rect 4909 2394 4943 2410
rect 5027 2786 5061 2802
rect 5027 2394 5061 2410
rect 5145 2786 5179 2839
rect 5145 2394 5179 2410
rect 5263 2786 5297 2802
rect 5263 2394 5297 2410
rect 5381 2786 5415 2839
rect 8091 2813 8107 2847
rect 8141 2813 8157 2847
rect 9760 2836 10030 2871
rect 5381 2394 5415 2410
rect 5499 2786 5533 2802
rect 9406 2783 9440 2799
rect 7695 2763 7729 2779
rect 5499 2394 5533 2410
rect 5628 2586 5662 2602
rect 5628 2394 5662 2410
rect 5746 2586 5780 2602
rect 5746 2394 5780 2410
rect 5864 2586 5898 2602
rect 5864 2394 5898 2410
rect 5982 2586 6016 2602
rect 5982 2394 6016 2410
rect 7695 2371 7729 2387
rect 7813 2763 7847 2779
rect 7813 2371 7847 2387
rect 7931 2763 7965 2779
rect 8048 2763 8082 2779
rect 8048 2571 8082 2587
rect 8166 2763 8200 2779
rect 8166 2571 8200 2587
rect 8922 2637 9192 2672
rect 8922 2583 8956 2637
rect 7931 2371 7965 2387
rect 8218 2437 8467 2480
rect 1225 2306 1241 2340
rect 1275 2306 1291 2340
rect 1343 2306 1359 2340
rect 1393 2306 1409 2340
rect 1705 2311 1954 2350
rect 8218 2347 8265 2437
rect 8428 2347 8467 2437
rect 8922 2391 8956 2407
rect 9040 2583 9074 2599
rect 9040 2391 9074 2407
rect 9158 2583 9192 2637
rect 9158 2391 9192 2407
rect 9276 2583 9310 2599
rect 9276 2391 9310 2407
rect 9406 2391 9440 2407
rect 9524 2783 9558 2799
rect 9524 2391 9558 2407
rect 9642 2783 9676 2799
rect 9642 2391 9676 2407
rect 9760 2783 9794 2836
rect 9760 2391 9794 2407
rect 9878 2783 9912 2799
rect 9878 2391 9912 2407
rect 9996 2783 10030 2836
rect 11658 2836 11928 2871
rect 9996 2391 10030 2407
rect 10114 2783 10148 2799
rect 11304 2783 11338 2799
rect 10820 2637 11090 2672
rect 10114 2391 10148 2407
rect 10243 2583 10277 2599
rect 10243 2391 10277 2407
rect 10361 2583 10395 2599
rect 10361 2391 10395 2407
rect 10479 2583 10513 2599
rect 10479 2391 10513 2407
rect 10597 2583 10631 2599
rect 10597 2391 10631 2407
rect 10820 2583 10854 2637
rect 10820 2391 10854 2407
rect 10938 2583 10972 2599
rect 10938 2391 10972 2407
rect 11056 2583 11090 2637
rect 11056 2391 11090 2407
rect 11174 2583 11208 2599
rect 11174 2391 11208 2407
rect 11304 2391 11338 2407
rect 11422 2783 11456 2799
rect 11422 2391 11456 2407
rect 11540 2783 11574 2799
rect 11540 2391 11574 2407
rect 11658 2783 11692 2836
rect 11658 2391 11692 2407
rect 11776 2783 11810 2799
rect 11776 2391 11810 2407
rect 11894 2783 11928 2836
rect 14625 2808 14641 2842
rect 14675 2808 14691 2842
rect 16294 2831 16564 2866
rect 11894 2391 11928 2407
rect 12012 2783 12046 2799
rect 15940 2778 15974 2794
rect 14229 2758 14263 2774
rect 12012 2391 12046 2407
rect 12141 2583 12175 2599
rect 12141 2391 12175 2407
rect 12259 2583 12293 2599
rect 12259 2391 12293 2407
rect 12377 2583 12411 2599
rect 12377 2391 12411 2407
rect 12495 2583 12529 2599
rect 12495 2391 12529 2407
rect 14229 2366 14263 2382
rect 14347 2758 14381 2774
rect 14347 2366 14381 2382
rect 14465 2758 14499 2774
rect 14582 2758 14616 2774
rect 14582 2566 14616 2582
rect 14700 2758 14734 2774
rect 14700 2566 14734 2582
rect 15456 2632 15726 2667
rect 15456 2578 15490 2632
rect 14465 2366 14499 2382
rect 14752 2432 15001 2475
rect 7738 2303 7754 2337
rect 7788 2303 7804 2337
rect 7856 2303 7872 2337
rect 7906 2303 7922 2337
rect 8218 2308 8467 2347
rect 14752 2342 14799 2432
rect 14962 2342 15001 2432
rect 15456 2386 15490 2402
rect 15574 2578 15608 2594
rect 15574 2386 15608 2402
rect 15692 2578 15726 2632
rect 15692 2386 15726 2402
rect 15810 2578 15844 2594
rect 15810 2386 15844 2402
rect 15940 2386 15974 2402
rect 16058 2778 16092 2794
rect 16058 2386 16092 2402
rect 16176 2778 16210 2794
rect 16176 2386 16210 2402
rect 16294 2778 16328 2831
rect 16294 2386 16328 2402
rect 16412 2778 16446 2794
rect 16412 2386 16446 2402
rect 16530 2778 16564 2831
rect 18192 2831 18462 2866
rect 16530 2386 16564 2402
rect 16648 2778 16682 2794
rect 17838 2778 17872 2794
rect 17354 2632 17624 2667
rect 16648 2386 16682 2402
rect 16777 2578 16811 2594
rect 16777 2386 16811 2402
rect 16895 2578 16929 2594
rect 16895 2386 16929 2402
rect 17013 2578 17047 2594
rect 17013 2386 17047 2402
rect 17131 2578 17165 2594
rect 17131 2386 17165 2402
rect 17354 2578 17388 2632
rect 17354 2386 17388 2402
rect 17472 2578 17506 2594
rect 17472 2386 17506 2402
rect 17590 2578 17624 2632
rect 17590 2386 17624 2402
rect 17708 2578 17742 2594
rect 17708 2386 17742 2402
rect 17838 2386 17872 2402
rect 17956 2778 17990 2794
rect 17956 2386 17990 2402
rect 18074 2778 18108 2794
rect 18074 2386 18108 2402
rect 18192 2778 18226 2831
rect 18192 2386 18226 2402
rect 18310 2778 18344 2794
rect 18310 2386 18344 2402
rect 18428 2778 18462 2831
rect 21183 2812 21199 2846
rect 21233 2812 21249 2846
rect 22852 2835 23122 2870
rect 18428 2386 18462 2402
rect 18546 2778 18580 2794
rect 22498 2782 22532 2798
rect 20787 2762 20821 2778
rect 18546 2386 18580 2402
rect 18675 2578 18709 2594
rect 18675 2386 18709 2402
rect 18793 2578 18827 2594
rect 18793 2386 18827 2402
rect 18911 2578 18945 2594
rect 18911 2386 18945 2402
rect 19029 2578 19063 2594
rect 19029 2386 19063 2402
rect 20787 2370 20821 2386
rect 20905 2762 20939 2778
rect 20905 2370 20939 2386
rect 21023 2762 21057 2778
rect 21140 2762 21174 2778
rect 21140 2570 21174 2586
rect 21258 2762 21292 2778
rect 21258 2570 21292 2586
rect 22014 2636 22284 2671
rect 22014 2582 22048 2636
rect 21023 2370 21057 2386
rect 21310 2436 21559 2479
rect 14272 2298 14288 2332
rect 14322 2298 14338 2332
rect 14390 2298 14406 2332
rect 14440 2298 14456 2332
rect 14752 2303 15001 2342
rect 21310 2346 21357 2436
rect 21520 2346 21559 2436
rect 22014 2390 22048 2406
rect 22132 2582 22166 2598
rect 22132 2390 22166 2406
rect 22250 2582 22284 2636
rect 22250 2390 22284 2406
rect 22368 2582 22402 2598
rect 22368 2390 22402 2406
rect 22498 2390 22532 2406
rect 22616 2782 22650 2798
rect 22616 2390 22650 2406
rect 22734 2782 22768 2798
rect 22734 2390 22768 2406
rect 22852 2782 22886 2835
rect 22852 2390 22886 2406
rect 22970 2782 23004 2798
rect 22970 2390 23004 2406
rect 23088 2782 23122 2835
rect 24750 2835 25020 2870
rect 23088 2390 23122 2406
rect 23206 2782 23240 2798
rect 24396 2782 24430 2798
rect 23912 2636 24182 2671
rect 23206 2390 23240 2406
rect 23335 2582 23369 2598
rect 23335 2390 23369 2406
rect 23453 2582 23487 2598
rect 23453 2390 23487 2406
rect 23571 2582 23605 2598
rect 23571 2390 23605 2406
rect 23689 2582 23723 2598
rect 23689 2390 23723 2406
rect 23912 2582 23946 2636
rect 23912 2390 23946 2406
rect 24030 2582 24064 2598
rect 24030 2390 24064 2406
rect 24148 2582 24182 2636
rect 24148 2390 24182 2406
rect 24266 2582 24300 2598
rect 24266 2390 24300 2406
rect 24396 2390 24430 2406
rect 24514 2782 24548 2798
rect 24514 2390 24548 2406
rect 24632 2782 24666 2798
rect 24632 2390 24666 2406
rect 24750 2782 24784 2835
rect 24750 2390 24784 2406
rect 24868 2782 24902 2798
rect 24868 2390 24902 2406
rect 24986 2782 25020 2835
rect 24986 2390 25020 2406
rect 25104 2782 25138 2798
rect 25104 2390 25138 2406
rect 25233 2582 25267 2598
rect 25233 2390 25267 2406
rect 25351 2582 25385 2598
rect 25351 2390 25385 2406
rect 25469 2582 25503 2598
rect 25469 2390 25503 2406
rect 25587 2582 25621 2598
rect 25587 2390 25621 2406
rect 20830 2302 20846 2336
rect 20880 2302 20896 2336
rect 20948 2302 20964 2336
rect 20998 2302 21014 2336
rect 21310 2307 21559 2346
rect 3873 2172 3907 2188
rect 10386 2169 10420 2185
rect 3873 2122 3907 2138
rect 5963 2151 6030 2167
rect 5963 2117 5980 2151
rect 6014 2117 6030 2151
rect 16920 2164 16954 2180
rect 10386 2119 10420 2135
rect 12476 2148 12543 2164
rect 2836 2093 2870 2109
rect 1335 2013 1558 2089
rect 1335 1864 1414 2013
rect 1481 1864 1558 2013
rect 1335 1758 1558 1864
rect 2954 2093 2988 2109
rect 2836 1701 2870 1717
rect 2953 1717 2954 1764
rect 3072 2093 3106 2109
rect 2988 1717 2989 1764
rect 1766 1649 2036 1683
rect 940 1599 974 1615
rect 940 1407 974 1423
rect 1058 1599 1092 1615
rect 1058 1407 1092 1423
rect 1176 1599 1210 1615
rect 1176 1407 1210 1423
rect 1294 1599 1328 1615
rect 1294 1407 1328 1423
rect 1412 1599 1446 1615
rect 1412 1407 1446 1423
rect 1530 1599 1564 1615
rect 1530 1407 1564 1423
rect 1648 1599 1682 1615
rect 1648 1407 1682 1423
rect 1766 1599 1800 1649
rect 1766 1407 1800 1423
rect 1884 1599 1918 1615
rect 1884 1407 1918 1423
rect 2002 1599 2036 1649
rect 2953 1659 2989 1717
rect 3190 2093 3224 2109
rect 3072 1701 3106 1717
rect 3188 1717 3190 1764
rect 3188 1659 3224 1717
rect 3308 2093 3342 2109
rect 3308 1701 3342 1717
rect 3426 2093 3460 2109
rect 3544 2093 3578 2109
rect 3460 1717 3462 1763
rect 3426 1659 3462 1717
rect 3544 1701 3578 1717
rect 4734 2093 4768 2109
rect 4852 2093 4886 2109
rect 4734 1701 4768 1717
rect 4851 1717 4852 1764
rect 4970 2093 5004 2109
rect 4886 1717 4887 1764
rect 4049 1659 4546 1677
rect 2953 1656 4546 1659
rect 2953 1622 4494 1656
rect 4528 1622 4546 1656
rect 2953 1619 4546 1622
rect 4851 1659 4887 1717
rect 5088 2093 5122 2109
rect 4970 1701 5004 1717
rect 5086 1717 5088 1764
rect 5086 1659 5122 1717
rect 5206 2093 5240 2109
rect 5206 1701 5240 1717
rect 5324 2093 5358 2109
rect 5442 2093 5476 2109
rect 5963 2101 6030 2117
rect 12476 2114 12493 2148
rect 12527 2114 12543 2148
rect 23478 2168 23512 2184
rect 16920 2114 16954 2130
rect 19010 2143 19077 2159
rect 5358 1717 5360 1763
rect 5324 1659 5360 1717
rect 9349 2090 9383 2106
rect 7848 2010 8071 2086
rect 7848 1861 7927 2010
rect 7994 1861 8071 2010
rect 7848 1755 8071 1861
rect 5442 1701 5476 1717
rect 9467 2090 9501 2106
rect 9349 1698 9383 1714
rect 9466 1714 9467 1761
rect 9585 2090 9619 2106
rect 9501 1714 9502 1761
rect 5947 1688 6047 1689
rect 5947 1659 6103 1688
rect 4851 1619 6103 1659
rect 2972 1618 4546 1619
rect 4870 1618 6103 1619
rect 2850 1529 2917 1545
rect 2850 1495 2866 1529
rect 2900 1495 2917 1529
rect 2850 1479 2917 1495
rect 2002 1407 2036 1423
rect 2681 1462 2715 1478
rect 2681 1412 2715 1428
rect 3027 1377 3061 1618
rect 4049 1601 4546 1618
rect 3497 1529 3564 1545
rect 3497 1495 3514 1529
rect 3548 1495 3564 1529
rect 3497 1479 3564 1495
rect 4748 1529 4815 1545
rect 4748 1495 4764 1529
rect 4798 1495 4815 1529
rect 4748 1479 4815 1495
rect 3804 1461 3838 1477
rect 3116 1411 3132 1445
rect 3166 1411 3182 1445
rect 3234 1412 3250 1446
rect 3284 1412 3300 1446
rect 3804 1411 3838 1427
rect 4579 1462 4613 1478
rect 4579 1412 4613 1428
rect 4925 1377 4959 1618
rect 5947 1590 6103 1618
rect 8279 1646 8549 1680
rect 7453 1596 7487 1612
rect 5947 1589 6047 1590
rect 5393 1530 5460 1546
rect 5393 1496 5410 1530
rect 5444 1496 5460 1530
rect 5393 1480 5460 1496
rect 5702 1461 5736 1477
rect 5014 1411 5030 1445
rect 5064 1411 5080 1445
rect 5132 1412 5148 1446
rect 5182 1412 5198 1446
rect 5702 1411 5736 1427
rect 7453 1404 7487 1420
rect 7571 1596 7605 1612
rect 7571 1404 7605 1420
rect 7689 1596 7723 1612
rect 7689 1404 7723 1420
rect 7807 1596 7841 1612
rect 7807 1404 7841 1420
rect 7925 1596 7959 1612
rect 7925 1404 7959 1420
rect 8043 1596 8077 1612
rect 8043 1404 8077 1420
rect 8161 1596 8195 1612
rect 8161 1404 8195 1420
rect 8279 1596 8313 1646
rect 8279 1404 8313 1420
rect 8397 1596 8431 1612
rect 8397 1404 8431 1420
rect 8515 1596 8549 1646
rect 9466 1656 9502 1714
rect 9703 2090 9737 2106
rect 9585 1698 9619 1714
rect 9701 1714 9703 1761
rect 9701 1656 9737 1714
rect 9821 2090 9855 2106
rect 9821 1698 9855 1714
rect 9939 2090 9973 2106
rect 10057 2090 10091 2106
rect 9973 1714 9975 1760
rect 9939 1656 9975 1714
rect 10057 1698 10091 1714
rect 11247 2090 11281 2106
rect 11365 2090 11399 2106
rect 11247 1698 11281 1714
rect 11364 1714 11365 1761
rect 11483 2090 11517 2106
rect 11399 1714 11400 1761
rect 10562 1656 11059 1674
rect 9466 1653 11059 1656
rect 9466 1619 11007 1653
rect 11041 1619 11059 1653
rect 9466 1616 11059 1619
rect 11364 1656 11400 1714
rect 11601 2090 11635 2106
rect 11483 1698 11517 1714
rect 11599 1714 11601 1761
rect 11599 1656 11635 1714
rect 11719 2090 11753 2106
rect 11719 1698 11753 1714
rect 11837 2090 11871 2106
rect 11955 2090 11989 2106
rect 12476 2098 12543 2114
rect 19010 2109 19027 2143
rect 19061 2109 19077 2143
rect 23478 2118 23512 2134
rect 25568 2147 25635 2163
rect 11871 1714 11873 1760
rect 11837 1656 11873 1714
rect 15883 2085 15917 2101
rect 14382 2005 14605 2081
rect 14382 1856 14461 2005
rect 14528 1856 14605 2005
rect 14382 1750 14605 1856
rect 11955 1698 11989 1714
rect 16001 2085 16035 2101
rect 15883 1693 15917 1709
rect 16000 1709 16001 1756
rect 16119 2085 16153 2101
rect 16035 1709 16036 1756
rect 12460 1685 12560 1686
rect 12460 1656 12616 1685
rect 11364 1616 12616 1656
rect 9485 1615 11059 1616
rect 11383 1615 12616 1616
rect 9363 1526 9430 1542
rect 9363 1492 9379 1526
rect 9413 1492 9430 1526
rect 9363 1476 9430 1492
rect 8515 1404 8549 1420
rect 9194 1459 9228 1475
rect 9194 1409 9228 1425
rect 1691 1329 1707 1363
rect 1741 1329 1757 1363
rect 2534 1361 2568 1377
rect 1573 1212 1589 1246
rect 1623 1212 1639 1246
rect 1177 1162 1211 1178
rect 1177 770 1211 786
rect 1295 1162 1329 1178
rect 1295 770 1329 786
rect 1413 1162 1447 1178
rect 1530 1162 1564 1178
rect 1530 970 1564 986
rect 1648 1162 1682 1178
rect 2534 1169 2568 1185
rect 2652 1361 2686 1377
rect 2652 1169 2686 1185
rect 2954 1361 2988 1377
rect 1648 970 1682 986
rect 3027 1361 3106 1377
rect 3027 1331 3072 1361
rect 2954 918 2989 985
rect 3072 969 3106 985
rect 3190 1361 3224 1377
rect 3190 969 3224 985
rect 3308 1361 3342 1377
rect 3426 1361 3460 1377
rect 3832 1361 3866 1377
rect 3832 1169 3866 1185
rect 3950 1361 3984 1377
rect 3950 1169 3984 1185
rect 4432 1361 4466 1377
rect 4432 1169 4466 1185
rect 4550 1361 4584 1377
rect 4550 1169 4584 1185
rect 4852 1361 4886 1377
rect 3308 969 3342 985
rect 3425 918 3460 985
rect 2954 883 3460 918
rect 4925 1361 5004 1377
rect 4925 1331 4970 1361
rect 4852 918 4887 985
rect 4970 969 5004 985
rect 5088 1361 5122 1377
rect 5088 969 5122 985
rect 5206 1361 5240 1377
rect 5324 1361 5358 1377
rect 5730 1361 5764 1377
rect 5730 1169 5764 1185
rect 5848 1361 5882 1377
rect 9540 1374 9574 1615
rect 10562 1598 11059 1615
rect 10010 1526 10077 1542
rect 10010 1492 10027 1526
rect 10061 1492 10077 1526
rect 10010 1476 10077 1492
rect 11261 1526 11328 1542
rect 11261 1492 11277 1526
rect 11311 1492 11328 1526
rect 11261 1476 11328 1492
rect 10317 1458 10351 1474
rect 9629 1408 9645 1442
rect 9679 1408 9695 1442
rect 9747 1409 9763 1443
rect 9797 1409 9813 1443
rect 10317 1408 10351 1424
rect 11092 1459 11126 1475
rect 11092 1409 11126 1425
rect 11438 1374 11472 1615
rect 12460 1587 12616 1615
rect 14813 1641 15083 1675
rect 13987 1591 14021 1607
rect 12460 1586 12560 1587
rect 11906 1527 11973 1543
rect 11906 1493 11923 1527
rect 11957 1493 11973 1527
rect 11906 1477 11973 1493
rect 12215 1458 12249 1474
rect 11527 1408 11543 1442
rect 11577 1408 11593 1442
rect 11645 1409 11661 1443
rect 11695 1409 11711 1443
rect 12215 1408 12249 1424
rect 13987 1399 14021 1415
rect 14105 1591 14139 1607
rect 14105 1399 14139 1415
rect 14223 1591 14257 1607
rect 14223 1399 14257 1415
rect 14341 1591 14375 1607
rect 14341 1399 14375 1415
rect 14459 1591 14493 1607
rect 14459 1399 14493 1415
rect 14577 1591 14611 1607
rect 14577 1399 14611 1415
rect 14695 1591 14729 1607
rect 14695 1399 14729 1415
rect 14813 1591 14847 1641
rect 14813 1399 14847 1415
rect 14931 1591 14965 1607
rect 14931 1399 14965 1415
rect 15049 1591 15083 1641
rect 16000 1651 16036 1709
rect 16237 2085 16271 2101
rect 16119 1693 16153 1709
rect 16235 1709 16237 1756
rect 16235 1651 16271 1709
rect 16355 2085 16389 2101
rect 16355 1693 16389 1709
rect 16473 2085 16507 2101
rect 16591 2085 16625 2101
rect 16507 1709 16509 1755
rect 16473 1651 16509 1709
rect 16591 1693 16625 1709
rect 17781 2085 17815 2101
rect 17899 2085 17933 2101
rect 17781 1693 17815 1709
rect 17898 1709 17899 1756
rect 18017 2085 18051 2101
rect 17933 1709 17934 1756
rect 17096 1651 17593 1669
rect 16000 1648 17593 1651
rect 16000 1614 17541 1648
rect 17575 1614 17593 1648
rect 16000 1611 17593 1614
rect 17898 1651 17934 1709
rect 18135 2085 18169 2101
rect 18017 1693 18051 1709
rect 18133 1709 18135 1756
rect 18133 1651 18169 1709
rect 18253 2085 18287 2101
rect 18253 1693 18287 1709
rect 18371 2085 18405 2101
rect 18489 2085 18523 2101
rect 19010 2093 19077 2109
rect 25568 2113 25585 2147
rect 25619 2113 25635 2147
rect 22441 2089 22475 2105
rect 18405 1709 18407 1755
rect 18371 1651 18407 1709
rect 20940 2009 21163 2085
rect 20940 1860 21019 2009
rect 21086 1860 21163 2009
rect 20940 1754 21163 1860
rect 18489 1693 18523 1709
rect 22559 2089 22593 2105
rect 22441 1697 22475 1713
rect 22558 1713 22559 1760
rect 22677 2089 22711 2105
rect 22593 1713 22594 1760
rect 18994 1680 19094 1681
rect 18994 1651 19150 1680
rect 17898 1611 19150 1651
rect 16019 1610 17593 1611
rect 17917 1610 19150 1611
rect 15897 1521 15964 1537
rect 15897 1487 15913 1521
rect 15947 1487 15964 1521
rect 15897 1471 15964 1487
rect 15049 1399 15083 1415
rect 15728 1454 15762 1470
rect 15728 1404 15762 1420
rect 8204 1326 8220 1360
rect 8254 1326 8270 1360
rect 9047 1358 9081 1374
rect 8086 1209 8102 1243
rect 8136 1209 8152 1243
rect 5848 1169 5882 1185
rect 5206 969 5240 985
rect 5323 918 5358 985
rect 4852 883 5358 918
rect 7690 1159 7724 1175
rect 1413 770 1447 786
rect 1700 836 1949 879
rect 1700 746 1747 836
rect 1910 746 1949 836
rect 7690 767 7724 783
rect 7808 1159 7842 1175
rect 7808 767 7842 783
rect 7926 1159 7960 1175
rect 8043 1159 8077 1175
rect 8043 967 8077 983
rect 8161 1159 8195 1175
rect 9047 1166 9081 1182
rect 9165 1358 9199 1374
rect 9165 1166 9199 1182
rect 9467 1358 9501 1374
rect 8161 967 8195 983
rect 9540 1358 9619 1374
rect 9540 1328 9585 1358
rect 9467 915 9502 982
rect 9585 966 9619 982
rect 9703 1358 9737 1374
rect 9703 966 9737 982
rect 9821 1358 9855 1374
rect 9939 1358 9973 1374
rect 10345 1358 10379 1374
rect 10345 1166 10379 1182
rect 10463 1358 10497 1374
rect 10463 1166 10497 1182
rect 10945 1358 10979 1374
rect 10945 1166 10979 1182
rect 11063 1358 11097 1374
rect 11063 1166 11097 1182
rect 11365 1358 11399 1374
rect 9821 966 9855 982
rect 9938 915 9973 982
rect 9467 880 9973 915
rect 11438 1358 11517 1374
rect 11438 1328 11483 1358
rect 11365 915 11400 982
rect 11483 966 11517 982
rect 11601 1358 11635 1374
rect 11601 966 11635 982
rect 11719 1358 11753 1374
rect 11837 1358 11871 1374
rect 12243 1358 12277 1374
rect 12243 1166 12277 1182
rect 12361 1358 12395 1374
rect 16074 1369 16108 1610
rect 17096 1593 17593 1610
rect 16544 1521 16611 1537
rect 16544 1487 16561 1521
rect 16595 1487 16611 1521
rect 16544 1471 16611 1487
rect 17795 1521 17862 1537
rect 17795 1487 17811 1521
rect 17845 1487 17862 1521
rect 17795 1471 17862 1487
rect 16851 1453 16885 1469
rect 16163 1403 16179 1437
rect 16213 1403 16229 1437
rect 16281 1404 16297 1438
rect 16331 1404 16347 1438
rect 16851 1403 16885 1419
rect 17626 1454 17660 1470
rect 17626 1404 17660 1420
rect 17972 1369 18006 1610
rect 18994 1582 19150 1610
rect 21371 1645 21641 1679
rect 20545 1595 20579 1611
rect 18994 1581 19094 1582
rect 18440 1522 18507 1538
rect 18440 1488 18457 1522
rect 18491 1488 18507 1522
rect 18440 1472 18507 1488
rect 18749 1453 18783 1469
rect 18061 1403 18077 1437
rect 18111 1403 18127 1437
rect 18179 1404 18195 1438
rect 18229 1404 18245 1438
rect 18749 1403 18783 1419
rect 20545 1403 20579 1419
rect 20663 1595 20697 1611
rect 20663 1403 20697 1419
rect 20781 1595 20815 1611
rect 20781 1403 20815 1419
rect 20899 1595 20933 1611
rect 20899 1403 20933 1419
rect 21017 1595 21051 1611
rect 21017 1403 21051 1419
rect 21135 1595 21169 1611
rect 21135 1403 21169 1419
rect 21253 1595 21287 1611
rect 21253 1403 21287 1419
rect 21371 1595 21405 1645
rect 21371 1403 21405 1419
rect 21489 1595 21523 1611
rect 21489 1403 21523 1419
rect 21607 1595 21641 1645
rect 22558 1655 22594 1713
rect 22795 2089 22829 2105
rect 22677 1697 22711 1713
rect 22793 1713 22795 1760
rect 22793 1655 22829 1713
rect 22913 2089 22947 2105
rect 22913 1697 22947 1713
rect 23031 2089 23065 2105
rect 23149 2089 23183 2105
rect 23065 1713 23067 1759
rect 23031 1655 23067 1713
rect 23149 1697 23183 1713
rect 24339 2089 24373 2105
rect 24457 2089 24491 2105
rect 24339 1697 24373 1713
rect 24456 1713 24457 1760
rect 24575 2089 24609 2105
rect 24491 1713 24492 1760
rect 23654 1655 24151 1673
rect 22558 1652 24151 1655
rect 22558 1618 24099 1652
rect 24133 1618 24151 1652
rect 22558 1615 24151 1618
rect 24456 1655 24492 1713
rect 24693 2089 24727 2105
rect 24575 1697 24609 1713
rect 24691 1713 24693 1760
rect 24691 1655 24727 1713
rect 24811 2089 24845 2105
rect 24811 1697 24845 1713
rect 24929 2089 24963 2105
rect 25047 2089 25081 2105
rect 25568 2097 25635 2113
rect 24963 1713 24965 1759
rect 24929 1655 24965 1713
rect 25047 1697 25081 1713
rect 25552 1684 25652 1685
rect 25552 1655 25708 1684
rect 24456 1615 25708 1655
rect 22577 1614 24151 1615
rect 24475 1614 25708 1615
rect 22455 1525 22522 1541
rect 22455 1491 22471 1525
rect 22505 1491 22522 1525
rect 22455 1475 22522 1491
rect 21607 1403 21641 1419
rect 22286 1458 22320 1474
rect 22286 1408 22320 1424
rect 22632 1373 22666 1614
rect 23654 1597 24151 1614
rect 23102 1525 23169 1541
rect 23102 1491 23119 1525
rect 23153 1491 23169 1525
rect 23102 1475 23169 1491
rect 24353 1525 24420 1541
rect 24353 1491 24369 1525
rect 24403 1491 24420 1525
rect 24353 1475 24420 1491
rect 23409 1457 23443 1473
rect 22721 1407 22737 1441
rect 22771 1407 22787 1441
rect 22839 1408 22855 1442
rect 22889 1408 22905 1442
rect 23409 1407 23443 1423
rect 24184 1458 24218 1474
rect 24184 1408 24218 1424
rect 24530 1373 24564 1614
rect 25552 1586 25708 1614
rect 25552 1585 25652 1586
rect 24998 1526 25065 1542
rect 24998 1492 25015 1526
rect 25049 1492 25065 1526
rect 24998 1476 25065 1492
rect 25307 1457 25341 1473
rect 24619 1407 24635 1441
rect 24669 1407 24685 1441
rect 24737 1408 24753 1442
rect 24787 1408 24803 1442
rect 25307 1407 25341 1423
rect 14738 1321 14754 1355
rect 14788 1321 14804 1355
rect 15581 1353 15615 1369
rect 14620 1204 14636 1238
rect 14670 1204 14686 1238
rect 12361 1166 12395 1182
rect 11719 966 11753 982
rect 11836 915 11871 982
rect 11365 880 11871 915
rect 14224 1154 14258 1170
rect 7926 767 7960 783
rect 8213 833 8462 876
rect 1220 702 1236 736
rect 1270 702 1286 736
rect 1338 702 1354 736
rect 1388 702 1404 736
rect 1700 707 1949 746
rect 8213 743 8260 833
rect 8423 743 8462 833
rect 14224 762 14258 778
rect 14342 1154 14376 1170
rect 14342 762 14376 778
rect 14460 1154 14494 1170
rect 14577 1154 14611 1170
rect 14577 962 14611 978
rect 14695 1154 14729 1170
rect 15581 1161 15615 1177
rect 15699 1353 15733 1369
rect 15699 1161 15733 1177
rect 16001 1353 16035 1369
rect 14695 962 14729 978
rect 16074 1353 16153 1369
rect 16074 1323 16119 1353
rect 16001 910 16036 977
rect 16119 961 16153 977
rect 16237 1353 16271 1369
rect 16237 961 16271 977
rect 16355 1353 16389 1369
rect 16473 1353 16507 1369
rect 16879 1353 16913 1369
rect 16879 1161 16913 1177
rect 16997 1353 17031 1369
rect 16997 1161 17031 1177
rect 17479 1353 17513 1369
rect 17479 1161 17513 1177
rect 17597 1353 17631 1369
rect 17597 1161 17631 1177
rect 17899 1353 17933 1369
rect 16355 961 16389 977
rect 16472 910 16507 977
rect 16001 875 16507 910
rect 17972 1353 18051 1369
rect 17972 1323 18017 1353
rect 17899 910 17934 977
rect 18017 961 18051 977
rect 18135 1353 18169 1369
rect 18135 961 18169 977
rect 18253 1353 18287 1369
rect 18371 1353 18405 1369
rect 18777 1353 18811 1369
rect 18777 1161 18811 1177
rect 18895 1353 18929 1369
rect 21296 1325 21312 1359
rect 21346 1325 21362 1359
rect 22139 1357 22173 1373
rect 21178 1208 21194 1242
rect 21228 1208 21244 1242
rect 18895 1161 18929 1177
rect 18253 961 18287 977
rect 18370 910 18405 977
rect 17899 875 18405 910
rect 20782 1158 20816 1174
rect 14460 762 14494 778
rect 14747 828 14996 871
rect 3125 676 3297 723
rect 7733 699 7749 733
rect 7783 699 7799 733
rect 7851 699 7867 733
rect 7901 699 7917 733
rect 8213 704 8462 743
rect 14747 738 14794 828
rect 14957 738 14996 828
rect 20782 766 20816 782
rect 20900 1158 20934 1174
rect 20900 766 20934 782
rect 21018 1158 21052 1174
rect 21135 1158 21169 1174
rect 21135 966 21169 982
rect 21253 1158 21287 1174
rect 22139 1165 22173 1181
rect 22257 1357 22291 1373
rect 22257 1165 22291 1181
rect 22559 1357 22593 1373
rect 21253 966 21287 982
rect 22632 1357 22711 1373
rect 22632 1327 22677 1357
rect 22559 914 22594 981
rect 22677 965 22711 981
rect 22795 1357 22829 1373
rect 22795 965 22829 981
rect 22913 1357 22947 1373
rect 23031 1357 23065 1373
rect 23437 1357 23471 1373
rect 23437 1165 23471 1181
rect 23555 1357 23589 1373
rect 23555 1165 23589 1181
rect 24037 1357 24071 1373
rect 24037 1165 24071 1181
rect 24155 1357 24189 1373
rect 24155 1165 24189 1181
rect 24457 1357 24491 1373
rect 22913 965 22947 981
rect 23030 914 23065 981
rect 22559 879 23065 914
rect 24530 1357 24609 1373
rect 24530 1327 24575 1357
rect 24457 914 24492 981
rect 24575 965 24609 981
rect 24693 1357 24727 1373
rect 24693 965 24727 981
rect 24811 1357 24845 1373
rect 24929 1357 24963 1373
rect 25335 1357 25369 1373
rect 25335 1165 25369 1181
rect 25453 1357 25487 1373
rect 25453 1165 25487 1181
rect 24811 965 24845 981
rect 24928 914 24963 981
rect 24457 879 24963 914
rect 21018 766 21052 782
rect 21305 832 21554 875
rect 3125 513 3164 676
rect 3254 513 3297 676
rect 3125 473 3297 513
rect 9638 673 9810 720
rect 14267 694 14283 728
rect 14317 694 14333 728
rect 14385 694 14401 728
rect 14435 694 14451 728
rect 14747 699 14996 738
rect 21305 742 21352 832
rect 21515 742 21554 832
rect 9638 510 9677 673
rect 9767 510 9810 673
rect 9638 470 9810 510
rect 16172 668 16344 715
rect 20825 698 20841 732
rect 20875 698 20891 732
rect 20943 698 20959 732
rect 20993 698 21009 732
rect 21305 703 21554 742
rect 16172 505 16211 668
rect 16301 505 16344 668
rect 16172 465 16344 505
rect 22730 672 22902 719
rect 22730 509 22769 672
rect 22859 509 22902 672
rect 22730 469 22902 509
rect 904 -287 1127 -211
rect 904 -436 981 -287
rect 1048 -436 1127 -287
rect 904 -542 1127 -436
rect 2051 -287 2274 -211
rect 2051 -436 2128 -287
rect 2195 -436 2274 -287
rect 1777 -501 1811 -485
rect 1777 -551 1811 -535
rect 2051 -542 2274 -436
rect 4533 -341 4756 -265
rect 4533 -490 4610 -341
rect 4677 -490 4756 -341
rect 2907 -507 2941 -491
rect 2907 -557 2941 -541
rect 4533 -596 4756 -490
rect 7462 -291 7685 -215
rect 7462 -440 7539 -291
rect 7606 -440 7685 -291
rect 7462 -546 7685 -440
rect 8609 -291 8832 -215
rect 8609 -440 8686 -291
rect 8753 -440 8832 -291
rect 8335 -505 8369 -489
rect 8335 -555 8369 -539
rect 8609 -546 8832 -440
rect 11091 -345 11314 -269
rect 11091 -494 11168 -345
rect 11235 -494 11314 -345
rect 9465 -511 9499 -495
rect 9465 -561 9499 -545
rect 11091 -600 11314 -494
rect 13996 -286 14219 -210
rect 13996 -435 14073 -286
rect 14140 -435 14219 -286
rect 13996 -541 14219 -435
rect 15143 -286 15366 -210
rect 15143 -435 15220 -286
rect 15287 -435 15366 -286
rect 14869 -500 14903 -484
rect 14869 -550 14903 -534
rect 15143 -541 15366 -435
rect 17625 -340 17848 -264
rect 17625 -489 17702 -340
rect 17769 -489 17848 -340
rect 15999 -506 16033 -490
rect 15999 -556 16033 -540
rect 17625 -595 17848 -489
rect 20509 -283 20732 -207
rect 20509 -432 20586 -283
rect 20653 -432 20732 -283
rect 20509 -538 20732 -432
rect 21656 -283 21879 -207
rect 21656 -432 21733 -283
rect 21800 -432 21879 -283
rect 21382 -497 21416 -481
rect 21382 -547 21416 -531
rect 21656 -538 21879 -432
rect 24138 -337 24361 -261
rect 24138 -486 24215 -337
rect 24282 -486 24361 -337
rect 22512 -503 22546 -487
rect 22512 -553 22546 -537
rect 24138 -592 24361 -486
rect 1777 -621 1811 -605
rect 942 -679 976 -663
rect 942 -1071 976 -1055
rect 1060 -679 1094 -663
rect 1060 -1071 1094 -1055
rect 1178 -679 1212 -663
rect 1178 -1071 1212 -1055
rect 1296 -679 1330 -663
rect 1296 -1071 1330 -1055
rect 1414 -679 1448 -663
rect 1414 -1071 1448 -1055
rect 1532 -679 1566 -663
rect 1532 -1071 1566 -1055
rect 1650 -679 1684 -663
rect 1777 -671 1811 -655
rect 2907 -625 2941 -609
rect 1650 -1071 1684 -1055
rect 2084 -683 2118 -667
rect 2084 -1075 2118 -1059
rect 2202 -683 2236 -667
rect 2202 -1075 2236 -1059
rect 2320 -683 2354 -667
rect 2320 -1075 2354 -1059
rect 2438 -683 2472 -667
rect 2438 -1075 2472 -1059
rect 2556 -683 2590 -667
rect 2556 -1075 2590 -1059
rect 2674 -683 2708 -667
rect 2674 -1075 2708 -1059
rect 2792 -683 2826 -667
rect 2907 -675 2941 -659
rect 8335 -625 8369 -609
rect 4055 -705 4325 -671
rect 4055 -755 4089 -705
rect 4055 -947 4089 -931
rect 4173 -755 4207 -739
rect 4173 -947 4207 -931
rect 4291 -755 4325 -705
rect 7500 -683 7534 -667
rect 4291 -947 4325 -931
rect 4409 -755 4443 -739
rect 4409 -947 4443 -931
rect 4527 -755 4561 -739
rect 4527 -947 4561 -931
rect 4645 -755 4679 -739
rect 4645 -947 4679 -931
rect 4763 -755 4797 -739
rect 4763 -947 4797 -931
rect 4881 -755 4915 -739
rect 4881 -947 4915 -931
rect 4999 -755 5033 -739
rect 4999 -947 5033 -931
rect 5117 -755 5151 -739
rect 5117 -947 5151 -931
rect 4334 -1025 4350 -991
rect 4384 -1025 4400 -991
rect 2792 -1075 2826 -1059
rect 7500 -1075 7534 -1059
rect 7618 -683 7652 -667
rect 7618 -1075 7652 -1059
rect 7736 -683 7770 -667
rect 7736 -1075 7770 -1059
rect 7854 -683 7888 -667
rect 7854 -1075 7888 -1059
rect 7972 -683 8006 -667
rect 7972 -1075 8006 -1059
rect 8090 -683 8124 -667
rect 8090 -1075 8124 -1059
rect 8208 -683 8242 -667
rect 8335 -675 8369 -659
rect 9465 -629 9499 -613
rect 14869 -620 14903 -604
rect 8208 -1075 8242 -1059
rect 8642 -687 8676 -671
rect 8642 -1079 8676 -1063
rect 8760 -687 8794 -671
rect 8760 -1079 8794 -1063
rect 8878 -687 8912 -671
rect 8878 -1079 8912 -1063
rect 8996 -687 9030 -671
rect 8996 -1079 9030 -1063
rect 9114 -687 9148 -671
rect 9114 -1079 9148 -1063
rect 9232 -687 9266 -671
rect 9232 -1079 9266 -1063
rect 9350 -687 9384 -671
rect 9465 -679 9499 -663
rect 10613 -709 10883 -675
rect 10613 -759 10647 -709
rect 10613 -951 10647 -935
rect 10731 -759 10765 -743
rect 10731 -951 10765 -935
rect 10849 -759 10883 -709
rect 14034 -678 14068 -662
rect 10849 -951 10883 -935
rect 10967 -759 11001 -743
rect 10967 -951 11001 -935
rect 11085 -759 11119 -743
rect 11085 -951 11119 -935
rect 11203 -759 11237 -743
rect 11203 -951 11237 -935
rect 11321 -759 11355 -743
rect 11321 -951 11355 -935
rect 11439 -759 11473 -743
rect 11439 -951 11473 -935
rect 11557 -759 11591 -743
rect 11557 -951 11591 -935
rect 11675 -759 11709 -743
rect 11675 -951 11709 -935
rect 10892 -1029 10908 -995
rect 10942 -1029 10958 -995
rect 9350 -1079 9384 -1063
rect 14034 -1070 14068 -1054
rect 14152 -678 14186 -662
rect 14152 -1070 14186 -1054
rect 14270 -678 14304 -662
rect 14270 -1070 14304 -1054
rect 14388 -678 14422 -662
rect 14388 -1070 14422 -1054
rect 14506 -678 14540 -662
rect 14506 -1070 14540 -1054
rect 14624 -678 14658 -662
rect 14624 -1070 14658 -1054
rect 14742 -678 14776 -662
rect 14869 -670 14903 -654
rect 15999 -624 16033 -608
rect 14742 -1070 14776 -1054
rect 15176 -682 15210 -666
rect 15176 -1074 15210 -1058
rect 15294 -682 15328 -666
rect 15294 -1074 15328 -1058
rect 15412 -682 15446 -666
rect 15412 -1074 15446 -1058
rect 15530 -682 15564 -666
rect 15530 -1074 15564 -1058
rect 15648 -682 15682 -666
rect 15648 -1074 15682 -1058
rect 15766 -682 15800 -666
rect 15766 -1074 15800 -1058
rect 15884 -682 15918 -666
rect 15999 -674 16033 -658
rect 21382 -617 21416 -601
rect 17147 -704 17417 -670
rect 17147 -754 17181 -704
rect 17147 -946 17181 -930
rect 17265 -754 17299 -738
rect 17265 -946 17299 -930
rect 17383 -754 17417 -704
rect 20547 -675 20581 -659
rect 17383 -946 17417 -930
rect 17501 -754 17535 -738
rect 17501 -946 17535 -930
rect 17619 -754 17653 -738
rect 17619 -946 17653 -930
rect 17737 -754 17771 -738
rect 17737 -946 17771 -930
rect 17855 -754 17889 -738
rect 17855 -946 17889 -930
rect 17973 -754 18007 -738
rect 17973 -946 18007 -930
rect 18091 -754 18125 -738
rect 18091 -946 18125 -930
rect 18209 -754 18243 -738
rect 18209 -946 18243 -930
rect 17426 -1024 17442 -990
rect 17476 -1024 17492 -990
rect 15884 -1074 15918 -1058
rect 20547 -1067 20581 -1051
rect 20665 -675 20699 -659
rect 20665 -1067 20699 -1051
rect 20783 -675 20817 -659
rect 20783 -1067 20817 -1051
rect 20901 -675 20935 -659
rect 20901 -1067 20935 -1051
rect 21019 -675 21053 -659
rect 21019 -1067 21053 -1051
rect 21137 -675 21171 -659
rect 21137 -1067 21171 -1051
rect 21255 -675 21289 -659
rect 21382 -667 21416 -651
rect 22512 -621 22546 -605
rect 21255 -1067 21289 -1051
rect 21689 -679 21723 -663
rect 21689 -1071 21723 -1055
rect 21807 -679 21841 -663
rect 21807 -1071 21841 -1055
rect 21925 -679 21959 -663
rect 21925 -1071 21959 -1055
rect 22043 -679 22077 -663
rect 22043 -1071 22077 -1055
rect 22161 -679 22195 -663
rect 22161 -1071 22195 -1055
rect 22279 -679 22313 -663
rect 22279 -1071 22313 -1055
rect 22397 -679 22431 -663
rect 22512 -671 22546 -655
rect 23660 -701 23930 -667
rect 23660 -751 23694 -701
rect 23660 -943 23694 -927
rect 23778 -751 23812 -735
rect 23778 -943 23812 -927
rect 23896 -751 23930 -701
rect 23896 -943 23930 -927
rect 24014 -751 24048 -735
rect 24014 -943 24048 -927
rect 24132 -751 24166 -735
rect 24132 -943 24166 -927
rect 24250 -751 24284 -735
rect 24250 -943 24284 -927
rect 24368 -751 24402 -735
rect 24368 -943 24402 -927
rect 24486 -751 24520 -735
rect 24486 -943 24520 -927
rect 24604 -751 24638 -735
rect 24604 -943 24638 -927
rect 24722 -751 24756 -735
rect 24722 -943 24756 -927
rect 23939 -1021 23955 -987
rect 23989 -1021 24005 -987
rect 22397 -1071 22431 -1055
rect 4452 -1142 4468 -1108
rect 4502 -1142 4518 -1108
rect 11010 -1146 11026 -1112
rect 11060 -1146 11076 -1112
rect 17544 -1141 17560 -1107
rect 17594 -1141 17610 -1107
rect 24057 -1138 24073 -1104
rect 24107 -1138 24123 -1104
rect 4409 -1192 4443 -1176
rect 1429 -1411 1445 -1377
rect 1479 -1411 1495 -1377
rect 2571 -1415 2587 -1381
rect 2621 -1415 2637 -1381
rect 4409 -1384 4443 -1368
rect 4527 -1192 4561 -1176
rect 4527 -1384 4561 -1368
rect 4644 -1192 4678 -1176
rect 867 -1462 901 -1446
rect 867 -1654 901 -1638
rect 985 -1462 1019 -1446
rect 985 -1654 1019 -1638
rect 1103 -1462 1137 -1446
rect 1103 -1654 1137 -1638
rect 1221 -1462 1255 -1446
rect 1221 -1654 1255 -1638
rect 1386 -1462 1420 -1446
rect 1386 -1654 1420 -1638
rect 1504 -1462 1538 -1446
rect 1504 -1654 1538 -1638
rect 1622 -1462 1656 -1446
rect 1622 -1654 1656 -1638
rect 1740 -1462 1774 -1446
rect 1740 -1654 1774 -1638
rect 2009 -1466 2043 -1450
rect 2009 -1658 2043 -1642
rect 2127 -1466 2161 -1450
rect 2127 -1658 2161 -1642
rect 2245 -1466 2279 -1450
rect 2245 -1658 2279 -1642
rect 2363 -1466 2397 -1450
rect 2363 -1658 2397 -1642
rect 2528 -1466 2562 -1450
rect 2528 -1658 2562 -1642
rect 2646 -1466 2680 -1450
rect 2646 -1658 2680 -1642
rect 2764 -1466 2798 -1450
rect 2764 -1658 2798 -1642
rect 2882 -1466 2916 -1450
rect 2882 -1658 2916 -1642
rect 4142 -1518 4391 -1475
rect 4142 -1608 4181 -1518
rect 4344 -1608 4391 -1518
rect 4644 -1584 4678 -1568
rect 4762 -1192 4796 -1176
rect 4762 -1584 4796 -1568
rect 4880 -1192 4914 -1176
rect 10967 -1196 11001 -1180
rect 7987 -1415 8003 -1381
rect 8037 -1415 8053 -1381
rect 9129 -1419 9145 -1385
rect 9179 -1419 9195 -1385
rect 10967 -1388 11001 -1372
rect 11085 -1196 11119 -1180
rect 11085 -1388 11119 -1372
rect 11202 -1196 11236 -1180
rect 4880 -1584 4914 -1568
rect 7425 -1466 7459 -1450
rect 4142 -1647 4391 -1608
rect 4687 -1652 4703 -1618
rect 4737 -1652 4753 -1618
rect 4805 -1652 4821 -1618
rect 4855 -1652 4871 -1618
rect 7425 -1658 7459 -1642
rect 7543 -1466 7577 -1450
rect 7543 -1658 7577 -1642
rect 7661 -1466 7695 -1450
rect 7661 -1658 7695 -1642
rect 7779 -1466 7813 -1450
rect 7779 -1658 7813 -1642
rect 7944 -1466 7978 -1450
rect 7944 -1658 7978 -1642
rect 8062 -1466 8096 -1450
rect 8062 -1658 8096 -1642
rect 8180 -1466 8214 -1450
rect 8180 -1658 8214 -1642
rect 8298 -1466 8332 -1450
rect 8298 -1658 8332 -1642
rect 8567 -1470 8601 -1454
rect 8567 -1662 8601 -1646
rect 8685 -1470 8719 -1454
rect 8685 -1662 8719 -1646
rect 8803 -1470 8837 -1454
rect 8803 -1662 8837 -1646
rect 8921 -1470 8955 -1454
rect 8921 -1662 8955 -1646
rect 9086 -1470 9120 -1454
rect 9086 -1662 9120 -1646
rect 9204 -1470 9238 -1454
rect 9204 -1662 9238 -1646
rect 9322 -1470 9356 -1454
rect 9322 -1662 9356 -1646
rect 9440 -1470 9474 -1454
rect 9440 -1662 9474 -1646
rect 10700 -1522 10949 -1479
rect 10700 -1612 10739 -1522
rect 10902 -1612 10949 -1522
rect 11202 -1588 11236 -1572
rect 11320 -1196 11354 -1180
rect 11320 -1588 11354 -1572
rect 11438 -1196 11472 -1180
rect 17501 -1191 17535 -1175
rect 14521 -1410 14537 -1376
rect 14571 -1410 14587 -1376
rect 15663 -1414 15679 -1380
rect 15713 -1414 15729 -1380
rect 17501 -1383 17535 -1367
rect 17619 -1191 17653 -1175
rect 17619 -1383 17653 -1367
rect 17736 -1191 17770 -1175
rect 11438 -1588 11472 -1572
rect 13959 -1461 13993 -1445
rect 10700 -1651 10949 -1612
rect 11245 -1656 11261 -1622
rect 11295 -1656 11311 -1622
rect 11363 -1656 11379 -1622
rect 11413 -1656 11429 -1622
rect 13959 -1653 13993 -1637
rect 14077 -1461 14111 -1445
rect 14077 -1653 14111 -1637
rect 14195 -1461 14229 -1445
rect 14195 -1653 14229 -1637
rect 14313 -1461 14347 -1445
rect 14313 -1653 14347 -1637
rect 14478 -1461 14512 -1445
rect 14478 -1653 14512 -1637
rect 14596 -1461 14630 -1445
rect 14596 -1653 14630 -1637
rect 14714 -1461 14748 -1445
rect 14714 -1653 14748 -1637
rect 14832 -1461 14866 -1445
rect 14832 -1653 14866 -1637
rect 15101 -1465 15135 -1449
rect 15101 -1657 15135 -1641
rect 15219 -1465 15253 -1449
rect 15219 -1657 15253 -1641
rect 15337 -1465 15371 -1449
rect 15337 -1657 15371 -1641
rect 15455 -1465 15489 -1449
rect 15455 -1657 15489 -1641
rect 15620 -1465 15654 -1449
rect 15620 -1657 15654 -1641
rect 15738 -1465 15772 -1449
rect 15738 -1657 15772 -1641
rect 15856 -1465 15890 -1449
rect 15856 -1657 15890 -1641
rect 15974 -1465 16008 -1449
rect 15974 -1657 16008 -1641
rect 17234 -1517 17483 -1474
rect 17234 -1607 17273 -1517
rect 17436 -1607 17483 -1517
rect 17736 -1583 17770 -1567
rect 17854 -1191 17888 -1175
rect 17854 -1583 17888 -1567
rect 17972 -1191 18006 -1175
rect 24014 -1188 24048 -1172
rect 21034 -1407 21050 -1373
rect 21084 -1407 21100 -1373
rect 22176 -1411 22192 -1377
rect 22226 -1411 22242 -1377
rect 24014 -1380 24048 -1364
rect 24132 -1188 24166 -1172
rect 24132 -1380 24166 -1364
rect 24249 -1188 24283 -1172
rect 17972 -1583 18006 -1567
rect 20472 -1458 20506 -1442
rect 17234 -1646 17483 -1607
rect 17779 -1651 17795 -1617
rect 17829 -1651 17845 -1617
rect 17897 -1651 17913 -1617
rect 17947 -1651 17963 -1617
rect 20472 -1650 20506 -1634
rect 20590 -1458 20624 -1442
rect 20590 -1650 20624 -1634
rect 20708 -1458 20742 -1442
rect 20708 -1650 20742 -1634
rect 20826 -1458 20860 -1442
rect 20826 -1650 20860 -1634
rect 20991 -1458 21025 -1442
rect 20991 -1650 21025 -1634
rect 21109 -1458 21143 -1442
rect 21109 -1650 21143 -1634
rect 21227 -1458 21261 -1442
rect 21227 -1650 21261 -1634
rect 21345 -1458 21379 -1442
rect 21345 -1650 21379 -1634
rect 21614 -1462 21648 -1446
rect 21614 -1654 21648 -1638
rect 21732 -1462 21766 -1446
rect 21732 -1654 21766 -1638
rect 21850 -1462 21884 -1446
rect 21850 -1654 21884 -1638
rect 21968 -1462 22002 -1446
rect 21968 -1654 22002 -1638
rect 22133 -1462 22167 -1446
rect 22133 -1654 22167 -1638
rect 22251 -1462 22285 -1446
rect 22251 -1654 22285 -1638
rect 22369 -1462 22403 -1446
rect 22369 -1654 22403 -1638
rect 22487 -1462 22521 -1446
rect 22487 -1654 22521 -1638
rect 23747 -1514 23996 -1471
rect 23747 -1604 23786 -1514
rect 23949 -1604 23996 -1514
rect 24249 -1580 24283 -1564
rect 24367 -1188 24401 -1172
rect 24367 -1580 24401 -1564
rect 24485 -1188 24519 -1172
rect 24485 -1580 24519 -1564
rect 23747 -1643 23996 -1604
rect 24292 -1648 24308 -1614
rect 24342 -1648 24358 -1614
rect 24410 -1648 24426 -1614
rect 24460 -1648 24476 -1614
rect 1587 -1891 1759 -1844
rect 1587 -2054 1630 -1891
rect 1720 -2054 1759 -1891
rect 1587 -2093 1759 -2054
rect 2729 -1889 2901 -1842
rect 2729 -2052 2772 -1889
rect 2862 -2052 2901 -1889
rect 8145 -1895 8317 -1848
rect 2729 -2091 2901 -2052
rect 4519 -1991 4742 -1915
rect 4519 -2140 4596 -1991
rect 4663 -2140 4742 -1991
rect 8145 -2058 8188 -1895
rect 8278 -2058 8317 -1895
rect 8145 -2097 8317 -2058
rect 9287 -1893 9459 -1846
rect 9287 -2056 9330 -1893
rect 9420 -2056 9459 -1893
rect 14679 -1890 14851 -1843
rect 9287 -2095 9459 -2056
rect 11077 -1995 11300 -1919
rect 4519 -2246 4742 -2140
rect 11077 -2144 11154 -1995
rect 11221 -2144 11300 -1995
rect 14679 -2053 14722 -1890
rect 14812 -2053 14851 -1890
rect 14679 -2092 14851 -2053
rect 15821 -1888 15993 -1841
rect 15821 -2051 15864 -1888
rect 15954 -2051 15993 -1888
rect 21192 -1887 21364 -1840
rect 15821 -2090 15993 -2051
rect 17611 -1990 17834 -1914
rect 11077 -2250 11300 -2144
rect 17611 -2139 17688 -1990
rect 17755 -2139 17834 -1990
rect 21192 -2050 21235 -1887
rect 21325 -2050 21364 -1887
rect 21192 -2089 21364 -2050
rect 22334 -1885 22506 -1838
rect 22334 -2048 22377 -1885
rect 22467 -2048 22506 -1885
rect 22334 -2087 22506 -2048
rect 24124 -1987 24347 -1911
rect 17611 -2245 17834 -2139
rect 24124 -2136 24201 -1987
rect 24268 -2136 24347 -1987
rect 24124 -2242 24347 -2136
rect 806 -2334 1031 -2258
rect 806 -2483 885 -2334
rect 952 -2483 1031 -2334
rect 806 -2589 1031 -2483
rect 4041 -2355 4311 -2321
rect 4041 -2405 4075 -2355
rect 4041 -2597 4075 -2581
rect 4159 -2405 4193 -2389
rect 4159 -2597 4193 -2581
rect 4277 -2405 4311 -2355
rect 7364 -2338 7589 -2262
rect 4277 -2597 4311 -2581
rect 4395 -2405 4429 -2389
rect 4395 -2597 4429 -2581
rect 4513 -2405 4547 -2389
rect 4513 -2597 4547 -2581
rect 4631 -2405 4665 -2389
rect 4631 -2597 4665 -2581
rect 4749 -2405 4783 -2389
rect 4749 -2597 4783 -2581
rect 4867 -2405 4901 -2389
rect 4867 -2597 4901 -2581
rect 4985 -2405 5019 -2389
rect 4985 -2597 5019 -2581
rect 5103 -2405 5137 -2389
rect 5103 -2597 5137 -2581
rect 7364 -2487 7443 -2338
rect 7510 -2487 7589 -2338
rect 7364 -2593 7589 -2487
rect 10599 -2359 10869 -2325
rect 10599 -2409 10633 -2359
rect 10599 -2601 10633 -2585
rect 10717 -2409 10751 -2393
rect 10717 -2601 10751 -2585
rect 10835 -2409 10869 -2359
rect 13898 -2333 14123 -2257
rect 10835 -2601 10869 -2585
rect 10953 -2409 10987 -2393
rect 10953 -2601 10987 -2585
rect 11071 -2409 11105 -2393
rect 11071 -2601 11105 -2585
rect 11189 -2409 11223 -2393
rect 11189 -2601 11223 -2585
rect 11307 -2409 11341 -2393
rect 11307 -2601 11341 -2585
rect 11425 -2409 11459 -2393
rect 11425 -2601 11459 -2585
rect 11543 -2409 11577 -2393
rect 11543 -2601 11577 -2585
rect 11661 -2409 11695 -2393
rect 11661 -2601 11695 -2585
rect 13898 -2482 13977 -2333
rect 14044 -2482 14123 -2333
rect 13898 -2588 14123 -2482
rect 17133 -2354 17403 -2320
rect 17133 -2404 17167 -2354
rect 17133 -2596 17167 -2580
rect 17251 -2404 17285 -2388
rect 17251 -2596 17285 -2580
rect 17369 -2404 17403 -2354
rect 20411 -2330 20636 -2254
rect 17369 -2596 17403 -2580
rect 17487 -2404 17521 -2388
rect 17487 -2596 17521 -2580
rect 17605 -2404 17639 -2388
rect 17605 -2596 17639 -2580
rect 17723 -2404 17757 -2388
rect 17723 -2596 17757 -2580
rect 17841 -2404 17875 -2388
rect 17841 -2596 17875 -2580
rect 17959 -2404 17993 -2388
rect 17959 -2596 17993 -2580
rect 18077 -2404 18111 -2388
rect 18077 -2596 18111 -2580
rect 18195 -2404 18229 -2388
rect 18195 -2596 18229 -2580
rect 20411 -2479 20490 -2330
rect 20557 -2479 20636 -2330
rect 20411 -2585 20636 -2479
rect 23646 -2351 23916 -2317
rect 23646 -2401 23680 -2351
rect 23646 -2593 23680 -2577
rect 23764 -2401 23798 -2385
rect 23764 -2593 23798 -2577
rect 23882 -2401 23916 -2351
rect 23882 -2593 23916 -2577
rect 24000 -2401 24034 -2385
rect 24000 -2593 24034 -2577
rect 24118 -2401 24152 -2385
rect 24118 -2593 24152 -2577
rect 24236 -2401 24270 -2385
rect 24236 -2593 24270 -2577
rect 24354 -2401 24388 -2385
rect 24354 -2593 24388 -2577
rect 24472 -2401 24506 -2385
rect 24472 -2593 24506 -2577
rect 24590 -2401 24624 -2385
rect 24590 -2593 24624 -2577
rect 24708 -2401 24742 -2385
rect 24708 -2593 24742 -2577
rect 4320 -2675 4336 -2641
rect 4370 -2675 4386 -2641
rect 10878 -2679 10894 -2645
rect 10928 -2679 10944 -2645
rect 17412 -2674 17428 -2640
rect 17462 -2674 17478 -2640
rect 23925 -2671 23941 -2637
rect 23975 -2671 23991 -2637
rect 667 -2769 937 -2734
rect 549 -2822 583 -2806
rect 66 -3022 100 -3006
rect 66 -3214 100 -3198
rect 184 -3022 218 -3006
rect 184 -3214 218 -3198
rect 302 -3022 336 -3006
rect 302 -3214 336 -3198
rect 420 -3022 454 -3006
rect 420 -3214 454 -3198
rect 549 -3214 583 -3198
rect 667 -2822 701 -2769
rect 667 -3214 701 -3198
rect 785 -2822 819 -2806
rect 785 -3214 819 -3198
rect 903 -2822 937 -2769
rect 2565 -2769 2835 -2734
rect 903 -3214 937 -3198
rect 1021 -2822 1055 -2806
rect 1021 -3214 1055 -3198
rect 1139 -2822 1173 -2806
rect 1139 -3214 1173 -3198
rect 1257 -2822 1291 -2806
rect 2447 -2822 2481 -2806
rect 1505 -2968 1775 -2933
rect 1257 -3214 1291 -3198
rect 1387 -3022 1421 -3006
rect 1387 -3214 1421 -3198
rect 1505 -3022 1539 -2968
rect 1505 -3214 1539 -3198
rect 1623 -3022 1657 -3006
rect 1623 -3214 1657 -3198
rect 1741 -3022 1775 -2968
rect 1741 -3214 1775 -3198
rect 1964 -3022 1998 -3006
rect 1964 -3214 1998 -3198
rect 2082 -3022 2116 -3006
rect 2082 -3214 2116 -3198
rect 2200 -3022 2234 -3006
rect 2200 -3214 2234 -3198
rect 2318 -3022 2352 -3006
rect 2318 -3214 2352 -3198
rect 2447 -3214 2481 -3198
rect 2565 -2822 2599 -2769
rect 2565 -3214 2599 -3198
rect 2683 -2822 2717 -2806
rect 2683 -3214 2717 -3198
rect 2801 -2822 2835 -2769
rect 4438 -2792 4454 -2758
rect 4488 -2792 4504 -2758
rect 7225 -2773 7495 -2738
rect 2801 -3214 2835 -3198
rect 2919 -2822 2953 -2806
rect 2919 -3214 2953 -3198
rect 3037 -2822 3071 -2806
rect 3037 -3214 3071 -3198
rect 3155 -2822 3189 -2806
rect 7107 -2826 7141 -2810
rect 4395 -2842 4429 -2826
rect 3403 -2968 3673 -2933
rect 3155 -3214 3189 -3198
rect 3285 -3022 3319 -3006
rect 3285 -3214 3319 -3198
rect 3403 -3022 3437 -2968
rect 3403 -3214 3437 -3198
rect 3521 -3022 3555 -3006
rect 3521 -3214 3555 -3198
rect 3639 -3022 3673 -2968
rect 4395 -3034 4429 -3018
rect 4513 -2842 4547 -2826
rect 4513 -3034 4547 -3018
rect 4630 -2842 4664 -2826
rect 3639 -3214 3673 -3198
rect 4128 -3168 4377 -3125
rect 4128 -3258 4167 -3168
rect 4330 -3258 4377 -3168
rect 4630 -3234 4664 -3218
rect 4748 -2842 4782 -2826
rect 4748 -3234 4782 -3218
rect 4866 -2842 4900 -2826
rect 6624 -3026 6658 -3010
rect 6624 -3218 6658 -3202
rect 6742 -3026 6776 -3010
rect 6742 -3218 6776 -3202
rect 6860 -3026 6894 -3010
rect 6860 -3218 6894 -3202
rect 6978 -3026 7012 -3010
rect 6978 -3218 7012 -3202
rect 7107 -3218 7141 -3202
rect 7225 -2826 7259 -2773
rect 7225 -3218 7259 -3202
rect 7343 -2826 7377 -2810
rect 7343 -3218 7377 -3202
rect 7461 -2826 7495 -2773
rect 9123 -2773 9393 -2738
rect 7461 -3218 7495 -3202
rect 7579 -2826 7613 -2810
rect 7579 -3218 7613 -3202
rect 7697 -2826 7731 -2810
rect 7697 -3218 7731 -3202
rect 7815 -2826 7849 -2810
rect 9005 -2826 9039 -2810
rect 8063 -2972 8333 -2937
rect 7815 -3218 7849 -3202
rect 7945 -3026 7979 -3010
rect 7945 -3218 7979 -3202
rect 8063 -3026 8097 -2972
rect 8063 -3218 8097 -3202
rect 8181 -3026 8215 -3010
rect 8181 -3218 8215 -3202
rect 8299 -3026 8333 -2972
rect 8299 -3218 8333 -3202
rect 8522 -3026 8556 -3010
rect 8522 -3218 8556 -3202
rect 8640 -3026 8674 -3010
rect 8640 -3218 8674 -3202
rect 8758 -3026 8792 -3010
rect 8758 -3218 8792 -3202
rect 8876 -3026 8910 -3010
rect 8876 -3218 8910 -3202
rect 9005 -3218 9039 -3202
rect 9123 -2826 9157 -2773
rect 9123 -3218 9157 -3202
rect 9241 -2826 9275 -2810
rect 9241 -3218 9275 -3202
rect 9359 -2826 9393 -2773
rect 10996 -2796 11012 -2762
rect 11046 -2796 11062 -2762
rect 13759 -2768 14029 -2733
rect 9359 -3218 9393 -3202
rect 9477 -2826 9511 -2810
rect 9477 -3218 9511 -3202
rect 9595 -2826 9629 -2810
rect 9595 -3218 9629 -3202
rect 9713 -2826 9747 -2810
rect 13641 -2821 13675 -2805
rect 10953 -2846 10987 -2830
rect 9961 -2972 10231 -2937
rect 9713 -3218 9747 -3202
rect 9843 -3026 9877 -3010
rect 9843 -3218 9877 -3202
rect 9961 -3026 9995 -2972
rect 9961 -3218 9995 -3202
rect 10079 -3026 10113 -3010
rect 10079 -3218 10113 -3202
rect 10197 -3026 10231 -2972
rect 10953 -3038 10987 -3022
rect 11071 -2846 11105 -2830
rect 11071 -3038 11105 -3022
rect 11188 -2846 11222 -2830
rect 10197 -3218 10231 -3202
rect 10686 -3172 10935 -3129
rect 4866 -3234 4900 -3218
rect 4128 -3297 4377 -3258
rect 10686 -3262 10725 -3172
rect 10888 -3262 10935 -3172
rect 11188 -3238 11222 -3222
rect 11306 -2846 11340 -2830
rect 11306 -3238 11340 -3222
rect 11424 -2846 11458 -2830
rect 13158 -3021 13192 -3005
rect 13158 -3213 13192 -3197
rect 13276 -3021 13310 -3005
rect 13276 -3213 13310 -3197
rect 13394 -3021 13428 -3005
rect 13394 -3213 13428 -3197
rect 13512 -3021 13546 -3005
rect 13512 -3213 13546 -3197
rect 13641 -3213 13675 -3197
rect 13759 -2821 13793 -2768
rect 13759 -3213 13793 -3197
rect 13877 -2821 13911 -2805
rect 13877 -3213 13911 -3197
rect 13995 -2821 14029 -2768
rect 15657 -2768 15927 -2733
rect 13995 -3213 14029 -3197
rect 14113 -2821 14147 -2805
rect 14113 -3213 14147 -3197
rect 14231 -2821 14265 -2805
rect 14231 -3213 14265 -3197
rect 14349 -2821 14383 -2805
rect 15539 -2821 15573 -2805
rect 14597 -2967 14867 -2932
rect 14349 -3213 14383 -3197
rect 14479 -3021 14513 -3005
rect 14479 -3213 14513 -3197
rect 14597 -3021 14631 -2967
rect 14597 -3213 14631 -3197
rect 14715 -3021 14749 -3005
rect 14715 -3213 14749 -3197
rect 14833 -3021 14867 -2967
rect 14833 -3213 14867 -3197
rect 15056 -3021 15090 -3005
rect 15056 -3213 15090 -3197
rect 15174 -3021 15208 -3005
rect 15174 -3213 15208 -3197
rect 15292 -3021 15326 -3005
rect 15292 -3213 15326 -3197
rect 15410 -3021 15444 -3005
rect 15410 -3213 15444 -3197
rect 15539 -3213 15573 -3197
rect 15657 -2821 15691 -2768
rect 15657 -3213 15691 -3197
rect 15775 -2821 15809 -2805
rect 15775 -3213 15809 -3197
rect 15893 -2821 15927 -2768
rect 17530 -2791 17546 -2757
rect 17580 -2791 17596 -2757
rect 20272 -2765 20542 -2730
rect 15893 -3213 15927 -3197
rect 16011 -2821 16045 -2805
rect 16011 -3213 16045 -3197
rect 16129 -2821 16163 -2805
rect 16129 -3213 16163 -3197
rect 16247 -2821 16281 -2805
rect 20154 -2818 20188 -2802
rect 17487 -2841 17521 -2825
rect 16495 -2967 16765 -2932
rect 16247 -3213 16281 -3197
rect 16377 -3021 16411 -3005
rect 16377 -3213 16411 -3197
rect 16495 -3021 16529 -2967
rect 16495 -3213 16529 -3197
rect 16613 -3021 16647 -3005
rect 16613 -3213 16647 -3197
rect 16731 -3021 16765 -2967
rect 17487 -3033 17521 -3017
rect 17605 -2841 17639 -2825
rect 17605 -3033 17639 -3017
rect 17722 -2841 17756 -2825
rect 16731 -3213 16765 -3197
rect 17220 -3167 17469 -3124
rect 11424 -3238 11458 -3222
rect 4673 -3302 4689 -3268
rect 4723 -3302 4739 -3268
rect 4791 -3302 4807 -3268
rect 4841 -3302 4857 -3268
rect 10686 -3301 10935 -3262
rect 17220 -3257 17259 -3167
rect 17422 -3257 17469 -3167
rect 17722 -3233 17756 -3217
rect 17840 -2841 17874 -2825
rect 17840 -3233 17874 -3217
rect 17958 -2841 17992 -2825
rect 19671 -3018 19705 -3002
rect 19671 -3210 19705 -3194
rect 19789 -3018 19823 -3002
rect 19789 -3210 19823 -3194
rect 19907 -3018 19941 -3002
rect 19907 -3210 19941 -3194
rect 20025 -3018 20059 -3002
rect 20025 -3210 20059 -3194
rect 20154 -3210 20188 -3194
rect 20272 -2818 20306 -2765
rect 20272 -3210 20306 -3194
rect 20390 -2818 20424 -2802
rect 20390 -3210 20424 -3194
rect 20508 -2818 20542 -2765
rect 22170 -2765 22440 -2730
rect 20508 -3210 20542 -3194
rect 20626 -2818 20660 -2802
rect 20626 -3210 20660 -3194
rect 20744 -2818 20778 -2802
rect 20744 -3210 20778 -3194
rect 20862 -2818 20896 -2802
rect 22052 -2818 22086 -2802
rect 21110 -2964 21380 -2929
rect 20862 -3210 20896 -3194
rect 20992 -3018 21026 -3002
rect 20992 -3210 21026 -3194
rect 21110 -3018 21144 -2964
rect 21110 -3210 21144 -3194
rect 21228 -3018 21262 -3002
rect 21228 -3210 21262 -3194
rect 21346 -3018 21380 -2964
rect 21346 -3210 21380 -3194
rect 21569 -3018 21603 -3002
rect 21569 -3210 21603 -3194
rect 21687 -3018 21721 -3002
rect 21687 -3210 21721 -3194
rect 21805 -3018 21839 -3002
rect 21805 -3210 21839 -3194
rect 21923 -3018 21957 -3002
rect 21923 -3210 21957 -3194
rect 22052 -3210 22086 -3194
rect 22170 -2818 22204 -2765
rect 22170 -3210 22204 -3194
rect 22288 -2818 22322 -2802
rect 22288 -3210 22322 -3194
rect 22406 -2818 22440 -2765
rect 24043 -2788 24059 -2754
rect 24093 -2788 24109 -2754
rect 22406 -3210 22440 -3194
rect 22524 -2818 22558 -2802
rect 22524 -3210 22558 -3194
rect 22642 -2818 22676 -2802
rect 22642 -3210 22676 -3194
rect 22760 -2818 22794 -2802
rect 24000 -2838 24034 -2822
rect 23008 -2964 23278 -2929
rect 22760 -3210 22794 -3194
rect 22890 -3018 22924 -3002
rect 22890 -3210 22924 -3194
rect 23008 -3018 23042 -2964
rect 23008 -3210 23042 -3194
rect 23126 -3018 23160 -3002
rect 23126 -3210 23160 -3194
rect 23244 -3018 23278 -2964
rect 24000 -3030 24034 -3014
rect 24118 -2838 24152 -2822
rect 24118 -3030 24152 -3014
rect 24235 -2838 24269 -2822
rect 23244 -3210 23278 -3194
rect 23733 -3164 23982 -3121
rect 17958 -3233 17992 -3217
rect 11231 -3306 11247 -3272
rect 11281 -3306 11297 -3272
rect 11349 -3306 11365 -3272
rect 11399 -3306 11415 -3272
rect 17220 -3296 17469 -3257
rect 23733 -3254 23772 -3164
rect 23935 -3254 23982 -3164
rect 24235 -3230 24269 -3214
rect 24353 -2838 24387 -2822
rect 24353 -3230 24387 -3214
rect 24471 -2838 24505 -2822
rect 24471 -3230 24505 -3214
rect 17765 -3301 17781 -3267
rect 17815 -3301 17831 -3267
rect 17883 -3301 17899 -3267
rect 17933 -3301 17949 -3267
rect 23733 -3293 23982 -3254
rect 24278 -3298 24294 -3264
rect 24328 -3298 24344 -3264
rect 24396 -3298 24412 -3264
rect 24446 -3298 24462 -3264
rect 2175 -3436 2209 -3420
rect 52 -3457 119 -3441
rect 52 -3491 68 -3457
rect 102 -3491 119 -3457
rect 8733 -3440 8767 -3424
rect 15267 -3435 15301 -3419
rect 2175 -3486 2209 -3470
rect 6610 -3461 6677 -3445
rect 52 -3507 119 -3491
rect 6610 -3495 6626 -3461
rect 6660 -3495 6677 -3461
rect 8733 -3490 8767 -3474
rect 13144 -3456 13211 -3440
rect 13144 -3490 13160 -3456
rect 13194 -3490 13211 -3456
rect 21780 -3432 21814 -3416
rect 15267 -3485 15301 -3469
rect 19657 -3453 19724 -3437
rect 606 -3515 640 -3499
rect 724 -3515 758 -3499
rect 606 -3907 640 -3891
rect 722 -3891 724 -3845
rect 35 -3920 135 -3919
rect -21 -3949 135 -3920
rect 722 -3949 758 -3891
rect 842 -3515 876 -3499
rect 842 -3907 876 -3891
rect 960 -3515 994 -3499
rect 1078 -3515 1112 -3499
rect 994 -3891 996 -3844
rect 960 -3949 996 -3891
rect 1196 -3515 1230 -3499
rect 1078 -3907 1112 -3891
rect 1195 -3891 1196 -3844
rect 1314 -3515 1348 -3499
rect 1230 -3891 1231 -3844
rect 1195 -3949 1231 -3891
rect 1314 -3907 1348 -3891
rect 2504 -3515 2538 -3499
rect 2622 -3515 2656 -3499
rect 2504 -3907 2538 -3891
rect 2620 -3891 2622 -3845
rect -21 -3989 1231 -3949
rect 1536 -3949 2033 -3931
rect 2620 -3949 2656 -3891
rect 2740 -3515 2774 -3499
rect 2740 -3907 2774 -3891
rect 2858 -3515 2892 -3499
rect 2976 -3515 3010 -3499
rect 2892 -3891 2894 -3844
rect 2858 -3949 2894 -3891
rect 3094 -3515 3128 -3499
rect 2976 -3907 3010 -3891
rect 3093 -3891 3094 -3844
rect 3212 -3515 3246 -3499
rect 6610 -3511 6677 -3495
rect 3128 -3891 3129 -3844
rect 3093 -3949 3129 -3891
rect 7164 -3519 7198 -3503
rect 4524 -3595 4747 -3519
rect 4524 -3744 4601 -3595
rect 4668 -3744 4747 -3595
rect 4524 -3850 4747 -3744
rect 3212 -3907 3246 -3891
rect 7282 -3519 7316 -3503
rect 7164 -3911 7198 -3895
rect 7280 -3895 7282 -3849
rect 6593 -3924 6693 -3923
rect 1536 -3952 3129 -3949
rect 1536 -3986 1554 -3952
rect 1588 -3986 3129 -3952
rect 1536 -3989 3129 -3986
rect 4046 -3959 4316 -3925
rect -21 -3990 1212 -3989
rect 1536 -3990 3110 -3989
rect -21 -4018 135 -3990
rect 35 -4019 135 -4018
rect 622 -4078 689 -4062
rect 622 -4112 638 -4078
rect 672 -4112 689 -4078
rect 622 -4128 689 -4112
rect 346 -4147 380 -4131
rect 346 -4197 380 -4181
rect 884 -4196 900 -4162
rect 934 -4196 950 -4162
rect 1002 -4197 1018 -4163
rect 1052 -4197 1068 -4163
rect 1123 -4231 1157 -3990
rect 1536 -4007 2033 -3990
rect 1267 -4079 1334 -4063
rect 1267 -4113 1284 -4079
rect 1318 -4113 1334 -4079
rect 1267 -4129 1334 -4113
rect 2518 -4079 2585 -4063
rect 2518 -4113 2534 -4079
rect 2568 -4113 2585 -4079
rect 2518 -4129 2585 -4113
rect 1469 -4146 1503 -4130
rect 1469 -4196 1503 -4180
rect 2244 -4147 2278 -4131
rect 2244 -4197 2278 -4181
rect 2782 -4196 2798 -4162
rect 2832 -4196 2848 -4162
rect 2900 -4197 2916 -4163
rect 2950 -4197 2966 -4163
rect 3021 -4231 3055 -3990
rect 4046 -4009 4080 -3959
rect 3165 -4079 3232 -4063
rect 3165 -4113 3182 -4079
rect 3216 -4113 3232 -4079
rect 3165 -4129 3232 -4113
rect 3367 -4146 3401 -4130
rect 3367 -4196 3401 -4180
rect 4046 -4201 4080 -4185
rect 4164 -4009 4198 -3993
rect 4164 -4201 4198 -4185
rect 4282 -4009 4316 -3959
rect 4282 -4201 4316 -4185
rect 4400 -4009 4434 -3993
rect 4400 -4201 4434 -4185
rect 4518 -4009 4552 -3993
rect 4518 -4201 4552 -4185
rect 4636 -4009 4670 -3993
rect 4636 -4201 4670 -4185
rect 4754 -4009 4788 -3993
rect 4754 -4201 4788 -4185
rect 4872 -4009 4906 -3993
rect 4872 -4201 4906 -4185
rect 4990 -4009 5024 -3993
rect 4990 -4201 5024 -4185
rect 5108 -4009 5142 -3993
rect 6537 -3953 6693 -3924
rect 7280 -3953 7316 -3895
rect 7400 -3519 7434 -3503
rect 7400 -3911 7434 -3895
rect 7518 -3519 7552 -3503
rect 7636 -3519 7670 -3503
rect 7552 -3895 7554 -3848
rect 7518 -3953 7554 -3895
rect 7754 -3519 7788 -3503
rect 7636 -3911 7670 -3895
rect 7753 -3895 7754 -3848
rect 7872 -3519 7906 -3503
rect 7788 -3895 7789 -3848
rect 7753 -3953 7789 -3895
rect 7872 -3911 7906 -3895
rect 9062 -3519 9096 -3503
rect 9180 -3519 9214 -3503
rect 9062 -3911 9096 -3895
rect 9178 -3895 9180 -3849
rect 6537 -3993 7789 -3953
rect 8094 -3953 8591 -3935
rect 9178 -3953 9214 -3895
rect 9298 -3519 9332 -3503
rect 9298 -3911 9332 -3895
rect 9416 -3519 9450 -3503
rect 9534 -3519 9568 -3503
rect 9450 -3895 9452 -3848
rect 9416 -3953 9452 -3895
rect 9652 -3519 9686 -3503
rect 9534 -3911 9568 -3895
rect 9651 -3895 9652 -3848
rect 9770 -3519 9804 -3503
rect 13144 -3506 13211 -3490
rect 19657 -3487 19673 -3453
rect 19707 -3487 19724 -3453
rect 21780 -3482 21814 -3466
rect 9686 -3895 9687 -3848
rect 9651 -3953 9687 -3895
rect 13698 -3514 13732 -3498
rect 11082 -3599 11305 -3523
rect 11082 -3748 11159 -3599
rect 11226 -3748 11305 -3599
rect 11082 -3854 11305 -3748
rect 9770 -3911 9804 -3895
rect 13816 -3514 13850 -3498
rect 13698 -3906 13732 -3890
rect 13814 -3890 13816 -3844
rect 13127 -3919 13227 -3918
rect 8094 -3956 9687 -3953
rect 8094 -3990 8112 -3956
rect 8146 -3990 9687 -3956
rect 8094 -3993 9687 -3990
rect 10604 -3963 10874 -3929
rect 6537 -3994 7770 -3993
rect 8094 -3994 9668 -3993
rect 6537 -4022 6693 -3994
rect 6593 -4023 6693 -4022
rect 7180 -4082 7247 -4066
rect 7180 -4116 7196 -4082
rect 7230 -4116 7247 -4082
rect 7180 -4132 7247 -4116
rect 5108 -4201 5142 -4185
rect 6904 -4151 6938 -4135
rect 6904 -4201 6938 -4185
rect 7442 -4200 7458 -4166
rect 7492 -4200 7508 -4166
rect 7560 -4201 7576 -4167
rect 7610 -4201 7626 -4167
rect 200 -4247 234 -4231
rect 200 -4439 234 -4423
rect 318 -4247 352 -4231
rect 318 -4439 352 -4423
rect 724 -4247 758 -4231
rect 842 -4247 876 -4231
rect 724 -4690 759 -4623
rect 842 -4639 876 -4623
rect 960 -4247 994 -4231
rect 960 -4639 994 -4623
rect 1078 -4247 1157 -4231
rect 1112 -4277 1157 -4247
rect 1196 -4247 1230 -4231
rect 1498 -4247 1532 -4231
rect 1498 -4439 1532 -4423
rect 1616 -4247 1650 -4231
rect 1616 -4439 1650 -4423
rect 2098 -4247 2132 -4231
rect 2098 -4439 2132 -4423
rect 2216 -4247 2250 -4231
rect 2216 -4439 2250 -4423
rect 2622 -4247 2656 -4231
rect 1078 -4639 1112 -4623
rect 1195 -4690 1230 -4623
rect 724 -4725 1230 -4690
rect 2740 -4247 2774 -4231
rect 2622 -4690 2657 -4623
rect 2740 -4639 2774 -4623
rect 2858 -4247 2892 -4231
rect 2858 -4639 2892 -4623
rect 2976 -4247 3055 -4231
rect 3010 -4277 3055 -4247
rect 3094 -4247 3128 -4231
rect 3396 -4247 3430 -4231
rect 3396 -4439 3430 -4423
rect 3514 -4247 3548 -4231
rect 7681 -4235 7715 -3994
rect 8094 -4011 8591 -3994
rect 7825 -4083 7892 -4067
rect 7825 -4117 7842 -4083
rect 7876 -4117 7892 -4083
rect 7825 -4133 7892 -4117
rect 9076 -4083 9143 -4067
rect 9076 -4117 9092 -4083
rect 9126 -4117 9143 -4083
rect 9076 -4133 9143 -4117
rect 8027 -4150 8061 -4134
rect 8027 -4200 8061 -4184
rect 8802 -4151 8836 -4135
rect 8802 -4201 8836 -4185
rect 9340 -4200 9356 -4166
rect 9390 -4200 9406 -4166
rect 9458 -4201 9474 -4167
rect 9508 -4201 9524 -4167
rect 9579 -4235 9613 -3994
rect 10604 -4013 10638 -3963
rect 9723 -4083 9790 -4067
rect 9723 -4117 9740 -4083
rect 9774 -4117 9790 -4083
rect 9723 -4133 9790 -4117
rect 9925 -4150 9959 -4134
rect 9925 -4200 9959 -4184
rect 10604 -4205 10638 -4189
rect 10722 -4013 10756 -3997
rect 10722 -4205 10756 -4189
rect 10840 -4013 10874 -3963
rect 10840 -4205 10874 -4189
rect 10958 -4013 10992 -3997
rect 10958 -4205 10992 -4189
rect 11076 -4013 11110 -3997
rect 11076 -4205 11110 -4189
rect 11194 -4013 11228 -3997
rect 11194 -4205 11228 -4189
rect 11312 -4013 11346 -3997
rect 11312 -4205 11346 -4189
rect 11430 -4013 11464 -3997
rect 11430 -4205 11464 -4189
rect 11548 -4013 11582 -3997
rect 11548 -4205 11582 -4189
rect 11666 -4013 11700 -3997
rect 13071 -3948 13227 -3919
rect 13814 -3948 13850 -3890
rect 13934 -3514 13968 -3498
rect 13934 -3906 13968 -3890
rect 14052 -3514 14086 -3498
rect 14170 -3514 14204 -3498
rect 14086 -3890 14088 -3843
rect 14052 -3948 14088 -3890
rect 14288 -3514 14322 -3498
rect 14170 -3906 14204 -3890
rect 14287 -3890 14288 -3843
rect 14406 -3514 14440 -3498
rect 14322 -3890 14323 -3843
rect 14287 -3948 14323 -3890
rect 14406 -3906 14440 -3890
rect 15596 -3514 15630 -3498
rect 15714 -3514 15748 -3498
rect 15596 -3906 15630 -3890
rect 15712 -3890 15714 -3844
rect 13071 -3988 14323 -3948
rect 14628 -3948 15125 -3930
rect 15712 -3948 15748 -3890
rect 15832 -3514 15866 -3498
rect 15832 -3906 15866 -3890
rect 15950 -3514 15984 -3498
rect 16068 -3514 16102 -3498
rect 15984 -3890 15986 -3843
rect 15950 -3948 15986 -3890
rect 16186 -3514 16220 -3498
rect 16068 -3906 16102 -3890
rect 16185 -3890 16186 -3843
rect 16304 -3514 16338 -3498
rect 19657 -3503 19724 -3487
rect 16220 -3890 16221 -3843
rect 16185 -3948 16221 -3890
rect 20211 -3511 20245 -3495
rect 17616 -3594 17839 -3518
rect 17616 -3743 17693 -3594
rect 17760 -3743 17839 -3594
rect 17616 -3849 17839 -3743
rect 16304 -3906 16338 -3890
rect 20329 -3511 20363 -3495
rect 20211 -3903 20245 -3887
rect 20327 -3887 20329 -3841
rect 19640 -3916 19740 -3915
rect 14628 -3951 16221 -3948
rect 14628 -3985 14646 -3951
rect 14680 -3985 16221 -3951
rect 14628 -3988 16221 -3985
rect 17138 -3958 17408 -3924
rect 13071 -3989 14304 -3988
rect 14628 -3989 16202 -3988
rect 13071 -4017 13227 -3989
rect 13127 -4018 13227 -4017
rect 13714 -4077 13781 -4061
rect 13714 -4111 13730 -4077
rect 13764 -4111 13781 -4077
rect 13714 -4127 13781 -4111
rect 11666 -4205 11700 -4189
rect 13438 -4146 13472 -4130
rect 13438 -4196 13472 -4180
rect 13976 -4195 13992 -4161
rect 14026 -4195 14042 -4161
rect 14094 -4196 14110 -4162
rect 14144 -4196 14160 -4162
rect 14215 -4230 14249 -3989
rect 14628 -4006 15125 -3989
rect 14359 -4078 14426 -4062
rect 14359 -4112 14376 -4078
rect 14410 -4112 14426 -4078
rect 14359 -4128 14426 -4112
rect 15610 -4078 15677 -4062
rect 15610 -4112 15626 -4078
rect 15660 -4112 15677 -4078
rect 15610 -4128 15677 -4112
rect 14561 -4145 14595 -4129
rect 14561 -4195 14595 -4179
rect 15336 -4146 15370 -4130
rect 15336 -4196 15370 -4180
rect 15874 -4195 15890 -4161
rect 15924 -4195 15940 -4161
rect 15992 -4196 16008 -4162
rect 16042 -4196 16058 -4162
rect 16113 -4230 16147 -3989
rect 17138 -4008 17172 -3958
rect 16257 -4078 16324 -4062
rect 16257 -4112 16274 -4078
rect 16308 -4112 16324 -4078
rect 16257 -4128 16324 -4112
rect 16459 -4145 16493 -4129
rect 16459 -4195 16493 -4179
rect 17138 -4200 17172 -4184
rect 17256 -4008 17290 -3992
rect 17256 -4200 17290 -4184
rect 17374 -4008 17408 -3958
rect 17374 -4200 17408 -4184
rect 17492 -4008 17526 -3992
rect 17492 -4200 17526 -4184
rect 17610 -4008 17644 -3992
rect 17610 -4200 17644 -4184
rect 17728 -4008 17762 -3992
rect 17728 -4200 17762 -4184
rect 17846 -4008 17880 -3992
rect 17846 -4200 17880 -4184
rect 17964 -4008 17998 -3992
rect 17964 -4200 17998 -4184
rect 18082 -4008 18116 -3992
rect 18082 -4200 18116 -4184
rect 18200 -4008 18234 -3992
rect 19584 -3945 19740 -3916
rect 20327 -3945 20363 -3887
rect 20447 -3511 20481 -3495
rect 20447 -3903 20481 -3887
rect 20565 -3511 20599 -3495
rect 20683 -3511 20717 -3495
rect 20599 -3887 20601 -3840
rect 20565 -3945 20601 -3887
rect 20801 -3511 20835 -3495
rect 20683 -3903 20717 -3887
rect 20800 -3887 20801 -3840
rect 20919 -3511 20953 -3495
rect 20835 -3887 20836 -3840
rect 20800 -3945 20836 -3887
rect 20919 -3903 20953 -3887
rect 22109 -3511 22143 -3495
rect 22227 -3511 22261 -3495
rect 22109 -3903 22143 -3887
rect 22225 -3887 22227 -3841
rect 19584 -3985 20836 -3945
rect 21141 -3945 21638 -3927
rect 22225 -3945 22261 -3887
rect 22345 -3511 22379 -3495
rect 22345 -3903 22379 -3887
rect 22463 -3511 22497 -3495
rect 22581 -3511 22615 -3495
rect 22497 -3887 22499 -3840
rect 22463 -3945 22499 -3887
rect 22699 -3511 22733 -3495
rect 22581 -3903 22615 -3887
rect 22698 -3887 22699 -3840
rect 22817 -3511 22851 -3495
rect 22733 -3887 22734 -3840
rect 22698 -3945 22734 -3887
rect 24129 -3591 24352 -3515
rect 24129 -3740 24206 -3591
rect 24273 -3740 24352 -3591
rect 24129 -3846 24352 -3740
rect 22817 -3903 22851 -3887
rect 21141 -3948 22734 -3945
rect 21141 -3982 21159 -3948
rect 21193 -3982 22734 -3948
rect 21141 -3985 22734 -3982
rect 23651 -3955 23921 -3921
rect 19584 -3986 20817 -3985
rect 21141 -3986 22715 -3985
rect 19584 -4014 19740 -3986
rect 19640 -4015 19740 -4014
rect 20227 -4074 20294 -4058
rect 20227 -4108 20243 -4074
rect 20277 -4108 20294 -4074
rect 20227 -4124 20294 -4108
rect 18200 -4200 18234 -4184
rect 19951 -4143 19985 -4127
rect 19951 -4193 19985 -4177
rect 20489 -4192 20505 -4158
rect 20539 -4192 20555 -4158
rect 20607 -4193 20623 -4159
rect 20657 -4193 20673 -4159
rect 20728 -4227 20762 -3986
rect 21141 -4003 21638 -3986
rect 20872 -4075 20939 -4059
rect 20872 -4109 20889 -4075
rect 20923 -4109 20939 -4075
rect 20872 -4125 20939 -4109
rect 22123 -4075 22190 -4059
rect 22123 -4109 22139 -4075
rect 22173 -4109 22190 -4075
rect 22123 -4125 22190 -4109
rect 21074 -4142 21108 -4126
rect 21074 -4192 21108 -4176
rect 21849 -4143 21883 -4127
rect 21849 -4193 21883 -4177
rect 22387 -4192 22403 -4158
rect 22437 -4192 22453 -4158
rect 22505 -4193 22521 -4159
rect 22555 -4193 22571 -4159
rect 22626 -4227 22660 -3986
rect 23651 -4005 23685 -3955
rect 22770 -4075 22837 -4059
rect 22770 -4109 22787 -4075
rect 22821 -4109 22837 -4075
rect 22770 -4125 22837 -4109
rect 22972 -4142 23006 -4126
rect 22972 -4192 23006 -4176
rect 23651 -4197 23685 -4181
rect 23769 -4005 23803 -3989
rect 23769 -4197 23803 -4181
rect 23887 -4005 23921 -3955
rect 23887 -4197 23921 -4181
rect 24005 -4005 24039 -3989
rect 24005 -4197 24039 -4181
rect 24123 -4005 24157 -3989
rect 24123 -4197 24157 -4181
rect 24241 -4005 24275 -3989
rect 24241 -4197 24275 -4181
rect 24359 -4005 24393 -3989
rect 24359 -4197 24393 -4181
rect 24477 -4005 24511 -3989
rect 24477 -4197 24511 -4181
rect 24595 -4005 24629 -3989
rect 24595 -4197 24629 -4181
rect 24713 -4005 24747 -3989
rect 24713 -4197 24747 -4181
rect 4325 -4279 4341 -4245
rect 4375 -4279 4391 -4245
rect 6758 -4251 6792 -4235
rect 4443 -4396 4459 -4362
rect 4493 -4396 4509 -4362
rect 3514 -4439 3548 -4423
rect 2976 -4639 3010 -4623
rect 3093 -4690 3128 -4623
rect 4400 -4446 4434 -4430
rect 4400 -4638 4434 -4622
rect 4518 -4446 4552 -4430
rect 4518 -4638 4552 -4622
rect 4635 -4446 4669 -4430
rect 2622 -4725 3128 -4690
rect 4133 -4772 4382 -4729
rect 4133 -4862 4172 -4772
rect 4335 -4862 4382 -4772
rect 4635 -4838 4669 -4822
rect 4753 -4446 4787 -4430
rect 4753 -4838 4787 -4822
rect 4871 -4446 4905 -4430
rect 6758 -4443 6792 -4427
rect 6876 -4251 6910 -4235
rect 6876 -4443 6910 -4427
rect 7282 -4251 7316 -4235
rect 7400 -4251 7434 -4235
rect 7282 -4694 7317 -4627
rect 7400 -4643 7434 -4627
rect 7518 -4251 7552 -4235
rect 7518 -4643 7552 -4627
rect 7636 -4251 7715 -4235
rect 7670 -4281 7715 -4251
rect 7754 -4251 7788 -4235
rect 8056 -4251 8090 -4235
rect 8056 -4443 8090 -4427
rect 8174 -4251 8208 -4235
rect 8174 -4443 8208 -4427
rect 8656 -4251 8690 -4235
rect 8656 -4443 8690 -4427
rect 8774 -4251 8808 -4235
rect 8774 -4443 8808 -4427
rect 9180 -4251 9214 -4235
rect 7636 -4643 7670 -4627
rect 7753 -4694 7788 -4627
rect 7282 -4729 7788 -4694
rect 9298 -4251 9332 -4235
rect 9180 -4694 9215 -4627
rect 9298 -4643 9332 -4627
rect 9416 -4251 9450 -4235
rect 9416 -4643 9450 -4627
rect 9534 -4251 9613 -4235
rect 9568 -4281 9613 -4251
rect 9652 -4251 9686 -4235
rect 9954 -4251 9988 -4235
rect 9954 -4443 9988 -4427
rect 10072 -4251 10106 -4235
rect 13292 -4246 13326 -4230
rect 10883 -4283 10899 -4249
rect 10933 -4283 10949 -4249
rect 11001 -4400 11017 -4366
rect 11051 -4400 11067 -4366
rect 10072 -4443 10106 -4427
rect 9534 -4643 9568 -4627
rect 9651 -4694 9686 -4627
rect 10958 -4450 10992 -4434
rect 10958 -4642 10992 -4626
rect 11076 -4450 11110 -4434
rect 11076 -4642 11110 -4626
rect 11193 -4450 11227 -4434
rect 9180 -4729 9686 -4694
rect 4871 -4838 4905 -4822
rect 10691 -4776 10940 -4733
rect 2785 -4932 2957 -4885
rect 4133 -4901 4382 -4862
rect 10691 -4866 10730 -4776
rect 10893 -4866 10940 -4776
rect 11193 -4842 11227 -4826
rect 11311 -4450 11345 -4434
rect 11311 -4842 11345 -4826
rect 11429 -4450 11463 -4434
rect 13292 -4438 13326 -4422
rect 13410 -4246 13444 -4230
rect 13410 -4438 13444 -4422
rect 13816 -4246 13850 -4230
rect 13934 -4246 13968 -4230
rect 13816 -4689 13851 -4622
rect 13934 -4638 13968 -4622
rect 14052 -4246 14086 -4230
rect 14052 -4638 14086 -4622
rect 14170 -4246 14249 -4230
rect 14204 -4276 14249 -4246
rect 14288 -4246 14322 -4230
rect 14590 -4246 14624 -4230
rect 14590 -4438 14624 -4422
rect 14708 -4246 14742 -4230
rect 14708 -4438 14742 -4422
rect 15190 -4246 15224 -4230
rect 15190 -4438 15224 -4422
rect 15308 -4246 15342 -4230
rect 15308 -4438 15342 -4422
rect 15714 -4246 15748 -4230
rect 14170 -4638 14204 -4622
rect 14287 -4689 14322 -4622
rect 13816 -4724 14322 -4689
rect 15832 -4246 15866 -4230
rect 15714 -4689 15749 -4622
rect 15832 -4638 15866 -4622
rect 15950 -4246 15984 -4230
rect 15950 -4638 15984 -4622
rect 16068 -4246 16147 -4230
rect 16102 -4276 16147 -4246
rect 16186 -4246 16220 -4230
rect 16488 -4246 16522 -4230
rect 16488 -4438 16522 -4422
rect 16606 -4246 16640 -4230
rect 19805 -4243 19839 -4227
rect 17417 -4278 17433 -4244
rect 17467 -4278 17483 -4244
rect 17535 -4395 17551 -4361
rect 17585 -4395 17601 -4361
rect 16606 -4438 16640 -4422
rect 16068 -4638 16102 -4622
rect 16185 -4689 16220 -4622
rect 17492 -4445 17526 -4429
rect 17492 -4637 17526 -4621
rect 17610 -4445 17644 -4429
rect 17610 -4637 17644 -4621
rect 17727 -4445 17761 -4429
rect 15714 -4724 16220 -4689
rect 11429 -4842 11463 -4826
rect 17225 -4771 17474 -4728
rect 4678 -4906 4694 -4872
rect 4728 -4906 4744 -4872
rect 4796 -4906 4812 -4872
rect 4846 -4906 4862 -4872
rect 2785 -5095 2828 -4932
rect 2918 -5095 2957 -4932
rect 2785 -5135 2957 -5095
rect 9343 -4936 9515 -4889
rect 10691 -4905 10940 -4866
rect 17225 -4861 17264 -4771
rect 17427 -4861 17474 -4771
rect 17727 -4837 17761 -4821
rect 17845 -4445 17879 -4429
rect 17845 -4837 17879 -4821
rect 17963 -4445 17997 -4429
rect 19805 -4435 19839 -4419
rect 19923 -4243 19957 -4227
rect 19923 -4435 19957 -4419
rect 20329 -4243 20363 -4227
rect 20447 -4243 20481 -4227
rect 20329 -4686 20364 -4619
rect 20447 -4635 20481 -4619
rect 20565 -4243 20599 -4227
rect 20565 -4635 20599 -4619
rect 20683 -4243 20762 -4227
rect 20717 -4273 20762 -4243
rect 20801 -4243 20835 -4227
rect 21103 -4243 21137 -4227
rect 21103 -4435 21137 -4419
rect 21221 -4243 21255 -4227
rect 21221 -4435 21255 -4419
rect 21703 -4243 21737 -4227
rect 21703 -4435 21737 -4419
rect 21821 -4243 21855 -4227
rect 21821 -4435 21855 -4419
rect 22227 -4243 22261 -4227
rect 20683 -4635 20717 -4619
rect 20800 -4686 20835 -4619
rect 20329 -4721 20835 -4686
rect 22345 -4243 22379 -4227
rect 22227 -4686 22262 -4619
rect 22345 -4635 22379 -4619
rect 22463 -4243 22497 -4227
rect 22463 -4635 22497 -4619
rect 22581 -4243 22660 -4227
rect 22615 -4273 22660 -4243
rect 22699 -4243 22733 -4227
rect 23001 -4243 23035 -4227
rect 23001 -4435 23035 -4419
rect 23119 -4243 23153 -4227
rect 23930 -4275 23946 -4241
rect 23980 -4275 23996 -4241
rect 24048 -4392 24064 -4358
rect 24098 -4392 24114 -4358
rect 23119 -4435 23153 -4419
rect 22581 -4635 22615 -4619
rect 22698 -4686 22733 -4619
rect 24005 -4442 24039 -4426
rect 24005 -4634 24039 -4618
rect 24123 -4442 24157 -4426
rect 24123 -4634 24157 -4618
rect 24240 -4442 24274 -4426
rect 22227 -4721 22733 -4686
rect 17963 -4837 17997 -4821
rect 23738 -4768 23987 -4725
rect 11236 -4910 11252 -4876
rect 11286 -4910 11302 -4876
rect 11354 -4910 11370 -4876
rect 11404 -4910 11420 -4876
rect 9343 -5099 9386 -4936
rect 9476 -5099 9515 -4936
rect 9343 -5139 9515 -5099
rect 15877 -4931 16049 -4884
rect 17225 -4900 17474 -4861
rect 23738 -4858 23777 -4768
rect 23940 -4858 23987 -4768
rect 24240 -4834 24274 -4818
rect 24358 -4442 24392 -4426
rect 24358 -4834 24392 -4818
rect 24476 -4442 24510 -4426
rect 24476 -4834 24510 -4818
rect 17770 -4905 17786 -4871
rect 17820 -4905 17836 -4871
rect 17888 -4905 17904 -4871
rect 17938 -4905 17954 -4871
rect 15877 -5094 15920 -4931
rect 16010 -5094 16049 -4931
rect 15877 -5134 16049 -5094
rect 22390 -4928 22562 -4881
rect 23738 -4897 23987 -4858
rect 24283 -4902 24299 -4868
rect 24333 -4902 24349 -4868
rect 24401 -4902 24417 -4868
rect 24451 -4902 24467 -4868
rect 22390 -5091 22433 -4928
rect 22523 -5091 22562 -4928
rect 22390 -5131 22562 -5091
<< viali >>
rect 3141 5067 3175 5101
rect 4271 5073 4305 5107
rect 9654 5064 9688 5098
rect 10784 5070 10818 5104
rect 16188 5059 16222 5093
rect 17318 5065 17352 5099
rect 22746 5063 22780 5097
rect 23876 5069 23910 5103
rect 3141 4949 3175 4983
rect 4271 4953 4305 4987
rect 931 4677 965 4853
rect 1049 4677 1083 4853
rect 1167 4677 1201 4853
rect 1285 4677 1319 4853
rect 1403 4677 1437 4853
rect 1521 4677 1555 4853
rect 1639 4677 1673 4853
rect 1757 4677 1791 4853
rect 1875 4677 1909 4853
rect 1993 4677 2027 4853
rect 1698 4583 1732 4617
rect 3256 4549 3290 4925
rect 3374 4549 3408 4925
rect 3492 4549 3526 4925
rect 3610 4549 3644 4925
rect 3728 4549 3762 4925
rect 3846 4549 3880 4925
rect 9654 4946 9688 4980
rect 3964 4549 3998 4925
rect 4398 4553 4432 4929
rect 4516 4553 4550 4929
rect 4634 4553 4668 4929
rect 4752 4553 4786 4929
rect 4870 4553 4904 4929
rect 4988 4553 5022 4929
rect 5106 4553 5140 4929
rect 10784 4950 10818 4984
rect 7444 4674 7478 4850
rect 7562 4674 7596 4850
rect 7680 4674 7714 4850
rect 7798 4674 7832 4850
rect 7916 4674 7950 4850
rect 8034 4674 8068 4850
rect 8152 4674 8186 4850
rect 8270 4674 8304 4850
rect 8388 4674 8422 4850
rect 8506 4674 8540 4850
rect 8211 4580 8245 4614
rect 9769 4546 9803 4922
rect 9887 4546 9921 4922
rect 10005 4546 10039 4922
rect 10123 4546 10157 4922
rect 10241 4546 10275 4922
rect 10359 4546 10393 4922
rect 10477 4546 10511 4922
rect 10911 4550 10945 4926
rect 11029 4550 11063 4926
rect 11147 4550 11181 4926
rect 11265 4550 11299 4926
rect 11383 4550 11417 4926
rect 11501 4550 11535 4926
rect 16188 4941 16222 4975
rect 11619 4550 11653 4926
rect 17318 4945 17352 4979
rect 13978 4669 14012 4845
rect 14096 4669 14130 4845
rect 14214 4669 14248 4845
rect 14332 4669 14366 4845
rect 14450 4669 14484 4845
rect 14568 4669 14602 4845
rect 14686 4669 14720 4845
rect 14804 4669 14838 4845
rect 14922 4669 14956 4845
rect 15040 4669 15074 4845
rect 14745 4575 14779 4609
rect 16303 4541 16337 4917
rect 16421 4541 16455 4917
rect 16539 4541 16573 4917
rect 16657 4541 16691 4917
rect 16775 4541 16809 4917
rect 16893 4541 16927 4917
rect 22746 4945 22780 4979
rect 17011 4541 17045 4917
rect 17445 4545 17479 4921
rect 17563 4545 17597 4921
rect 17681 4545 17715 4921
rect 17799 4545 17833 4921
rect 17917 4545 17951 4921
rect 18035 4545 18069 4921
rect 18153 4545 18187 4921
rect 23876 4949 23910 4983
rect 20536 4673 20570 4849
rect 20654 4673 20688 4849
rect 20772 4673 20806 4849
rect 20890 4673 20924 4849
rect 21008 4673 21042 4849
rect 21126 4673 21160 4849
rect 21244 4673 21278 4849
rect 21362 4673 21396 4849
rect 21480 4673 21514 4849
rect 21598 4673 21632 4849
rect 21303 4579 21337 4613
rect 22861 4545 22895 4921
rect 22979 4545 23013 4921
rect 23097 4545 23131 4921
rect 23215 4545 23249 4921
rect 23333 4545 23367 4921
rect 23451 4545 23485 4921
rect 23569 4545 23603 4921
rect 24003 4549 24037 4925
rect 24121 4549 24155 4925
rect 24239 4549 24273 4925
rect 24357 4549 24391 4925
rect 24475 4549 24509 4925
rect 24593 4549 24627 4925
rect 24711 4549 24745 4925
rect 1580 4466 1614 4500
rect 8093 4463 8127 4497
rect 14627 4458 14661 4492
rect 21185 4462 21219 4496
rect 1168 4040 1202 4416
rect 1286 4040 1320 4416
rect 1404 4040 1438 4416
rect 1521 4240 1555 4416
rect 1639 4240 1673 4416
rect 3461 4193 3495 4227
rect 4603 4197 4637 4231
rect 1227 3956 1261 3990
rect 1345 3956 1379 3990
rect 3166 3966 3200 4142
rect 3284 3966 3318 4142
rect 3402 3966 3436 4142
rect 3520 3966 3554 4142
rect 3685 3966 3719 4142
rect 3803 3966 3837 4142
rect 3921 3966 3955 4142
rect 4039 3966 4073 4142
rect 4308 3970 4342 4146
rect 4426 3970 4460 4146
rect 4544 3970 4578 4146
rect 4662 3970 4696 4146
rect 4827 3970 4861 4146
rect 4945 3970 4979 4146
rect 5063 3970 5097 4146
rect 5181 3970 5215 4146
rect 7681 4037 7715 4413
rect 7799 4037 7833 4413
rect 7917 4037 7951 4413
rect 8034 4237 8068 4413
rect 8152 4237 8186 4413
rect 9974 4190 10008 4224
rect 11116 4194 11150 4228
rect 7740 3953 7774 3987
rect 7858 3953 7892 3987
rect 9679 3963 9713 4139
rect 9797 3963 9831 4139
rect 9915 3963 9949 4139
rect 10033 3963 10067 4139
rect 10198 3963 10232 4139
rect 10316 3963 10350 4139
rect 10434 3963 10468 4139
rect 10552 3963 10586 4139
rect 10821 3967 10855 4143
rect 10939 3967 10973 4143
rect 11057 3967 11091 4143
rect 11175 3967 11209 4143
rect 11340 3967 11374 4143
rect 11458 3967 11492 4143
rect 11576 3967 11610 4143
rect 11694 3967 11728 4143
rect 14215 4032 14249 4408
rect 14333 4032 14367 4408
rect 14451 4032 14485 4408
rect 14568 4232 14602 4408
rect 14686 4232 14720 4408
rect 16508 4185 16542 4219
rect 17650 4189 17684 4223
rect 14274 3948 14308 3982
rect 14392 3948 14426 3982
rect 16213 3958 16247 4134
rect 16331 3958 16365 4134
rect 16449 3958 16483 4134
rect 16567 3958 16601 4134
rect 16732 3958 16766 4134
rect 16850 3958 16884 4134
rect 16968 3958 17002 4134
rect 17086 3958 17120 4134
rect 17355 3962 17389 4138
rect 17473 3962 17507 4138
rect 17591 3962 17625 4138
rect 17709 3962 17743 4138
rect 17874 3962 17908 4138
rect 17992 3962 18026 4138
rect 18110 3962 18144 4138
rect 18228 3962 18262 4138
rect 20773 4036 20807 4412
rect 20891 4036 20925 4412
rect 21009 4036 21043 4412
rect 21126 4236 21160 4412
rect 21244 4236 21278 4412
rect 23066 4189 23100 4223
rect 24208 4193 24242 4227
rect 20832 3952 20866 3986
rect 20950 3952 20984 3986
rect 22771 3962 22805 4138
rect 22889 3962 22923 4138
rect 23007 3962 23041 4138
rect 23125 3962 23159 4138
rect 23290 3962 23324 4138
rect 23408 3962 23442 4138
rect 23526 3962 23560 4138
rect 23644 3962 23678 4138
rect 23913 3966 23947 4142
rect 24031 3966 24065 4142
rect 24149 3966 24183 4142
rect 24267 3966 24301 4142
rect 24432 3966 24466 4142
rect 24550 3966 24584 4142
rect 24668 3966 24702 4142
rect 24786 3966 24820 4142
rect 945 3027 979 3203
rect 1063 3027 1097 3203
rect 1181 3027 1215 3203
rect 1299 3027 1333 3203
rect 1417 3027 1451 3203
rect 1535 3027 1569 3203
rect 1653 3027 1687 3203
rect 1771 3027 1805 3203
rect 1889 3027 1923 3203
rect 2007 3027 2041 3203
rect 7458 3024 7492 3200
rect 7576 3024 7610 3200
rect 7694 3024 7728 3200
rect 7812 3024 7846 3200
rect 7930 3024 7964 3200
rect 8048 3024 8082 3200
rect 8166 3024 8200 3200
rect 8284 3024 8318 3200
rect 8402 3024 8436 3200
rect 8520 3024 8554 3200
rect 13992 3019 14026 3195
rect 14110 3019 14144 3195
rect 14228 3019 14262 3195
rect 14346 3019 14380 3195
rect 14464 3019 14498 3195
rect 14582 3019 14616 3195
rect 14700 3019 14734 3195
rect 14818 3019 14852 3195
rect 14936 3019 14970 3195
rect 15054 3019 15088 3195
rect 20550 3023 20584 3199
rect 20668 3023 20702 3199
rect 20786 3023 20820 3199
rect 20904 3023 20938 3199
rect 21022 3023 21056 3199
rect 21140 3023 21174 3199
rect 21258 3023 21292 3199
rect 21376 3023 21410 3199
rect 21494 3023 21528 3199
rect 21612 3023 21646 3199
rect 1712 2933 1746 2967
rect 8225 2930 8259 2964
rect 14759 2925 14793 2959
rect 21317 2929 21351 2963
rect 1594 2816 1628 2850
rect 1182 2390 1216 2766
rect 1300 2390 1334 2766
rect 1418 2390 1452 2766
rect 1535 2590 1569 2766
rect 1653 2590 1687 2766
rect 2409 2410 2443 2586
rect 2527 2410 2561 2586
rect 2645 2410 2679 2586
rect 2763 2410 2797 2586
rect 2893 2410 2927 2786
rect 3011 2410 3045 2786
rect 3129 2410 3163 2786
rect 3247 2410 3281 2786
rect 3365 2410 3399 2786
rect 3483 2410 3517 2786
rect 3601 2410 3635 2786
rect 3730 2410 3764 2586
rect 3848 2410 3882 2586
rect 3966 2410 4000 2586
rect 4084 2410 4118 2586
rect 4307 2410 4341 2586
rect 4425 2410 4459 2586
rect 4543 2410 4577 2586
rect 4661 2410 4695 2586
rect 4791 2410 4825 2786
rect 4909 2410 4943 2786
rect 5027 2410 5061 2786
rect 5145 2410 5179 2786
rect 5263 2410 5297 2786
rect 8107 2813 8141 2847
rect 5381 2410 5415 2786
rect 5499 2410 5533 2786
rect 5628 2410 5662 2586
rect 5746 2410 5780 2586
rect 5864 2410 5898 2586
rect 5982 2410 6016 2586
rect 7695 2387 7729 2763
rect 7813 2387 7847 2763
rect 7931 2387 7965 2763
rect 8048 2587 8082 2763
rect 8166 2587 8200 2763
rect 1241 2306 1275 2340
rect 1359 2306 1393 2340
rect 8922 2407 8956 2583
rect 9040 2407 9074 2583
rect 9158 2407 9192 2583
rect 9276 2407 9310 2583
rect 9406 2407 9440 2783
rect 9524 2407 9558 2783
rect 9642 2407 9676 2783
rect 9760 2407 9794 2783
rect 9878 2407 9912 2783
rect 9996 2407 10030 2783
rect 10114 2407 10148 2783
rect 10243 2407 10277 2583
rect 10361 2407 10395 2583
rect 10479 2407 10513 2583
rect 10597 2407 10631 2583
rect 10820 2407 10854 2583
rect 10938 2407 10972 2583
rect 11056 2407 11090 2583
rect 11174 2407 11208 2583
rect 11304 2407 11338 2783
rect 11422 2407 11456 2783
rect 11540 2407 11574 2783
rect 11658 2407 11692 2783
rect 11776 2407 11810 2783
rect 14641 2808 14675 2842
rect 11894 2407 11928 2783
rect 12012 2407 12046 2783
rect 12141 2407 12175 2583
rect 12259 2407 12293 2583
rect 12377 2407 12411 2583
rect 12495 2407 12529 2583
rect 14229 2382 14263 2758
rect 14347 2382 14381 2758
rect 14465 2382 14499 2758
rect 14582 2582 14616 2758
rect 14700 2582 14734 2758
rect 7754 2303 7788 2337
rect 7872 2303 7906 2337
rect 15456 2402 15490 2578
rect 15574 2402 15608 2578
rect 15692 2402 15726 2578
rect 15810 2402 15844 2578
rect 15940 2402 15974 2778
rect 16058 2402 16092 2778
rect 16176 2402 16210 2778
rect 16294 2402 16328 2778
rect 16412 2402 16446 2778
rect 16530 2402 16564 2778
rect 16648 2402 16682 2778
rect 16777 2402 16811 2578
rect 16895 2402 16929 2578
rect 17013 2402 17047 2578
rect 17131 2402 17165 2578
rect 17354 2402 17388 2578
rect 17472 2402 17506 2578
rect 17590 2402 17624 2578
rect 17708 2402 17742 2578
rect 17838 2402 17872 2778
rect 17956 2402 17990 2778
rect 18074 2402 18108 2778
rect 18192 2402 18226 2778
rect 18310 2402 18344 2778
rect 21199 2812 21233 2846
rect 18428 2402 18462 2778
rect 18546 2402 18580 2778
rect 18675 2402 18709 2578
rect 18793 2402 18827 2578
rect 18911 2402 18945 2578
rect 19029 2402 19063 2578
rect 20787 2386 20821 2762
rect 20905 2386 20939 2762
rect 21023 2386 21057 2762
rect 21140 2586 21174 2762
rect 21258 2586 21292 2762
rect 14288 2298 14322 2332
rect 14406 2298 14440 2332
rect 22014 2406 22048 2582
rect 22132 2406 22166 2582
rect 22250 2406 22284 2582
rect 22368 2406 22402 2582
rect 22498 2406 22532 2782
rect 22616 2406 22650 2782
rect 22734 2406 22768 2782
rect 22852 2406 22886 2782
rect 22970 2406 23004 2782
rect 23088 2406 23122 2782
rect 23206 2406 23240 2782
rect 23335 2406 23369 2582
rect 23453 2406 23487 2582
rect 23571 2406 23605 2582
rect 23689 2406 23723 2582
rect 23912 2406 23946 2582
rect 24030 2406 24064 2582
rect 24148 2406 24182 2582
rect 24266 2406 24300 2582
rect 24396 2406 24430 2782
rect 24514 2406 24548 2782
rect 24632 2406 24666 2782
rect 24750 2406 24784 2782
rect 24868 2406 24902 2782
rect 24986 2406 25020 2782
rect 25104 2406 25138 2782
rect 25233 2406 25267 2582
rect 25351 2406 25385 2582
rect 25469 2406 25503 2582
rect 25587 2406 25621 2582
rect 20846 2302 20880 2336
rect 20964 2302 20998 2336
rect 3873 2138 3907 2172
rect 5980 2117 6014 2151
rect 10386 2135 10420 2169
rect 2836 1717 2870 2093
rect 2954 1717 2988 2093
rect 940 1423 974 1599
rect 1058 1423 1092 1599
rect 1176 1423 1210 1599
rect 1294 1423 1328 1599
rect 1412 1423 1446 1599
rect 1530 1423 1564 1599
rect 1648 1423 1682 1599
rect 1766 1423 1800 1599
rect 1884 1423 1918 1599
rect 3072 1717 3106 2093
rect 3190 1717 3224 2093
rect 3308 1717 3342 2093
rect 3426 1717 3460 2093
rect 3544 1717 3578 2093
rect 4734 1717 4768 2093
rect 4852 1717 4886 2093
rect 4970 1717 5004 2093
rect 5088 1717 5122 2093
rect 5206 1717 5240 2093
rect 5324 1717 5358 2093
rect 12493 2114 12527 2148
rect 16920 2130 16954 2164
rect 5442 1717 5476 2093
rect 9349 1714 9383 2090
rect 9467 1714 9501 2090
rect 2002 1423 2036 1599
rect 2866 1495 2900 1529
rect 2681 1428 2715 1462
rect 3514 1495 3548 1529
rect 4764 1495 4798 1529
rect 3132 1411 3166 1445
rect 3250 1412 3284 1446
rect 3804 1427 3838 1461
rect 4579 1428 4613 1462
rect 6103 1590 6235 1688
rect 5410 1496 5444 1530
rect 5030 1411 5064 1445
rect 5148 1412 5182 1446
rect 5702 1427 5736 1461
rect 7453 1420 7487 1596
rect 7571 1420 7605 1596
rect 7689 1420 7723 1596
rect 7807 1420 7841 1596
rect 7925 1420 7959 1596
rect 8043 1420 8077 1596
rect 8161 1420 8195 1596
rect 8279 1420 8313 1596
rect 8397 1420 8431 1596
rect 9585 1714 9619 2090
rect 9703 1714 9737 2090
rect 9821 1714 9855 2090
rect 9939 1714 9973 2090
rect 10057 1714 10091 2090
rect 11247 1714 11281 2090
rect 11365 1714 11399 2090
rect 11483 1714 11517 2090
rect 11601 1714 11635 2090
rect 11719 1714 11753 2090
rect 11837 1714 11871 2090
rect 19027 2109 19061 2143
rect 23478 2134 23512 2168
rect 11955 1714 11989 2090
rect 15883 1709 15917 2085
rect 16001 1709 16035 2085
rect 8515 1420 8549 1596
rect 9379 1492 9413 1526
rect 9194 1425 9228 1459
rect 1707 1329 1741 1363
rect 1589 1212 1623 1246
rect 2534 1185 2568 1361
rect 1177 786 1211 1162
rect 1295 786 1329 1162
rect 1413 786 1447 1162
rect 1530 986 1564 1162
rect 2652 1185 2686 1361
rect 1648 986 1682 1162
rect 2954 985 2988 1361
rect 3072 985 3106 1361
rect 3190 985 3224 1361
rect 3308 985 3342 1361
rect 3426 985 3460 1361
rect 3832 1185 3866 1361
rect 3950 1185 3984 1361
rect 4432 1185 4466 1361
rect 4550 1185 4584 1361
rect 4852 985 4886 1361
rect 4970 985 5004 1361
rect 5088 985 5122 1361
rect 5206 985 5240 1361
rect 5324 985 5358 1361
rect 5730 1185 5764 1361
rect 10027 1492 10061 1526
rect 11277 1492 11311 1526
rect 9645 1408 9679 1442
rect 9763 1409 9797 1443
rect 10317 1424 10351 1458
rect 11092 1425 11126 1459
rect 12616 1587 12748 1685
rect 11923 1493 11957 1527
rect 11543 1408 11577 1442
rect 11661 1409 11695 1443
rect 12215 1424 12249 1458
rect 13987 1415 14021 1591
rect 14105 1415 14139 1591
rect 14223 1415 14257 1591
rect 14341 1415 14375 1591
rect 14459 1415 14493 1591
rect 14577 1415 14611 1591
rect 14695 1415 14729 1591
rect 14813 1415 14847 1591
rect 14931 1415 14965 1591
rect 16119 1709 16153 2085
rect 16237 1709 16271 2085
rect 16355 1709 16389 2085
rect 16473 1709 16507 2085
rect 16591 1709 16625 2085
rect 17781 1709 17815 2085
rect 17899 1709 17933 2085
rect 18017 1709 18051 2085
rect 18135 1709 18169 2085
rect 18253 1709 18287 2085
rect 18371 1709 18405 2085
rect 25585 2113 25619 2147
rect 18489 1709 18523 2085
rect 22441 1713 22475 2089
rect 22559 1713 22593 2089
rect 15049 1415 15083 1591
rect 15913 1487 15947 1521
rect 15728 1420 15762 1454
rect 5848 1185 5882 1361
rect 8220 1326 8254 1360
rect 8102 1209 8136 1243
rect 9047 1182 9081 1358
rect 7690 783 7724 1159
rect 7808 783 7842 1159
rect 7926 783 7960 1159
rect 8043 983 8077 1159
rect 9165 1182 9199 1358
rect 8161 983 8195 1159
rect 9467 982 9501 1358
rect 9585 982 9619 1358
rect 9703 982 9737 1358
rect 9821 982 9855 1358
rect 9939 982 9973 1358
rect 10345 1182 10379 1358
rect 10463 1182 10497 1358
rect 10945 1182 10979 1358
rect 11063 1182 11097 1358
rect 11365 982 11399 1358
rect 11483 982 11517 1358
rect 11601 982 11635 1358
rect 11719 982 11753 1358
rect 11837 982 11871 1358
rect 12243 1182 12277 1358
rect 16561 1487 16595 1521
rect 17811 1487 17845 1521
rect 16179 1403 16213 1437
rect 16297 1404 16331 1438
rect 16851 1419 16885 1453
rect 17626 1420 17660 1454
rect 19150 1582 19282 1680
rect 18457 1488 18491 1522
rect 18077 1403 18111 1437
rect 18195 1404 18229 1438
rect 18749 1419 18783 1453
rect 20545 1419 20579 1595
rect 20663 1419 20697 1595
rect 20781 1419 20815 1595
rect 20899 1419 20933 1595
rect 21017 1419 21051 1595
rect 21135 1419 21169 1595
rect 21253 1419 21287 1595
rect 21371 1419 21405 1595
rect 21489 1419 21523 1595
rect 22677 1713 22711 2089
rect 22795 1713 22829 2089
rect 22913 1713 22947 2089
rect 23031 1713 23065 2089
rect 23149 1713 23183 2089
rect 24339 1713 24373 2089
rect 24457 1713 24491 2089
rect 24575 1713 24609 2089
rect 24693 1713 24727 2089
rect 24811 1713 24845 2089
rect 24929 1713 24963 2089
rect 25047 1713 25081 2089
rect 21607 1419 21641 1595
rect 22471 1491 22505 1525
rect 22286 1424 22320 1458
rect 23119 1491 23153 1525
rect 24369 1491 24403 1525
rect 22737 1407 22771 1441
rect 22855 1408 22889 1442
rect 23409 1423 23443 1457
rect 24184 1424 24218 1458
rect 25708 1586 25840 1684
rect 25015 1492 25049 1526
rect 24635 1407 24669 1441
rect 24753 1408 24787 1442
rect 25307 1423 25341 1457
rect 12361 1182 12395 1358
rect 14754 1321 14788 1355
rect 14636 1204 14670 1238
rect 15581 1177 15615 1353
rect 1236 702 1270 736
rect 1354 702 1388 736
rect 14224 778 14258 1154
rect 14342 778 14376 1154
rect 14460 778 14494 1154
rect 14577 978 14611 1154
rect 15699 1177 15733 1353
rect 14695 978 14729 1154
rect 16001 977 16035 1353
rect 16119 977 16153 1353
rect 16237 977 16271 1353
rect 16355 977 16389 1353
rect 16473 977 16507 1353
rect 16879 1177 16913 1353
rect 16997 1177 17031 1353
rect 17479 1177 17513 1353
rect 17597 1177 17631 1353
rect 17899 977 17933 1353
rect 18017 977 18051 1353
rect 18135 977 18169 1353
rect 18253 977 18287 1353
rect 18371 977 18405 1353
rect 18777 1177 18811 1353
rect 18895 1177 18929 1353
rect 21312 1325 21346 1359
rect 21194 1208 21228 1242
rect 22139 1181 22173 1357
rect 7749 699 7783 733
rect 7867 699 7901 733
rect 20782 782 20816 1158
rect 20900 782 20934 1158
rect 21018 782 21052 1158
rect 21135 982 21169 1158
rect 22257 1181 22291 1357
rect 21253 982 21287 1158
rect 22559 981 22593 1357
rect 22677 981 22711 1357
rect 22795 981 22829 1357
rect 22913 981 22947 1357
rect 23031 981 23065 1357
rect 23437 1181 23471 1357
rect 23555 1181 23589 1357
rect 24037 1181 24071 1357
rect 24155 1181 24189 1357
rect 24457 981 24491 1357
rect 24575 981 24609 1357
rect 24693 981 24727 1357
rect 24811 981 24845 1357
rect 24929 981 24963 1357
rect 25335 1181 25369 1357
rect 25453 1181 25487 1357
rect 14283 694 14317 728
rect 14401 694 14435 728
rect 20841 698 20875 732
rect 20959 698 20993 732
rect 1777 -535 1811 -501
rect 2907 -541 2941 -507
rect 8335 -539 8369 -505
rect 9465 -545 9499 -511
rect 14869 -534 14903 -500
rect 15999 -540 16033 -506
rect 21382 -531 21416 -497
rect 22512 -537 22546 -503
rect 1777 -655 1811 -621
rect 942 -1055 976 -679
rect 1060 -1055 1094 -679
rect 1178 -1055 1212 -679
rect 1296 -1055 1330 -679
rect 1414 -1055 1448 -679
rect 1532 -1055 1566 -679
rect 2907 -659 2941 -625
rect 1650 -1055 1684 -679
rect 2084 -1059 2118 -683
rect 2202 -1059 2236 -683
rect 2320 -1059 2354 -683
rect 2438 -1059 2472 -683
rect 2556 -1059 2590 -683
rect 2674 -1059 2708 -683
rect 8335 -659 8369 -625
rect 2792 -1059 2826 -683
rect 4055 -931 4089 -755
rect 4173 -931 4207 -755
rect 4291 -931 4325 -755
rect 4409 -931 4443 -755
rect 4527 -931 4561 -755
rect 4645 -931 4679 -755
rect 4763 -931 4797 -755
rect 4881 -931 4915 -755
rect 4999 -931 5033 -755
rect 5117 -931 5151 -755
rect 4350 -1025 4384 -991
rect 7500 -1059 7534 -683
rect 7618 -1059 7652 -683
rect 7736 -1059 7770 -683
rect 7854 -1059 7888 -683
rect 7972 -1059 8006 -683
rect 8090 -1059 8124 -683
rect 9465 -663 9499 -629
rect 14869 -654 14903 -620
rect 8208 -1059 8242 -683
rect 8642 -1063 8676 -687
rect 8760 -1063 8794 -687
rect 8878 -1063 8912 -687
rect 8996 -1063 9030 -687
rect 9114 -1063 9148 -687
rect 9232 -1063 9266 -687
rect 9350 -1063 9384 -687
rect 10613 -935 10647 -759
rect 10731 -935 10765 -759
rect 10849 -935 10883 -759
rect 10967 -935 11001 -759
rect 11085 -935 11119 -759
rect 11203 -935 11237 -759
rect 11321 -935 11355 -759
rect 11439 -935 11473 -759
rect 11557 -935 11591 -759
rect 11675 -935 11709 -759
rect 10908 -1029 10942 -995
rect 14034 -1054 14068 -678
rect 14152 -1054 14186 -678
rect 14270 -1054 14304 -678
rect 14388 -1054 14422 -678
rect 14506 -1054 14540 -678
rect 14624 -1054 14658 -678
rect 15999 -658 16033 -624
rect 14742 -1054 14776 -678
rect 15176 -1058 15210 -682
rect 15294 -1058 15328 -682
rect 15412 -1058 15446 -682
rect 15530 -1058 15564 -682
rect 15648 -1058 15682 -682
rect 15766 -1058 15800 -682
rect 21382 -651 21416 -617
rect 15884 -1058 15918 -682
rect 17147 -930 17181 -754
rect 17265 -930 17299 -754
rect 17383 -930 17417 -754
rect 17501 -930 17535 -754
rect 17619 -930 17653 -754
rect 17737 -930 17771 -754
rect 17855 -930 17889 -754
rect 17973 -930 18007 -754
rect 18091 -930 18125 -754
rect 18209 -930 18243 -754
rect 17442 -1024 17476 -990
rect 20547 -1051 20581 -675
rect 20665 -1051 20699 -675
rect 20783 -1051 20817 -675
rect 20901 -1051 20935 -675
rect 21019 -1051 21053 -675
rect 21137 -1051 21171 -675
rect 22512 -655 22546 -621
rect 21255 -1051 21289 -675
rect 21689 -1055 21723 -679
rect 21807 -1055 21841 -679
rect 21925 -1055 21959 -679
rect 22043 -1055 22077 -679
rect 22161 -1055 22195 -679
rect 22279 -1055 22313 -679
rect 22397 -1055 22431 -679
rect 23660 -927 23694 -751
rect 23778 -927 23812 -751
rect 23896 -927 23930 -751
rect 24014 -927 24048 -751
rect 24132 -927 24166 -751
rect 24250 -927 24284 -751
rect 24368 -927 24402 -751
rect 24486 -927 24520 -751
rect 24604 -927 24638 -751
rect 24722 -927 24756 -751
rect 23955 -1021 23989 -987
rect 4468 -1142 4502 -1108
rect 11026 -1146 11060 -1112
rect 17560 -1141 17594 -1107
rect 24073 -1138 24107 -1104
rect 4409 -1368 4443 -1192
rect 1445 -1411 1479 -1377
rect 2587 -1415 2621 -1381
rect 4527 -1368 4561 -1192
rect 867 -1638 901 -1462
rect 985 -1638 1019 -1462
rect 1103 -1638 1137 -1462
rect 1221 -1638 1255 -1462
rect 1386 -1638 1420 -1462
rect 1504 -1638 1538 -1462
rect 1622 -1638 1656 -1462
rect 1740 -1638 1774 -1462
rect 2009 -1642 2043 -1466
rect 2127 -1642 2161 -1466
rect 2245 -1642 2279 -1466
rect 2363 -1642 2397 -1466
rect 2528 -1642 2562 -1466
rect 2646 -1642 2680 -1466
rect 2764 -1642 2798 -1466
rect 2882 -1642 2916 -1466
rect 4644 -1568 4678 -1192
rect 4762 -1568 4796 -1192
rect 4880 -1568 4914 -1192
rect 10967 -1372 11001 -1196
rect 8003 -1415 8037 -1381
rect 9145 -1419 9179 -1385
rect 11085 -1372 11119 -1196
rect 4703 -1652 4737 -1618
rect 4821 -1652 4855 -1618
rect 7425 -1642 7459 -1466
rect 7543 -1642 7577 -1466
rect 7661 -1642 7695 -1466
rect 7779 -1642 7813 -1466
rect 7944 -1642 7978 -1466
rect 8062 -1642 8096 -1466
rect 8180 -1642 8214 -1466
rect 8298 -1642 8332 -1466
rect 8567 -1646 8601 -1470
rect 8685 -1646 8719 -1470
rect 8803 -1646 8837 -1470
rect 8921 -1646 8955 -1470
rect 9086 -1646 9120 -1470
rect 9204 -1646 9238 -1470
rect 9322 -1646 9356 -1470
rect 9440 -1646 9474 -1470
rect 11202 -1572 11236 -1196
rect 11320 -1572 11354 -1196
rect 11438 -1572 11472 -1196
rect 17501 -1367 17535 -1191
rect 14537 -1410 14571 -1376
rect 15679 -1414 15713 -1380
rect 17619 -1367 17653 -1191
rect 11261 -1656 11295 -1622
rect 11379 -1656 11413 -1622
rect 13959 -1637 13993 -1461
rect 14077 -1637 14111 -1461
rect 14195 -1637 14229 -1461
rect 14313 -1637 14347 -1461
rect 14478 -1637 14512 -1461
rect 14596 -1637 14630 -1461
rect 14714 -1637 14748 -1461
rect 14832 -1637 14866 -1461
rect 15101 -1641 15135 -1465
rect 15219 -1641 15253 -1465
rect 15337 -1641 15371 -1465
rect 15455 -1641 15489 -1465
rect 15620 -1641 15654 -1465
rect 15738 -1641 15772 -1465
rect 15856 -1641 15890 -1465
rect 15974 -1641 16008 -1465
rect 17736 -1567 17770 -1191
rect 17854 -1567 17888 -1191
rect 17972 -1567 18006 -1191
rect 24014 -1364 24048 -1188
rect 21050 -1407 21084 -1373
rect 22192 -1411 22226 -1377
rect 24132 -1364 24166 -1188
rect 17795 -1651 17829 -1617
rect 17913 -1651 17947 -1617
rect 20472 -1634 20506 -1458
rect 20590 -1634 20624 -1458
rect 20708 -1634 20742 -1458
rect 20826 -1634 20860 -1458
rect 20991 -1634 21025 -1458
rect 21109 -1634 21143 -1458
rect 21227 -1634 21261 -1458
rect 21345 -1634 21379 -1458
rect 21614 -1638 21648 -1462
rect 21732 -1638 21766 -1462
rect 21850 -1638 21884 -1462
rect 21968 -1638 22002 -1462
rect 22133 -1638 22167 -1462
rect 22251 -1638 22285 -1462
rect 22369 -1638 22403 -1462
rect 22487 -1638 22521 -1462
rect 24249 -1564 24283 -1188
rect 24367 -1564 24401 -1188
rect 24485 -1564 24519 -1188
rect 24308 -1648 24342 -1614
rect 24426 -1648 24460 -1614
rect 4041 -2581 4075 -2405
rect 4159 -2581 4193 -2405
rect 4277 -2581 4311 -2405
rect 4395 -2581 4429 -2405
rect 4513 -2581 4547 -2405
rect 4631 -2581 4665 -2405
rect 4749 -2581 4783 -2405
rect 4867 -2581 4901 -2405
rect 4985 -2581 5019 -2405
rect 5103 -2581 5137 -2405
rect 10599 -2585 10633 -2409
rect 10717 -2585 10751 -2409
rect 10835 -2585 10869 -2409
rect 10953 -2585 10987 -2409
rect 11071 -2585 11105 -2409
rect 11189 -2585 11223 -2409
rect 11307 -2585 11341 -2409
rect 11425 -2585 11459 -2409
rect 11543 -2585 11577 -2409
rect 11661 -2585 11695 -2409
rect 17133 -2580 17167 -2404
rect 17251 -2580 17285 -2404
rect 17369 -2580 17403 -2404
rect 17487 -2580 17521 -2404
rect 17605 -2580 17639 -2404
rect 17723 -2580 17757 -2404
rect 17841 -2580 17875 -2404
rect 17959 -2580 17993 -2404
rect 18077 -2580 18111 -2404
rect 18195 -2580 18229 -2404
rect 23646 -2577 23680 -2401
rect 23764 -2577 23798 -2401
rect 23882 -2577 23916 -2401
rect 24000 -2577 24034 -2401
rect 24118 -2577 24152 -2401
rect 24236 -2577 24270 -2401
rect 24354 -2577 24388 -2401
rect 24472 -2577 24506 -2401
rect 24590 -2577 24624 -2401
rect 24708 -2577 24742 -2401
rect 4336 -2675 4370 -2641
rect 10894 -2679 10928 -2645
rect 17428 -2674 17462 -2640
rect 23941 -2671 23975 -2637
rect 66 -3198 100 -3022
rect 184 -3198 218 -3022
rect 302 -3198 336 -3022
rect 420 -3198 454 -3022
rect 549 -3198 583 -2822
rect 667 -3198 701 -2822
rect 785 -3198 819 -2822
rect 903 -3198 937 -2822
rect 1021 -3198 1055 -2822
rect 1139 -3198 1173 -2822
rect 1257 -3198 1291 -2822
rect 1387 -3198 1421 -3022
rect 1505 -3198 1539 -3022
rect 1623 -3198 1657 -3022
rect 1741 -3198 1775 -3022
rect 1964 -3198 1998 -3022
rect 2082 -3198 2116 -3022
rect 2200 -3198 2234 -3022
rect 2318 -3198 2352 -3022
rect 2447 -3198 2481 -2822
rect 2565 -3198 2599 -2822
rect 2683 -3198 2717 -2822
rect 4454 -2792 4488 -2758
rect 2801 -3198 2835 -2822
rect 2919 -3198 2953 -2822
rect 3037 -3198 3071 -2822
rect 3155 -3198 3189 -2822
rect 3285 -3198 3319 -3022
rect 3403 -3198 3437 -3022
rect 3521 -3198 3555 -3022
rect 3639 -3198 3673 -3022
rect 4395 -3018 4429 -2842
rect 4513 -3018 4547 -2842
rect 4630 -3218 4664 -2842
rect 4748 -3218 4782 -2842
rect 4866 -3218 4900 -2842
rect 6624 -3202 6658 -3026
rect 6742 -3202 6776 -3026
rect 6860 -3202 6894 -3026
rect 6978 -3202 7012 -3026
rect 7107 -3202 7141 -2826
rect 7225 -3202 7259 -2826
rect 7343 -3202 7377 -2826
rect 7461 -3202 7495 -2826
rect 7579 -3202 7613 -2826
rect 7697 -3202 7731 -2826
rect 7815 -3202 7849 -2826
rect 7945 -3202 7979 -3026
rect 8063 -3202 8097 -3026
rect 8181 -3202 8215 -3026
rect 8299 -3202 8333 -3026
rect 8522 -3202 8556 -3026
rect 8640 -3202 8674 -3026
rect 8758 -3202 8792 -3026
rect 8876 -3202 8910 -3026
rect 9005 -3202 9039 -2826
rect 9123 -3202 9157 -2826
rect 9241 -3202 9275 -2826
rect 11012 -2796 11046 -2762
rect 9359 -3202 9393 -2826
rect 9477 -3202 9511 -2826
rect 9595 -3202 9629 -2826
rect 9713 -3202 9747 -2826
rect 9843 -3202 9877 -3026
rect 9961 -3202 9995 -3026
rect 10079 -3202 10113 -3026
rect 10197 -3202 10231 -3026
rect 10953 -3022 10987 -2846
rect 11071 -3022 11105 -2846
rect 11188 -3222 11222 -2846
rect 11306 -3222 11340 -2846
rect 11424 -3222 11458 -2846
rect 13158 -3197 13192 -3021
rect 13276 -3197 13310 -3021
rect 13394 -3197 13428 -3021
rect 13512 -3197 13546 -3021
rect 13641 -3197 13675 -2821
rect 13759 -3197 13793 -2821
rect 13877 -3197 13911 -2821
rect 13995 -3197 14029 -2821
rect 14113 -3197 14147 -2821
rect 14231 -3197 14265 -2821
rect 14349 -3197 14383 -2821
rect 14479 -3197 14513 -3021
rect 14597 -3197 14631 -3021
rect 14715 -3197 14749 -3021
rect 14833 -3197 14867 -3021
rect 15056 -3197 15090 -3021
rect 15174 -3197 15208 -3021
rect 15292 -3197 15326 -3021
rect 15410 -3197 15444 -3021
rect 15539 -3197 15573 -2821
rect 15657 -3197 15691 -2821
rect 15775 -3197 15809 -2821
rect 17546 -2791 17580 -2757
rect 15893 -3197 15927 -2821
rect 16011 -3197 16045 -2821
rect 16129 -3197 16163 -2821
rect 16247 -3197 16281 -2821
rect 16377 -3197 16411 -3021
rect 16495 -3197 16529 -3021
rect 16613 -3197 16647 -3021
rect 16731 -3197 16765 -3021
rect 17487 -3017 17521 -2841
rect 17605 -3017 17639 -2841
rect 4689 -3302 4723 -3268
rect 4807 -3302 4841 -3268
rect 17722 -3217 17756 -2841
rect 17840 -3217 17874 -2841
rect 17958 -3217 17992 -2841
rect 19671 -3194 19705 -3018
rect 19789 -3194 19823 -3018
rect 19907 -3194 19941 -3018
rect 20025 -3194 20059 -3018
rect 20154 -3194 20188 -2818
rect 20272 -3194 20306 -2818
rect 20390 -3194 20424 -2818
rect 20508 -3194 20542 -2818
rect 20626 -3194 20660 -2818
rect 20744 -3194 20778 -2818
rect 20862 -3194 20896 -2818
rect 20992 -3194 21026 -3018
rect 21110 -3194 21144 -3018
rect 21228 -3194 21262 -3018
rect 21346 -3194 21380 -3018
rect 21569 -3194 21603 -3018
rect 21687 -3194 21721 -3018
rect 21805 -3194 21839 -3018
rect 21923 -3194 21957 -3018
rect 22052 -3194 22086 -2818
rect 22170 -3194 22204 -2818
rect 22288 -3194 22322 -2818
rect 24059 -2788 24093 -2754
rect 22406 -3194 22440 -2818
rect 22524 -3194 22558 -2818
rect 22642 -3194 22676 -2818
rect 22760 -3194 22794 -2818
rect 22890 -3194 22924 -3018
rect 23008 -3194 23042 -3018
rect 23126 -3194 23160 -3018
rect 23244 -3194 23278 -3018
rect 24000 -3014 24034 -2838
rect 24118 -3014 24152 -2838
rect 11247 -3306 11281 -3272
rect 11365 -3306 11399 -3272
rect 24235 -3214 24269 -2838
rect 24353 -3214 24387 -2838
rect 24471 -3214 24505 -2838
rect 17781 -3301 17815 -3267
rect 17899 -3301 17933 -3267
rect 24294 -3298 24328 -3264
rect 24412 -3298 24446 -3264
rect 68 -3491 102 -3457
rect 2175 -3470 2209 -3436
rect 6626 -3495 6660 -3461
rect 8733 -3474 8767 -3440
rect 13160 -3490 13194 -3456
rect 15267 -3469 15301 -3435
rect 606 -3891 640 -3515
rect 724 -3891 758 -3515
rect -153 -4018 -21 -3920
rect 842 -3891 876 -3515
rect 960 -3891 994 -3515
rect 1078 -3891 1112 -3515
rect 1196 -3891 1230 -3515
rect 1314 -3891 1348 -3515
rect 2504 -3891 2538 -3515
rect 2622 -3891 2656 -3515
rect 2740 -3891 2774 -3515
rect 2858 -3891 2892 -3515
rect 2976 -3891 3010 -3515
rect 3094 -3891 3128 -3515
rect 3212 -3891 3246 -3515
rect 7164 -3895 7198 -3519
rect 7282 -3895 7316 -3519
rect 638 -4112 672 -4078
rect 346 -4181 380 -4147
rect 900 -4196 934 -4162
rect 1018 -4197 1052 -4163
rect 1284 -4113 1318 -4079
rect 2534 -4113 2568 -4079
rect 1469 -4180 1503 -4146
rect 2244 -4181 2278 -4147
rect 2798 -4196 2832 -4162
rect 2916 -4197 2950 -4163
rect 3182 -4113 3216 -4079
rect 3367 -4180 3401 -4146
rect 4046 -4185 4080 -4009
rect 4164 -4185 4198 -4009
rect 4282 -4185 4316 -4009
rect 4400 -4185 4434 -4009
rect 4518 -4185 4552 -4009
rect 4636 -4185 4670 -4009
rect 4754 -4185 4788 -4009
rect 4872 -4185 4906 -4009
rect 4990 -4185 5024 -4009
rect 5108 -4185 5142 -4009
rect 6405 -4022 6537 -3924
rect 7400 -3895 7434 -3519
rect 7518 -3895 7552 -3519
rect 7636 -3895 7670 -3519
rect 7754 -3895 7788 -3519
rect 7872 -3895 7906 -3519
rect 9062 -3895 9096 -3519
rect 9180 -3895 9214 -3519
rect 9298 -3895 9332 -3519
rect 9416 -3895 9450 -3519
rect 9534 -3895 9568 -3519
rect 9652 -3895 9686 -3519
rect 19673 -3487 19707 -3453
rect 21780 -3466 21814 -3432
rect 9770 -3895 9804 -3519
rect 13698 -3890 13732 -3514
rect 13816 -3890 13850 -3514
rect 7196 -4116 7230 -4082
rect 6904 -4185 6938 -4151
rect 7458 -4200 7492 -4166
rect 7576 -4201 7610 -4167
rect 200 -4423 234 -4247
rect 318 -4423 352 -4247
rect 724 -4623 758 -4247
rect 842 -4623 876 -4247
rect 960 -4623 994 -4247
rect 1078 -4623 1112 -4247
rect 1196 -4623 1230 -4247
rect 1498 -4423 1532 -4247
rect 1616 -4423 1650 -4247
rect 2098 -4423 2132 -4247
rect 2216 -4423 2250 -4247
rect 2622 -4623 2656 -4247
rect 2740 -4623 2774 -4247
rect 2858 -4623 2892 -4247
rect 2976 -4623 3010 -4247
rect 3094 -4623 3128 -4247
rect 3396 -4423 3430 -4247
rect 7842 -4117 7876 -4083
rect 9092 -4117 9126 -4083
rect 8027 -4184 8061 -4150
rect 8802 -4185 8836 -4151
rect 9356 -4200 9390 -4166
rect 9474 -4201 9508 -4167
rect 9740 -4117 9774 -4083
rect 9925 -4184 9959 -4150
rect 10604 -4189 10638 -4013
rect 10722 -4189 10756 -4013
rect 10840 -4189 10874 -4013
rect 10958 -4189 10992 -4013
rect 11076 -4189 11110 -4013
rect 11194 -4189 11228 -4013
rect 11312 -4189 11346 -4013
rect 11430 -4189 11464 -4013
rect 11548 -4189 11582 -4013
rect 11666 -4189 11700 -4013
rect 12939 -4017 13071 -3919
rect 13934 -3890 13968 -3514
rect 14052 -3890 14086 -3514
rect 14170 -3890 14204 -3514
rect 14288 -3890 14322 -3514
rect 14406 -3890 14440 -3514
rect 15596 -3890 15630 -3514
rect 15714 -3890 15748 -3514
rect 15832 -3890 15866 -3514
rect 15950 -3890 15984 -3514
rect 16068 -3890 16102 -3514
rect 16186 -3890 16220 -3514
rect 16304 -3890 16338 -3514
rect 20211 -3887 20245 -3511
rect 20329 -3887 20363 -3511
rect 13730 -4111 13764 -4077
rect 13438 -4180 13472 -4146
rect 13992 -4195 14026 -4161
rect 14110 -4196 14144 -4162
rect 14376 -4112 14410 -4078
rect 15626 -4112 15660 -4078
rect 14561 -4179 14595 -4145
rect 15336 -4180 15370 -4146
rect 15890 -4195 15924 -4161
rect 16008 -4196 16042 -4162
rect 16274 -4112 16308 -4078
rect 16459 -4179 16493 -4145
rect 17138 -4184 17172 -4008
rect 17256 -4184 17290 -4008
rect 17374 -4184 17408 -4008
rect 17492 -4184 17526 -4008
rect 17610 -4184 17644 -4008
rect 17728 -4184 17762 -4008
rect 17846 -4184 17880 -4008
rect 17964 -4184 17998 -4008
rect 18082 -4184 18116 -4008
rect 18200 -4184 18234 -4008
rect 19452 -4014 19584 -3916
rect 20447 -3887 20481 -3511
rect 20565 -3887 20599 -3511
rect 20683 -3887 20717 -3511
rect 20801 -3887 20835 -3511
rect 20919 -3887 20953 -3511
rect 22109 -3887 22143 -3511
rect 22227 -3887 22261 -3511
rect 22345 -3887 22379 -3511
rect 22463 -3887 22497 -3511
rect 22581 -3887 22615 -3511
rect 22699 -3887 22733 -3511
rect 22817 -3887 22851 -3511
rect 20243 -4108 20277 -4074
rect 19951 -4177 19985 -4143
rect 20505 -4192 20539 -4158
rect 20623 -4193 20657 -4159
rect 20889 -4109 20923 -4075
rect 22139 -4109 22173 -4075
rect 21074 -4176 21108 -4142
rect 21849 -4177 21883 -4143
rect 22403 -4192 22437 -4158
rect 22521 -4193 22555 -4159
rect 22787 -4109 22821 -4075
rect 22972 -4176 23006 -4142
rect 23651 -4181 23685 -4005
rect 23769 -4181 23803 -4005
rect 23887 -4181 23921 -4005
rect 24005 -4181 24039 -4005
rect 24123 -4181 24157 -4005
rect 24241 -4181 24275 -4005
rect 24359 -4181 24393 -4005
rect 24477 -4181 24511 -4005
rect 24595 -4181 24629 -4005
rect 24713 -4181 24747 -4005
rect 3514 -4423 3548 -4247
rect 4341 -4279 4375 -4245
rect 4459 -4396 4493 -4362
rect 6758 -4427 6792 -4251
rect 4400 -4622 4434 -4446
rect 4518 -4622 4552 -4446
rect 4635 -4822 4669 -4446
rect 4753 -4822 4787 -4446
rect 6876 -4427 6910 -4251
rect 4871 -4822 4905 -4446
rect 7282 -4627 7316 -4251
rect 7400 -4627 7434 -4251
rect 7518 -4627 7552 -4251
rect 7636 -4627 7670 -4251
rect 7754 -4627 7788 -4251
rect 8056 -4427 8090 -4251
rect 8174 -4427 8208 -4251
rect 8656 -4427 8690 -4251
rect 8774 -4427 8808 -4251
rect 9180 -4627 9214 -4251
rect 9298 -4627 9332 -4251
rect 9416 -4627 9450 -4251
rect 9534 -4627 9568 -4251
rect 9652 -4627 9686 -4251
rect 9954 -4427 9988 -4251
rect 10072 -4427 10106 -4251
rect 10899 -4283 10933 -4249
rect 11017 -4400 11051 -4366
rect 13292 -4422 13326 -4246
rect 10958 -4626 10992 -4450
rect 11076 -4626 11110 -4450
rect 11193 -4826 11227 -4450
rect 11311 -4826 11345 -4450
rect 13410 -4422 13444 -4246
rect 11429 -4826 11463 -4450
rect 13816 -4622 13850 -4246
rect 13934 -4622 13968 -4246
rect 14052 -4622 14086 -4246
rect 14170 -4622 14204 -4246
rect 14288 -4622 14322 -4246
rect 14590 -4422 14624 -4246
rect 14708 -4422 14742 -4246
rect 15190 -4422 15224 -4246
rect 15308 -4422 15342 -4246
rect 15714 -4622 15748 -4246
rect 15832 -4622 15866 -4246
rect 15950 -4622 15984 -4246
rect 16068 -4622 16102 -4246
rect 16186 -4622 16220 -4246
rect 16488 -4422 16522 -4246
rect 16606 -4422 16640 -4246
rect 17433 -4278 17467 -4244
rect 17551 -4395 17585 -4361
rect 19805 -4419 19839 -4243
rect 17492 -4621 17526 -4445
rect 17610 -4621 17644 -4445
rect 4694 -4906 4728 -4872
rect 4812 -4906 4846 -4872
rect 17727 -4821 17761 -4445
rect 17845 -4821 17879 -4445
rect 19923 -4419 19957 -4243
rect 17963 -4821 17997 -4445
rect 20329 -4619 20363 -4243
rect 20447 -4619 20481 -4243
rect 20565 -4619 20599 -4243
rect 20683 -4619 20717 -4243
rect 20801 -4619 20835 -4243
rect 21103 -4419 21137 -4243
rect 21221 -4419 21255 -4243
rect 21703 -4419 21737 -4243
rect 21821 -4419 21855 -4243
rect 22227 -4619 22261 -4243
rect 22345 -4619 22379 -4243
rect 22463 -4619 22497 -4243
rect 22581 -4619 22615 -4243
rect 22699 -4619 22733 -4243
rect 23001 -4419 23035 -4243
rect 23119 -4419 23153 -4243
rect 23946 -4275 23980 -4241
rect 24064 -4392 24098 -4358
rect 24005 -4618 24039 -4442
rect 24123 -4618 24157 -4442
rect 11252 -4910 11286 -4876
rect 11370 -4910 11404 -4876
rect 24240 -4818 24274 -4442
rect 24358 -4818 24392 -4442
rect 24476 -4818 24510 -4442
rect 17786 -4905 17820 -4871
rect 17904 -4905 17938 -4871
rect 24299 -4902 24333 -4868
rect 24417 -4902 24451 -4868
<< metal1 >>
rect 1328 5151 1548 5171
rect 1328 5043 1372 5151
rect 1504 5043 1548 5151
rect 3125 5109 3181 5117
rect 1328 5001 1548 5043
rect 2199 5101 3181 5109
rect 2199 5067 3141 5101
rect 3175 5067 3181 5101
rect 3844 5097 3854 5205
rect 3986 5142 3996 5205
rect 3986 5131 3998 5142
rect 3986 5097 3999 5131
rect 4255 5121 4311 5123
rect 2199 5051 3181 5067
rect 3854 5059 3999 5097
rect 2199 5050 3178 5051
rect 932 4971 1909 5001
rect 932 4865 964 4971
rect 1168 4865 1200 4971
rect 1404 4865 1436 4971
rect 1640 4865 1672 4971
rect 1875 4865 1909 4971
rect 925 4853 971 4865
rect 925 4677 931 4853
rect 965 4677 971 4853
rect 925 4665 971 4677
rect 1043 4853 1089 4865
rect 1043 4677 1049 4853
rect 1083 4677 1089 4853
rect 1043 4665 1089 4677
rect 1161 4853 1207 4865
rect 1161 4677 1167 4853
rect 1201 4677 1207 4853
rect 1161 4665 1207 4677
rect 1279 4853 1325 4865
rect 1279 4677 1285 4853
rect 1319 4677 1325 4853
rect 1279 4665 1325 4677
rect 1397 4853 1443 4865
rect 1397 4677 1403 4853
rect 1437 4677 1443 4853
rect 1397 4665 1443 4677
rect 1515 4853 1561 4865
rect 1515 4677 1521 4853
rect 1555 4677 1561 4853
rect 1515 4665 1561 4677
rect 1633 4853 1679 4865
rect 1633 4677 1639 4853
rect 1673 4677 1679 4853
rect 1633 4665 1679 4677
rect 1751 4853 1797 4865
rect 1751 4677 1757 4853
rect 1791 4677 1797 4853
rect 1751 4665 1797 4677
rect 1869 4853 1915 4865
rect 1869 4677 1875 4853
rect 1909 4677 1915 4853
rect 1869 4665 1915 4677
rect 1987 4853 2033 4865
rect 1987 4677 1993 4853
rect 2027 4677 2033 4853
rect 1987 4665 2033 4677
rect 1048 4571 1084 4665
rect 1284 4571 1320 4665
rect 1520 4572 1556 4665
rect 1682 4617 1748 4624
rect 1682 4583 1698 4617
rect 1732 4583 1748 4617
rect 1682 4572 1748 4583
rect 1520 4571 1748 4572
rect 1048 4542 1748 4571
rect 1048 4541 1630 4542
rect 1168 4428 1202 4541
rect 1564 4500 1630 4541
rect 1564 4466 1580 4500
rect 1614 4466 1630 4500
rect 1564 4459 1630 4466
rect 1992 4460 2027 4665
rect 2199 4460 2266 5050
rect 3958 5027 3999 5059
rect 4245 5055 4255 5121
rect 4311 5055 4321 5121
rect 4991 5097 5001 5205
rect 5133 5142 5143 5205
rect 7841 5148 8061 5168
rect 5133 5131 5145 5142
rect 5133 5097 5146 5131
rect 5001 5059 5146 5097
rect 5105 5031 5146 5059
rect 3374 4999 3644 5027
rect 3115 4933 3125 4999
rect 3191 4933 3201 4999
rect 3374 4937 3408 4999
rect 3610 4937 3644 4999
rect 3728 4999 3999 5027
rect 4516 5003 4786 5031
rect 3728 4937 3762 4999
rect 3964 4937 3999 4999
rect 4140 4987 4311 5003
rect 4140 4953 4271 4987
rect 4305 4953 4311 4987
rect 4140 4937 4311 4953
rect 4516 4941 4550 5003
rect 4752 4941 4786 5003
rect 4870 5003 5146 5031
rect 4870 4941 4904 5003
rect 5106 4941 5146 5003
rect 7841 5040 7885 5148
rect 8017 5040 8061 5148
rect 9638 5106 9694 5114
rect 7841 4998 8061 5040
rect 8712 5098 9694 5106
rect 8712 5064 9654 5098
rect 9688 5064 9694 5098
rect 10357 5094 10367 5202
rect 10499 5139 10509 5202
rect 10499 5128 10511 5139
rect 10499 5094 10512 5128
rect 10768 5118 10824 5120
rect 8712 5048 9694 5064
rect 10367 5056 10512 5094
rect 8712 5047 9691 5048
rect 3250 4925 3296 4937
rect 3250 4549 3256 4925
rect 3290 4549 3296 4925
rect 3250 4537 3296 4549
rect 3368 4925 3414 4937
rect 3368 4549 3374 4925
rect 3408 4549 3414 4925
rect 3368 4537 3414 4549
rect 3486 4925 3532 4937
rect 3486 4549 3492 4925
rect 3526 4549 3532 4925
rect 3486 4537 3532 4549
rect 3604 4925 3650 4937
rect 3604 4549 3610 4925
rect 3644 4549 3650 4925
rect 3604 4537 3650 4549
rect 3722 4925 3768 4937
rect 3722 4549 3728 4925
rect 3762 4549 3768 4925
rect 3722 4537 3768 4549
rect 3840 4925 3886 4937
rect 3840 4549 3846 4925
rect 3880 4549 3886 4925
rect 3840 4537 3886 4549
rect 3958 4925 4004 4937
rect 3958 4549 3964 4925
rect 3998 4549 4004 4925
rect 3958 4537 4004 4549
rect 1992 4432 2266 4460
rect 1638 4428 2266 4432
rect 1162 4416 1208 4428
rect -10 4023 279 4198
rect 1162 4040 1168 4416
rect 1202 4040 1208 4416
rect 1162 4028 1208 4040
rect 1280 4416 1326 4428
rect 1280 4040 1286 4416
rect 1320 4040 1326 4416
rect 1280 4028 1326 4040
rect 1398 4416 1444 4428
rect 1398 4040 1404 4416
rect 1438 4064 1444 4416
rect 1515 4416 1561 4428
rect 1515 4240 1521 4416
rect 1555 4240 1561 4416
rect 1515 4228 1561 4240
rect 1633 4416 2266 4428
rect 1633 4240 1639 4416
rect 1673 4403 2266 4416
rect 3256 4495 3290 4537
rect 3492 4495 3526 4537
rect 3256 4467 3526 4495
rect 3610 4496 3644 4537
rect 3846 4496 3880 4537
rect 3610 4467 3880 4496
rect 3256 4419 3290 4467
rect 1673 4240 1679 4403
rect 3256 4389 3319 4419
rect 1633 4228 1679 4240
rect 3284 4297 3319 4389
rect 3284 4261 3511 4297
rect 3781 4286 3791 4383
rect 3890 4286 3900 4383
rect 3964 4354 3998 4537
rect 3964 4300 4073 4354
rect 1521 4112 1556 4228
rect 3284 4154 3319 4261
rect 3445 4227 3511 4261
rect 3445 4193 3461 4227
rect 3495 4193 3511 4227
rect 3792 4285 3889 4286
rect 3792 4218 3849 4285
rect 3445 4187 3511 4193
rect 3686 4182 3955 4218
rect 3686 4154 3719 4182
rect 3922 4154 3955 4182
rect 4039 4154 4073 4300
rect 3160 4142 3206 4154
rect 1652 4112 1760 4122
rect 1521 4064 1652 4112
rect 1438 4040 1652 4064
rect 1398 4028 1652 4040
rect 1404 4024 1652 4028
rect -10 3996 1040 4023
rect -10 3990 1277 3996
rect -10 3956 1227 3990
rect 1261 3956 1277 3990
rect -10 3940 1277 3956
rect 1329 3990 1395 3996
rect 1329 3956 1345 3990
rect 1379 3956 1395 3990
rect 1578 3980 1652 4024
rect 1652 3970 1760 3980
rect -10 3924 1040 3940
rect -10 3923 977 3924
rect -10 3919 512 3923
rect -10 3918 279 3919
rect 7 3508 296 3670
rect 7 3402 144 3508
rect 256 3495 296 3508
rect 256 3402 298 3495
rect 7 3391 298 3402
rect 7 3390 296 3391
rect 7 2396 295 2558
rect 7 2290 143 2396
rect 255 2394 295 2396
rect 261 2383 295 2394
rect 7 2288 149 2290
rect 261 2288 296 2383
rect 7 2279 296 2288
rect 7 2278 295 2279
rect 7 2277 263 2278
rect 419 2025 512 3919
rect 575 3860 1041 3882
rect 1329 3860 1395 3956
rect 3160 3966 3166 4142
rect 3200 3966 3206 4142
rect 3160 3954 3206 3966
rect 3278 4142 3324 4154
rect 3278 3966 3284 4142
rect 3318 3966 3324 4142
rect 3278 3954 3324 3966
rect 3396 4142 3442 4154
rect 3396 3966 3402 4142
rect 3436 3966 3442 4142
rect 3396 3954 3442 3966
rect 3514 4142 3560 4154
rect 3514 3966 3520 4142
rect 3554 4087 3560 4142
rect 3679 4142 3725 4154
rect 3679 4087 3685 4142
rect 3554 3999 3685 4087
rect 3554 3966 3560 3999
rect 3514 3954 3560 3966
rect 3679 3966 3685 3999
rect 3719 3966 3725 4142
rect 3679 3954 3725 3966
rect 3797 4142 3843 4154
rect 3797 3966 3803 4142
rect 3837 3966 3843 4142
rect 3797 3954 3843 3966
rect 3915 4142 3961 4154
rect 3915 3966 3921 4142
rect 3955 3966 3961 4142
rect 3915 3954 3961 3966
rect 4033 4142 4079 4154
rect 4033 3966 4039 4142
rect 4073 3966 4079 4142
rect 4033 3954 4079 3966
rect 3166 3915 3200 3954
rect 3402 3915 3436 3954
rect 3166 3880 3436 3915
rect 3803 3916 3836 3954
rect 4039 3916 4072 3954
rect 3803 3880 4072 3916
rect 575 3812 1395 3860
rect 3200 3879 3436 3880
rect 575 3781 1041 3812
rect 3200 3805 3332 3879
rect 575 3525 680 3781
rect 3190 3697 3200 3805
rect 3332 3697 3342 3805
rect 575 3419 638 3525
rect 750 3419 760 3525
rect 1342 3501 1562 3521
rect 575 3408 724 3419
rect 575 2231 680 3408
rect 1342 3393 1386 3501
rect 1518 3393 1562 3501
rect 1342 3351 1562 3393
rect 4140 3366 4202 4937
rect 4392 4929 4438 4941
rect 4392 4553 4398 4929
rect 4432 4553 4438 4929
rect 4392 4541 4438 4553
rect 4510 4929 4556 4941
rect 4510 4553 4516 4929
rect 4550 4553 4556 4929
rect 4510 4541 4556 4553
rect 4628 4929 4674 4941
rect 4628 4553 4634 4929
rect 4668 4553 4674 4929
rect 4628 4541 4674 4553
rect 4746 4929 4792 4941
rect 4746 4553 4752 4929
rect 4786 4553 4792 4929
rect 4746 4541 4792 4553
rect 4864 4929 4910 4941
rect 4864 4553 4870 4929
rect 4904 4553 4910 4929
rect 4864 4541 4910 4553
rect 4982 4929 5028 4941
rect 4982 4553 4988 4929
rect 5022 4553 5028 4929
rect 4982 4541 5028 4553
rect 5100 4929 5146 4941
rect 5100 4553 5106 4929
rect 5140 4553 5146 4929
rect 7445 4968 8422 4998
rect 7445 4862 7477 4968
rect 7681 4862 7713 4968
rect 7917 4862 7949 4968
rect 8153 4862 8185 4968
rect 8388 4862 8422 4968
rect 7438 4850 7484 4862
rect 7438 4674 7444 4850
rect 7478 4674 7484 4850
rect 7438 4662 7484 4674
rect 7556 4850 7602 4862
rect 7556 4674 7562 4850
rect 7596 4674 7602 4850
rect 7556 4662 7602 4674
rect 7674 4850 7720 4862
rect 7674 4674 7680 4850
rect 7714 4674 7720 4850
rect 7674 4662 7720 4674
rect 7792 4850 7838 4862
rect 7792 4674 7798 4850
rect 7832 4674 7838 4850
rect 7792 4662 7838 4674
rect 7910 4850 7956 4862
rect 7910 4674 7916 4850
rect 7950 4674 7956 4850
rect 7910 4662 7956 4674
rect 8028 4850 8074 4862
rect 8028 4674 8034 4850
rect 8068 4674 8074 4850
rect 8028 4662 8074 4674
rect 8146 4850 8192 4862
rect 8146 4674 8152 4850
rect 8186 4674 8192 4850
rect 8146 4662 8192 4674
rect 8264 4850 8310 4862
rect 8264 4674 8270 4850
rect 8304 4674 8310 4850
rect 8264 4662 8310 4674
rect 8382 4850 8428 4862
rect 8382 4674 8388 4850
rect 8422 4674 8428 4850
rect 8382 4662 8428 4674
rect 8500 4850 8546 4862
rect 8500 4674 8506 4850
rect 8540 4674 8546 4850
rect 8500 4662 8546 4674
rect 5100 4541 5146 4553
rect 7561 4568 7597 4662
rect 7797 4568 7833 4662
rect 8033 4569 8069 4662
rect 8195 4614 8261 4621
rect 8195 4580 8211 4614
rect 8245 4580 8261 4614
rect 8195 4569 8261 4580
rect 8033 4568 8261 4569
rect 4398 4499 4432 4541
rect 4634 4499 4668 4541
rect 4398 4471 4668 4499
rect 4752 4500 4786 4541
rect 4988 4500 5022 4541
rect 4752 4471 5022 4500
rect 4398 4423 4432 4471
rect 4398 4393 4461 4423
rect 4426 4301 4461 4393
rect 4933 4363 5033 4384
rect 4933 4309 4947 4363
rect 5012 4309 5033 4363
rect 4933 4304 5033 4309
rect 5106 4358 5140 4541
rect 7561 4539 8261 4568
rect 7561 4538 8143 4539
rect 7681 4425 7715 4538
rect 8077 4497 8143 4538
rect 8077 4463 8093 4497
rect 8127 4463 8143 4497
rect 8077 4456 8143 4463
rect 8505 4457 8540 4662
rect 8712 4457 8779 5047
rect 10471 5024 10512 5056
rect 10758 5052 10768 5118
rect 10824 5052 10834 5118
rect 11504 5094 11514 5202
rect 11646 5139 11656 5202
rect 14375 5143 14595 5163
rect 11646 5128 11658 5139
rect 11646 5094 11659 5128
rect 11514 5056 11659 5094
rect 11618 5028 11659 5056
rect 9887 4996 10157 5024
rect 9628 4930 9638 4996
rect 9704 4930 9714 4996
rect 9887 4934 9921 4996
rect 10123 4934 10157 4996
rect 10241 4996 10512 5024
rect 11029 5000 11299 5028
rect 10241 4934 10275 4996
rect 10477 4934 10512 4996
rect 10653 4984 10824 5000
rect 10653 4950 10784 4984
rect 10818 4950 10824 4984
rect 10653 4934 10824 4950
rect 11029 4938 11063 5000
rect 11265 4938 11299 5000
rect 11383 5000 11659 5028
rect 11383 4938 11417 5000
rect 11619 4938 11659 5000
rect 14375 5035 14419 5143
rect 14551 5035 14595 5143
rect 16172 5101 16228 5109
rect 14375 4993 14595 5035
rect 15246 5093 16228 5101
rect 15246 5059 16188 5093
rect 16222 5059 16228 5093
rect 16891 5089 16901 5197
rect 17033 5134 17043 5197
rect 17033 5123 17045 5134
rect 17033 5089 17046 5123
rect 17302 5113 17358 5115
rect 15246 5043 16228 5059
rect 16901 5051 17046 5089
rect 15246 5042 16225 5043
rect 9763 4922 9809 4934
rect 9763 4546 9769 4922
rect 9803 4546 9809 4922
rect 9763 4534 9809 4546
rect 9881 4922 9927 4934
rect 9881 4546 9887 4922
rect 9921 4546 9927 4922
rect 9881 4534 9927 4546
rect 9999 4922 10045 4934
rect 9999 4546 10005 4922
rect 10039 4546 10045 4922
rect 9999 4534 10045 4546
rect 10117 4922 10163 4934
rect 10117 4546 10123 4922
rect 10157 4546 10163 4922
rect 10117 4534 10163 4546
rect 10235 4922 10281 4934
rect 10235 4546 10241 4922
rect 10275 4546 10281 4922
rect 10235 4534 10281 4546
rect 10353 4922 10399 4934
rect 10353 4546 10359 4922
rect 10393 4546 10399 4922
rect 10353 4534 10399 4546
rect 10471 4922 10517 4934
rect 10471 4546 10477 4922
rect 10511 4546 10517 4922
rect 10471 4534 10517 4546
rect 8505 4429 8779 4457
rect 8151 4425 8779 4429
rect 7675 4413 7721 4425
rect 6108 4372 6215 4374
rect 5106 4304 5215 4358
rect 4426 4265 4653 4301
rect 4426 4158 4461 4265
rect 4587 4231 4653 4265
rect 4587 4197 4603 4231
rect 4637 4197 4653 4231
rect 4934 4289 5031 4304
rect 4934 4222 4991 4289
rect 4587 4191 4653 4197
rect 4828 4186 5097 4222
rect 4828 4158 4861 4186
rect 5064 4158 5097 4186
rect 5181 4158 5215 4304
rect 6032 4297 6042 4372
rect 6110 4297 6215 4372
rect 6059 4296 6215 4297
rect 4302 4146 4348 4158
rect 4302 3970 4308 4146
rect 4342 3970 4348 4146
rect 4302 3958 4348 3970
rect 4420 4146 4466 4158
rect 4420 3970 4426 4146
rect 4460 3970 4466 4146
rect 4420 3958 4466 3970
rect 4538 4146 4584 4158
rect 4538 3970 4544 4146
rect 4578 3970 4584 4146
rect 4538 3958 4584 3970
rect 4656 4146 4702 4158
rect 4656 3970 4662 4146
rect 4696 4091 4702 4146
rect 4821 4146 4867 4158
rect 4821 4091 4827 4146
rect 4696 4003 4827 4091
rect 4696 3970 4702 4003
rect 4656 3958 4702 3970
rect 4821 3970 4827 4003
rect 4861 3970 4867 4146
rect 4821 3958 4867 3970
rect 4939 4146 4985 4158
rect 4939 3970 4945 4146
rect 4979 3970 4985 4146
rect 4939 3958 4985 3970
rect 5057 4146 5103 4158
rect 5057 3970 5063 4146
rect 5097 3970 5103 4146
rect 5057 3958 5103 3970
rect 5175 4146 5221 4158
rect 5175 3970 5181 4146
rect 5215 3970 5221 4146
rect 5175 3958 5221 3970
rect 4308 3919 4342 3958
rect 4544 3919 4578 3958
rect 4308 3883 4578 3919
rect 4945 3920 4978 3958
rect 5181 3920 5214 3958
rect 4945 3884 5214 3920
rect 4308 3882 4474 3883
rect 4342 3803 4474 3882
rect 4332 3695 4342 3803
rect 4474 3695 4484 3803
rect 946 3321 1923 3351
rect 4140 3349 4203 3366
rect 4065 3345 4203 3349
rect 946 3215 978 3321
rect 1182 3215 1214 3321
rect 1418 3215 1450 3321
rect 1654 3215 1686 3321
rect 1889 3215 1923 3321
rect 2233 3311 4203 3345
rect 2231 3282 4203 3311
rect 2231 3266 2277 3282
rect 4065 3280 4203 3282
rect 939 3203 985 3215
rect 939 3027 945 3203
rect 979 3027 985 3203
rect 939 3015 985 3027
rect 1057 3203 1103 3215
rect 1057 3027 1063 3203
rect 1097 3027 1103 3203
rect 1057 3015 1103 3027
rect 1175 3203 1221 3215
rect 1175 3027 1181 3203
rect 1215 3027 1221 3203
rect 1175 3015 1221 3027
rect 1293 3203 1339 3215
rect 1293 3027 1299 3203
rect 1333 3027 1339 3203
rect 1293 3015 1339 3027
rect 1411 3203 1457 3215
rect 1411 3027 1417 3203
rect 1451 3027 1457 3203
rect 1411 3015 1457 3027
rect 1529 3203 1575 3215
rect 1529 3027 1535 3203
rect 1569 3027 1575 3203
rect 1529 3015 1575 3027
rect 1647 3203 1693 3215
rect 1647 3027 1653 3203
rect 1687 3027 1693 3203
rect 1647 3015 1693 3027
rect 1765 3203 1811 3215
rect 1765 3027 1771 3203
rect 1805 3027 1811 3203
rect 1765 3015 1811 3027
rect 1883 3203 1929 3215
rect 1883 3027 1889 3203
rect 1923 3027 1929 3203
rect 1883 3015 1929 3027
rect 2001 3203 2047 3215
rect 2001 3027 2007 3203
rect 2041 3027 2047 3203
rect 2001 3015 2047 3027
rect 1062 2921 1098 3015
rect 1298 2921 1334 3015
rect 1534 2922 1570 3015
rect 1696 2967 1762 2974
rect 1696 2933 1712 2967
rect 1746 2933 1762 2967
rect 1696 2922 1762 2933
rect 1534 2921 1762 2922
rect 1062 2892 1762 2921
rect 1062 2891 1644 2892
rect 1182 2778 1216 2891
rect 1578 2850 1644 2891
rect 1578 2816 1594 2850
rect 1628 2816 1644 2850
rect 1578 2809 1644 2816
rect 2006 2797 2041 3015
rect 2230 2814 2277 3266
rect 3189 3050 3199 3158
rect 3331 3050 3341 3158
rect 5087 3050 5097 3158
rect 5229 3050 5239 3158
rect 3199 3010 3331 3050
rect 5097 3010 5229 3050
rect 3198 2944 3331 3010
rect 5096 2944 5229 3010
rect 2527 2901 4000 2944
rect 2230 2798 2276 2814
rect 2195 2797 2276 2798
rect 2006 2782 2276 2797
rect 1652 2778 2276 2782
rect 1176 2766 1222 2778
rect 911 2288 921 2406
rect 1039 2374 1049 2406
rect 1176 2390 1182 2766
rect 1216 2390 1222 2766
rect 1176 2378 1222 2390
rect 1294 2766 1340 2778
rect 1294 2390 1300 2766
rect 1334 2390 1340 2766
rect 1294 2378 1340 2390
rect 1412 2766 1458 2778
rect 1412 2390 1418 2766
rect 1452 2414 1458 2766
rect 1529 2766 1575 2778
rect 1529 2590 1535 2766
rect 1569 2590 1575 2766
rect 1529 2578 1575 2590
rect 1647 2766 2276 2778
rect 1647 2590 1653 2766
rect 1687 2754 2276 2766
rect 1687 2753 1929 2754
rect 1687 2590 1693 2753
rect 2195 2752 2276 2754
rect 2527 2598 2561 2901
rect 2893 2798 2927 2901
rect 3129 2798 3163 2901
rect 3365 2798 3399 2901
rect 3601 2798 3635 2901
rect 2887 2786 2933 2798
rect 1647 2578 1693 2590
rect 2403 2586 2449 2598
rect 1535 2462 1570 2578
rect 1666 2462 1774 2472
rect 1535 2414 1666 2462
rect 1452 2390 1666 2414
rect 1412 2378 1666 2390
rect 1418 2374 1666 2378
rect 1039 2346 1054 2374
rect 1039 2340 1291 2346
rect 1039 2306 1241 2340
rect 1275 2306 1291 2340
rect 1039 2290 1291 2306
rect 1343 2340 1409 2346
rect 1343 2306 1359 2340
rect 1393 2306 1409 2340
rect 1592 2330 1666 2374
rect 2403 2410 2409 2586
rect 2443 2410 2449 2586
rect 2403 2398 2449 2410
rect 2521 2586 2567 2598
rect 2521 2410 2527 2586
rect 2561 2410 2567 2586
rect 2521 2398 2567 2410
rect 2639 2586 2685 2598
rect 2639 2410 2645 2586
rect 2679 2410 2685 2586
rect 2639 2398 2685 2410
rect 2757 2586 2803 2598
rect 2887 2586 2893 2786
rect 2757 2410 2763 2586
rect 2797 2410 2893 2586
rect 2927 2410 2933 2786
rect 2757 2398 2803 2410
rect 2887 2398 2933 2410
rect 3005 2786 3051 2798
rect 3005 2410 3011 2786
rect 3045 2410 3051 2786
rect 3005 2398 3051 2410
rect 3123 2786 3169 2798
rect 3123 2410 3129 2786
rect 3163 2410 3169 2786
rect 3123 2398 3169 2410
rect 3241 2786 3287 2798
rect 3241 2410 3247 2786
rect 3281 2410 3287 2786
rect 3241 2398 3287 2410
rect 3359 2786 3405 2798
rect 3359 2410 3365 2786
rect 3399 2410 3405 2786
rect 3359 2398 3405 2410
rect 3477 2786 3523 2798
rect 3477 2410 3483 2786
rect 3517 2410 3523 2786
rect 3477 2398 3523 2410
rect 3595 2786 3641 2798
rect 3595 2410 3601 2786
rect 3635 2586 3641 2786
rect 3966 2598 4000 2901
rect 4425 2901 5898 2944
rect 4425 2598 4459 2901
rect 4791 2798 4825 2901
rect 5027 2798 5061 2901
rect 5263 2798 5297 2901
rect 5499 2798 5533 2901
rect 4785 2786 4831 2798
rect 3724 2586 3770 2598
rect 3635 2410 3730 2586
rect 3764 2410 3770 2586
rect 3595 2398 3641 2410
rect 3724 2398 3770 2410
rect 3842 2586 3888 2598
rect 3842 2410 3848 2586
rect 3882 2410 3888 2586
rect 3842 2398 3888 2410
rect 3960 2586 4006 2598
rect 3960 2410 3966 2586
rect 4000 2410 4006 2586
rect 3960 2398 4006 2410
rect 4078 2586 4124 2598
rect 4078 2410 4084 2586
rect 4118 2410 4124 2586
rect 4078 2398 4124 2410
rect 4301 2586 4347 2598
rect 4301 2410 4307 2586
rect 4341 2410 4347 2586
rect 4301 2398 4347 2410
rect 4419 2586 4465 2598
rect 4419 2410 4425 2586
rect 4459 2410 4465 2586
rect 4419 2398 4465 2410
rect 4537 2586 4583 2598
rect 4537 2410 4543 2586
rect 4577 2410 4583 2586
rect 4537 2398 4583 2410
rect 4655 2586 4701 2598
rect 4785 2586 4791 2786
rect 4655 2410 4661 2586
rect 4695 2410 4791 2586
rect 4825 2410 4831 2786
rect 4655 2398 4701 2410
rect 4785 2398 4831 2410
rect 4903 2786 4949 2798
rect 4903 2410 4909 2786
rect 4943 2410 4949 2786
rect 4903 2398 4949 2410
rect 5021 2786 5067 2798
rect 5021 2410 5027 2786
rect 5061 2410 5067 2786
rect 5021 2398 5067 2410
rect 5139 2786 5185 2798
rect 5139 2410 5145 2786
rect 5179 2410 5185 2786
rect 5139 2398 5185 2410
rect 5257 2786 5303 2798
rect 5257 2410 5263 2786
rect 5297 2410 5303 2786
rect 5257 2398 5303 2410
rect 5375 2786 5421 2798
rect 5375 2410 5381 2786
rect 5415 2410 5421 2786
rect 5375 2398 5421 2410
rect 5493 2786 5539 2798
rect 5493 2410 5499 2786
rect 5533 2586 5539 2786
rect 5864 2598 5898 2901
rect 5622 2586 5668 2598
rect 5533 2410 5628 2586
rect 5662 2410 5668 2586
rect 5493 2398 5539 2410
rect 5622 2398 5668 2410
rect 5740 2586 5786 2598
rect 5740 2410 5746 2586
rect 5780 2410 5786 2586
rect 5740 2398 5786 2410
rect 5858 2586 5904 2598
rect 5858 2410 5864 2586
rect 5898 2410 5904 2586
rect 5858 2398 5904 2410
rect 5976 2586 6022 2598
rect 5976 2410 5982 2586
rect 6016 2410 6022 2586
rect 6108 2552 6215 4296
rect 6503 4020 6792 4195
rect 7675 4037 7681 4413
rect 7715 4037 7721 4413
rect 7675 4025 7721 4037
rect 7793 4413 7839 4425
rect 7793 4037 7799 4413
rect 7833 4037 7839 4413
rect 7793 4025 7839 4037
rect 7911 4413 7957 4425
rect 7911 4037 7917 4413
rect 7951 4061 7957 4413
rect 8028 4413 8074 4425
rect 8028 4237 8034 4413
rect 8068 4237 8074 4413
rect 8028 4225 8074 4237
rect 8146 4413 8779 4425
rect 8146 4237 8152 4413
rect 8186 4400 8779 4413
rect 9769 4492 9803 4534
rect 10005 4492 10039 4534
rect 9769 4464 10039 4492
rect 10123 4493 10157 4534
rect 10359 4493 10393 4534
rect 10123 4464 10393 4493
rect 9769 4416 9803 4464
rect 8186 4237 8192 4400
rect 9769 4386 9832 4416
rect 8146 4225 8192 4237
rect 9797 4294 9832 4386
rect 9797 4258 10024 4294
rect 10294 4283 10304 4380
rect 10403 4283 10413 4380
rect 10477 4351 10511 4534
rect 10477 4297 10586 4351
rect 8034 4109 8069 4225
rect 9797 4151 9832 4258
rect 9958 4224 10024 4258
rect 9958 4190 9974 4224
rect 10008 4190 10024 4224
rect 10305 4282 10402 4283
rect 10305 4215 10362 4282
rect 9958 4184 10024 4190
rect 10199 4179 10468 4215
rect 10199 4151 10232 4179
rect 10435 4151 10468 4179
rect 10552 4151 10586 4297
rect 9673 4139 9719 4151
rect 8165 4109 8273 4119
rect 8034 4061 8165 4109
rect 7951 4037 8165 4061
rect 7911 4025 8165 4037
rect 7917 4021 8165 4025
rect 6503 3993 7553 4020
rect 6503 3987 7790 3993
rect 6503 3953 7740 3987
rect 7774 3953 7790 3987
rect 6503 3937 7790 3953
rect 7842 3987 7908 3993
rect 7842 3953 7858 3987
rect 7892 3953 7908 3987
rect 8091 3977 8165 4021
rect 8165 3967 8273 3977
rect 6503 3921 7553 3937
rect 6503 3920 7490 3921
rect 6503 3916 7025 3920
rect 6503 3915 6792 3916
rect 6520 3505 6809 3667
rect 6520 3399 6657 3505
rect 6769 3492 6809 3505
rect 6769 3399 6811 3492
rect 6520 3388 6811 3399
rect 6520 3387 6809 3388
rect 6520 2552 6808 2555
rect 6108 2436 6808 2552
rect 6108 2433 6215 2436
rect 5976 2398 6022 2410
rect 1666 2320 1774 2330
rect 2409 2364 2443 2398
rect 3011 2364 3045 2398
rect 3247 2364 3281 2398
rect 2409 2329 2568 2364
rect 3011 2329 3281 2364
rect 3848 2364 3882 2398
rect 4084 2364 4118 2398
rect 3848 2329 4118 2364
rect 4307 2364 4341 2398
rect 4909 2364 4943 2398
rect 5145 2364 5179 2398
rect 4307 2329 4466 2364
rect 4909 2329 5179 2364
rect 5746 2364 5780 2398
rect 5982 2364 6016 2398
rect 5746 2329 6016 2364
rect 6520 2393 6808 2436
rect 1039 2288 1054 2290
rect 954 2274 1054 2288
rect 954 2231 1054 2232
rect 575 2210 1054 2231
rect 1343 2210 1409 2306
rect 575 2162 1409 2210
rect 575 2133 1054 2162
rect 575 2131 680 2133
rect 954 2132 1054 2133
rect 408 1946 418 2025
rect 511 1946 521 2025
rect 419 772 512 1946
rect 1337 1897 1557 1917
rect 1337 1789 1381 1897
rect 1513 1789 1557 1897
rect 1337 1747 1557 1789
rect 941 1717 1918 1747
rect 941 1611 973 1717
rect 1177 1611 1209 1717
rect 1413 1611 1445 1717
rect 1649 1611 1681 1717
rect 1884 1611 1918 1717
rect 934 1599 980 1611
rect 934 1423 940 1599
rect 974 1423 980 1599
rect 934 1411 980 1423
rect 1052 1599 1098 1611
rect 1052 1423 1058 1599
rect 1092 1423 1098 1599
rect 1052 1411 1098 1423
rect 1170 1599 1216 1611
rect 1170 1423 1176 1599
rect 1210 1423 1216 1599
rect 1170 1411 1216 1423
rect 1288 1599 1334 1611
rect 1288 1423 1294 1599
rect 1328 1423 1334 1599
rect 1288 1411 1334 1423
rect 1406 1599 1452 1611
rect 1406 1423 1412 1599
rect 1446 1423 1452 1599
rect 1406 1411 1452 1423
rect 1524 1599 1570 1611
rect 1524 1423 1530 1599
rect 1564 1423 1570 1599
rect 1524 1411 1570 1423
rect 1642 1599 1688 1611
rect 1642 1423 1648 1599
rect 1682 1423 1688 1599
rect 1642 1411 1688 1423
rect 1760 1599 1806 1611
rect 1760 1423 1766 1599
rect 1800 1423 1806 1599
rect 1760 1411 1806 1423
rect 1878 1599 1924 1611
rect 1878 1423 1884 1599
rect 1918 1423 1924 1599
rect 1878 1411 1924 1423
rect 1996 1599 2042 1611
rect 1996 1423 2002 1599
rect 2036 1423 2042 1599
rect 1996 1411 2042 1423
rect 2534 1545 2568 2329
rect 3247 2267 3281 2329
rect 2836 2229 3578 2267
rect 2836 2105 2870 2229
rect 3072 2105 3106 2229
rect 3308 2105 3342 2229
rect 3544 2105 3578 2229
rect 3834 2122 3844 2188
rect 3907 2122 3917 2188
rect 2830 2093 2876 2105
rect 2830 1717 2836 2093
rect 2870 1717 2876 2093
rect 2830 1705 2876 1717
rect 2948 2093 2994 2105
rect 2948 1717 2954 2093
rect 2988 1717 2994 2093
rect 2948 1705 2994 1717
rect 3066 2093 3112 2105
rect 3066 1717 3072 2093
rect 3106 1717 3112 2093
rect 3066 1705 3112 1717
rect 3184 2093 3230 2105
rect 3184 1717 3190 2093
rect 3224 1717 3230 2093
rect 3184 1705 3230 1717
rect 3302 2093 3348 2105
rect 3302 1717 3308 2093
rect 3342 1717 3348 2093
rect 3302 1705 3348 1717
rect 3420 2093 3466 2105
rect 3420 1717 3426 2093
rect 3460 1717 3466 2093
rect 3420 1705 3466 1717
rect 3538 2093 3584 2105
rect 3538 1717 3544 2093
rect 3578 1717 3584 2093
rect 3538 1705 3584 1717
rect 3950 1546 3984 2329
rect 3677 1545 3984 1546
rect 2534 1540 2850 1545
rect 3564 1540 3984 1545
rect 2534 1529 2917 1540
rect 2534 1502 2866 1529
rect 1057 1317 1093 1411
rect 1293 1317 1329 1411
rect 1529 1318 1565 1411
rect 1691 1363 1757 1370
rect 1691 1329 1707 1363
rect 1741 1329 1757 1363
rect 1691 1318 1757 1329
rect 1529 1317 1757 1318
rect 1057 1288 1757 1317
rect 1057 1287 1639 1288
rect 1177 1174 1211 1287
rect 1573 1246 1639 1287
rect 1573 1212 1589 1246
rect 1623 1212 1639 1246
rect 1573 1205 1639 1212
rect 2001 1178 2036 1411
rect 2534 1373 2568 1502
rect 2850 1495 2866 1502
rect 2900 1495 2917 1529
rect 2850 1489 2917 1495
rect 3497 1529 3984 1540
rect 3497 1495 3514 1529
rect 3548 1502 3984 1529
rect 3548 1495 3564 1502
rect 3677 1501 3984 1502
rect 3497 1489 3564 1495
rect 2675 1462 2731 1474
rect 2675 1428 2681 1462
rect 2715 1461 2731 1462
rect 3788 1461 3844 1473
rect 2715 1445 3182 1461
rect 2715 1428 3132 1445
rect 2675 1412 3132 1428
rect 3116 1411 3132 1412
rect 3166 1411 3182 1445
rect 3116 1404 3182 1411
rect 3234 1446 3804 1461
rect 3234 1412 3250 1446
rect 3284 1427 3804 1446
rect 3838 1427 3844 1461
rect 3284 1412 3844 1427
rect 3234 1402 3301 1412
rect 3788 1411 3844 1412
rect 3950 1373 3984 1501
rect 4432 1545 4466 2329
rect 5145 2267 5179 2329
rect 4734 2229 5476 2267
rect 4734 2105 4768 2229
rect 4970 2105 5004 2229
rect 5206 2105 5240 2229
rect 5442 2105 5476 2229
rect 4728 2093 4774 2105
rect 4728 1717 4734 2093
rect 4768 1717 4774 2093
rect 4728 1705 4774 1717
rect 4846 2093 4892 2105
rect 4846 1717 4852 2093
rect 4886 1717 4892 2093
rect 4846 1705 4892 1717
rect 4964 2093 5010 2105
rect 4964 1717 4970 2093
rect 5004 1717 5010 2093
rect 4964 1705 5010 1717
rect 5082 2093 5128 2105
rect 5082 1717 5088 2093
rect 5122 1717 5128 2093
rect 5082 1705 5128 1717
rect 5200 2093 5246 2105
rect 5200 1717 5206 2093
rect 5240 1717 5246 2093
rect 5200 1705 5246 1717
rect 5318 2093 5364 2105
rect 5318 1717 5324 2093
rect 5358 1717 5364 2093
rect 5318 1705 5364 1717
rect 5436 2093 5482 2105
rect 5436 1717 5442 2093
rect 5476 1717 5482 2093
rect 5436 1705 5482 1717
rect 5848 1546 5882 2329
rect 6520 2287 6656 2393
rect 6768 2391 6808 2393
rect 6774 2380 6808 2391
rect 6520 2285 6662 2287
rect 6774 2285 6809 2380
rect 6520 2276 6809 2285
rect 6520 2275 6808 2276
rect 6520 2274 6776 2275
rect 5460 1545 5529 1546
rect 5575 1545 5882 1546
rect 4432 1540 4748 1545
rect 5460 1541 5882 1545
rect 4432 1529 4815 1540
rect 4432 1502 4764 1529
rect 4432 1373 4466 1502
rect 4748 1495 4764 1502
rect 4798 1495 4815 1529
rect 4748 1489 4815 1495
rect 5393 1530 5882 1541
rect 5393 1496 5410 1530
rect 5444 1502 5882 1530
rect 5444 1496 5460 1502
rect 5575 1501 5882 1502
rect 5393 1490 5460 1496
rect 4573 1462 4629 1474
rect 4573 1428 4579 1462
rect 4613 1461 4629 1462
rect 5686 1461 5742 1473
rect 4613 1445 5080 1461
rect 4613 1428 5030 1445
rect 4573 1412 5030 1428
rect 5014 1411 5030 1412
rect 5064 1411 5080 1445
rect 5014 1404 5080 1411
rect 5132 1446 5702 1461
rect 5132 1412 5148 1446
rect 5182 1427 5702 1446
rect 5736 1427 5742 1461
rect 5182 1412 5742 1427
rect 5132 1402 5199 1412
rect 5686 1411 5742 1412
rect 5848 1373 5882 1501
rect 5963 2151 6030 2175
rect 5963 2117 5980 2151
rect 6014 2117 6030 2151
rect 1647 1174 2036 1178
rect 1171 1162 1217 1174
rect 1171 786 1177 1162
rect 1211 786 1217 1162
rect 1171 774 1217 786
rect 1289 1162 1335 1174
rect 1289 786 1295 1162
rect 1329 786 1335 1162
rect 1289 774 1335 786
rect 1407 1162 1453 1174
rect 1407 786 1413 1162
rect 1447 810 1453 1162
rect 1524 1162 1570 1174
rect 1524 986 1530 1162
rect 1564 986 1570 1162
rect 1524 974 1570 986
rect 1642 1162 2036 1174
rect 2528 1361 2574 1373
rect 2528 1185 2534 1361
rect 2568 1185 2574 1361
rect 2528 1173 2574 1185
rect 2646 1361 2692 1373
rect 2646 1185 2652 1361
rect 2686 1185 2692 1361
rect 2646 1173 2692 1185
rect 2948 1361 2994 1373
rect 1642 986 1648 1162
rect 1682 1149 2036 1162
rect 1682 986 1688 1149
rect 1958 1146 2036 1149
rect 1958 1094 1968 1146
rect 2031 1094 2041 1146
rect 1963 1088 2036 1094
rect 1642 974 1688 986
rect 1530 858 1565 974
rect 2651 879 2685 1173
rect 2948 985 2954 1361
rect 2988 985 2994 1361
rect 2948 973 2994 985
rect 3066 1361 3112 1373
rect 3066 985 3072 1361
rect 3106 985 3112 1361
rect 3066 973 3112 985
rect 3184 1361 3230 1373
rect 3184 985 3190 1361
rect 3224 985 3230 1361
rect 3184 973 3230 985
rect 3302 1361 3348 1373
rect 3302 985 3308 1361
rect 3342 985 3348 1361
rect 3302 973 3348 985
rect 3420 1361 3466 1373
rect 3420 985 3426 1361
rect 3460 985 3466 1361
rect 3826 1361 3872 1373
rect 3826 1185 3832 1361
rect 3866 1185 3872 1361
rect 3826 1173 3872 1185
rect 3944 1361 3990 1373
rect 3944 1185 3950 1361
rect 3984 1185 3990 1361
rect 3944 1173 3990 1185
rect 4426 1361 4472 1373
rect 4426 1185 4432 1361
rect 4466 1185 4472 1361
rect 4426 1173 4472 1185
rect 4544 1361 4590 1373
rect 4544 1185 4550 1361
rect 4584 1185 4590 1361
rect 4544 1173 4590 1185
rect 4846 1361 4892 1373
rect 3420 973 3466 985
rect 3308 879 3342 973
rect 3832 879 3865 1173
rect 1661 858 1769 868
rect 1530 810 1661 858
rect 1447 786 1661 810
rect 1407 774 1661 786
rect 419 770 1004 772
rect 1413 770 1661 774
rect 419 742 1049 770
rect 419 736 1286 742
rect 419 702 1236 736
rect 1270 702 1286 736
rect 419 686 1286 702
rect 1338 736 1404 742
rect 1338 702 1354 736
rect 1388 702 1404 736
rect 1587 726 1661 770
rect 2651 847 3865 879
rect 4549 879 4583 1173
rect 4846 985 4852 1361
rect 4886 985 4892 1361
rect 4846 973 4892 985
rect 4964 1361 5010 1373
rect 4964 985 4970 1361
rect 5004 985 5010 1361
rect 4964 973 5010 985
rect 5082 1361 5128 1373
rect 5082 985 5088 1361
rect 5122 985 5128 1361
rect 5082 973 5128 985
rect 5200 1361 5246 1373
rect 5200 985 5206 1361
rect 5240 985 5246 1361
rect 5200 973 5246 985
rect 5318 1361 5364 1373
rect 5318 985 5324 1361
rect 5358 985 5364 1361
rect 5724 1361 5770 1373
rect 5724 1185 5730 1361
rect 5764 1185 5770 1361
rect 5724 1173 5770 1185
rect 5842 1361 5888 1373
rect 5842 1185 5848 1361
rect 5882 1185 5888 1361
rect 5842 1173 5888 1185
rect 5318 973 5364 985
rect 5206 879 5240 973
rect 5730 879 5763 1173
rect 4549 847 5763 879
rect 3144 762 3276 847
rect 5042 762 5174 847
rect 1661 716 1769 726
rect 419 670 1049 686
rect 419 666 1004 670
rect 419 665 520 666
rect 949 617 1049 628
rect 913 511 923 617
rect 1035 606 1049 617
rect 1338 606 1404 702
rect 3134 654 3144 762
rect 3276 654 3286 762
rect 5032 654 5042 762
rect 5174 654 5184 762
rect 5963 734 6030 2117
rect 6932 2022 7025 3916
rect 7088 3857 7554 3879
rect 7842 3857 7908 3953
rect 9673 3963 9679 4139
rect 9713 3963 9719 4139
rect 9673 3951 9719 3963
rect 9791 4139 9837 4151
rect 9791 3963 9797 4139
rect 9831 3963 9837 4139
rect 9791 3951 9837 3963
rect 9909 4139 9955 4151
rect 9909 3963 9915 4139
rect 9949 3963 9955 4139
rect 9909 3951 9955 3963
rect 10027 4139 10073 4151
rect 10027 3963 10033 4139
rect 10067 4084 10073 4139
rect 10192 4139 10238 4151
rect 10192 4084 10198 4139
rect 10067 3996 10198 4084
rect 10067 3963 10073 3996
rect 10027 3951 10073 3963
rect 10192 3963 10198 3996
rect 10232 3963 10238 4139
rect 10192 3951 10238 3963
rect 10310 4139 10356 4151
rect 10310 3963 10316 4139
rect 10350 3963 10356 4139
rect 10310 3951 10356 3963
rect 10428 4139 10474 4151
rect 10428 3963 10434 4139
rect 10468 3963 10474 4139
rect 10428 3951 10474 3963
rect 10546 4139 10592 4151
rect 10546 3963 10552 4139
rect 10586 3963 10592 4139
rect 10546 3951 10592 3963
rect 9679 3912 9713 3951
rect 9915 3912 9949 3951
rect 9679 3877 9949 3912
rect 10316 3913 10349 3951
rect 10552 3913 10585 3951
rect 10316 3877 10585 3913
rect 7088 3809 7908 3857
rect 9713 3876 9949 3877
rect 7088 3778 7554 3809
rect 9713 3802 9845 3876
rect 7088 3522 7193 3778
rect 9703 3694 9713 3802
rect 9845 3694 9855 3802
rect 7088 3416 7151 3522
rect 7263 3416 7273 3522
rect 7855 3498 8075 3518
rect 7088 3405 7237 3416
rect 7088 2228 7193 3405
rect 7855 3390 7899 3498
rect 8031 3390 8075 3498
rect 7855 3348 8075 3390
rect 10653 3363 10715 4934
rect 10905 4926 10951 4938
rect 10905 4550 10911 4926
rect 10945 4550 10951 4926
rect 10905 4538 10951 4550
rect 11023 4926 11069 4938
rect 11023 4550 11029 4926
rect 11063 4550 11069 4926
rect 11023 4538 11069 4550
rect 11141 4926 11187 4938
rect 11141 4550 11147 4926
rect 11181 4550 11187 4926
rect 11141 4538 11187 4550
rect 11259 4926 11305 4938
rect 11259 4550 11265 4926
rect 11299 4550 11305 4926
rect 11259 4538 11305 4550
rect 11377 4926 11423 4938
rect 11377 4550 11383 4926
rect 11417 4550 11423 4926
rect 11377 4538 11423 4550
rect 11495 4926 11541 4938
rect 11495 4550 11501 4926
rect 11535 4550 11541 4926
rect 11495 4538 11541 4550
rect 11613 4926 11659 4938
rect 11613 4550 11619 4926
rect 11653 4550 11659 4926
rect 13979 4963 14956 4993
rect 13979 4857 14011 4963
rect 14215 4857 14247 4963
rect 14451 4857 14483 4963
rect 14687 4857 14719 4963
rect 14922 4857 14956 4963
rect 13972 4845 14018 4857
rect 13972 4669 13978 4845
rect 14012 4669 14018 4845
rect 13972 4657 14018 4669
rect 14090 4845 14136 4857
rect 14090 4669 14096 4845
rect 14130 4669 14136 4845
rect 14090 4657 14136 4669
rect 14208 4845 14254 4857
rect 14208 4669 14214 4845
rect 14248 4669 14254 4845
rect 14208 4657 14254 4669
rect 14326 4845 14372 4857
rect 14326 4669 14332 4845
rect 14366 4669 14372 4845
rect 14326 4657 14372 4669
rect 14444 4845 14490 4857
rect 14444 4669 14450 4845
rect 14484 4669 14490 4845
rect 14444 4657 14490 4669
rect 14562 4845 14608 4857
rect 14562 4669 14568 4845
rect 14602 4669 14608 4845
rect 14562 4657 14608 4669
rect 14680 4845 14726 4857
rect 14680 4669 14686 4845
rect 14720 4669 14726 4845
rect 14680 4657 14726 4669
rect 14798 4845 14844 4857
rect 14798 4669 14804 4845
rect 14838 4669 14844 4845
rect 14798 4657 14844 4669
rect 14916 4845 14962 4857
rect 14916 4669 14922 4845
rect 14956 4669 14962 4845
rect 14916 4657 14962 4669
rect 15034 4845 15080 4857
rect 15034 4669 15040 4845
rect 15074 4669 15080 4845
rect 15034 4657 15080 4669
rect 11613 4538 11659 4550
rect 14095 4563 14131 4657
rect 14331 4563 14367 4657
rect 14567 4564 14603 4657
rect 14729 4609 14795 4616
rect 14729 4575 14745 4609
rect 14779 4575 14795 4609
rect 14729 4564 14795 4575
rect 14567 4563 14795 4564
rect 10911 4496 10945 4538
rect 11147 4496 11181 4538
rect 10911 4468 11181 4496
rect 11265 4497 11299 4538
rect 11501 4497 11535 4538
rect 11265 4468 11535 4497
rect 10911 4420 10945 4468
rect 10911 4390 10974 4420
rect 10939 4298 10974 4390
rect 11446 4360 11546 4381
rect 11446 4306 11460 4360
rect 11525 4306 11546 4360
rect 11446 4301 11546 4306
rect 11619 4355 11653 4538
rect 14095 4534 14795 4563
rect 14095 4533 14677 4534
rect 14215 4420 14249 4533
rect 14611 4492 14677 4533
rect 14611 4458 14627 4492
rect 14661 4458 14677 4492
rect 14611 4451 14677 4458
rect 15039 4452 15074 4657
rect 15246 4452 15313 5042
rect 17005 5019 17046 5051
rect 17292 5047 17302 5113
rect 17358 5047 17368 5113
rect 18038 5089 18048 5197
rect 18180 5134 18190 5197
rect 20933 5147 21153 5167
rect 18180 5123 18192 5134
rect 18180 5089 18193 5123
rect 18048 5051 18193 5089
rect 18152 5023 18193 5051
rect 16421 4991 16691 5019
rect 16162 4925 16172 4991
rect 16238 4925 16248 4991
rect 16421 4929 16455 4991
rect 16657 4929 16691 4991
rect 16775 4991 17046 5019
rect 17563 4995 17833 5023
rect 16775 4929 16809 4991
rect 17011 4929 17046 4991
rect 17187 4979 17358 4995
rect 17187 4945 17318 4979
rect 17352 4945 17358 4979
rect 17187 4929 17358 4945
rect 17563 4933 17597 4995
rect 17799 4933 17833 4995
rect 17917 4995 18193 5023
rect 20933 5039 20977 5147
rect 21109 5039 21153 5147
rect 22730 5105 22786 5113
rect 20933 4997 21153 5039
rect 21804 5097 22786 5105
rect 21804 5063 22746 5097
rect 22780 5063 22786 5097
rect 23449 5093 23459 5201
rect 23591 5138 23601 5201
rect 23591 5127 23603 5138
rect 23591 5093 23604 5127
rect 23860 5117 23916 5119
rect 21804 5047 22786 5063
rect 23459 5055 23604 5093
rect 21804 5046 22783 5047
rect 17917 4933 17951 4995
rect 18153 4933 18193 4995
rect 16297 4917 16343 4929
rect 16297 4541 16303 4917
rect 16337 4541 16343 4917
rect 16297 4529 16343 4541
rect 16415 4917 16461 4929
rect 16415 4541 16421 4917
rect 16455 4541 16461 4917
rect 16415 4529 16461 4541
rect 16533 4917 16579 4929
rect 16533 4541 16539 4917
rect 16573 4541 16579 4917
rect 16533 4529 16579 4541
rect 16651 4917 16697 4929
rect 16651 4541 16657 4917
rect 16691 4541 16697 4917
rect 16651 4529 16697 4541
rect 16769 4917 16815 4929
rect 16769 4541 16775 4917
rect 16809 4541 16815 4917
rect 16769 4529 16815 4541
rect 16887 4917 16933 4929
rect 16887 4541 16893 4917
rect 16927 4541 16933 4917
rect 16887 4529 16933 4541
rect 17005 4917 17051 4929
rect 17005 4541 17011 4917
rect 17045 4541 17051 4917
rect 17005 4529 17051 4541
rect 15039 4424 15313 4452
rect 14685 4420 15313 4424
rect 14209 4408 14255 4420
rect 12628 4369 12727 4373
rect 11619 4301 11728 4355
rect 10939 4262 11166 4298
rect 10939 4155 10974 4262
rect 11100 4228 11166 4262
rect 11100 4194 11116 4228
rect 11150 4194 11166 4228
rect 11447 4286 11544 4301
rect 11447 4219 11504 4286
rect 11100 4188 11166 4194
rect 11341 4183 11610 4219
rect 11341 4155 11374 4183
rect 11577 4155 11610 4183
rect 11694 4155 11728 4301
rect 12545 4294 12555 4369
rect 12623 4294 12727 4369
rect 12572 4293 12727 4294
rect 10815 4143 10861 4155
rect 10815 3967 10821 4143
rect 10855 3967 10861 4143
rect 10815 3955 10861 3967
rect 10933 4143 10979 4155
rect 10933 3967 10939 4143
rect 10973 3967 10979 4143
rect 10933 3955 10979 3967
rect 11051 4143 11097 4155
rect 11051 3967 11057 4143
rect 11091 3967 11097 4143
rect 11051 3955 11097 3967
rect 11169 4143 11215 4155
rect 11169 3967 11175 4143
rect 11209 4088 11215 4143
rect 11334 4143 11380 4155
rect 11334 4088 11340 4143
rect 11209 4000 11340 4088
rect 11209 3967 11215 4000
rect 11169 3955 11215 3967
rect 11334 3967 11340 4000
rect 11374 3967 11380 4143
rect 11334 3955 11380 3967
rect 11452 4143 11498 4155
rect 11452 3967 11458 4143
rect 11492 3967 11498 4143
rect 11452 3955 11498 3967
rect 11570 4143 11616 4155
rect 11570 3967 11576 4143
rect 11610 3967 11616 4143
rect 11570 3955 11616 3967
rect 11688 4143 11734 4155
rect 11688 3967 11694 4143
rect 11728 3967 11734 4143
rect 11688 3955 11734 3967
rect 10821 3916 10855 3955
rect 11057 3916 11091 3955
rect 10821 3880 11091 3916
rect 11458 3917 11491 3955
rect 11694 3917 11727 3955
rect 11458 3881 11727 3917
rect 10821 3879 10987 3880
rect 10855 3800 10987 3879
rect 10845 3692 10855 3800
rect 10987 3692 10997 3800
rect 7459 3318 8436 3348
rect 10653 3346 10716 3363
rect 10578 3342 10716 3346
rect 7459 3212 7491 3318
rect 7695 3212 7727 3318
rect 7931 3212 7963 3318
rect 8167 3212 8199 3318
rect 8402 3212 8436 3318
rect 8746 3308 10716 3342
rect 8744 3279 10716 3308
rect 8744 3263 8790 3279
rect 10578 3277 10716 3279
rect 7452 3200 7498 3212
rect 7452 3024 7458 3200
rect 7492 3024 7498 3200
rect 7452 3012 7498 3024
rect 7570 3200 7616 3212
rect 7570 3024 7576 3200
rect 7610 3024 7616 3200
rect 7570 3012 7616 3024
rect 7688 3200 7734 3212
rect 7688 3024 7694 3200
rect 7728 3024 7734 3200
rect 7688 3012 7734 3024
rect 7806 3200 7852 3212
rect 7806 3024 7812 3200
rect 7846 3024 7852 3200
rect 7806 3012 7852 3024
rect 7924 3200 7970 3212
rect 7924 3024 7930 3200
rect 7964 3024 7970 3200
rect 7924 3012 7970 3024
rect 8042 3200 8088 3212
rect 8042 3024 8048 3200
rect 8082 3024 8088 3200
rect 8042 3012 8088 3024
rect 8160 3200 8206 3212
rect 8160 3024 8166 3200
rect 8200 3024 8206 3200
rect 8160 3012 8206 3024
rect 8278 3200 8324 3212
rect 8278 3024 8284 3200
rect 8318 3024 8324 3200
rect 8278 3012 8324 3024
rect 8396 3200 8442 3212
rect 8396 3024 8402 3200
rect 8436 3024 8442 3200
rect 8396 3012 8442 3024
rect 8514 3200 8560 3212
rect 8514 3024 8520 3200
rect 8554 3024 8560 3200
rect 8514 3012 8560 3024
rect 7575 2918 7611 3012
rect 7811 2918 7847 3012
rect 8047 2919 8083 3012
rect 8209 2964 8275 2971
rect 8209 2930 8225 2964
rect 8259 2930 8275 2964
rect 8209 2919 8275 2930
rect 8047 2918 8275 2919
rect 7575 2889 8275 2918
rect 7575 2888 8157 2889
rect 7695 2775 7729 2888
rect 8091 2847 8157 2888
rect 8091 2813 8107 2847
rect 8141 2813 8157 2847
rect 8091 2806 8157 2813
rect 8519 2794 8554 3012
rect 8743 2811 8790 3263
rect 9702 3047 9712 3155
rect 9844 3047 9854 3155
rect 11600 3047 11610 3155
rect 11742 3047 11752 3155
rect 9712 3007 9844 3047
rect 11610 3007 11742 3047
rect 9711 2941 9844 3007
rect 11609 2941 11742 3007
rect 9040 2898 10513 2941
rect 8743 2795 8789 2811
rect 8708 2794 8789 2795
rect 8519 2779 8789 2794
rect 8165 2775 8789 2779
rect 7689 2763 7735 2775
rect 7424 2285 7434 2403
rect 7552 2371 7562 2403
rect 7689 2387 7695 2763
rect 7729 2387 7735 2763
rect 7689 2375 7735 2387
rect 7807 2763 7853 2775
rect 7807 2387 7813 2763
rect 7847 2387 7853 2763
rect 7807 2375 7853 2387
rect 7925 2763 7971 2775
rect 7925 2387 7931 2763
rect 7965 2411 7971 2763
rect 8042 2763 8088 2775
rect 8042 2587 8048 2763
rect 8082 2587 8088 2763
rect 8042 2575 8088 2587
rect 8160 2763 8789 2775
rect 8160 2587 8166 2763
rect 8200 2751 8789 2763
rect 8200 2750 8442 2751
rect 8200 2587 8206 2750
rect 8708 2749 8789 2751
rect 9040 2595 9074 2898
rect 9406 2795 9440 2898
rect 9642 2795 9676 2898
rect 9878 2795 9912 2898
rect 10114 2795 10148 2898
rect 9400 2783 9446 2795
rect 8160 2575 8206 2587
rect 8916 2583 8962 2595
rect 8048 2459 8083 2575
rect 8179 2459 8287 2469
rect 8048 2411 8179 2459
rect 7965 2387 8179 2411
rect 7925 2375 8179 2387
rect 7931 2371 8179 2375
rect 7552 2343 7567 2371
rect 7552 2337 7804 2343
rect 7552 2303 7754 2337
rect 7788 2303 7804 2337
rect 7552 2287 7804 2303
rect 7856 2337 7922 2343
rect 7856 2303 7872 2337
rect 7906 2303 7922 2337
rect 8105 2327 8179 2371
rect 8916 2407 8922 2583
rect 8956 2407 8962 2583
rect 8916 2395 8962 2407
rect 9034 2583 9080 2595
rect 9034 2407 9040 2583
rect 9074 2407 9080 2583
rect 9034 2395 9080 2407
rect 9152 2583 9198 2595
rect 9152 2407 9158 2583
rect 9192 2407 9198 2583
rect 9152 2395 9198 2407
rect 9270 2583 9316 2595
rect 9400 2583 9406 2783
rect 9270 2407 9276 2583
rect 9310 2407 9406 2583
rect 9440 2407 9446 2783
rect 9270 2395 9316 2407
rect 9400 2395 9446 2407
rect 9518 2783 9564 2795
rect 9518 2407 9524 2783
rect 9558 2407 9564 2783
rect 9518 2395 9564 2407
rect 9636 2783 9682 2795
rect 9636 2407 9642 2783
rect 9676 2407 9682 2783
rect 9636 2395 9682 2407
rect 9754 2783 9800 2795
rect 9754 2407 9760 2783
rect 9794 2407 9800 2783
rect 9754 2395 9800 2407
rect 9872 2783 9918 2795
rect 9872 2407 9878 2783
rect 9912 2407 9918 2783
rect 9872 2395 9918 2407
rect 9990 2783 10036 2795
rect 9990 2407 9996 2783
rect 10030 2407 10036 2783
rect 9990 2395 10036 2407
rect 10108 2783 10154 2795
rect 10108 2407 10114 2783
rect 10148 2583 10154 2783
rect 10479 2595 10513 2898
rect 10938 2898 12411 2941
rect 10938 2595 10972 2898
rect 11304 2795 11338 2898
rect 11540 2795 11574 2898
rect 11776 2795 11810 2898
rect 12012 2795 12046 2898
rect 11298 2783 11344 2795
rect 10237 2583 10283 2595
rect 10148 2407 10243 2583
rect 10277 2407 10283 2583
rect 10108 2395 10154 2407
rect 10237 2395 10283 2407
rect 10355 2583 10401 2595
rect 10355 2407 10361 2583
rect 10395 2407 10401 2583
rect 10355 2395 10401 2407
rect 10473 2583 10519 2595
rect 10473 2407 10479 2583
rect 10513 2407 10519 2583
rect 10473 2395 10519 2407
rect 10591 2583 10637 2595
rect 10591 2407 10597 2583
rect 10631 2407 10637 2583
rect 10591 2395 10637 2407
rect 10814 2583 10860 2595
rect 10814 2407 10820 2583
rect 10854 2407 10860 2583
rect 10814 2395 10860 2407
rect 10932 2583 10978 2595
rect 10932 2407 10938 2583
rect 10972 2407 10978 2583
rect 10932 2395 10978 2407
rect 11050 2583 11096 2595
rect 11050 2407 11056 2583
rect 11090 2407 11096 2583
rect 11050 2395 11096 2407
rect 11168 2583 11214 2595
rect 11298 2583 11304 2783
rect 11168 2407 11174 2583
rect 11208 2407 11304 2583
rect 11338 2407 11344 2783
rect 11168 2395 11214 2407
rect 11298 2395 11344 2407
rect 11416 2783 11462 2795
rect 11416 2407 11422 2783
rect 11456 2407 11462 2783
rect 11416 2395 11462 2407
rect 11534 2783 11580 2795
rect 11534 2407 11540 2783
rect 11574 2407 11580 2783
rect 11534 2395 11580 2407
rect 11652 2783 11698 2795
rect 11652 2407 11658 2783
rect 11692 2407 11698 2783
rect 11652 2395 11698 2407
rect 11770 2783 11816 2795
rect 11770 2407 11776 2783
rect 11810 2407 11816 2783
rect 11770 2395 11816 2407
rect 11888 2783 11934 2795
rect 11888 2407 11894 2783
rect 11928 2407 11934 2783
rect 11888 2395 11934 2407
rect 12006 2783 12052 2795
rect 12006 2407 12012 2783
rect 12046 2583 12052 2783
rect 12377 2595 12411 2898
rect 12135 2583 12181 2595
rect 12046 2407 12141 2583
rect 12175 2407 12181 2583
rect 12006 2395 12052 2407
rect 12135 2395 12181 2407
rect 12253 2583 12299 2595
rect 12253 2407 12259 2583
rect 12293 2407 12299 2583
rect 12253 2395 12299 2407
rect 12371 2583 12417 2595
rect 12371 2407 12377 2583
rect 12411 2407 12417 2583
rect 12371 2395 12417 2407
rect 12489 2583 12535 2595
rect 12489 2407 12495 2583
rect 12529 2407 12535 2583
rect 12628 2547 12727 4293
rect 13037 4015 13326 4190
rect 14209 4032 14215 4408
rect 14249 4032 14255 4408
rect 14209 4020 14255 4032
rect 14327 4408 14373 4420
rect 14327 4032 14333 4408
rect 14367 4032 14373 4408
rect 14327 4020 14373 4032
rect 14445 4408 14491 4420
rect 14445 4032 14451 4408
rect 14485 4056 14491 4408
rect 14562 4408 14608 4420
rect 14562 4232 14568 4408
rect 14602 4232 14608 4408
rect 14562 4220 14608 4232
rect 14680 4408 15313 4420
rect 14680 4232 14686 4408
rect 14720 4395 15313 4408
rect 16303 4487 16337 4529
rect 16539 4487 16573 4529
rect 16303 4459 16573 4487
rect 16657 4488 16691 4529
rect 16893 4488 16927 4529
rect 16657 4459 16927 4488
rect 16303 4411 16337 4459
rect 14720 4232 14726 4395
rect 16303 4381 16366 4411
rect 14680 4220 14726 4232
rect 16331 4289 16366 4381
rect 16331 4253 16558 4289
rect 16828 4278 16838 4375
rect 16937 4278 16947 4375
rect 17011 4346 17045 4529
rect 17011 4292 17120 4346
rect 14568 4104 14603 4220
rect 16331 4146 16366 4253
rect 16492 4219 16558 4253
rect 16492 4185 16508 4219
rect 16542 4185 16558 4219
rect 16839 4277 16936 4278
rect 16839 4210 16896 4277
rect 16492 4179 16558 4185
rect 16733 4174 17002 4210
rect 16733 4146 16766 4174
rect 16969 4146 17002 4174
rect 17086 4146 17120 4292
rect 16207 4134 16253 4146
rect 14699 4104 14807 4114
rect 14568 4056 14699 4104
rect 14485 4032 14699 4056
rect 14445 4020 14699 4032
rect 14451 4016 14699 4020
rect 13037 3988 14087 4015
rect 13037 3982 14324 3988
rect 13037 3948 14274 3982
rect 14308 3948 14324 3982
rect 13037 3932 14324 3948
rect 14376 3982 14442 3988
rect 14376 3948 14392 3982
rect 14426 3948 14442 3982
rect 14625 3972 14699 4016
rect 14699 3962 14807 3972
rect 13037 3916 14087 3932
rect 13037 3915 14024 3916
rect 13037 3911 13559 3915
rect 13037 3910 13326 3911
rect 13054 3500 13343 3662
rect 13054 3394 13191 3500
rect 13303 3487 13343 3500
rect 13303 3394 13345 3487
rect 13054 3383 13345 3394
rect 13054 3382 13343 3383
rect 13054 2547 13342 2550
rect 12628 2437 13342 2547
rect 12489 2395 12535 2407
rect 8179 2317 8287 2327
rect 8922 2361 8956 2395
rect 9524 2361 9558 2395
rect 9760 2361 9794 2395
rect 8922 2326 9081 2361
rect 9524 2326 9794 2361
rect 10361 2361 10395 2395
rect 10597 2361 10631 2395
rect 10361 2326 10631 2361
rect 10820 2361 10854 2395
rect 11422 2361 11456 2395
rect 11658 2361 11692 2395
rect 10820 2326 10979 2361
rect 11422 2326 11692 2361
rect 12259 2361 12293 2395
rect 12495 2361 12529 2395
rect 12259 2326 12529 2361
rect 13054 2388 13342 2437
rect 7552 2285 7567 2287
rect 7467 2271 7567 2285
rect 7467 2228 7567 2229
rect 7088 2207 7567 2228
rect 7856 2207 7922 2303
rect 7088 2159 7922 2207
rect 7088 2130 7567 2159
rect 7088 2128 7193 2130
rect 7467 2129 7567 2130
rect 6921 1943 6931 2022
rect 7024 1943 7034 2022
rect 6091 1688 6247 1694
rect 6091 1590 6103 1688
rect 6235 1590 6247 1688
rect 6091 1584 6247 1590
rect 6932 769 7025 1943
rect 7850 1894 8070 1914
rect 7850 1786 7894 1894
rect 8026 1786 8070 1894
rect 7850 1744 8070 1786
rect 7454 1714 8431 1744
rect 7454 1608 7486 1714
rect 7690 1608 7722 1714
rect 7926 1608 7958 1714
rect 8162 1608 8194 1714
rect 8397 1608 8431 1714
rect 7447 1596 7493 1608
rect 7447 1420 7453 1596
rect 7487 1420 7493 1596
rect 7447 1408 7493 1420
rect 7565 1596 7611 1608
rect 7565 1420 7571 1596
rect 7605 1420 7611 1596
rect 7565 1408 7611 1420
rect 7683 1596 7729 1608
rect 7683 1420 7689 1596
rect 7723 1420 7729 1596
rect 7683 1408 7729 1420
rect 7801 1596 7847 1608
rect 7801 1420 7807 1596
rect 7841 1420 7847 1596
rect 7801 1408 7847 1420
rect 7919 1596 7965 1608
rect 7919 1420 7925 1596
rect 7959 1420 7965 1596
rect 7919 1408 7965 1420
rect 8037 1596 8083 1608
rect 8037 1420 8043 1596
rect 8077 1420 8083 1596
rect 8037 1408 8083 1420
rect 8155 1596 8201 1608
rect 8155 1420 8161 1596
rect 8195 1420 8201 1596
rect 8155 1408 8201 1420
rect 8273 1596 8319 1608
rect 8273 1420 8279 1596
rect 8313 1420 8319 1596
rect 8273 1408 8319 1420
rect 8391 1596 8437 1608
rect 8391 1420 8397 1596
rect 8431 1420 8437 1596
rect 8391 1408 8437 1420
rect 8509 1596 8555 1608
rect 8509 1420 8515 1596
rect 8549 1420 8555 1596
rect 8509 1408 8555 1420
rect 9047 1542 9081 2326
rect 9760 2264 9794 2326
rect 9349 2226 10091 2264
rect 9349 2102 9383 2226
rect 9585 2102 9619 2226
rect 9821 2102 9855 2226
rect 10057 2102 10091 2226
rect 10347 2119 10357 2185
rect 10420 2119 10430 2185
rect 9343 2090 9389 2102
rect 9343 1714 9349 2090
rect 9383 1714 9389 2090
rect 9343 1702 9389 1714
rect 9461 2090 9507 2102
rect 9461 1714 9467 2090
rect 9501 1714 9507 2090
rect 9461 1702 9507 1714
rect 9579 2090 9625 2102
rect 9579 1714 9585 2090
rect 9619 1714 9625 2090
rect 9579 1702 9625 1714
rect 9697 2090 9743 2102
rect 9697 1714 9703 2090
rect 9737 1714 9743 2090
rect 9697 1702 9743 1714
rect 9815 2090 9861 2102
rect 9815 1714 9821 2090
rect 9855 1714 9861 2090
rect 9815 1702 9861 1714
rect 9933 2090 9979 2102
rect 9933 1714 9939 2090
rect 9973 1714 9979 2090
rect 9933 1702 9979 1714
rect 10051 2090 10097 2102
rect 10051 1714 10057 2090
rect 10091 1714 10097 2090
rect 10051 1702 10097 1714
rect 10463 1543 10497 2326
rect 10190 1542 10497 1543
rect 9047 1537 9363 1542
rect 10077 1537 10497 1542
rect 9047 1526 9430 1537
rect 9047 1499 9379 1526
rect 7570 1314 7606 1408
rect 7806 1314 7842 1408
rect 8042 1315 8078 1408
rect 8204 1360 8270 1367
rect 8204 1326 8220 1360
rect 8254 1326 8270 1360
rect 8204 1315 8270 1326
rect 8042 1314 8270 1315
rect 7570 1285 8270 1314
rect 7570 1284 8152 1285
rect 7690 1171 7724 1284
rect 8086 1243 8152 1284
rect 8086 1209 8102 1243
rect 8136 1209 8152 1243
rect 8086 1202 8152 1209
rect 8514 1175 8549 1408
rect 9047 1370 9081 1499
rect 9363 1492 9379 1499
rect 9413 1492 9430 1526
rect 9363 1486 9430 1492
rect 10010 1526 10497 1537
rect 10010 1492 10027 1526
rect 10061 1499 10497 1526
rect 10061 1492 10077 1499
rect 10190 1498 10497 1499
rect 10010 1486 10077 1492
rect 9188 1459 9244 1471
rect 9188 1425 9194 1459
rect 9228 1458 9244 1459
rect 10301 1458 10357 1470
rect 9228 1442 9695 1458
rect 9228 1425 9645 1442
rect 9188 1409 9645 1425
rect 9629 1408 9645 1409
rect 9679 1408 9695 1442
rect 9629 1401 9695 1408
rect 9747 1443 10317 1458
rect 9747 1409 9763 1443
rect 9797 1424 10317 1443
rect 10351 1424 10357 1458
rect 9797 1409 10357 1424
rect 9747 1399 9814 1409
rect 10301 1408 10357 1409
rect 10463 1370 10497 1498
rect 10945 1542 10979 2326
rect 11658 2264 11692 2326
rect 11247 2226 11989 2264
rect 11247 2102 11281 2226
rect 11483 2102 11517 2226
rect 11719 2102 11753 2226
rect 11955 2102 11989 2226
rect 11241 2090 11287 2102
rect 11241 1714 11247 2090
rect 11281 1714 11287 2090
rect 11241 1702 11287 1714
rect 11359 2090 11405 2102
rect 11359 1714 11365 2090
rect 11399 1714 11405 2090
rect 11359 1702 11405 1714
rect 11477 2090 11523 2102
rect 11477 1714 11483 2090
rect 11517 1714 11523 2090
rect 11477 1702 11523 1714
rect 11595 2090 11641 2102
rect 11595 1714 11601 2090
rect 11635 1714 11641 2090
rect 11595 1702 11641 1714
rect 11713 2090 11759 2102
rect 11713 1714 11719 2090
rect 11753 1714 11759 2090
rect 11713 1702 11759 1714
rect 11831 2090 11877 2102
rect 11831 1714 11837 2090
rect 11871 1714 11877 2090
rect 11831 1702 11877 1714
rect 11949 2090 11995 2102
rect 11949 1714 11955 2090
rect 11989 1714 11995 2090
rect 11949 1702 11995 1714
rect 12361 1543 12395 2326
rect 13054 2282 13190 2388
rect 13302 2386 13342 2388
rect 13308 2375 13342 2386
rect 13054 2280 13196 2282
rect 13308 2280 13343 2375
rect 13054 2271 13343 2280
rect 13054 2270 13342 2271
rect 13054 2269 13310 2270
rect 11973 1542 12042 1543
rect 12088 1542 12395 1543
rect 10945 1537 11261 1542
rect 11973 1538 12395 1542
rect 10945 1526 11328 1537
rect 10945 1499 11277 1526
rect 10945 1370 10979 1499
rect 11261 1492 11277 1499
rect 11311 1492 11328 1526
rect 11261 1486 11328 1492
rect 11906 1527 12395 1538
rect 11906 1493 11923 1527
rect 11957 1499 12395 1527
rect 11957 1493 11973 1499
rect 12088 1498 12395 1499
rect 11906 1487 11973 1493
rect 11086 1459 11142 1471
rect 11086 1425 11092 1459
rect 11126 1458 11142 1459
rect 12199 1458 12255 1470
rect 11126 1442 11593 1458
rect 11126 1425 11543 1442
rect 11086 1409 11543 1425
rect 11527 1408 11543 1409
rect 11577 1408 11593 1442
rect 11527 1401 11593 1408
rect 11645 1443 12215 1458
rect 11645 1409 11661 1443
rect 11695 1424 12215 1443
rect 12249 1424 12255 1458
rect 11695 1409 12255 1424
rect 11645 1399 11712 1409
rect 12199 1408 12255 1409
rect 12361 1370 12395 1498
rect 12476 2148 12543 2172
rect 12476 2114 12493 2148
rect 12527 2114 12543 2148
rect 8160 1171 8549 1175
rect 7684 1159 7730 1171
rect 7684 783 7690 1159
rect 7724 783 7730 1159
rect 7684 771 7730 783
rect 7802 1159 7848 1171
rect 7802 783 7808 1159
rect 7842 783 7848 1159
rect 7802 771 7848 783
rect 7920 1159 7966 1171
rect 7920 783 7926 1159
rect 7960 807 7966 1159
rect 8037 1159 8083 1171
rect 8037 983 8043 1159
rect 8077 983 8083 1159
rect 8037 971 8083 983
rect 8155 1159 8549 1171
rect 9041 1358 9087 1370
rect 9041 1182 9047 1358
rect 9081 1182 9087 1358
rect 9041 1170 9087 1182
rect 9159 1358 9205 1370
rect 9159 1182 9165 1358
rect 9199 1182 9205 1358
rect 9159 1170 9205 1182
rect 9461 1358 9507 1370
rect 8155 983 8161 1159
rect 8195 1146 8549 1159
rect 8195 983 8201 1146
rect 8471 1143 8549 1146
rect 8471 1091 8481 1143
rect 8544 1091 8554 1143
rect 8476 1085 8549 1091
rect 8155 971 8201 983
rect 8043 855 8078 971
rect 9164 876 9198 1170
rect 9461 982 9467 1358
rect 9501 982 9507 1358
rect 9461 970 9507 982
rect 9579 1358 9625 1370
rect 9579 982 9585 1358
rect 9619 982 9625 1358
rect 9579 970 9625 982
rect 9697 1358 9743 1370
rect 9697 982 9703 1358
rect 9737 982 9743 1358
rect 9697 970 9743 982
rect 9815 1358 9861 1370
rect 9815 982 9821 1358
rect 9855 982 9861 1358
rect 9815 970 9861 982
rect 9933 1358 9979 1370
rect 9933 982 9939 1358
rect 9973 982 9979 1358
rect 10339 1358 10385 1370
rect 10339 1182 10345 1358
rect 10379 1182 10385 1358
rect 10339 1170 10385 1182
rect 10457 1358 10503 1370
rect 10457 1182 10463 1358
rect 10497 1182 10503 1358
rect 10457 1170 10503 1182
rect 10939 1358 10985 1370
rect 10939 1182 10945 1358
rect 10979 1182 10985 1358
rect 10939 1170 10985 1182
rect 11057 1358 11103 1370
rect 11057 1182 11063 1358
rect 11097 1182 11103 1358
rect 11057 1170 11103 1182
rect 11359 1358 11405 1370
rect 9933 970 9979 982
rect 9821 876 9855 970
rect 10345 876 10378 1170
rect 8174 855 8282 865
rect 8043 807 8174 855
rect 7960 783 8174 807
rect 7920 771 8174 783
rect 6932 767 7517 769
rect 7926 767 8174 771
rect 6932 739 7562 767
rect 1035 558 1404 606
rect 1035 528 1049 558
rect 1035 511 1045 528
rect 1337 455 1403 558
rect 5963 455 6029 734
rect 6932 733 7799 739
rect 6932 699 7749 733
rect 7783 699 7799 733
rect 6932 683 7799 699
rect 7851 733 7917 739
rect 7851 699 7867 733
rect 7901 699 7917 733
rect 8100 723 8174 767
rect 9164 844 10378 876
rect 11062 876 11096 1170
rect 11359 982 11365 1358
rect 11399 982 11405 1358
rect 11359 970 11405 982
rect 11477 1358 11523 1370
rect 11477 982 11483 1358
rect 11517 982 11523 1358
rect 11477 970 11523 982
rect 11595 1358 11641 1370
rect 11595 982 11601 1358
rect 11635 982 11641 1358
rect 11595 970 11641 982
rect 11713 1358 11759 1370
rect 11713 982 11719 1358
rect 11753 982 11759 1358
rect 11713 970 11759 982
rect 11831 1358 11877 1370
rect 11831 982 11837 1358
rect 11871 982 11877 1358
rect 12237 1358 12283 1370
rect 12237 1182 12243 1358
rect 12277 1182 12283 1358
rect 12237 1170 12283 1182
rect 12355 1358 12401 1370
rect 12355 1182 12361 1358
rect 12395 1182 12401 1358
rect 12355 1170 12401 1182
rect 11831 970 11877 982
rect 11719 876 11753 970
rect 12243 876 12276 1170
rect 11062 844 12276 876
rect 9657 759 9789 844
rect 11555 759 11687 844
rect 8174 713 8282 723
rect 6932 667 7562 683
rect 6932 663 7517 667
rect 6932 662 7033 663
rect 7462 614 7562 625
rect 7426 508 7436 614
rect 7548 603 7562 614
rect 7851 603 7917 699
rect 9647 651 9657 759
rect 9789 651 9799 759
rect 11545 651 11555 759
rect 11687 651 11697 759
rect 12476 731 12543 2114
rect 13466 2017 13559 3911
rect 13622 3852 14088 3874
rect 14376 3852 14442 3948
rect 16207 3958 16213 4134
rect 16247 3958 16253 4134
rect 16207 3946 16253 3958
rect 16325 4134 16371 4146
rect 16325 3958 16331 4134
rect 16365 3958 16371 4134
rect 16325 3946 16371 3958
rect 16443 4134 16489 4146
rect 16443 3958 16449 4134
rect 16483 3958 16489 4134
rect 16443 3946 16489 3958
rect 16561 4134 16607 4146
rect 16561 3958 16567 4134
rect 16601 4079 16607 4134
rect 16726 4134 16772 4146
rect 16726 4079 16732 4134
rect 16601 3991 16732 4079
rect 16601 3958 16607 3991
rect 16561 3946 16607 3958
rect 16726 3958 16732 3991
rect 16766 3958 16772 4134
rect 16726 3946 16772 3958
rect 16844 4134 16890 4146
rect 16844 3958 16850 4134
rect 16884 3958 16890 4134
rect 16844 3946 16890 3958
rect 16962 4134 17008 4146
rect 16962 3958 16968 4134
rect 17002 3958 17008 4134
rect 16962 3946 17008 3958
rect 17080 4134 17126 4146
rect 17080 3958 17086 4134
rect 17120 3958 17126 4134
rect 17080 3946 17126 3958
rect 16213 3907 16247 3946
rect 16449 3907 16483 3946
rect 16213 3872 16483 3907
rect 16850 3908 16883 3946
rect 17086 3908 17119 3946
rect 16850 3872 17119 3908
rect 13622 3804 14442 3852
rect 16247 3871 16483 3872
rect 13622 3773 14088 3804
rect 16247 3797 16379 3871
rect 13622 3517 13727 3773
rect 16237 3689 16247 3797
rect 16379 3689 16389 3797
rect 13622 3411 13685 3517
rect 13797 3411 13807 3517
rect 14389 3493 14609 3513
rect 13622 3400 13771 3411
rect 13622 2223 13727 3400
rect 14389 3385 14433 3493
rect 14565 3385 14609 3493
rect 14389 3343 14609 3385
rect 17187 3358 17249 4929
rect 17439 4921 17485 4933
rect 17439 4545 17445 4921
rect 17479 4545 17485 4921
rect 17439 4533 17485 4545
rect 17557 4921 17603 4933
rect 17557 4545 17563 4921
rect 17597 4545 17603 4921
rect 17557 4533 17603 4545
rect 17675 4921 17721 4933
rect 17675 4545 17681 4921
rect 17715 4545 17721 4921
rect 17675 4533 17721 4545
rect 17793 4921 17839 4933
rect 17793 4545 17799 4921
rect 17833 4545 17839 4921
rect 17793 4533 17839 4545
rect 17911 4921 17957 4933
rect 17911 4545 17917 4921
rect 17951 4545 17957 4921
rect 17911 4533 17957 4545
rect 18029 4921 18075 4933
rect 18029 4545 18035 4921
rect 18069 4545 18075 4921
rect 18029 4533 18075 4545
rect 18147 4921 18193 4933
rect 18147 4545 18153 4921
rect 18187 4545 18193 4921
rect 20537 4967 21514 4997
rect 20537 4861 20569 4967
rect 20773 4861 20805 4967
rect 21009 4861 21041 4967
rect 21245 4861 21277 4967
rect 21480 4861 21514 4967
rect 20530 4849 20576 4861
rect 20530 4673 20536 4849
rect 20570 4673 20576 4849
rect 20530 4661 20576 4673
rect 20648 4849 20694 4861
rect 20648 4673 20654 4849
rect 20688 4673 20694 4849
rect 20648 4661 20694 4673
rect 20766 4849 20812 4861
rect 20766 4673 20772 4849
rect 20806 4673 20812 4849
rect 20766 4661 20812 4673
rect 20884 4849 20930 4861
rect 20884 4673 20890 4849
rect 20924 4673 20930 4849
rect 20884 4661 20930 4673
rect 21002 4849 21048 4861
rect 21002 4673 21008 4849
rect 21042 4673 21048 4849
rect 21002 4661 21048 4673
rect 21120 4849 21166 4861
rect 21120 4673 21126 4849
rect 21160 4673 21166 4849
rect 21120 4661 21166 4673
rect 21238 4849 21284 4861
rect 21238 4673 21244 4849
rect 21278 4673 21284 4849
rect 21238 4661 21284 4673
rect 21356 4849 21402 4861
rect 21356 4673 21362 4849
rect 21396 4673 21402 4849
rect 21356 4661 21402 4673
rect 21474 4849 21520 4861
rect 21474 4673 21480 4849
rect 21514 4673 21520 4849
rect 21474 4661 21520 4673
rect 21592 4849 21638 4861
rect 21592 4673 21598 4849
rect 21632 4673 21638 4849
rect 21592 4661 21638 4673
rect 18147 4533 18193 4545
rect 20653 4567 20689 4661
rect 20889 4567 20925 4661
rect 21125 4568 21161 4661
rect 21287 4613 21353 4620
rect 21287 4579 21303 4613
rect 21337 4579 21353 4613
rect 21287 4568 21353 4579
rect 21125 4567 21353 4568
rect 20653 4538 21353 4567
rect 20653 4537 21235 4538
rect 17445 4491 17479 4533
rect 17681 4491 17715 4533
rect 17445 4463 17715 4491
rect 17799 4492 17833 4533
rect 18035 4492 18069 4533
rect 17799 4463 18069 4492
rect 17445 4415 17479 4463
rect 17445 4385 17508 4415
rect 17473 4293 17508 4385
rect 17980 4355 18080 4376
rect 17980 4301 17994 4355
rect 18059 4301 18080 4355
rect 17980 4296 18080 4301
rect 18153 4350 18187 4533
rect 20773 4424 20807 4537
rect 21169 4496 21235 4537
rect 21169 4462 21185 4496
rect 21219 4462 21235 4496
rect 21169 4455 21235 4462
rect 21597 4456 21632 4661
rect 21804 4456 21871 5046
rect 23563 5023 23604 5055
rect 23850 5051 23860 5117
rect 23916 5051 23926 5117
rect 24596 5093 24606 5201
rect 24738 5138 24748 5201
rect 24738 5127 24750 5138
rect 24738 5093 24751 5127
rect 24606 5055 24751 5093
rect 24710 5027 24751 5055
rect 22979 4995 23249 5023
rect 22720 4929 22730 4995
rect 22796 4929 22806 4995
rect 22979 4933 23013 4995
rect 23215 4933 23249 4995
rect 23333 4995 23604 5023
rect 24121 4999 24391 5027
rect 23333 4933 23367 4995
rect 23569 4933 23604 4995
rect 23745 4983 23916 4999
rect 23745 4949 23876 4983
rect 23910 4949 23916 4983
rect 23745 4933 23916 4949
rect 24121 4937 24155 4999
rect 24357 4937 24391 4999
rect 24475 4999 24751 5027
rect 24475 4937 24509 4999
rect 24711 4937 24751 4999
rect 22855 4921 22901 4933
rect 22855 4545 22861 4921
rect 22895 4545 22901 4921
rect 22855 4533 22901 4545
rect 22973 4921 23019 4933
rect 22973 4545 22979 4921
rect 23013 4545 23019 4921
rect 22973 4533 23019 4545
rect 23091 4921 23137 4933
rect 23091 4545 23097 4921
rect 23131 4545 23137 4921
rect 23091 4533 23137 4545
rect 23209 4921 23255 4933
rect 23209 4545 23215 4921
rect 23249 4545 23255 4921
rect 23209 4533 23255 4545
rect 23327 4921 23373 4933
rect 23327 4545 23333 4921
rect 23367 4545 23373 4921
rect 23327 4533 23373 4545
rect 23445 4921 23491 4933
rect 23445 4545 23451 4921
rect 23485 4545 23491 4921
rect 23445 4533 23491 4545
rect 23563 4921 23609 4933
rect 23563 4545 23569 4921
rect 23603 4545 23609 4921
rect 23563 4533 23609 4545
rect 21597 4428 21871 4456
rect 21243 4424 21871 4428
rect 20767 4412 20813 4424
rect 19165 4364 19257 4367
rect 18153 4296 18262 4350
rect 17473 4257 17700 4293
rect 17473 4150 17508 4257
rect 17634 4223 17700 4257
rect 17634 4189 17650 4223
rect 17684 4189 17700 4223
rect 17981 4281 18078 4296
rect 17981 4214 18038 4281
rect 17634 4183 17700 4189
rect 17875 4178 18144 4214
rect 17875 4150 17908 4178
rect 18111 4150 18144 4178
rect 18228 4150 18262 4296
rect 19079 4289 19089 4364
rect 19157 4289 19257 4364
rect 19106 4288 19257 4289
rect 17349 4138 17395 4150
rect 17349 3962 17355 4138
rect 17389 3962 17395 4138
rect 17349 3950 17395 3962
rect 17467 4138 17513 4150
rect 17467 3962 17473 4138
rect 17507 3962 17513 4138
rect 17467 3950 17513 3962
rect 17585 4138 17631 4150
rect 17585 3962 17591 4138
rect 17625 3962 17631 4138
rect 17585 3950 17631 3962
rect 17703 4138 17749 4150
rect 17703 3962 17709 4138
rect 17743 4083 17749 4138
rect 17868 4138 17914 4150
rect 17868 4083 17874 4138
rect 17743 3995 17874 4083
rect 17743 3962 17749 3995
rect 17703 3950 17749 3962
rect 17868 3962 17874 3995
rect 17908 3962 17914 4138
rect 17868 3950 17914 3962
rect 17986 4138 18032 4150
rect 17986 3962 17992 4138
rect 18026 3962 18032 4138
rect 17986 3950 18032 3962
rect 18104 4138 18150 4150
rect 18104 3962 18110 4138
rect 18144 3962 18150 4138
rect 18104 3950 18150 3962
rect 18222 4138 18268 4150
rect 18222 3962 18228 4138
rect 18262 3962 18268 4138
rect 18222 3950 18268 3962
rect 17355 3911 17389 3950
rect 17591 3911 17625 3950
rect 17355 3875 17625 3911
rect 17992 3912 18025 3950
rect 18228 3912 18261 3950
rect 17992 3876 18261 3912
rect 17355 3874 17521 3875
rect 17389 3795 17521 3874
rect 17379 3687 17389 3795
rect 17521 3687 17531 3795
rect 13993 3313 14970 3343
rect 17187 3341 17250 3358
rect 17112 3337 17250 3341
rect 13993 3207 14025 3313
rect 14229 3207 14261 3313
rect 14465 3207 14497 3313
rect 14701 3207 14733 3313
rect 14936 3207 14970 3313
rect 15280 3303 17250 3337
rect 15278 3274 17250 3303
rect 15278 3258 15324 3274
rect 17112 3272 17250 3274
rect 13986 3195 14032 3207
rect 13986 3019 13992 3195
rect 14026 3019 14032 3195
rect 13986 3007 14032 3019
rect 14104 3195 14150 3207
rect 14104 3019 14110 3195
rect 14144 3019 14150 3195
rect 14104 3007 14150 3019
rect 14222 3195 14268 3207
rect 14222 3019 14228 3195
rect 14262 3019 14268 3195
rect 14222 3007 14268 3019
rect 14340 3195 14386 3207
rect 14340 3019 14346 3195
rect 14380 3019 14386 3195
rect 14340 3007 14386 3019
rect 14458 3195 14504 3207
rect 14458 3019 14464 3195
rect 14498 3019 14504 3195
rect 14458 3007 14504 3019
rect 14576 3195 14622 3207
rect 14576 3019 14582 3195
rect 14616 3019 14622 3195
rect 14576 3007 14622 3019
rect 14694 3195 14740 3207
rect 14694 3019 14700 3195
rect 14734 3019 14740 3195
rect 14694 3007 14740 3019
rect 14812 3195 14858 3207
rect 14812 3019 14818 3195
rect 14852 3019 14858 3195
rect 14812 3007 14858 3019
rect 14930 3195 14976 3207
rect 14930 3019 14936 3195
rect 14970 3019 14976 3195
rect 14930 3007 14976 3019
rect 15048 3195 15094 3207
rect 15048 3019 15054 3195
rect 15088 3019 15094 3195
rect 15048 3007 15094 3019
rect 14109 2913 14145 3007
rect 14345 2913 14381 3007
rect 14581 2914 14617 3007
rect 14743 2959 14809 2966
rect 14743 2925 14759 2959
rect 14793 2925 14809 2959
rect 14743 2914 14809 2925
rect 14581 2913 14809 2914
rect 14109 2884 14809 2913
rect 14109 2883 14691 2884
rect 14229 2770 14263 2883
rect 14625 2842 14691 2883
rect 14625 2808 14641 2842
rect 14675 2808 14691 2842
rect 14625 2801 14691 2808
rect 15053 2789 15088 3007
rect 15277 2806 15324 3258
rect 16236 3042 16246 3150
rect 16378 3042 16388 3150
rect 18134 3042 18144 3150
rect 18276 3042 18286 3150
rect 16246 3002 16378 3042
rect 18144 3002 18276 3042
rect 16245 2936 16378 3002
rect 18143 2936 18276 3002
rect 15574 2893 17047 2936
rect 15277 2790 15323 2806
rect 15242 2789 15323 2790
rect 15053 2774 15323 2789
rect 14699 2770 15323 2774
rect 14223 2758 14269 2770
rect 13958 2280 13968 2398
rect 14086 2366 14096 2398
rect 14223 2382 14229 2758
rect 14263 2382 14269 2758
rect 14223 2370 14269 2382
rect 14341 2758 14387 2770
rect 14341 2382 14347 2758
rect 14381 2382 14387 2758
rect 14341 2370 14387 2382
rect 14459 2758 14505 2770
rect 14459 2382 14465 2758
rect 14499 2406 14505 2758
rect 14576 2758 14622 2770
rect 14576 2582 14582 2758
rect 14616 2582 14622 2758
rect 14576 2570 14622 2582
rect 14694 2758 15323 2770
rect 14694 2582 14700 2758
rect 14734 2746 15323 2758
rect 14734 2745 14976 2746
rect 14734 2582 14740 2745
rect 15242 2744 15323 2746
rect 15574 2590 15608 2893
rect 15940 2790 15974 2893
rect 16176 2790 16210 2893
rect 16412 2790 16446 2893
rect 16648 2790 16682 2893
rect 15934 2778 15980 2790
rect 14694 2570 14740 2582
rect 15450 2578 15496 2590
rect 14582 2454 14617 2570
rect 14713 2454 14821 2464
rect 14582 2406 14713 2454
rect 14499 2382 14713 2406
rect 14459 2370 14713 2382
rect 14465 2366 14713 2370
rect 14086 2338 14101 2366
rect 14086 2332 14338 2338
rect 14086 2298 14288 2332
rect 14322 2298 14338 2332
rect 14086 2282 14338 2298
rect 14390 2332 14456 2338
rect 14390 2298 14406 2332
rect 14440 2298 14456 2332
rect 14639 2322 14713 2366
rect 15450 2402 15456 2578
rect 15490 2402 15496 2578
rect 15450 2390 15496 2402
rect 15568 2578 15614 2590
rect 15568 2402 15574 2578
rect 15608 2402 15614 2578
rect 15568 2390 15614 2402
rect 15686 2578 15732 2590
rect 15686 2402 15692 2578
rect 15726 2402 15732 2578
rect 15686 2390 15732 2402
rect 15804 2578 15850 2590
rect 15934 2578 15940 2778
rect 15804 2402 15810 2578
rect 15844 2402 15940 2578
rect 15974 2402 15980 2778
rect 15804 2390 15850 2402
rect 15934 2390 15980 2402
rect 16052 2778 16098 2790
rect 16052 2402 16058 2778
rect 16092 2402 16098 2778
rect 16052 2390 16098 2402
rect 16170 2778 16216 2790
rect 16170 2402 16176 2778
rect 16210 2402 16216 2778
rect 16170 2390 16216 2402
rect 16288 2778 16334 2790
rect 16288 2402 16294 2778
rect 16328 2402 16334 2778
rect 16288 2390 16334 2402
rect 16406 2778 16452 2790
rect 16406 2402 16412 2778
rect 16446 2402 16452 2778
rect 16406 2390 16452 2402
rect 16524 2778 16570 2790
rect 16524 2402 16530 2778
rect 16564 2402 16570 2778
rect 16524 2390 16570 2402
rect 16642 2778 16688 2790
rect 16642 2402 16648 2778
rect 16682 2578 16688 2778
rect 17013 2590 17047 2893
rect 17472 2893 18945 2936
rect 17472 2590 17506 2893
rect 17838 2790 17872 2893
rect 18074 2790 18108 2893
rect 18310 2790 18344 2893
rect 18546 2790 18580 2893
rect 17832 2778 17878 2790
rect 16771 2578 16817 2590
rect 16682 2402 16777 2578
rect 16811 2402 16817 2578
rect 16642 2390 16688 2402
rect 16771 2390 16817 2402
rect 16889 2578 16935 2590
rect 16889 2402 16895 2578
rect 16929 2402 16935 2578
rect 16889 2390 16935 2402
rect 17007 2578 17053 2590
rect 17007 2402 17013 2578
rect 17047 2402 17053 2578
rect 17007 2390 17053 2402
rect 17125 2578 17171 2590
rect 17125 2402 17131 2578
rect 17165 2402 17171 2578
rect 17125 2390 17171 2402
rect 17348 2578 17394 2590
rect 17348 2402 17354 2578
rect 17388 2402 17394 2578
rect 17348 2390 17394 2402
rect 17466 2578 17512 2590
rect 17466 2402 17472 2578
rect 17506 2402 17512 2578
rect 17466 2390 17512 2402
rect 17584 2578 17630 2590
rect 17584 2402 17590 2578
rect 17624 2402 17630 2578
rect 17584 2390 17630 2402
rect 17702 2578 17748 2590
rect 17832 2578 17838 2778
rect 17702 2402 17708 2578
rect 17742 2402 17838 2578
rect 17872 2402 17878 2778
rect 17702 2390 17748 2402
rect 17832 2390 17878 2402
rect 17950 2778 17996 2790
rect 17950 2402 17956 2778
rect 17990 2402 17996 2778
rect 17950 2390 17996 2402
rect 18068 2778 18114 2790
rect 18068 2402 18074 2778
rect 18108 2402 18114 2778
rect 18068 2390 18114 2402
rect 18186 2778 18232 2790
rect 18186 2402 18192 2778
rect 18226 2402 18232 2778
rect 18186 2390 18232 2402
rect 18304 2778 18350 2790
rect 18304 2402 18310 2778
rect 18344 2402 18350 2778
rect 18304 2390 18350 2402
rect 18422 2778 18468 2790
rect 18422 2402 18428 2778
rect 18462 2402 18468 2778
rect 18422 2390 18468 2402
rect 18540 2778 18586 2790
rect 18540 2402 18546 2778
rect 18580 2578 18586 2778
rect 18911 2590 18945 2893
rect 18669 2578 18715 2590
rect 18580 2402 18675 2578
rect 18709 2402 18715 2578
rect 18540 2390 18586 2402
rect 18669 2390 18715 2402
rect 18787 2578 18833 2590
rect 18787 2402 18793 2578
rect 18827 2402 18833 2578
rect 18787 2390 18833 2402
rect 18905 2578 18951 2590
rect 18905 2402 18911 2578
rect 18945 2402 18951 2578
rect 18905 2390 18951 2402
rect 19023 2578 19069 2590
rect 19023 2402 19029 2578
rect 19063 2402 19069 2578
rect 19165 2552 19257 4288
rect 19595 4019 19884 4194
rect 20767 4036 20773 4412
rect 20807 4036 20813 4412
rect 20767 4024 20813 4036
rect 20885 4412 20931 4424
rect 20885 4036 20891 4412
rect 20925 4036 20931 4412
rect 20885 4024 20931 4036
rect 21003 4412 21049 4424
rect 21003 4036 21009 4412
rect 21043 4060 21049 4412
rect 21120 4412 21166 4424
rect 21120 4236 21126 4412
rect 21160 4236 21166 4412
rect 21120 4224 21166 4236
rect 21238 4412 21871 4424
rect 21238 4236 21244 4412
rect 21278 4399 21871 4412
rect 22861 4491 22895 4533
rect 23097 4491 23131 4533
rect 22861 4463 23131 4491
rect 23215 4492 23249 4533
rect 23451 4492 23485 4533
rect 23215 4463 23485 4492
rect 22861 4415 22895 4463
rect 21278 4236 21284 4399
rect 22861 4385 22924 4415
rect 21238 4224 21284 4236
rect 22889 4293 22924 4385
rect 22889 4257 23116 4293
rect 23386 4282 23396 4379
rect 23495 4282 23505 4379
rect 23569 4350 23603 4533
rect 23569 4296 23678 4350
rect 21126 4108 21161 4224
rect 22889 4150 22924 4257
rect 23050 4223 23116 4257
rect 23050 4189 23066 4223
rect 23100 4189 23116 4223
rect 23397 4281 23494 4282
rect 23397 4214 23454 4281
rect 23050 4183 23116 4189
rect 23291 4178 23560 4214
rect 23291 4150 23324 4178
rect 23527 4150 23560 4178
rect 23644 4150 23678 4296
rect 22765 4138 22811 4150
rect 21257 4108 21365 4118
rect 21126 4060 21257 4108
rect 21043 4036 21257 4060
rect 21003 4024 21257 4036
rect 21009 4020 21257 4024
rect 19595 3992 20645 4019
rect 19595 3986 20882 3992
rect 19595 3952 20832 3986
rect 20866 3952 20882 3986
rect 19595 3936 20882 3952
rect 20934 3986 21000 3992
rect 20934 3952 20950 3986
rect 20984 3952 21000 3986
rect 21183 3976 21257 4020
rect 21257 3966 21365 3976
rect 19595 3920 20645 3936
rect 19595 3919 20582 3920
rect 19595 3915 20117 3919
rect 19595 3914 19884 3915
rect 19612 3504 19901 3666
rect 19612 3398 19749 3504
rect 19861 3491 19901 3504
rect 19861 3398 19903 3491
rect 19612 3387 19903 3398
rect 19612 3386 19901 3387
rect 19612 2552 19900 2554
rect 19165 2436 19900 2552
rect 19023 2390 19069 2402
rect 19612 2392 19900 2436
rect 14713 2312 14821 2322
rect 15456 2356 15490 2390
rect 16058 2356 16092 2390
rect 16294 2356 16328 2390
rect 15456 2321 15615 2356
rect 16058 2321 16328 2356
rect 16895 2356 16929 2390
rect 17131 2356 17165 2390
rect 16895 2321 17165 2356
rect 17354 2356 17388 2390
rect 17956 2356 17990 2390
rect 18192 2356 18226 2390
rect 17354 2321 17513 2356
rect 17956 2321 18226 2356
rect 18793 2356 18827 2390
rect 19029 2356 19063 2390
rect 18793 2321 19063 2356
rect 14086 2280 14101 2282
rect 14001 2266 14101 2280
rect 14001 2223 14101 2224
rect 13622 2202 14101 2223
rect 14390 2202 14456 2298
rect 13622 2154 14456 2202
rect 13622 2125 14101 2154
rect 13622 2123 13727 2125
rect 14001 2124 14101 2125
rect 13455 1938 13465 2017
rect 13558 1938 13568 2017
rect 12604 1685 12760 1691
rect 12604 1587 12616 1685
rect 12748 1587 12760 1685
rect 12604 1581 12760 1587
rect 13466 764 13559 1938
rect 14384 1889 14604 1909
rect 14384 1781 14428 1889
rect 14560 1781 14604 1889
rect 14384 1739 14604 1781
rect 13988 1709 14965 1739
rect 13988 1603 14020 1709
rect 14224 1603 14256 1709
rect 14460 1603 14492 1709
rect 14696 1603 14728 1709
rect 14931 1603 14965 1709
rect 13981 1591 14027 1603
rect 13981 1415 13987 1591
rect 14021 1415 14027 1591
rect 13981 1403 14027 1415
rect 14099 1591 14145 1603
rect 14099 1415 14105 1591
rect 14139 1415 14145 1591
rect 14099 1403 14145 1415
rect 14217 1591 14263 1603
rect 14217 1415 14223 1591
rect 14257 1415 14263 1591
rect 14217 1403 14263 1415
rect 14335 1591 14381 1603
rect 14335 1415 14341 1591
rect 14375 1415 14381 1591
rect 14335 1403 14381 1415
rect 14453 1591 14499 1603
rect 14453 1415 14459 1591
rect 14493 1415 14499 1591
rect 14453 1403 14499 1415
rect 14571 1591 14617 1603
rect 14571 1415 14577 1591
rect 14611 1415 14617 1591
rect 14571 1403 14617 1415
rect 14689 1591 14735 1603
rect 14689 1415 14695 1591
rect 14729 1415 14735 1591
rect 14689 1403 14735 1415
rect 14807 1591 14853 1603
rect 14807 1415 14813 1591
rect 14847 1415 14853 1591
rect 14807 1403 14853 1415
rect 14925 1591 14971 1603
rect 14925 1415 14931 1591
rect 14965 1415 14971 1591
rect 14925 1403 14971 1415
rect 15043 1591 15089 1603
rect 15043 1415 15049 1591
rect 15083 1415 15089 1591
rect 15043 1403 15089 1415
rect 15581 1537 15615 2321
rect 16294 2259 16328 2321
rect 15883 2221 16625 2259
rect 15883 2097 15917 2221
rect 16119 2097 16153 2221
rect 16355 2097 16389 2221
rect 16591 2097 16625 2221
rect 16881 2114 16891 2180
rect 16954 2114 16964 2180
rect 15877 2085 15923 2097
rect 15877 1709 15883 2085
rect 15917 1709 15923 2085
rect 15877 1697 15923 1709
rect 15995 2085 16041 2097
rect 15995 1709 16001 2085
rect 16035 1709 16041 2085
rect 15995 1697 16041 1709
rect 16113 2085 16159 2097
rect 16113 1709 16119 2085
rect 16153 1709 16159 2085
rect 16113 1697 16159 1709
rect 16231 2085 16277 2097
rect 16231 1709 16237 2085
rect 16271 1709 16277 2085
rect 16231 1697 16277 1709
rect 16349 2085 16395 2097
rect 16349 1709 16355 2085
rect 16389 1709 16395 2085
rect 16349 1697 16395 1709
rect 16467 2085 16513 2097
rect 16467 1709 16473 2085
rect 16507 1709 16513 2085
rect 16467 1697 16513 1709
rect 16585 2085 16631 2097
rect 16585 1709 16591 2085
rect 16625 1709 16631 2085
rect 16585 1697 16631 1709
rect 16997 1538 17031 2321
rect 16724 1537 17031 1538
rect 15581 1532 15897 1537
rect 16611 1532 17031 1537
rect 15581 1521 15964 1532
rect 15581 1494 15913 1521
rect 14104 1309 14140 1403
rect 14340 1309 14376 1403
rect 14576 1310 14612 1403
rect 14738 1355 14804 1362
rect 14738 1321 14754 1355
rect 14788 1321 14804 1355
rect 14738 1310 14804 1321
rect 14576 1309 14804 1310
rect 14104 1280 14804 1309
rect 14104 1279 14686 1280
rect 14224 1166 14258 1279
rect 14620 1238 14686 1279
rect 14620 1204 14636 1238
rect 14670 1204 14686 1238
rect 14620 1197 14686 1204
rect 15048 1170 15083 1403
rect 15581 1365 15615 1494
rect 15897 1487 15913 1494
rect 15947 1487 15964 1521
rect 15897 1481 15964 1487
rect 16544 1521 17031 1532
rect 16544 1487 16561 1521
rect 16595 1494 17031 1521
rect 16595 1487 16611 1494
rect 16724 1493 17031 1494
rect 16544 1481 16611 1487
rect 15722 1454 15778 1466
rect 15722 1420 15728 1454
rect 15762 1453 15778 1454
rect 16835 1453 16891 1465
rect 15762 1437 16229 1453
rect 15762 1420 16179 1437
rect 15722 1404 16179 1420
rect 16163 1403 16179 1404
rect 16213 1403 16229 1437
rect 16163 1396 16229 1403
rect 16281 1438 16851 1453
rect 16281 1404 16297 1438
rect 16331 1419 16851 1438
rect 16885 1419 16891 1453
rect 16331 1404 16891 1419
rect 16281 1394 16348 1404
rect 16835 1403 16891 1404
rect 16997 1365 17031 1493
rect 17479 1537 17513 2321
rect 18192 2259 18226 2321
rect 17781 2221 18523 2259
rect 17781 2097 17815 2221
rect 18017 2097 18051 2221
rect 18253 2097 18287 2221
rect 18489 2097 18523 2221
rect 17775 2085 17821 2097
rect 17775 1709 17781 2085
rect 17815 1709 17821 2085
rect 17775 1697 17821 1709
rect 17893 2085 17939 2097
rect 17893 1709 17899 2085
rect 17933 1709 17939 2085
rect 17893 1697 17939 1709
rect 18011 2085 18057 2097
rect 18011 1709 18017 2085
rect 18051 1709 18057 2085
rect 18011 1697 18057 1709
rect 18129 2085 18175 2097
rect 18129 1709 18135 2085
rect 18169 1709 18175 2085
rect 18129 1697 18175 1709
rect 18247 2085 18293 2097
rect 18247 1709 18253 2085
rect 18287 1709 18293 2085
rect 18247 1697 18293 1709
rect 18365 2085 18411 2097
rect 18365 1709 18371 2085
rect 18405 1709 18411 2085
rect 18365 1697 18411 1709
rect 18483 2085 18529 2097
rect 18483 1709 18489 2085
rect 18523 1709 18529 2085
rect 18483 1697 18529 1709
rect 18895 1538 18929 2321
rect 19612 2286 19748 2392
rect 19860 2390 19900 2392
rect 19866 2379 19900 2390
rect 19612 2284 19754 2286
rect 19866 2284 19901 2379
rect 19612 2275 19901 2284
rect 19612 2274 19900 2275
rect 19612 2273 19868 2274
rect 18507 1537 18576 1538
rect 18622 1537 18929 1538
rect 17479 1532 17795 1537
rect 18507 1533 18929 1537
rect 17479 1521 17862 1532
rect 17479 1494 17811 1521
rect 17479 1365 17513 1494
rect 17795 1487 17811 1494
rect 17845 1487 17862 1521
rect 17795 1481 17862 1487
rect 18440 1522 18929 1533
rect 18440 1488 18457 1522
rect 18491 1494 18929 1522
rect 18491 1488 18507 1494
rect 18622 1493 18929 1494
rect 18440 1482 18507 1488
rect 17620 1454 17676 1466
rect 17620 1420 17626 1454
rect 17660 1453 17676 1454
rect 18733 1453 18789 1465
rect 17660 1437 18127 1453
rect 17660 1420 18077 1437
rect 17620 1404 18077 1420
rect 18061 1403 18077 1404
rect 18111 1403 18127 1437
rect 18061 1396 18127 1403
rect 18179 1438 18749 1453
rect 18179 1404 18195 1438
rect 18229 1419 18749 1438
rect 18783 1419 18789 1453
rect 18229 1404 18789 1419
rect 18179 1394 18246 1404
rect 18733 1403 18789 1404
rect 18895 1365 18929 1493
rect 19010 2143 19077 2167
rect 19010 2109 19027 2143
rect 19061 2109 19077 2143
rect 14694 1166 15083 1170
rect 14218 1154 14264 1166
rect 14218 778 14224 1154
rect 14258 778 14264 1154
rect 14218 766 14264 778
rect 14336 1154 14382 1166
rect 14336 778 14342 1154
rect 14376 778 14382 1154
rect 14336 766 14382 778
rect 14454 1154 14500 1166
rect 14454 778 14460 1154
rect 14494 802 14500 1154
rect 14571 1154 14617 1166
rect 14571 978 14577 1154
rect 14611 978 14617 1154
rect 14571 966 14617 978
rect 14689 1154 15083 1166
rect 15575 1353 15621 1365
rect 15575 1177 15581 1353
rect 15615 1177 15621 1353
rect 15575 1165 15621 1177
rect 15693 1353 15739 1365
rect 15693 1177 15699 1353
rect 15733 1177 15739 1353
rect 15693 1165 15739 1177
rect 15995 1353 16041 1365
rect 14689 978 14695 1154
rect 14729 1141 15083 1154
rect 14729 978 14735 1141
rect 15005 1138 15083 1141
rect 15005 1086 15015 1138
rect 15078 1086 15088 1138
rect 15010 1080 15083 1086
rect 14689 966 14735 978
rect 14577 850 14612 966
rect 15698 871 15732 1165
rect 15995 977 16001 1353
rect 16035 977 16041 1353
rect 15995 965 16041 977
rect 16113 1353 16159 1365
rect 16113 977 16119 1353
rect 16153 977 16159 1353
rect 16113 965 16159 977
rect 16231 1353 16277 1365
rect 16231 977 16237 1353
rect 16271 977 16277 1353
rect 16231 965 16277 977
rect 16349 1353 16395 1365
rect 16349 977 16355 1353
rect 16389 977 16395 1353
rect 16349 965 16395 977
rect 16467 1353 16513 1365
rect 16467 977 16473 1353
rect 16507 977 16513 1353
rect 16873 1353 16919 1365
rect 16873 1177 16879 1353
rect 16913 1177 16919 1353
rect 16873 1165 16919 1177
rect 16991 1353 17037 1365
rect 16991 1177 16997 1353
rect 17031 1177 17037 1353
rect 16991 1165 17037 1177
rect 17473 1353 17519 1365
rect 17473 1177 17479 1353
rect 17513 1177 17519 1353
rect 17473 1165 17519 1177
rect 17591 1353 17637 1365
rect 17591 1177 17597 1353
rect 17631 1177 17637 1353
rect 17591 1165 17637 1177
rect 17893 1353 17939 1365
rect 16467 965 16513 977
rect 16355 871 16389 965
rect 16879 871 16912 1165
rect 14708 850 14816 860
rect 14577 802 14708 850
rect 14494 778 14708 802
rect 14454 766 14708 778
rect 13466 762 14051 764
rect 14460 762 14708 766
rect 13466 734 14096 762
rect 7548 555 7917 603
rect 7548 525 7562 555
rect 7548 508 7558 525
rect 1335 375 6029 455
rect 7850 452 7916 555
rect 12476 452 12542 731
rect 13466 728 14333 734
rect 13466 694 14283 728
rect 14317 694 14333 728
rect 13466 678 14333 694
rect 14385 728 14451 734
rect 14385 694 14401 728
rect 14435 694 14451 728
rect 14634 718 14708 762
rect 15698 839 16912 871
rect 17596 871 17630 1165
rect 17893 977 17899 1353
rect 17933 977 17939 1353
rect 17893 965 17939 977
rect 18011 1353 18057 1365
rect 18011 977 18017 1353
rect 18051 977 18057 1353
rect 18011 965 18057 977
rect 18129 1353 18175 1365
rect 18129 977 18135 1353
rect 18169 977 18175 1353
rect 18129 965 18175 977
rect 18247 1353 18293 1365
rect 18247 977 18253 1353
rect 18287 977 18293 1353
rect 18247 965 18293 977
rect 18365 1353 18411 1365
rect 18365 977 18371 1353
rect 18405 977 18411 1353
rect 18771 1353 18817 1365
rect 18771 1177 18777 1353
rect 18811 1177 18817 1353
rect 18771 1165 18817 1177
rect 18889 1353 18935 1365
rect 18889 1177 18895 1353
rect 18929 1177 18935 1353
rect 18889 1165 18935 1177
rect 18365 965 18411 977
rect 18253 871 18287 965
rect 18777 871 18810 1165
rect 17596 839 18810 871
rect 16191 754 16323 839
rect 18089 754 18221 839
rect 14708 708 14816 718
rect 13466 662 14096 678
rect 13466 658 14051 662
rect 13466 657 13567 658
rect 13996 609 14096 620
rect 13960 503 13970 609
rect 14082 598 14096 609
rect 14385 598 14451 694
rect 16181 646 16191 754
rect 16323 646 16333 754
rect 18079 646 18089 754
rect 18221 646 18231 754
rect 19010 726 19077 2109
rect 20024 2021 20117 3915
rect 20180 3856 20646 3878
rect 20934 3856 21000 3952
rect 22765 3962 22771 4138
rect 22805 3962 22811 4138
rect 22765 3950 22811 3962
rect 22883 4138 22929 4150
rect 22883 3962 22889 4138
rect 22923 3962 22929 4138
rect 22883 3950 22929 3962
rect 23001 4138 23047 4150
rect 23001 3962 23007 4138
rect 23041 3962 23047 4138
rect 23001 3950 23047 3962
rect 23119 4138 23165 4150
rect 23119 3962 23125 4138
rect 23159 4083 23165 4138
rect 23284 4138 23330 4150
rect 23284 4083 23290 4138
rect 23159 3995 23290 4083
rect 23159 3962 23165 3995
rect 23119 3950 23165 3962
rect 23284 3962 23290 3995
rect 23324 3962 23330 4138
rect 23284 3950 23330 3962
rect 23402 4138 23448 4150
rect 23402 3962 23408 4138
rect 23442 3962 23448 4138
rect 23402 3950 23448 3962
rect 23520 4138 23566 4150
rect 23520 3962 23526 4138
rect 23560 3962 23566 4138
rect 23520 3950 23566 3962
rect 23638 4138 23684 4150
rect 23638 3962 23644 4138
rect 23678 3962 23684 4138
rect 23638 3950 23684 3962
rect 22771 3911 22805 3950
rect 23007 3911 23041 3950
rect 22771 3876 23041 3911
rect 23408 3912 23441 3950
rect 23644 3912 23677 3950
rect 23408 3876 23677 3912
rect 20180 3808 21000 3856
rect 22805 3875 23041 3876
rect 20180 3777 20646 3808
rect 22805 3801 22937 3875
rect 20180 3521 20285 3777
rect 22795 3693 22805 3801
rect 22937 3693 22947 3801
rect 20180 3415 20243 3521
rect 20355 3415 20365 3521
rect 20947 3497 21167 3517
rect 20180 3404 20329 3415
rect 20180 2227 20285 3404
rect 20947 3389 20991 3497
rect 21123 3389 21167 3497
rect 20947 3347 21167 3389
rect 23745 3362 23807 4933
rect 23997 4925 24043 4937
rect 23997 4549 24003 4925
rect 24037 4549 24043 4925
rect 23997 4537 24043 4549
rect 24115 4925 24161 4937
rect 24115 4549 24121 4925
rect 24155 4549 24161 4925
rect 24115 4537 24161 4549
rect 24233 4925 24279 4937
rect 24233 4549 24239 4925
rect 24273 4549 24279 4925
rect 24233 4537 24279 4549
rect 24351 4925 24397 4937
rect 24351 4549 24357 4925
rect 24391 4549 24397 4925
rect 24351 4537 24397 4549
rect 24469 4925 24515 4937
rect 24469 4549 24475 4925
rect 24509 4549 24515 4925
rect 24469 4537 24515 4549
rect 24587 4925 24633 4937
rect 24587 4549 24593 4925
rect 24627 4549 24633 4925
rect 24587 4537 24633 4549
rect 24705 4925 24751 4937
rect 24705 4549 24711 4925
rect 24745 4549 24751 4925
rect 24705 4537 24751 4549
rect 24003 4495 24037 4537
rect 24239 4495 24273 4537
rect 24003 4467 24273 4495
rect 24357 4496 24391 4537
rect 24593 4496 24627 4537
rect 24357 4467 24627 4496
rect 24003 4419 24037 4467
rect 24003 4389 24066 4419
rect 24031 4297 24066 4389
rect 24538 4359 24638 4380
rect 24538 4305 24552 4359
rect 24617 4305 24638 4359
rect 24538 4300 24638 4305
rect 24711 4354 24745 4537
rect 25745 4368 26111 4370
rect 24711 4300 24820 4354
rect 24031 4261 24258 4297
rect 24031 4154 24066 4261
rect 24192 4227 24258 4261
rect 24192 4193 24208 4227
rect 24242 4193 24258 4227
rect 24539 4285 24636 4300
rect 24539 4218 24596 4285
rect 24192 4187 24258 4193
rect 24433 4182 24702 4218
rect 24433 4154 24466 4182
rect 24669 4154 24702 4182
rect 24786 4154 24820 4300
rect 25637 4293 25647 4368
rect 25715 4293 26111 4368
rect 25664 4292 26111 4293
rect 25710 4288 26111 4292
rect 23907 4142 23953 4154
rect 23907 3966 23913 4142
rect 23947 3966 23953 4142
rect 23907 3954 23953 3966
rect 24025 4142 24071 4154
rect 24025 3966 24031 4142
rect 24065 3966 24071 4142
rect 24025 3954 24071 3966
rect 24143 4142 24189 4154
rect 24143 3966 24149 4142
rect 24183 3966 24189 4142
rect 24143 3954 24189 3966
rect 24261 4142 24307 4154
rect 24261 3966 24267 4142
rect 24301 4087 24307 4142
rect 24426 4142 24472 4154
rect 24426 4087 24432 4142
rect 24301 3999 24432 4087
rect 24301 3966 24307 3999
rect 24261 3954 24307 3966
rect 24426 3966 24432 3999
rect 24466 3966 24472 4142
rect 24426 3954 24472 3966
rect 24544 4142 24590 4154
rect 24544 3966 24550 4142
rect 24584 3966 24590 4142
rect 24544 3954 24590 3966
rect 24662 4142 24708 4154
rect 24662 3966 24668 4142
rect 24702 3966 24708 4142
rect 24662 3954 24708 3966
rect 24780 4142 24826 4154
rect 24780 3966 24786 4142
rect 24820 3966 24826 4142
rect 24780 3954 24826 3966
rect 23913 3915 23947 3954
rect 24149 3915 24183 3954
rect 23913 3879 24183 3915
rect 24550 3916 24583 3954
rect 24786 3916 24819 3954
rect 24550 3880 24819 3916
rect 23913 3878 24079 3879
rect 23947 3799 24079 3878
rect 23937 3691 23947 3799
rect 24079 3691 24089 3799
rect 25984 3370 26111 4288
rect 20551 3317 21528 3347
rect 23745 3345 23808 3362
rect 23670 3341 23808 3345
rect 20551 3211 20583 3317
rect 20787 3211 20819 3317
rect 21023 3211 21055 3317
rect 21259 3211 21291 3317
rect 21494 3211 21528 3317
rect 21838 3307 23808 3341
rect 21836 3278 23808 3307
rect 21836 3262 21882 3278
rect 23670 3276 23808 3278
rect 25986 3263 26109 3370
rect 20544 3199 20590 3211
rect 20544 3023 20550 3199
rect 20584 3023 20590 3199
rect 20544 3011 20590 3023
rect 20662 3199 20708 3211
rect 20662 3023 20668 3199
rect 20702 3023 20708 3199
rect 20662 3011 20708 3023
rect 20780 3199 20826 3211
rect 20780 3023 20786 3199
rect 20820 3023 20826 3199
rect 20780 3011 20826 3023
rect 20898 3199 20944 3211
rect 20898 3023 20904 3199
rect 20938 3023 20944 3199
rect 20898 3011 20944 3023
rect 21016 3199 21062 3211
rect 21016 3023 21022 3199
rect 21056 3023 21062 3199
rect 21016 3011 21062 3023
rect 21134 3199 21180 3211
rect 21134 3023 21140 3199
rect 21174 3023 21180 3199
rect 21134 3011 21180 3023
rect 21252 3199 21298 3211
rect 21252 3023 21258 3199
rect 21292 3023 21298 3199
rect 21252 3011 21298 3023
rect 21370 3199 21416 3211
rect 21370 3023 21376 3199
rect 21410 3023 21416 3199
rect 21370 3011 21416 3023
rect 21488 3199 21534 3211
rect 21488 3023 21494 3199
rect 21528 3023 21534 3199
rect 21488 3011 21534 3023
rect 21606 3199 21652 3211
rect 21606 3023 21612 3199
rect 21646 3023 21652 3199
rect 21606 3011 21652 3023
rect 20667 2917 20703 3011
rect 20903 2917 20939 3011
rect 21139 2918 21175 3011
rect 21301 2963 21367 2970
rect 21301 2929 21317 2963
rect 21351 2929 21367 2963
rect 21301 2918 21367 2929
rect 21139 2917 21367 2918
rect 20667 2888 21367 2917
rect 20667 2887 21249 2888
rect 20787 2774 20821 2887
rect 21183 2846 21249 2887
rect 21183 2812 21199 2846
rect 21233 2812 21249 2846
rect 21183 2805 21249 2812
rect 21611 2793 21646 3011
rect 21835 2810 21882 3262
rect 22794 3046 22804 3154
rect 22936 3046 22946 3154
rect 24692 3046 24702 3154
rect 24834 3046 24844 3154
rect 22804 3006 22936 3046
rect 24702 3006 24834 3046
rect 22803 2940 22936 3006
rect 24701 2940 24834 3006
rect 22132 2897 23605 2940
rect 21835 2794 21881 2810
rect 21800 2793 21881 2794
rect 21611 2778 21881 2793
rect 21257 2774 21881 2778
rect 20781 2762 20827 2774
rect 20516 2284 20526 2402
rect 20644 2370 20654 2402
rect 20781 2386 20787 2762
rect 20821 2386 20827 2762
rect 20781 2374 20827 2386
rect 20899 2762 20945 2774
rect 20899 2386 20905 2762
rect 20939 2386 20945 2762
rect 20899 2374 20945 2386
rect 21017 2762 21063 2774
rect 21017 2386 21023 2762
rect 21057 2410 21063 2762
rect 21134 2762 21180 2774
rect 21134 2586 21140 2762
rect 21174 2586 21180 2762
rect 21134 2574 21180 2586
rect 21252 2762 21881 2774
rect 21252 2586 21258 2762
rect 21292 2750 21881 2762
rect 21292 2749 21534 2750
rect 21292 2586 21298 2749
rect 21800 2748 21881 2750
rect 22132 2594 22166 2897
rect 22498 2794 22532 2897
rect 22734 2794 22768 2897
rect 22970 2794 23004 2897
rect 23206 2794 23240 2897
rect 22492 2782 22538 2794
rect 21252 2574 21298 2586
rect 22008 2582 22054 2594
rect 21140 2458 21175 2574
rect 21271 2458 21379 2468
rect 21140 2410 21271 2458
rect 21057 2386 21271 2410
rect 21017 2374 21271 2386
rect 21023 2370 21271 2374
rect 20644 2342 20659 2370
rect 20644 2336 20896 2342
rect 20644 2302 20846 2336
rect 20880 2302 20896 2336
rect 20644 2286 20896 2302
rect 20948 2336 21014 2342
rect 20948 2302 20964 2336
rect 20998 2302 21014 2336
rect 21197 2326 21271 2370
rect 22008 2406 22014 2582
rect 22048 2406 22054 2582
rect 22008 2394 22054 2406
rect 22126 2582 22172 2594
rect 22126 2406 22132 2582
rect 22166 2406 22172 2582
rect 22126 2394 22172 2406
rect 22244 2582 22290 2594
rect 22244 2406 22250 2582
rect 22284 2406 22290 2582
rect 22244 2394 22290 2406
rect 22362 2582 22408 2594
rect 22492 2582 22498 2782
rect 22362 2406 22368 2582
rect 22402 2406 22498 2582
rect 22532 2406 22538 2782
rect 22362 2394 22408 2406
rect 22492 2394 22538 2406
rect 22610 2782 22656 2794
rect 22610 2406 22616 2782
rect 22650 2406 22656 2782
rect 22610 2394 22656 2406
rect 22728 2782 22774 2794
rect 22728 2406 22734 2782
rect 22768 2406 22774 2782
rect 22728 2394 22774 2406
rect 22846 2782 22892 2794
rect 22846 2406 22852 2782
rect 22886 2406 22892 2782
rect 22846 2394 22892 2406
rect 22964 2782 23010 2794
rect 22964 2406 22970 2782
rect 23004 2406 23010 2782
rect 22964 2394 23010 2406
rect 23082 2782 23128 2794
rect 23082 2406 23088 2782
rect 23122 2406 23128 2782
rect 23082 2394 23128 2406
rect 23200 2782 23246 2794
rect 23200 2406 23206 2782
rect 23240 2582 23246 2782
rect 23571 2594 23605 2897
rect 24030 2897 25503 2940
rect 24030 2594 24064 2897
rect 24396 2794 24430 2897
rect 24632 2794 24666 2897
rect 24868 2794 24902 2897
rect 25104 2794 25138 2897
rect 24390 2782 24436 2794
rect 23329 2582 23375 2594
rect 23240 2406 23335 2582
rect 23369 2406 23375 2582
rect 23200 2394 23246 2406
rect 23329 2394 23375 2406
rect 23447 2582 23493 2594
rect 23447 2406 23453 2582
rect 23487 2406 23493 2582
rect 23447 2394 23493 2406
rect 23565 2582 23611 2594
rect 23565 2406 23571 2582
rect 23605 2406 23611 2582
rect 23565 2394 23611 2406
rect 23683 2582 23729 2594
rect 23683 2406 23689 2582
rect 23723 2406 23729 2582
rect 23683 2394 23729 2406
rect 23906 2582 23952 2594
rect 23906 2406 23912 2582
rect 23946 2406 23952 2582
rect 23906 2394 23952 2406
rect 24024 2582 24070 2594
rect 24024 2406 24030 2582
rect 24064 2406 24070 2582
rect 24024 2394 24070 2406
rect 24142 2582 24188 2594
rect 24142 2406 24148 2582
rect 24182 2406 24188 2582
rect 24142 2394 24188 2406
rect 24260 2582 24306 2594
rect 24390 2582 24396 2782
rect 24260 2406 24266 2582
rect 24300 2406 24396 2582
rect 24430 2406 24436 2782
rect 24260 2394 24306 2406
rect 24390 2394 24436 2406
rect 24508 2782 24554 2794
rect 24508 2406 24514 2782
rect 24548 2406 24554 2782
rect 24508 2394 24554 2406
rect 24626 2782 24672 2794
rect 24626 2406 24632 2782
rect 24666 2406 24672 2782
rect 24626 2394 24672 2406
rect 24744 2782 24790 2794
rect 24744 2406 24750 2782
rect 24784 2406 24790 2782
rect 24744 2394 24790 2406
rect 24862 2782 24908 2794
rect 24862 2406 24868 2782
rect 24902 2406 24908 2782
rect 24862 2394 24908 2406
rect 24980 2782 25026 2794
rect 24980 2406 24986 2782
rect 25020 2406 25026 2782
rect 24980 2394 25026 2406
rect 25098 2782 25144 2794
rect 25098 2406 25104 2782
rect 25138 2582 25144 2782
rect 25469 2594 25503 2897
rect 25227 2582 25273 2594
rect 25138 2406 25233 2582
rect 25267 2406 25273 2582
rect 25098 2394 25144 2406
rect 25227 2394 25273 2406
rect 25345 2582 25391 2594
rect 25345 2406 25351 2582
rect 25385 2406 25391 2582
rect 25345 2394 25391 2406
rect 25463 2582 25509 2594
rect 25463 2406 25469 2582
rect 25503 2406 25509 2582
rect 25463 2394 25509 2406
rect 25581 2582 25627 2594
rect 25581 2406 25587 2582
rect 25621 2406 25627 2582
rect 25581 2394 25627 2406
rect 21271 2316 21379 2326
rect 22014 2360 22048 2394
rect 22616 2360 22650 2394
rect 22852 2360 22886 2394
rect 22014 2325 22173 2360
rect 22616 2325 22886 2360
rect 23453 2360 23487 2394
rect 23689 2360 23723 2394
rect 23453 2325 23723 2360
rect 23912 2360 23946 2394
rect 24514 2360 24548 2394
rect 24750 2360 24784 2394
rect 23912 2325 24071 2360
rect 24514 2325 24784 2360
rect 25351 2360 25385 2394
rect 25587 2360 25621 2394
rect 25351 2325 25621 2360
rect 20644 2284 20659 2286
rect 20559 2270 20659 2284
rect 20559 2227 20659 2228
rect 20180 2206 20659 2227
rect 20948 2206 21014 2302
rect 20180 2158 21014 2206
rect 20180 2129 20659 2158
rect 20180 2127 20285 2129
rect 20559 2128 20659 2129
rect 20013 1942 20023 2021
rect 20116 1942 20126 2021
rect 19138 1680 19294 1686
rect 19138 1582 19150 1680
rect 19282 1582 19294 1680
rect 19138 1576 19294 1582
rect 20024 768 20117 1942
rect 20942 1893 21162 1913
rect 20942 1785 20986 1893
rect 21118 1785 21162 1893
rect 20942 1743 21162 1785
rect 20546 1713 21523 1743
rect 20546 1607 20578 1713
rect 20782 1607 20814 1713
rect 21018 1607 21050 1713
rect 21254 1607 21286 1713
rect 21489 1607 21523 1713
rect 20539 1595 20585 1607
rect 20539 1419 20545 1595
rect 20579 1419 20585 1595
rect 20539 1407 20585 1419
rect 20657 1595 20703 1607
rect 20657 1419 20663 1595
rect 20697 1419 20703 1595
rect 20657 1407 20703 1419
rect 20775 1595 20821 1607
rect 20775 1419 20781 1595
rect 20815 1419 20821 1595
rect 20775 1407 20821 1419
rect 20893 1595 20939 1607
rect 20893 1419 20899 1595
rect 20933 1419 20939 1595
rect 20893 1407 20939 1419
rect 21011 1595 21057 1607
rect 21011 1419 21017 1595
rect 21051 1419 21057 1595
rect 21011 1407 21057 1419
rect 21129 1595 21175 1607
rect 21129 1419 21135 1595
rect 21169 1419 21175 1595
rect 21129 1407 21175 1419
rect 21247 1595 21293 1607
rect 21247 1419 21253 1595
rect 21287 1419 21293 1595
rect 21247 1407 21293 1419
rect 21365 1595 21411 1607
rect 21365 1419 21371 1595
rect 21405 1419 21411 1595
rect 21365 1407 21411 1419
rect 21483 1595 21529 1607
rect 21483 1419 21489 1595
rect 21523 1419 21529 1595
rect 21483 1407 21529 1419
rect 21601 1595 21647 1607
rect 21601 1419 21607 1595
rect 21641 1419 21647 1595
rect 21601 1407 21647 1419
rect 22139 1541 22173 2325
rect 22852 2263 22886 2325
rect 22441 2225 23183 2263
rect 22441 2101 22475 2225
rect 22677 2101 22711 2225
rect 22913 2101 22947 2225
rect 23149 2101 23183 2225
rect 23439 2118 23449 2184
rect 23512 2118 23522 2184
rect 22435 2089 22481 2101
rect 22435 1713 22441 2089
rect 22475 1713 22481 2089
rect 22435 1701 22481 1713
rect 22553 2089 22599 2101
rect 22553 1713 22559 2089
rect 22593 1713 22599 2089
rect 22553 1701 22599 1713
rect 22671 2089 22717 2101
rect 22671 1713 22677 2089
rect 22711 1713 22717 2089
rect 22671 1701 22717 1713
rect 22789 2089 22835 2101
rect 22789 1713 22795 2089
rect 22829 1713 22835 2089
rect 22789 1701 22835 1713
rect 22907 2089 22953 2101
rect 22907 1713 22913 2089
rect 22947 1713 22953 2089
rect 22907 1701 22953 1713
rect 23025 2089 23071 2101
rect 23025 1713 23031 2089
rect 23065 1713 23071 2089
rect 23025 1701 23071 1713
rect 23143 2089 23189 2101
rect 23143 1713 23149 2089
rect 23183 1713 23189 2089
rect 23143 1701 23189 1713
rect 23555 1542 23589 2325
rect 23282 1541 23589 1542
rect 22139 1536 22455 1541
rect 23169 1536 23589 1541
rect 22139 1525 22522 1536
rect 22139 1498 22471 1525
rect 20662 1313 20698 1407
rect 20898 1313 20934 1407
rect 21134 1314 21170 1407
rect 21296 1359 21362 1366
rect 21296 1325 21312 1359
rect 21346 1325 21362 1359
rect 21296 1314 21362 1325
rect 21134 1313 21362 1314
rect 20662 1284 21362 1313
rect 20662 1283 21244 1284
rect 20782 1170 20816 1283
rect 21178 1242 21244 1283
rect 21178 1208 21194 1242
rect 21228 1208 21244 1242
rect 21178 1201 21244 1208
rect 21606 1174 21641 1407
rect 22139 1369 22173 1498
rect 22455 1491 22471 1498
rect 22505 1491 22522 1525
rect 22455 1485 22522 1491
rect 23102 1525 23589 1536
rect 23102 1491 23119 1525
rect 23153 1498 23589 1525
rect 23153 1491 23169 1498
rect 23282 1497 23589 1498
rect 23102 1485 23169 1491
rect 22280 1458 22336 1470
rect 22280 1424 22286 1458
rect 22320 1457 22336 1458
rect 23393 1457 23449 1469
rect 22320 1441 22787 1457
rect 22320 1424 22737 1441
rect 22280 1408 22737 1424
rect 22721 1407 22737 1408
rect 22771 1407 22787 1441
rect 22721 1400 22787 1407
rect 22839 1442 23409 1457
rect 22839 1408 22855 1442
rect 22889 1423 23409 1442
rect 23443 1423 23449 1457
rect 22889 1408 23449 1423
rect 22839 1398 22906 1408
rect 23393 1407 23449 1408
rect 23555 1369 23589 1497
rect 24037 1541 24071 2325
rect 24750 2263 24784 2325
rect 24339 2225 25081 2263
rect 24339 2101 24373 2225
rect 24575 2101 24609 2225
rect 24811 2101 24845 2225
rect 25047 2101 25081 2225
rect 24333 2089 24379 2101
rect 24333 1713 24339 2089
rect 24373 1713 24379 2089
rect 24333 1701 24379 1713
rect 24451 2089 24497 2101
rect 24451 1713 24457 2089
rect 24491 1713 24497 2089
rect 24451 1701 24497 1713
rect 24569 2089 24615 2101
rect 24569 1713 24575 2089
rect 24609 1713 24615 2089
rect 24569 1701 24615 1713
rect 24687 2089 24733 2101
rect 24687 1713 24693 2089
rect 24727 1713 24733 2089
rect 24687 1701 24733 1713
rect 24805 2089 24851 2101
rect 24805 1713 24811 2089
rect 24845 1713 24851 2089
rect 24805 1701 24851 1713
rect 24923 2089 24969 2101
rect 24923 1713 24929 2089
rect 24963 1713 24969 2089
rect 24923 1701 24969 1713
rect 25041 2089 25087 2101
rect 25041 1713 25047 2089
rect 25081 1713 25087 2089
rect 25041 1701 25087 1713
rect 25453 1542 25487 2325
rect 25065 1541 25134 1542
rect 25180 1541 25487 1542
rect 24037 1536 24353 1541
rect 25065 1537 25487 1541
rect 24037 1525 24420 1536
rect 24037 1498 24369 1525
rect 24037 1369 24071 1498
rect 24353 1491 24369 1498
rect 24403 1491 24420 1525
rect 24353 1485 24420 1491
rect 24998 1526 25487 1537
rect 24998 1492 25015 1526
rect 25049 1498 25487 1526
rect 25049 1492 25065 1498
rect 25180 1497 25487 1498
rect 24998 1486 25065 1492
rect 24178 1458 24234 1470
rect 24178 1424 24184 1458
rect 24218 1457 24234 1458
rect 25291 1457 25347 1469
rect 24218 1441 24685 1457
rect 24218 1424 24635 1441
rect 24178 1408 24635 1424
rect 24619 1407 24635 1408
rect 24669 1407 24685 1441
rect 24619 1400 24685 1407
rect 24737 1442 25307 1457
rect 24737 1408 24753 1442
rect 24787 1423 25307 1442
rect 25341 1423 25347 1457
rect 24787 1408 25347 1423
rect 24737 1398 24804 1408
rect 25291 1407 25347 1408
rect 25453 1369 25487 1497
rect 25568 2147 25635 2171
rect 25568 2113 25585 2147
rect 25619 2113 25635 2147
rect 21252 1170 21641 1174
rect 20776 1158 20822 1170
rect 20776 782 20782 1158
rect 20816 782 20822 1158
rect 20776 770 20822 782
rect 20894 1158 20940 1170
rect 20894 782 20900 1158
rect 20934 782 20940 1158
rect 20894 770 20940 782
rect 21012 1158 21058 1170
rect 21012 782 21018 1158
rect 21052 806 21058 1158
rect 21129 1158 21175 1170
rect 21129 982 21135 1158
rect 21169 982 21175 1158
rect 21129 970 21175 982
rect 21247 1158 21641 1170
rect 22133 1357 22179 1369
rect 22133 1181 22139 1357
rect 22173 1181 22179 1357
rect 22133 1169 22179 1181
rect 22251 1357 22297 1369
rect 22251 1181 22257 1357
rect 22291 1181 22297 1357
rect 22251 1169 22297 1181
rect 22553 1357 22599 1369
rect 21247 982 21253 1158
rect 21287 1145 21641 1158
rect 21287 982 21293 1145
rect 21563 1142 21641 1145
rect 21563 1090 21573 1142
rect 21636 1090 21646 1142
rect 21568 1084 21641 1090
rect 21247 970 21293 982
rect 21135 854 21170 970
rect 22256 875 22290 1169
rect 22553 981 22559 1357
rect 22593 981 22599 1357
rect 22553 969 22599 981
rect 22671 1357 22717 1369
rect 22671 981 22677 1357
rect 22711 981 22717 1357
rect 22671 969 22717 981
rect 22789 1357 22835 1369
rect 22789 981 22795 1357
rect 22829 981 22835 1357
rect 22789 969 22835 981
rect 22907 1357 22953 1369
rect 22907 981 22913 1357
rect 22947 981 22953 1357
rect 22907 969 22953 981
rect 23025 1357 23071 1369
rect 23025 981 23031 1357
rect 23065 981 23071 1357
rect 23431 1357 23477 1369
rect 23431 1181 23437 1357
rect 23471 1181 23477 1357
rect 23431 1169 23477 1181
rect 23549 1357 23595 1369
rect 23549 1181 23555 1357
rect 23589 1181 23595 1357
rect 23549 1169 23595 1181
rect 24031 1357 24077 1369
rect 24031 1181 24037 1357
rect 24071 1181 24077 1357
rect 24031 1169 24077 1181
rect 24149 1357 24195 1369
rect 24149 1181 24155 1357
rect 24189 1181 24195 1357
rect 24149 1169 24195 1181
rect 24451 1357 24497 1369
rect 23025 969 23071 981
rect 22913 875 22947 969
rect 23437 875 23470 1169
rect 21266 854 21374 864
rect 21135 806 21266 854
rect 21052 782 21266 806
rect 21012 770 21266 782
rect 20024 766 20609 768
rect 21018 766 21266 770
rect 20024 738 20654 766
rect 20024 732 20891 738
rect 14082 550 14451 598
rect 14082 520 14096 550
rect 14082 503 14092 520
rect 7848 372 12542 452
rect 14384 447 14450 550
rect 19010 447 19076 726
rect 20024 698 20841 732
rect 20875 698 20891 732
rect 20024 682 20891 698
rect 20943 732 21009 738
rect 20943 698 20959 732
rect 20993 698 21009 732
rect 21192 722 21266 766
rect 22256 843 23470 875
rect 24154 875 24188 1169
rect 24451 981 24457 1357
rect 24491 981 24497 1357
rect 24451 969 24497 981
rect 24569 1357 24615 1369
rect 24569 981 24575 1357
rect 24609 981 24615 1357
rect 24569 969 24615 981
rect 24687 1357 24733 1369
rect 24687 981 24693 1357
rect 24727 981 24733 1357
rect 24687 969 24733 981
rect 24805 1357 24851 1369
rect 24805 981 24811 1357
rect 24845 981 24851 1357
rect 24805 969 24851 981
rect 24923 1357 24969 1369
rect 24923 981 24929 1357
rect 24963 981 24969 1357
rect 25329 1357 25375 1369
rect 25329 1181 25335 1357
rect 25369 1181 25375 1357
rect 25329 1169 25375 1181
rect 25447 1357 25493 1369
rect 25447 1181 25453 1357
rect 25487 1181 25493 1357
rect 25447 1169 25493 1181
rect 24923 969 24969 981
rect 24811 875 24845 969
rect 25335 875 25368 1169
rect 24154 843 25368 875
rect 22749 758 22881 843
rect 24647 758 24779 843
rect 21266 712 21374 722
rect 20024 666 20654 682
rect 20024 662 20609 666
rect 20024 661 20125 662
rect 20554 613 20654 624
rect 20518 507 20528 613
rect 20640 602 20654 613
rect 20943 602 21009 698
rect 22739 650 22749 758
rect 22881 650 22891 758
rect 24637 650 24647 758
rect 24779 650 24789 758
rect 25568 730 25635 2113
rect 25696 1684 25852 1690
rect 25696 1586 25708 1684
rect 25840 1586 25852 1684
rect 25696 1580 25852 1586
rect 20640 554 21009 602
rect 20640 524 20654 554
rect 20640 507 20650 524
rect 20942 451 21008 554
rect 25568 451 25634 730
rect 14382 367 19076 447
rect 20940 371 25634 451
rect 939 -466 949 -403
rect 937 -477 949 -466
rect 936 -511 949 -477
rect 1081 -511 1091 -403
rect 2086 -466 2096 -403
rect 2084 -477 2096 -466
rect 1771 -487 1827 -485
rect 936 -549 1081 -511
rect 936 -577 977 -549
rect 1761 -553 1771 -487
rect 1827 -553 1837 -487
rect 2083 -511 2096 -477
rect 2228 -511 2238 -403
rect 4534 -457 4754 -437
rect 2901 -499 2957 -491
rect 2901 -507 3883 -499
rect 2083 -549 2228 -511
rect 2901 -541 2907 -507
rect 2941 -541 3883 -507
rect 936 -605 1212 -577
rect 936 -667 976 -605
rect 1178 -667 1212 -605
rect 1296 -605 1566 -577
rect 2083 -581 2124 -549
rect 2901 -557 3883 -541
rect 2904 -558 3883 -557
rect 1296 -667 1330 -605
rect 1532 -667 1566 -605
rect 1771 -621 1942 -605
rect 1771 -655 1777 -621
rect 1811 -655 1942 -621
rect 936 -679 982 -667
rect 936 -1055 942 -679
rect 976 -1055 982 -679
rect 936 -1067 982 -1055
rect 1054 -679 1100 -667
rect 1054 -1055 1060 -679
rect 1094 -1055 1100 -679
rect 1054 -1067 1100 -1055
rect 1172 -679 1218 -667
rect 1172 -1055 1178 -679
rect 1212 -1055 1218 -679
rect 1172 -1067 1218 -1055
rect 1290 -679 1336 -667
rect 1290 -1055 1296 -679
rect 1330 -1055 1336 -679
rect 1290 -1067 1336 -1055
rect 1408 -679 1454 -667
rect 1408 -1055 1414 -679
rect 1448 -1055 1454 -679
rect 1408 -1067 1454 -1055
rect 1526 -679 1572 -667
rect 1526 -1055 1532 -679
rect 1566 -1055 1572 -679
rect 1526 -1067 1572 -1055
rect 1644 -679 1690 -667
rect 1771 -671 1942 -655
rect 2083 -609 2354 -581
rect 2083 -671 2118 -609
rect 2320 -671 2354 -609
rect 2438 -609 2708 -581
rect 2438 -671 2472 -609
rect 2674 -671 2708 -609
rect 1644 -1055 1650 -679
rect 1684 -1055 1690 -679
rect 1644 -1067 1690 -1055
rect -128 -1311 -28 -1236
rect 40 -1311 50 -1236
rect 942 -1250 976 -1067
rect 1060 -1108 1094 -1067
rect 1296 -1108 1330 -1067
rect 1060 -1137 1330 -1108
rect 1414 -1109 1448 -1067
rect 1650 -1109 1684 -1067
rect 1414 -1137 1684 -1109
rect 1650 -1185 1684 -1137
rect 1621 -1215 1684 -1185
rect 867 -1304 976 -1250
rect 1049 -1245 1149 -1224
rect 1049 -1299 1070 -1245
rect 1135 -1299 1149 -1245
rect 1049 -1304 1149 -1299
rect -128 -1312 23 -1311
rect 867 -1450 901 -1304
rect 1051 -1319 1148 -1304
rect 1621 -1307 1656 -1215
rect 1091 -1386 1148 -1319
rect 1429 -1343 1656 -1307
rect 1429 -1377 1495 -1343
rect 985 -1422 1254 -1386
rect 1429 -1411 1445 -1377
rect 1479 -1411 1495 -1377
rect 1429 -1417 1495 -1411
rect 985 -1450 1018 -1422
rect 1221 -1450 1254 -1422
rect 1621 -1450 1656 -1343
rect 861 -1462 907 -1450
rect 861 -1638 867 -1462
rect 901 -1638 907 -1462
rect 861 -1650 907 -1638
rect 979 -1462 1025 -1450
rect 979 -1638 985 -1462
rect 1019 -1638 1025 -1462
rect 979 -1650 1025 -1638
rect 1097 -1462 1143 -1450
rect 1097 -1638 1103 -1462
rect 1137 -1638 1143 -1462
rect 1097 -1650 1143 -1638
rect 1215 -1462 1261 -1450
rect 1215 -1638 1221 -1462
rect 1255 -1517 1261 -1462
rect 1380 -1462 1426 -1450
rect 1380 -1517 1386 -1462
rect 1255 -1605 1386 -1517
rect 1255 -1638 1261 -1605
rect 1215 -1650 1261 -1638
rect 1380 -1638 1386 -1605
rect 1420 -1638 1426 -1462
rect 1380 -1650 1426 -1638
rect 1498 -1462 1544 -1450
rect 1498 -1638 1504 -1462
rect 1538 -1638 1544 -1462
rect 1498 -1650 1544 -1638
rect 1616 -1462 1662 -1450
rect 1616 -1638 1622 -1462
rect 1656 -1638 1662 -1462
rect 1616 -1650 1662 -1638
rect 1734 -1462 1780 -1450
rect 1734 -1638 1740 -1462
rect 1774 -1638 1780 -1462
rect 1734 -1650 1780 -1638
rect 868 -1688 901 -1650
rect 1104 -1688 1137 -1650
rect 868 -1724 1137 -1688
rect 1504 -1689 1538 -1650
rect 1740 -1689 1774 -1650
rect 1504 -1725 1774 -1689
rect 1608 -1726 1774 -1725
rect 1608 -1805 1740 -1726
rect 1598 -1913 1608 -1805
rect 1740 -1913 1750 -1805
rect 1880 -2242 1942 -671
rect 2078 -683 2124 -671
rect 2078 -1059 2084 -683
rect 2118 -1059 2124 -683
rect 2078 -1071 2124 -1059
rect 2196 -683 2242 -671
rect 2196 -1059 2202 -683
rect 2236 -1059 2242 -683
rect 2196 -1071 2242 -1059
rect 2314 -683 2360 -671
rect 2314 -1059 2320 -683
rect 2354 -1059 2360 -683
rect 2314 -1071 2360 -1059
rect 2432 -683 2478 -671
rect 2432 -1059 2438 -683
rect 2472 -1059 2478 -683
rect 2432 -1071 2478 -1059
rect 2550 -683 2596 -671
rect 2550 -1059 2556 -683
rect 2590 -1059 2596 -683
rect 2550 -1071 2596 -1059
rect 2668 -683 2714 -671
rect 2668 -1059 2674 -683
rect 2708 -1059 2714 -683
rect 2668 -1071 2714 -1059
rect 2786 -683 2832 -671
rect 2881 -675 2891 -609
rect 2957 -675 2967 -609
rect 2786 -1059 2792 -683
rect 2826 -1059 2832 -683
rect 2786 -1071 2832 -1059
rect 2084 -1254 2118 -1071
rect 2202 -1112 2236 -1071
rect 2438 -1112 2472 -1071
rect 2202 -1141 2472 -1112
rect 2556 -1113 2590 -1071
rect 2792 -1113 2826 -1071
rect 2556 -1141 2826 -1113
rect 2792 -1189 2826 -1141
rect 2763 -1219 2826 -1189
rect 3816 -1148 3883 -558
rect 4534 -565 4578 -457
rect 4710 -565 4754 -457
rect 7497 -470 7507 -407
rect 7495 -481 7507 -470
rect 4534 -607 4754 -565
rect 7494 -515 7507 -481
rect 7639 -515 7649 -407
rect 8644 -470 8654 -407
rect 8642 -481 8654 -470
rect 8329 -491 8385 -489
rect 7494 -553 7639 -515
rect 7494 -581 7535 -553
rect 8319 -557 8329 -491
rect 8385 -557 8395 -491
rect 8641 -515 8654 -481
rect 8786 -515 8796 -407
rect 11092 -461 11312 -441
rect 9459 -503 9515 -495
rect 9459 -511 10441 -503
rect 8641 -553 8786 -515
rect 9459 -545 9465 -511
rect 9499 -545 10441 -511
rect 4173 -637 5150 -607
rect 4173 -743 4207 -637
rect 4410 -743 4442 -637
rect 4646 -743 4678 -637
rect 4882 -743 4914 -637
rect 5118 -743 5150 -637
rect 7494 -609 7770 -581
rect 7494 -671 7534 -609
rect 7736 -671 7770 -609
rect 7854 -609 8124 -581
rect 8641 -585 8682 -553
rect 9459 -561 10441 -545
rect 9462 -562 10441 -561
rect 7854 -671 7888 -609
rect 8090 -671 8124 -609
rect 8329 -625 8500 -609
rect 8329 -659 8335 -625
rect 8369 -659 8500 -625
rect 7494 -683 7540 -671
rect 4049 -755 4095 -743
rect 4049 -931 4055 -755
rect 4089 -931 4095 -755
rect 4049 -943 4095 -931
rect 4167 -755 4213 -743
rect 4167 -931 4173 -755
rect 4207 -931 4213 -755
rect 4167 -943 4213 -931
rect 4285 -755 4331 -743
rect 4285 -931 4291 -755
rect 4325 -931 4331 -755
rect 4285 -943 4331 -931
rect 4403 -755 4449 -743
rect 4403 -931 4409 -755
rect 4443 -931 4449 -755
rect 4403 -943 4449 -931
rect 4521 -755 4567 -743
rect 4521 -931 4527 -755
rect 4561 -931 4567 -755
rect 4521 -943 4567 -931
rect 4639 -755 4685 -743
rect 4639 -931 4645 -755
rect 4679 -931 4685 -755
rect 4639 -943 4685 -931
rect 4757 -755 4803 -743
rect 4757 -931 4763 -755
rect 4797 -931 4803 -755
rect 4757 -943 4803 -931
rect 4875 -755 4921 -743
rect 4875 -931 4881 -755
rect 4915 -931 4921 -755
rect 4875 -943 4921 -931
rect 4993 -755 5039 -743
rect 4993 -931 4999 -755
rect 5033 -931 5039 -755
rect 4993 -943 5039 -931
rect 5111 -755 5157 -743
rect 5111 -931 5117 -755
rect 5151 -931 5157 -755
rect 5111 -943 5157 -931
rect 4055 -1148 4090 -943
rect 4334 -991 4400 -984
rect 4334 -1025 4350 -991
rect 4384 -1025 4400 -991
rect 4334 -1036 4400 -1025
rect 4526 -1036 4562 -943
rect 4334 -1037 4562 -1036
rect 4762 -1037 4798 -943
rect 4998 -1037 5034 -943
rect 4334 -1066 5034 -1037
rect 3816 -1176 4090 -1148
rect 4452 -1067 5034 -1066
rect 7494 -1059 7500 -683
rect 7534 -1059 7540 -683
rect 4452 -1108 4518 -1067
rect 4452 -1142 4468 -1108
rect 4502 -1142 4518 -1108
rect 4452 -1149 4518 -1142
rect 3816 -1180 4444 -1176
rect 4880 -1180 4914 -1067
rect 7494 -1071 7540 -1059
rect 7612 -683 7658 -671
rect 7612 -1059 7618 -683
rect 7652 -1059 7658 -683
rect 7612 -1071 7658 -1059
rect 7730 -683 7776 -671
rect 7730 -1059 7736 -683
rect 7770 -1059 7776 -683
rect 7730 -1071 7776 -1059
rect 7848 -683 7894 -671
rect 7848 -1059 7854 -683
rect 7888 -1059 7894 -683
rect 7848 -1071 7894 -1059
rect 7966 -683 8012 -671
rect 7966 -1059 7972 -683
rect 8006 -1059 8012 -683
rect 7966 -1071 8012 -1059
rect 8084 -683 8130 -671
rect 8084 -1059 8090 -683
rect 8124 -1059 8130 -683
rect 8084 -1071 8130 -1059
rect 8202 -683 8248 -671
rect 8329 -675 8500 -659
rect 8641 -613 8912 -585
rect 8641 -675 8676 -613
rect 8878 -675 8912 -613
rect 8996 -613 9266 -585
rect 8996 -675 9030 -613
rect 9232 -675 9266 -613
rect 8202 -1059 8208 -683
rect 8242 -1059 8248 -683
rect 8202 -1071 8248 -1059
rect 3816 -1192 4449 -1180
rect 3816 -1205 4409 -1192
rect 2009 -1308 2118 -1254
rect 2009 -1454 2043 -1308
rect 2182 -1322 2192 -1225
rect 2291 -1322 2301 -1225
rect 2763 -1311 2798 -1219
rect 2193 -1323 2290 -1322
rect 2233 -1390 2290 -1323
rect 2571 -1347 2798 -1311
rect 2571 -1381 2637 -1347
rect 2127 -1426 2396 -1390
rect 2571 -1415 2587 -1381
rect 2621 -1415 2637 -1381
rect 2571 -1421 2637 -1415
rect 2127 -1454 2160 -1426
rect 2363 -1454 2396 -1426
rect 2763 -1454 2798 -1347
rect 4403 -1368 4409 -1205
rect 4443 -1368 4449 -1192
rect 4403 -1380 4449 -1368
rect 4521 -1192 4567 -1180
rect 4521 -1368 4527 -1192
rect 4561 -1368 4567 -1192
rect 4521 -1380 4567 -1368
rect 4638 -1192 4684 -1180
rect 2003 -1466 2049 -1454
rect 2003 -1642 2009 -1466
rect 2043 -1642 2049 -1466
rect 2003 -1654 2049 -1642
rect 2121 -1466 2167 -1454
rect 2121 -1642 2127 -1466
rect 2161 -1642 2167 -1466
rect 2121 -1654 2167 -1642
rect 2239 -1466 2285 -1454
rect 2239 -1642 2245 -1466
rect 2279 -1642 2285 -1466
rect 2239 -1654 2285 -1642
rect 2357 -1466 2403 -1454
rect 2357 -1642 2363 -1466
rect 2397 -1521 2403 -1466
rect 2522 -1466 2568 -1454
rect 2522 -1521 2528 -1466
rect 2397 -1609 2528 -1521
rect 2397 -1642 2403 -1609
rect 2357 -1654 2403 -1642
rect 2522 -1642 2528 -1609
rect 2562 -1642 2568 -1466
rect 2522 -1654 2568 -1642
rect 2640 -1466 2686 -1454
rect 2640 -1642 2646 -1466
rect 2680 -1642 2686 -1466
rect 2640 -1654 2686 -1642
rect 2758 -1466 2804 -1454
rect 2758 -1642 2764 -1466
rect 2798 -1642 2804 -1466
rect 2758 -1654 2804 -1642
rect 2876 -1466 2922 -1454
rect 2876 -1642 2882 -1466
rect 2916 -1642 2922 -1466
rect 4322 -1496 4430 -1486
rect 4526 -1496 4561 -1380
rect 4430 -1544 4561 -1496
rect 4638 -1544 4644 -1192
rect 4430 -1568 4644 -1544
rect 4678 -1568 4684 -1192
rect 4430 -1580 4684 -1568
rect 4756 -1192 4802 -1180
rect 4756 -1568 4762 -1192
rect 4796 -1568 4802 -1192
rect 4756 -1580 4802 -1568
rect 4874 -1192 4920 -1180
rect 4874 -1568 4880 -1192
rect 4914 -1568 4920 -1192
rect 6430 -1240 6529 -1238
rect 6430 -1315 6530 -1240
rect 6598 -1315 6608 -1240
rect 7500 -1254 7534 -1071
rect 7618 -1112 7652 -1071
rect 7854 -1112 7888 -1071
rect 7618 -1141 7888 -1112
rect 7972 -1113 8006 -1071
rect 8208 -1113 8242 -1071
rect 7972 -1141 8242 -1113
rect 8208 -1189 8242 -1141
rect 8179 -1219 8242 -1189
rect 7425 -1308 7534 -1254
rect 7607 -1249 7707 -1228
rect 7607 -1303 7628 -1249
rect 7693 -1303 7707 -1249
rect 7607 -1308 7707 -1303
rect 6430 -1316 6581 -1315
rect 4874 -1580 4920 -1568
rect 4430 -1584 4678 -1580
rect 4430 -1628 4504 -1584
rect 5803 -1585 6092 -1410
rect 5042 -1612 6092 -1585
rect 4687 -1618 4753 -1612
rect 4322 -1638 4430 -1628
rect 2876 -1654 2922 -1642
rect 4687 -1652 4703 -1618
rect 4737 -1652 4753 -1618
rect 2010 -1692 2043 -1654
rect 2246 -1692 2279 -1654
rect 2010 -1728 2279 -1692
rect 2646 -1693 2680 -1654
rect 2882 -1693 2916 -1654
rect 2646 -1728 2916 -1693
rect 2646 -1729 2882 -1728
rect 2750 -1803 2882 -1729
rect 4687 -1748 4753 -1652
rect 4805 -1618 6092 -1612
rect 4805 -1652 4821 -1618
rect 4855 -1652 6092 -1618
rect 4805 -1668 6092 -1652
rect 5042 -1684 6092 -1668
rect 5105 -1685 6092 -1684
rect 5570 -1689 6092 -1685
rect 5041 -1748 5507 -1726
rect 4687 -1796 5507 -1748
rect 2740 -1911 2750 -1803
rect 2882 -1911 2892 -1803
rect 5041 -1827 5507 -1796
rect 5402 -2083 5507 -1827
rect 1879 -2259 1942 -2242
rect 4520 -2107 4740 -2087
rect 4520 -2215 4564 -2107
rect 4696 -2215 4740 -2107
rect 5322 -2189 5332 -2083
rect 5444 -2189 5507 -2083
rect 5358 -2200 5507 -2189
rect 4520 -2257 4740 -2215
rect 1879 -2263 2017 -2259
rect 1879 -2297 3849 -2263
rect 4159 -2287 5136 -2257
rect 1879 -2326 3851 -2297
rect 1879 -2328 2017 -2326
rect 3805 -2342 3851 -2326
rect 843 -2558 853 -2450
rect 985 -2558 995 -2450
rect 2741 -2558 2751 -2450
rect 2883 -2558 2893 -2450
rect 853 -2598 985 -2558
rect 2751 -2598 2883 -2558
rect 853 -2664 986 -2598
rect 2751 -2664 2884 -2598
rect 184 -2707 1657 -2664
rect 184 -3010 218 -2707
rect 549 -2810 583 -2707
rect 785 -2810 819 -2707
rect 1021 -2810 1055 -2707
rect 1257 -2810 1291 -2707
rect 543 -2822 589 -2810
rect 60 -3022 106 -3010
rect 60 -3198 66 -3022
rect 100 -3198 106 -3022
rect 60 -3210 106 -3198
rect 178 -3022 224 -3010
rect 178 -3198 184 -3022
rect 218 -3198 224 -3022
rect 178 -3210 224 -3198
rect 296 -3022 342 -3010
rect 296 -3198 302 -3022
rect 336 -3198 342 -3022
rect 296 -3210 342 -3198
rect 414 -3022 460 -3010
rect 543 -3022 549 -2822
rect 414 -3198 420 -3022
rect 454 -3198 549 -3022
rect 583 -3198 589 -2822
rect 414 -3210 460 -3198
rect 543 -3210 589 -3198
rect 661 -2822 707 -2810
rect 661 -3198 667 -2822
rect 701 -3198 707 -2822
rect 661 -3210 707 -3198
rect 779 -2822 825 -2810
rect 779 -3198 785 -2822
rect 819 -3198 825 -2822
rect 779 -3210 825 -3198
rect 897 -2822 943 -2810
rect 897 -3198 903 -2822
rect 937 -3198 943 -2822
rect 897 -3210 943 -3198
rect 1015 -2822 1061 -2810
rect 1015 -3198 1021 -2822
rect 1055 -3198 1061 -2822
rect 1015 -3210 1061 -3198
rect 1133 -2822 1179 -2810
rect 1133 -3198 1139 -2822
rect 1173 -3198 1179 -2822
rect 1133 -3210 1179 -3198
rect 1251 -2822 1297 -2810
rect 1251 -3198 1257 -2822
rect 1291 -3022 1297 -2822
rect 1623 -3010 1657 -2707
rect 2082 -2707 3555 -2664
rect 2082 -3010 2116 -2707
rect 2447 -2810 2481 -2707
rect 2683 -2810 2717 -2707
rect 2919 -2810 2953 -2707
rect 3155 -2810 3189 -2707
rect 2441 -2822 2487 -2810
rect 1381 -3022 1427 -3010
rect 1291 -3198 1387 -3022
rect 1421 -3198 1427 -3022
rect 1251 -3210 1297 -3198
rect 1381 -3210 1427 -3198
rect 1499 -3022 1545 -3010
rect 1499 -3198 1505 -3022
rect 1539 -3198 1545 -3022
rect 1499 -3210 1545 -3198
rect 1617 -3022 1663 -3010
rect 1617 -3198 1623 -3022
rect 1657 -3198 1663 -3022
rect 1617 -3210 1663 -3198
rect 1735 -3022 1781 -3010
rect 1735 -3198 1741 -3022
rect 1775 -3198 1781 -3022
rect 1735 -3210 1781 -3198
rect 1958 -3022 2004 -3010
rect 1958 -3198 1964 -3022
rect 1998 -3198 2004 -3022
rect 1958 -3210 2004 -3198
rect 2076 -3022 2122 -3010
rect 2076 -3198 2082 -3022
rect 2116 -3198 2122 -3022
rect 2076 -3210 2122 -3198
rect 2194 -3022 2240 -3010
rect 2194 -3198 2200 -3022
rect 2234 -3198 2240 -3022
rect 2194 -3210 2240 -3198
rect 2312 -3022 2358 -3010
rect 2441 -3022 2447 -2822
rect 2312 -3198 2318 -3022
rect 2352 -3198 2447 -3022
rect 2481 -3198 2487 -2822
rect 2312 -3210 2358 -3198
rect 2441 -3210 2487 -3198
rect 2559 -2822 2605 -2810
rect 2559 -3198 2565 -2822
rect 2599 -3198 2605 -2822
rect 2559 -3210 2605 -3198
rect 2677 -2822 2723 -2810
rect 2677 -3198 2683 -2822
rect 2717 -3198 2723 -2822
rect 2677 -3210 2723 -3198
rect 2795 -2822 2841 -2810
rect 2795 -3198 2801 -2822
rect 2835 -3198 2841 -2822
rect 2795 -3210 2841 -3198
rect 2913 -2822 2959 -2810
rect 2913 -3198 2919 -2822
rect 2953 -3198 2959 -2822
rect 2913 -3210 2959 -3198
rect 3031 -2822 3077 -2810
rect 3031 -3198 3037 -2822
rect 3071 -3198 3077 -2822
rect 3031 -3210 3077 -3198
rect 3149 -2822 3195 -2810
rect 3149 -3198 3155 -2822
rect 3189 -3022 3195 -2822
rect 3521 -3010 3555 -2707
rect 3805 -2794 3852 -2342
rect 4159 -2393 4193 -2287
rect 4396 -2393 4428 -2287
rect 4632 -2393 4664 -2287
rect 4868 -2393 4900 -2287
rect 5104 -2393 5136 -2287
rect 4035 -2405 4081 -2393
rect 4035 -2581 4041 -2405
rect 4075 -2581 4081 -2405
rect 4035 -2593 4081 -2581
rect 4153 -2405 4199 -2393
rect 4153 -2581 4159 -2405
rect 4193 -2581 4199 -2405
rect 4153 -2593 4199 -2581
rect 4271 -2405 4317 -2393
rect 4271 -2581 4277 -2405
rect 4311 -2581 4317 -2405
rect 4271 -2593 4317 -2581
rect 4389 -2405 4435 -2393
rect 4389 -2581 4395 -2405
rect 4429 -2581 4435 -2405
rect 4389 -2593 4435 -2581
rect 4507 -2405 4553 -2393
rect 4507 -2581 4513 -2405
rect 4547 -2581 4553 -2405
rect 4507 -2593 4553 -2581
rect 4625 -2405 4671 -2393
rect 4625 -2581 4631 -2405
rect 4665 -2581 4671 -2405
rect 4625 -2593 4671 -2581
rect 4743 -2405 4789 -2393
rect 4743 -2581 4749 -2405
rect 4783 -2581 4789 -2405
rect 4743 -2593 4789 -2581
rect 4861 -2405 4907 -2393
rect 4861 -2581 4867 -2405
rect 4901 -2581 4907 -2405
rect 4861 -2593 4907 -2581
rect 4979 -2405 5025 -2393
rect 4979 -2581 4985 -2405
rect 5019 -2581 5025 -2405
rect 4979 -2593 5025 -2581
rect 5097 -2405 5143 -2393
rect 5097 -2581 5103 -2405
rect 5137 -2581 5143 -2405
rect 5097 -2593 5143 -2581
rect 3806 -2810 3852 -2794
rect 3806 -2811 3887 -2810
rect 4041 -2811 4076 -2593
rect 4320 -2641 4386 -2634
rect 4320 -2675 4336 -2641
rect 4370 -2675 4386 -2641
rect 4320 -2686 4386 -2675
rect 4512 -2686 4548 -2593
rect 4320 -2687 4548 -2686
rect 4748 -2687 4784 -2593
rect 4984 -2687 5020 -2593
rect 4320 -2716 5020 -2687
rect 4438 -2717 5020 -2716
rect 4438 -2758 4504 -2717
rect 4438 -2792 4454 -2758
rect 4488 -2792 4504 -2758
rect 4438 -2799 4504 -2792
rect 3806 -2826 4076 -2811
rect 3806 -2830 4430 -2826
rect 4866 -2830 4900 -2717
rect 3806 -2842 4435 -2830
rect 3806 -2854 4395 -2842
rect 3806 -2856 3887 -2854
rect 4153 -2855 4395 -2854
rect 3279 -3022 3325 -3010
rect 3189 -3198 3285 -3022
rect 3319 -3198 3325 -3022
rect 3149 -3210 3195 -3198
rect 3279 -3210 3325 -3198
rect 3397 -3022 3443 -3010
rect 3397 -3198 3403 -3022
rect 3437 -3198 3443 -3022
rect 3397 -3210 3443 -3198
rect 3515 -3022 3561 -3010
rect 3515 -3198 3521 -3022
rect 3555 -3198 3561 -3022
rect 3515 -3210 3561 -3198
rect 3633 -3022 3679 -3010
rect 3633 -3198 3639 -3022
rect 3673 -3198 3679 -3022
rect 4389 -3018 4395 -2855
rect 4429 -3018 4435 -2842
rect 4389 -3030 4435 -3018
rect 4507 -2842 4553 -2830
rect 4507 -3018 4513 -2842
rect 4547 -3018 4553 -2842
rect 4507 -3030 4553 -3018
rect 4624 -2842 4670 -2830
rect 3633 -3210 3679 -3198
rect 4308 -3146 4416 -3136
rect 4512 -3146 4547 -3030
rect 66 -3244 100 -3210
rect 302 -3244 336 -3210
rect 66 -3279 336 -3244
rect 903 -3244 937 -3210
rect 1139 -3244 1173 -3210
rect 1741 -3244 1775 -3210
rect 903 -3279 1173 -3244
rect 1616 -3279 1775 -3244
rect 1964 -3244 1998 -3210
rect 2200 -3244 2234 -3210
rect 1964 -3279 2234 -3244
rect 2801 -3244 2835 -3210
rect 3037 -3244 3071 -3210
rect 3639 -3244 3673 -3210
rect 2801 -3279 3071 -3244
rect 3514 -3279 3673 -3244
rect 4416 -3194 4547 -3146
rect 4624 -3194 4630 -2842
rect 4416 -3218 4630 -3194
rect 4664 -3218 4670 -2842
rect 4416 -3230 4670 -3218
rect 4742 -2842 4788 -2830
rect 4742 -3218 4748 -2842
rect 4782 -3218 4788 -2842
rect 4742 -3230 4788 -3218
rect 4860 -2842 4906 -2830
rect 4860 -3218 4866 -2842
rect 4900 -3218 4906 -2842
rect 4860 -3230 4906 -3218
rect 4416 -3234 4664 -3230
rect 5033 -3234 5043 -3202
rect 4416 -3278 4490 -3234
rect 5028 -3262 5043 -3234
rect 4673 -3268 4739 -3262
rect 52 -3457 119 -3433
rect 52 -3491 68 -3457
rect 102 -3491 119 -3457
rect -165 -3920 -9 -3914
rect -165 -4018 -153 -3920
rect -21 -4018 -9 -3920
rect -165 -4024 -9 -4018
rect 52 -4874 119 -3491
rect 200 -4062 234 -3279
rect 903 -3341 937 -3279
rect 606 -3379 1348 -3341
rect 606 -3503 640 -3379
rect 842 -3503 876 -3379
rect 1078 -3503 1112 -3379
rect 1314 -3503 1348 -3379
rect 600 -3515 646 -3503
rect 600 -3891 606 -3515
rect 640 -3891 646 -3515
rect 600 -3903 646 -3891
rect 718 -3515 764 -3503
rect 718 -3891 724 -3515
rect 758 -3891 764 -3515
rect 718 -3903 764 -3891
rect 836 -3515 882 -3503
rect 836 -3891 842 -3515
rect 876 -3891 882 -3515
rect 836 -3903 882 -3891
rect 954 -3515 1000 -3503
rect 954 -3891 960 -3515
rect 994 -3891 1000 -3515
rect 954 -3903 1000 -3891
rect 1072 -3515 1118 -3503
rect 1072 -3891 1078 -3515
rect 1112 -3891 1118 -3515
rect 1072 -3903 1118 -3891
rect 1190 -3515 1236 -3503
rect 1190 -3891 1196 -3515
rect 1230 -3891 1236 -3515
rect 1190 -3903 1236 -3891
rect 1308 -3515 1354 -3503
rect 1308 -3891 1314 -3515
rect 1348 -3891 1354 -3515
rect 1308 -3903 1354 -3891
rect 200 -4063 507 -4062
rect 553 -4063 622 -4062
rect 1616 -4063 1650 -3279
rect 200 -4067 622 -4063
rect 200 -4078 689 -4067
rect 1334 -4068 1650 -4063
rect 200 -4106 638 -4078
rect 200 -4107 507 -4106
rect 200 -4235 234 -4107
rect 622 -4112 638 -4106
rect 672 -4112 689 -4078
rect 622 -4118 689 -4112
rect 1267 -4079 1650 -4068
rect 1267 -4113 1284 -4079
rect 1318 -4106 1650 -4079
rect 1318 -4113 1334 -4106
rect 1267 -4119 1334 -4113
rect 340 -4147 396 -4135
rect 1453 -4146 1509 -4134
rect 1453 -4147 1469 -4146
rect 340 -4181 346 -4147
rect 380 -4162 950 -4147
rect 380 -4181 900 -4162
rect 340 -4196 900 -4181
rect 934 -4196 950 -4162
rect 340 -4197 396 -4196
rect 883 -4206 950 -4196
rect 1002 -4163 1469 -4147
rect 1002 -4197 1018 -4163
rect 1052 -4180 1469 -4163
rect 1503 -4180 1509 -4146
rect 1052 -4196 1509 -4180
rect 1052 -4197 1068 -4196
rect 1002 -4204 1068 -4197
rect 1616 -4235 1650 -4106
rect 2098 -4062 2132 -3279
rect 2801 -3341 2835 -3279
rect 2504 -3379 3246 -3341
rect 2165 -3486 2175 -3420
rect 2238 -3486 2248 -3420
rect 2504 -3503 2538 -3379
rect 2740 -3503 2774 -3379
rect 2976 -3503 3010 -3379
rect 3212 -3503 3246 -3379
rect 2498 -3515 2544 -3503
rect 2498 -3891 2504 -3515
rect 2538 -3891 2544 -3515
rect 2498 -3903 2544 -3891
rect 2616 -3515 2662 -3503
rect 2616 -3891 2622 -3515
rect 2656 -3891 2662 -3515
rect 2616 -3903 2662 -3891
rect 2734 -3515 2780 -3503
rect 2734 -3891 2740 -3515
rect 2774 -3891 2780 -3515
rect 2734 -3903 2780 -3891
rect 2852 -3515 2898 -3503
rect 2852 -3891 2858 -3515
rect 2892 -3891 2898 -3515
rect 2852 -3903 2898 -3891
rect 2970 -3515 3016 -3503
rect 2970 -3891 2976 -3515
rect 3010 -3891 3016 -3515
rect 2970 -3903 3016 -3891
rect 3088 -3515 3134 -3503
rect 3088 -3891 3094 -3515
rect 3128 -3891 3134 -3515
rect 3088 -3903 3134 -3891
rect 3206 -3515 3252 -3503
rect 3206 -3891 3212 -3515
rect 3246 -3891 3252 -3515
rect 3206 -3903 3252 -3891
rect 2098 -4063 2405 -4062
rect 3514 -4063 3548 -3279
rect 4308 -3288 4416 -3278
rect 4673 -3302 4689 -3268
rect 4723 -3302 4739 -3268
rect 4673 -3398 4739 -3302
rect 4791 -3268 5043 -3262
rect 4791 -3302 4807 -3268
rect 4841 -3302 5043 -3268
rect 4791 -3318 5043 -3302
rect 5028 -3320 5043 -3318
rect 5161 -3320 5171 -3202
rect 5028 -3334 5128 -3320
rect 5028 -3377 5128 -3376
rect 5402 -3377 5507 -2200
rect 5028 -3398 5507 -3377
rect 4673 -3446 5507 -3398
rect 5028 -3475 5507 -3446
rect 5028 -3476 5128 -3475
rect 5402 -3477 5507 -3475
rect 5570 -3583 5663 -1689
rect 5803 -1690 6092 -1689
rect 5786 -2100 6075 -1938
rect 5786 -2113 5826 -2100
rect 5784 -2206 5826 -2113
rect 5938 -2206 6075 -2100
rect 5784 -2217 6075 -2206
rect 5786 -2218 6075 -2217
rect 6430 -3050 6529 -1316
rect 7425 -1454 7459 -1308
rect 7609 -1323 7706 -1308
rect 8179 -1311 8214 -1219
rect 7649 -1390 7706 -1323
rect 7987 -1347 8214 -1311
rect 7987 -1381 8053 -1347
rect 7543 -1426 7812 -1390
rect 7987 -1415 8003 -1381
rect 8037 -1415 8053 -1381
rect 7987 -1421 8053 -1415
rect 7543 -1454 7576 -1426
rect 7779 -1454 7812 -1426
rect 8179 -1454 8214 -1347
rect 7419 -1466 7465 -1454
rect 7419 -1642 7425 -1466
rect 7459 -1642 7465 -1466
rect 7419 -1654 7465 -1642
rect 7537 -1466 7583 -1454
rect 7537 -1642 7543 -1466
rect 7577 -1642 7583 -1466
rect 7537 -1654 7583 -1642
rect 7655 -1466 7701 -1454
rect 7655 -1642 7661 -1466
rect 7695 -1642 7701 -1466
rect 7655 -1654 7701 -1642
rect 7773 -1466 7819 -1454
rect 7773 -1642 7779 -1466
rect 7813 -1521 7819 -1466
rect 7938 -1466 7984 -1454
rect 7938 -1521 7944 -1466
rect 7813 -1609 7944 -1521
rect 7813 -1642 7819 -1609
rect 7773 -1654 7819 -1642
rect 7938 -1642 7944 -1609
rect 7978 -1642 7984 -1466
rect 7938 -1654 7984 -1642
rect 8056 -1466 8102 -1454
rect 8056 -1642 8062 -1466
rect 8096 -1642 8102 -1466
rect 8056 -1654 8102 -1642
rect 8174 -1466 8220 -1454
rect 8174 -1642 8180 -1466
rect 8214 -1642 8220 -1466
rect 8174 -1654 8220 -1642
rect 8292 -1466 8338 -1454
rect 8292 -1642 8298 -1466
rect 8332 -1642 8338 -1466
rect 8292 -1654 8338 -1642
rect 7426 -1692 7459 -1654
rect 7662 -1692 7695 -1654
rect 7426 -1728 7695 -1692
rect 8062 -1693 8096 -1654
rect 8298 -1693 8332 -1654
rect 8062 -1729 8332 -1693
rect 8166 -1730 8332 -1729
rect 8166 -1809 8298 -1730
rect 8156 -1917 8166 -1809
rect 8298 -1917 8308 -1809
rect 8438 -2246 8500 -675
rect 8636 -687 8682 -675
rect 8636 -1063 8642 -687
rect 8676 -1063 8682 -687
rect 8636 -1075 8682 -1063
rect 8754 -687 8800 -675
rect 8754 -1063 8760 -687
rect 8794 -1063 8800 -687
rect 8754 -1075 8800 -1063
rect 8872 -687 8918 -675
rect 8872 -1063 8878 -687
rect 8912 -1063 8918 -687
rect 8872 -1075 8918 -1063
rect 8990 -687 9036 -675
rect 8990 -1063 8996 -687
rect 9030 -1063 9036 -687
rect 8990 -1075 9036 -1063
rect 9108 -687 9154 -675
rect 9108 -1063 9114 -687
rect 9148 -1063 9154 -687
rect 9108 -1075 9154 -1063
rect 9226 -687 9272 -675
rect 9226 -1063 9232 -687
rect 9266 -1063 9272 -687
rect 9226 -1075 9272 -1063
rect 9344 -687 9390 -675
rect 9439 -679 9449 -613
rect 9515 -679 9525 -613
rect 9344 -1063 9350 -687
rect 9384 -1063 9390 -687
rect 9344 -1075 9390 -1063
rect 8642 -1258 8676 -1075
rect 8760 -1116 8794 -1075
rect 8996 -1116 9030 -1075
rect 8760 -1145 9030 -1116
rect 9114 -1117 9148 -1075
rect 9350 -1117 9384 -1075
rect 9114 -1145 9384 -1117
rect 9350 -1193 9384 -1145
rect 9321 -1223 9384 -1193
rect 10374 -1152 10441 -562
rect 11092 -569 11136 -461
rect 11268 -569 11312 -461
rect 14031 -465 14041 -402
rect 14029 -476 14041 -465
rect 11092 -611 11312 -569
rect 14028 -510 14041 -476
rect 14173 -510 14183 -402
rect 15178 -465 15188 -402
rect 15176 -476 15188 -465
rect 14863 -486 14919 -484
rect 14028 -548 14173 -510
rect 14028 -576 14069 -548
rect 14853 -552 14863 -486
rect 14919 -552 14929 -486
rect 15175 -510 15188 -476
rect 15320 -510 15330 -402
rect 17626 -456 17846 -436
rect 15993 -498 16049 -490
rect 15993 -506 16975 -498
rect 15175 -548 15320 -510
rect 15993 -540 15999 -506
rect 16033 -540 16975 -506
rect 14028 -604 14304 -576
rect 10731 -641 11708 -611
rect 10731 -747 10765 -641
rect 10968 -747 11000 -641
rect 11204 -747 11236 -641
rect 11440 -747 11472 -641
rect 11676 -747 11708 -641
rect 14028 -666 14068 -604
rect 14270 -666 14304 -604
rect 14388 -604 14658 -576
rect 15175 -580 15216 -548
rect 15993 -556 16975 -540
rect 15996 -557 16975 -556
rect 14388 -666 14422 -604
rect 14624 -666 14658 -604
rect 14863 -620 15034 -604
rect 14863 -654 14869 -620
rect 14903 -654 15034 -620
rect 14028 -678 14074 -666
rect 10607 -759 10653 -747
rect 10607 -935 10613 -759
rect 10647 -935 10653 -759
rect 10607 -947 10653 -935
rect 10725 -759 10771 -747
rect 10725 -935 10731 -759
rect 10765 -935 10771 -759
rect 10725 -947 10771 -935
rect 10843 -759 10889 -747
rect 10843 -935 10849 -759
rect 10883 -935 10889 -759
rect 10843 -947 10889 -935
rect 10961 -759 11007 -747
rect 10961 -935 10967 -759
rect 11001 -935 11007 -759
rect 10961 -947 11007 -935
rect 11079 -759 11125 -747
rect 11079 -935 11085 -759
rect 11119 -935 11125 -759
rect 11079 -947 11125 -935
rect 11197 -759 11243 -747
rect 11197 -935 11203 -759
rect 11237 -935 11243 -759
rect 11197 -947 11243 -935
rect 11315 -759 11361 -747
rect 11315 -935 11321 -759
rect 11355 -935 11361 -759
rect 11315 -947 11361 -935
rect 11433 -759 11479 -747
rect 11433 -935 11439 -759
rect 11473 -935 11479 -759
rect 11433 -947 11479 -935
rect 11551 -759 11597 -747
rect 11551 -935 11557 -759
rect 11591 -935 11597 -759
rect 11551 -947 11597 -935
rect 11669 -759 11715 -747
rect 11669 -935 11675 -759
rect 11709 -935 11715 -759
rect 11669 -947 11715 -935
rect 10613 -1152 10648 -947
rect 10892 -995 10958 -988
rect 10892 -1029 10908 -995
rect 10942 -1029 10958 -995
rect 10892 -1040 10958 -1029
rect 11084 -1040 11120 -947
rect 10892 -1041 11120 -1040
rect 11320 -1041 11356 -947
rect 11556 -1041 11592 -947
rect 10892 -1070 11592 -1041
rect 14028 -1054 14034 -678
rect 14068 -1054 14074 -678
rect 14028 -1066 14074 -1054
rect 14146 -678 14192 -666
rect 14146 -1054 14152 -678
rect 14186 -1054 14192 -678
rect 14146 -1066 14192 -1054
rect 14264 -678 14310 -666
rect 14264 -1054 14270 -678
rect 14304 -1054 14310 -678
rect 14264 -1066 14310 -1054
rect 14382 -678 14428 -666
rect 14382 -1054 14388 -678
rect 14422 -1054 14428 -678
rect 14382 -1066 14428 -1054
rect 14500 -678 14546 -666
rect 14500 -1054 14506 -678
rect 14540 -1054 14546 -678
rect 14500 -1066 14546 -1054
rect 14618 -678 14664 -666
rect 14618 -1054 14624 -678
rect 14658 -1054 14664 -678
rect 14618 -1066 14664 -1054
rect 14736 -678 14782 -666
rect 14863 -670 15034 -654
rect 15175 -608 15446 -580
rect 15175 -670 15210 -608
rect 15412 -670 15446 -608
rect 15530 -608 15800 -580
rect 15530 -670 15564 -608
rect 15766 -670 15800 -608
rect 14736 -1054 14742 -678
rect 14776 -1054 14782 -678
rect 14736 -1066 14782 -1054
rect 10374 -1180 10648 -1152
rect 11010 -1071 11592 -1070
rect 11010 -1112 11076 -1071
rect 11010 -1146 11026 -1112
rect 11060 -1146 11076 -1112
rect 11010 -1153 11076 -1146
rect 10374 -1184 11002 -1180
rect 11438 -1184 11472 -1071
rect 10374 -1196 11007 -1184
rect 10374 -1209 10967 -1196
rect 8567 -1312 8676 -1258
rect 8567 -1458 8601 -1312
rect 8740 -1326 8750 -1229
rect 8849 -1326 8859 -1229
rect 9321 -1315 9356 -1223
rect 8751 -1327 8848 -1326
rect 8791 -1394 8848 -1327
rect 9129 -1351 9356 -1315
rect 9129 -1385 9195 -1351
rect 8685 -1430 8954 -1394
rect 9129 -1419 9145 -1385
rect 9179 -1419 9195 -1385
rect 9129 -1425 9195 -1419
rect 8685 -1458 8718 -1430
rect 8921 -1458 8954 -1430
rect 9321 -1458 9356 -1351
rect 10961 -1372 10967 -1209
rect 11001 -1372 11007 -1196
rect 10961 -1384 11007 -1372
rect 11079 -1196 11125 -1184
rect 11079 -1372 11085 -1196
rect 11119 -1372 11125 -1196
rect 11079 -1384 11125 -1372
rect 11196 -1196 11242 -1184
rect 8561 -1470 8607 -1458
rect 8561 -1646 8567 -1470
rect 8601 -1646 8607 -1470
rect 8561 -1658 8607 -1646
rect 8679 -1470 8725 -1458
rect 8679 -1646 8685 -1470
rect 8719 -1646 8725 -1470
rect 8679 -1658 8725 -1646
rect 8797 -1470 8843 -1458
rect 8797 -1646 8803 -1470
rect 8837 -1646 8843 -1470
rect 8797 -1658 8843 -1646
rect 8915 -1470 8961 -1458
rect 8915 -1646 8921 -1470
rect 8955 -1525 8961 -1470
rect 9080 -1470 9126 -1458
rect 9080 -1525 9086 -1470
rect 8955 -1613 9086 -1525
rect 8955 -1646 8961 -1613
rect 8915 -1658 8961 -1646
rect 9080 -1646 9086 -1613
rect 9120 -1646 9126 -1470
rect 9080 -1658 9126 -1646
rect 9198 -1470 9244 -1458
rect 9198 -1646 9204 -1470
rect 9238 -1646 9244 -1470
rect 9198 -1658 9244 -1646
rect 9316 -1470 9362 -1458
rect 9316 -1646 9322 -1470
rect 9356 -1646 9362 -1470
rect 9316 -1658 9362 -1646
rect 9434 -1470 9480 -1458
rect 9434 -1646 9440 -1470
rect 9474 -1646 9480 -1470
rect 10880 -1500 10988 -1490
rect 11084 -1500 11119 -1384
rect 10988 -1548 11119 -1500
rect 11196 -1548 11202 -1196
rect 10988 -1572 11202 -1548
rect 11236 -1572 11242 -1196
rect 10988 -1584 11242 -1572
rect 11314 -1196 11360 -1184
rect 11314 -1572 11320 -1196
rect 11354 -1572 11360 -1196
rect 11314 -1584 11360 -1572
rect 11432 -1196 11478 -1184
rect 11432 -1572 11438 -1196
rect 11472 -1572 11478 -1196
rect 12964 -1252 13064 -1235
rect 12962 -1310 13064 -1252
rect 13132 -1310 13142 -1235
rect 14034 -1249 14068 -1066
rect 14152 -1107 14186 -1066
rect 14388 -1107 14422 -1066
rect 14152 -1136 14422 -1107
rect 14506 -1108 14540 -1066
rect 14742 -1108 14776 -1066
rect 14506 -1136 14776 -1108
rect 14742 -1184 14776 -1136
rect 14713 -1214 14776 -1184
rect 13959 -1303 14068 -1249
rect 14141 -1244 14241 -1223
rect 14141 -1298 14162 -1244
rect 14227 -1298 14241 -1244
rect 14141 -1303 14241 -1298
rect 12962 -1311 13115 -1310
rect 11432 -1584 11478 -1572
rect 10988 -1588 11236 -1584
rect 10988 -1632 11062 -1588
rect 12361 -1589 12650 -1414
rect 11600 -1616 12650 -1589
rect 11245 -1622 11311 -1616
rect 10880 -1642 10988 -1632
rect 9434 -1658 9480 -1646
rect 11245 -1656 11261 -1622
rect 11295 -1656 11311 -1622
rect 8568 -1696 8601 -1658
rect 8804 -1696 8837 -1658
rect 8568 -1732 8837 -1696
rect 9204 -1697 9238 -1658
rect 9440 -1697 9474 -1658
rect 9204 -1732 9474 -1697
rect 9204 -1733 9440 -1732
rect 9308 -1807 9440 -1733
rect 11245 -1752 11311 -1656
rect 11363 -1622 12650 -1616
rect 11363 -1656 11379 -1622
rect 11413 -1656 12650 -1622
rect 11363 -1672 12650 -1656
rect 11600 -1688 12650 -1672
rect 11663 -1689 12650 -1688
rect 12128 -1693 12650 -1689
rect 11599 -1752 12065 -1730
rect 11245 -1800 12065 -1752
rect 9298 -1915 9308 -1807
rect 9440 -1915 9450 -1807
rect 11599 -1831 12065 -1800
rect 11960 -2087 12065 -1831
rect 8437 -2263 8500 -2246
rect 11078 -2111 11298 -2091
rect 11078 -2219 11122 -2111
rect 11254 -2219 11298 -2111
rect 11880 -2193 11890 -2087
rect 12002 -2193 12065 -2087
rect 11916 -2204 12065 -2193
rect 11078 -2261 11298 -2219
rect 8437 -2267 8575 -2263
rect 8437 -2301 10407 -2267
rect 10717 -2291 11694 -2261
rect 8437 -2330 10409 -2301
rect 8437 -2332 8575 -2330
rect 10363 -2346 10409 -2330
rect 7401 -2562 7411 -2454
rect 7543 -2562 7553 -2454
rect 9299 -2562 9309 -2454
rect 9441 -2562 9451 -2454
rect 7411 -2602 7543 -2562
rect 9309 -2602 9441 -2562
rect 7411 -2668 7544 -2602
rect 9309 -2668 9442 -2602
rect 6742 -2711 8215 -2668
rect 6742 -3014 6776 -2711
rect 7107 -2814 7141 -2711
rect 7343 -2814 7377 -2711
rect 7579 -2814 7613 -2711
rect 7815 -2814 7849 -2711
rect 7101 -2826 7147 -2814
rect 5787 -3153 6529 -3050
rect 6618 -3026 6664 -3014
rect 5787 -3212 6075 -3153
rect 5787 -3214 5827 -3212
rect 5787 -3225 5821 -3214
rect 5786 -3320 5821 -3225
rect 5939 -3318 6075 -3212
rect 6618 -3202 6624 -3026
rect 6658 -3202 6664 -3026
rect 6618 -3214 6664 -3202
rect 6736 -3026 6782 -3014
rect 6736 -3202 6742 -3026
rect 6776 -3202 6782 -3026
rect 6736 -3214 6782 -3202
rect 6854 -3026 6900 -3014
rect 6854 -3202 6860 -3026
rect 6894 -3202 6900 -3026
rect 6854 -3214 6900 -3202
rect 6972 -3026 7018 -3014
rect 7101 -3026 7107 -2826
rect 6972 -3202 6978 -3026
rect 7012 -3202 7107 -3026
rect 7141 -3202 7147 -2826
rect 6972 -3214 7018 -3202
rect 7101 -3214 7147 -3202
rect 7219 -2826 7265 -2814
rect 7219 -3202 7225 -2826
rect 7259 -3202 7265 -2826
rect 7219 -3214 7265 -3202
rect 7337 -2826 7383 -2814
rect 7337 -3202 7343 -2826
rect 7377 -3202 7383 -2826
rect 7337 -3214 7383 -3202
rect 7455 -2826 7501 -2814
rect 7455 -3202 7461 -2826
rect 7495 -3202 7501 -2826
rect 7455 -3214 7501 -3202
rect 7573 -2826 7619 -2814
rect 7573 -3202 7579 -2826
rect 7613 -3202 7619 -2826
rect 7573 -3214 7619 -3202
rect 7691 -2826 7737 -2814
rect 7691 -3202 7697 -2826
rect 7731 -3202 7737 -2826
rect 7691 -3214 7737 -3202
rect 7809 -2826 7855 -2814
rect 7809 -3202 7815 -2826
rect 7849 -3026 7855 -2826
rect 8181 -3014 8215 -2711
rect 8640 -2711 10113 -2668
rect 8640 -3014 8674 -2711
rect 9005 -2814 9039 -2711
rect 9241 -2814 9275 -2711
rect 9477 -2814 9511 -2711
rect 9713 -2814 9747 -2711
rect 8999 -2826 9045 -2814
rect 7939 -3026 7985 -3014
rect 7849 -3202 7945 -3026
rect 7979 -3202 7985 -3026
rect 7809 -3214 7855 -3202
rect 7939 -3214 7985 -3202
rect 8057 -3026 8103 -3014
rect 8057 -3202 8063 -3026
rect 8097 -3202 8103 -3026
rect 8057 -3214 8103 -3202
rect 8175 -3026 8221 -3014
rect 8175 -3202 8181 -3026
rect 8215 -3202 8221 -3026
rect 8175 -3214 8221 -3202
rect 8293 -3026 8339 -3014
rect 8293 -3202 8299 -3026
rect 8333 -3202 8339 -3026
rect 8293 -3214 8339 -3202
rect 8516 -3026 8562 -3014
rect 8516 -3202 8522 -3026
rect 8556 -3202 8562 -3026
rect 8516 -3214 8562 -3202
rect 8634 -3026 8680 -3014
rect 8634 -3202 8640 -3026
rect 8674 -3202 8680 -3026
rect 8634 -3214 8680 -3202
rect 8752 -3026 8798 -3014
rect 8752 -3202 8758 -3026
rect 8792 -3202 8798 -3026
rect 8752 -3214 8798 -3202
rect 8870 -3026 8916 -3014
rect 8999 -3026 9005 -2826
rect 8870 -3202 8876 -3026
rect 8910 -3202 9005 -3026
rect 9039 -3202 9045 -2826
rect 8870 -3214 8916 -3202
rect 8999 -3214 9045 -3202
rect 9117 -2826 9163 -2814
rect 9117 -3202 9123 -2826
rect 9157 -3202 9163 -2826
rect 9117 -3214 9163 -3202
rect 9235 -2826 9281 -2814
rect 9235 -3202 9241 -2826
rect 9275 -3202 9281 -2826
rect 9235 -3214 9281 -3202
rect 9353 -2826 9399 -2814
rect 9353 -3202 9359 -2826
rect 9393 -3202 9399 -2826
rect 9353 -3214 9399 -3202
rect 9471 -2826 9517 -2814
rect 9471 -3202 9477 -2826
rect 9511 -3202 9517 -2826
rect 9471 -3214 9517 -3202
rect 9589 -2826 9635 -2814
rect 9589 -3202 9595 -2826
rect 9629 -3202 9635 -2826
rect 9589 -3214 9635 -3202
rect 9707 -2826 9753 -2814
rect 9707 -3202 9713 -2826
rect 9747 -3026 9753 -2826
rect 10079 -3014 10113 -2711
rect 10363 -2798 10410 -2346
rect 10717 -2397 10751 -2291
rect 10954 -2397 10986 -2291
rect 11190 -2397 11222 -2291
rect 11426 -2397 11458 -2291
rect 11662 -2397 11694 -2291
rect 10593 -2409 10639 -2397
rect 10593 -2585 10599 -2409
rect 10633 -2585 10639 -2409
rect 10593 -2597 10639 -2585
rect 10711 -2409 10757 -2397
rect 10711 -2585 10717 -2409
rect 10751 -2585 10757 -2409
rect 10711 -2597 10757 -2585
rect 10829 -2409 10875 -2397
rect 10829 -2585 10835 -2409
rect 10869 -2585 10875 -2409
rect 10829 -2597 10875 -2585
rect 10947 -2409 10993 -2397
rect 10947 -2585 10953 -2409
rect 10987 -2585 10993 -2409
rect 10947 -2597 10993 -2585
rect 11065 -2409 11111 -2397
rect 11065 -2585 11071 -2409
rect 11105 -2585 11111 -2409
rect 11065 -2597 11111 -2585
rect 11183 -2409 11229 -2397
rect 11183 -2585 11189 -2409
rect 11223 -2585 11229 -2409
rect 11183 -2597 11229 -2585
rect 11301 -2409 11347 -2397
rect 11301 -2585 11307 -2409
rect 11341 -2585 11347 -2409
rect 11301 -2597 11347 -2585
rect 11419 -2409 11465 -2397
rect 11419 -2585 11425 -2409
rect 11459 -2585 11465 -2409
rect 11419 -2597 11465 -2585
rect 11537 -2409 11583 -2397
rect 11537 -2585 11543 -2409
rect 11577 -2585 11583 -2409
rect 11537 -2597 11583 -2585
rect 11655 -2409 11701 -2397
rect 11655 -2585 11661 -2409
rect 11695 -2585 11701 -2409
rect 11655 -2597 11701 -2585
rect 10364 -2814 10410 -2798
rect 10364 -2815 10445 -2814
rect 10599 -2815 10634 -2597
rect 10878 -2645 10944 -2638
rect 10878 -2679 10894 -2645
rect 10928 -2679 10944 -2645
rect 10878 -2690 10944 -2679
rect 11070 -2690 11106 -2597
rect 10878 -2691 11106 -2690
rect 11306 -2691 11342 -2597
rect 11542 -2691 11578 -2597
rect 10878 -2720 11578 -2691
rect 10996 -2721 11578 -2720
rect 10996 -2762 11062 -2721
rect 10996 -2796 11012 -2762
rect 11046 -2796 11062 -2762
rect 10996 -2803 11062 -2796
rect 10364 -2830 10634 -2815
rect 10364 -2834 10988 -2830
rect 11424 -2834 11458 -2721
rect 10364 -2846 10993 -2834
rect 10364 -2858 10953 -2846
rect 10364 -2860 10445 -2858
rect 10711 -2859 10953 -2858
rect 9837 -3026 9883 -3014
rect 9747 -3202 9843 -3026
rect 9877 -3202 9883 -3026
rect 9707 -3214 9753 -3202
rect 9837 -3214 9883 -3202
rect 9955 -3026 10001 -3014
rect 9955 -3202 9961 -3026
rect 9995 -3202 10001 -3026
rect 9955 -3214 10001 -3202
rect 10073 -3026 10119 -3014
rect 10073 -3202 10079 -3026
rect 10113 -3202 10119 -3026
rect 10073 -3214 10119 -3202
rect 10191 -3026 10237 -3014
rect 10191 -3202 10197 -3026
rect 10231 -3202 10237 -3026
rect 10947 -3022 10953 -2859
rect 10987 -3022 10993 -2846
rect 10947 -3034 10993 -3022
rect 11065 -2846 11111 -2834
rect 11065 -3022 11071 -2846
rect 11105 -3022 11111 -2846
rect 11065 -3034 11111 -3022
rect 11182 -2846 11228 -2834
rect 10191 -3214 10237 -3202
rect 10866 -3150 10974 -3140
rect 11070 -3150 11105 -3034
rect 6624 -3248 6658 -3214
rect 6860 -3248 6894 -3214
rect 6624 -3283 6894 -3248
rect 7461 -3248 7495 -3214
rect 7697 -3248 7731 -3214
rect 8299 -3248 8333 -3214
rect 7461 -3283 7731 -3248
rect 8174 -3283 8333 -3248
rect 8522 -3248 8556 -3214
rect 8758 -3248 8792 -3214
rect 8522 -3283 8792 -3248
rect 9359 -3248 9393 -3214
rect 9595 -3248 9629 -3214
rect 10197 -3248 10231 -3214
rect 9359 -3283 9629 -3248
rect 10072 -3283 10231 -3248
rect 10974 -3198 11105 -3150
rect 11182 -3198 11188 -2846
rect 10974 -3222 11188 -3198
rect 11222 -3222 11228 -2846
rect 10974 -3234 11228 -3222
rect 11300 -2846 11346 -2834
rect 11300 -3222 11306 -2846
rect 11340 -3222 11346 -2846
rect 11300 -3234 11346 -3222
rect 11418 -2846 11464 -2834
rect 11418 -3222 11424 -2846
rect 11458 -3222 11464 -2846
rect 11418 -3234 11464 -3222
rect 10974 -3238 11222 -3234
rect 11591 -3238 11601 -3206
rect 10974 -3282 11048 -3238
rect 11586 -3266 11601 -3238
rect 11231 -3272 11297 -3266
rect 5933 -3320 6075 -3318
rect 5786 -3329 6075 -3320
rect 5787 -3330 6075 -3329
rect 5819 -3331 6075 -3330
rect 6610 -3461 6677 -3437
rect 6610 -3495 6626 -3461
rect 6660 -3495 6677 -3461
rect 5561 -3662 5571 -3583
rect 5664 -3662 5674 -3583
rect 4525 -3711 4745 -3691
rect 4525 -3819 4569 -3711
rect 4701 -3819 4745 -3711
rect 4525 -3861 4745 -3819
rect 4164 -3891 5141 -3861
rect 4164 -3997 4198 -3891
rect 4401 -3997 4433 -3891
rect 4637 -3997 4669 -3891
rect 4873 -3997 4905 -3891
rect 5109 -3997 5141 -3891
rect 2098 -4068 2518 -4063
rect 3232 -4068 3548 -4063
rect 2098 -4079 2585 -4068
rect 2098 -4106 2534 -4079
rect 2098 -4107 2405 -4106
rect 2098 -4235 2132 -4107
rect 2518 -4113 2534 -4106
rect 2568 -4113 2585 -4079
rect 2518 -4119 2585 -4113
rect 3165 -4079 3548 -4068
rect 3165 -4113 3182 -4079
rect 3216 -4106 3548 -4079
rect 3216 -4113 3232 -4106
rect 3165 -4119 3232 -4113
rect 2238 -4147 2294 -4135
rect 3351 -4146 3407 -4134
rect 3351 -4147 3367 -4146
rect 2238 -4181 2244 -4147
rect 2278 -4162 2848 -4147
rect 2278 -4181 2798 -4162
rect 2238 -4196 2798 -4181
rect 2832 -4196 2848 -4162
rect 2238 -4197 2294 -4196
rect 2781 -4206 2848 -4196
rect 2900 -4163 3367 -4147
rect 2900 -4197 2916 -4163
rect 2950 -4180 3367 -4163
rect 3401 -4180 3407 -4146
rect 2950 -4196 3407 -4180
rect 2950 -4197 2966 -4196
rect 2900 -4204 2966 -4197
rect 3514 -4235 3548 -4106
rect 4040 -4009 4086 -3997
rect 4040 -4185 4046 -4009
rect 4080 -4185 4086 -4009
rect 4040 -4197 4086 -4185
rect 4158 -4009 4204 -3997
rect 4158 -4185 4164 -4009
rect 4198 -4185 4204 -4009
rect 4158 -4197 4204 -4185
rect 4276 -4009 4322 -3997
rect 4276 -4185 4282 -4009
rect 4316 -4185 4322 -4009
rect 4276 -4197 4322 -4185
rect 4394 -4009 4440 -3997
rect 4394 -4185 4400 -4009
rect 4434 -4185 4440 -4009
rect 4394 -4197 4440 -4185
rect 4512 -4009 4558 -3997
rect 4512 -4185 4518 -4009
rect 4552 -4185 4558 -4009
rect 4512 -4197 4558 -4185
rect 4630 -4009 4676 -3997
rect 4630 -4185 4636 -4009
rect 4670 -4185 4676 -4009
rect 4630 -4197 4676 -4185
rect 4748 -4009 4794 -3997
rect 4748 -4185 4754 -4009
rect 4788 -4185 4794 -4009
rect 4748 -4197 4794 -4185
rect 4866 -4009 4912 -3997
rect 4866 -4185 4872 -4009
rect 4906 -4185 4912 -4009
rect 4866 -4197 4912 -4185
rect 4984 -4009 5030 -3997
rect 4984 -4185 4990 -4009
rect 5024 -4185 5030 -4009
rect 4984 -4197 5030 -4185
rect 5102 -4009 5148 -3997
rect 5102 -4185 5108 -4009
rect 5142 -4185 5148 -4009
rect 5102 -4197 5148 -4185
rect 194 -4247 240 -4235
rect 194 -4423 200 -4247
rect 234 -4423 240 -4247
rect 194 -4435 240 -4423
rect 312 -4247 358 -4235
rect 312 -4423 318 -4247
rect 352 -4423 358 -4247
rect 312 -4435 358 -4423
rect 718 -4247 764 -4235
rect 319 -4729 352 -4435
rect 718 -4623 724 -4247
rect 758 -4623 764 -4247
rect 718 -4635 764 -4623
rect 836 -4247 882 -4235
rect 836 -4623 842 -4247
rect 876 -4623 882 -4247
rect 836 -4635 882 -4623
rect 954 -4247 1000 -4235
rect 954 -4623 960 -4247
rect 994 -4623 1000 -4247
rect 954 -4635 1000 -4623
rect 1072 -4247 1118 -4235
rect 1072 -4623 1078 -4247
rect 1112 -4623 1118 -4247
rect 1072 -4635 1118 -4623
rect 1190 -4247 1236 -4235
rect 1190 -4623 1196 -4247
rect 1230 -4623 1236 -4247
rect 1492 -4247 1538 -4235
rect 1492 -4423 1498 -4247
rect 1532 -4423 1538 -4247
rect 1492 -4435 1538 -4423
rect 1610 -4247 1656 -4235
rect 1610 -4423 1616 -4247
rect 1650 -4423 1656 -4247
rect 1610 -4435 1656 -4423
rect 2092 -4247 2138 -4235
rect 2092 -4423 2098 -4247
rect 2132 -4423 2138 -4247
rect 2092 -4435 2138 -4423
rect 2210 -4247 2256 -4235
rect 2210 -4423 2216 -4247
rect 2250 -4423 2256 -4247
rect 2210 -4435 2256 -4423
rect 2616 -4247 2662 -4235
rect 1190 -4635 1236 -4623
rect 842 -4729 876 -4635
rect 1499 -4729 1533 -4435
rect 319 -4761 1533 -4729
rect 2217 -4729 2250 -4435
rect 2616 -4623 2622 -4247
rect 2656 -4623 2662 -4247
rect 2616 -4635 2662 -4623
rect 2734 -4247 2780 -4235
rect 2734 -4623 2740 -4247
rect 2774 -4623 2780 -4247
rect 2734 -4635 2780 -4623
rect 2852 -4247 2898 -4235
rect 2852 -4623 2858 -4247
rect 2892 -4623 2898 -4247
rect 2852 -4635 2898 -4623
rect 2970 -4247 3016 -4235
rect 2970 -4623 2976 -4247
rect 3010 -4623 3016 -4247
rect 2970 -4635 3016 -4623
rect 3088 -4247 3134 -4235
rect 3088 -4623 3094 -4247
rect 3128 -4623 3134 -4247
rect 3390 -4247 3436 -4235
rect 3390 -4423 3396 -4247
rect 3430 -4423 3436 -4247
rect 3390 -4435 3436 -4423
rect 3508 -4247 3554 -4235
rect 3508 -4423 3514 -4247
rect 3548 -4423 3554 -4247
rect 3508 -4435 3554 -4423
rect 4046 -4430 4081 -4197
rect 4325 -4245 4391 -4238
rect 4325 -4279 4341 -4245
rect 4375 -4279 4391 -4245
rect 4325 -4290 4391 -4279
rect 4517 -4290 4553 -4197
rect 4325 -4291 4553 -4290
rect 4753 -4291 4789 -4197
rect 4989 -4291 5025 -4197
rect 4325 -4320 5025 -4291
rect 4443 -4321 5025 -4320
rect 4443 -4362 4509 -4321
rect 4443 -4396 4459 -4362
rect 4493 -4396 4509 -4362
rect 4443 -4403 4509 -4396
rect 4046 -4434 4435 -4430
rect 4871 -4434 4905 -4321
rect 3088 -4635 3134 -4623
rect 2740 -4729 2774 -4635
rect 3397 -4729 3431 -4435
rect 4046 -4446 4440 -4434
rect 4046 -4459 4400 -4446
rect 4046 -4462 4124 -4459
rect 4041 -4514 4051 -4462
rect 4114 -4514 4124 -4462
rect 4046 -4520 4119 -4514
rect 4394 -4622 4400 -4459
rect 4434 -4622 4440 -4446
rect 4394 -4634 4440 -4622
rect 4512 -4446 4558 -4434
rect 4512 -4622 4518 -4446
rect 4552 -4622 4558 -4446
rect 4512 -4634 4558 -4622
rect 4629 -4446 4675 -4434
rect 2217 -4761 3431 -4729
rect 4313 -4750 4421 -4740
rect 4517 -4750 4552 -4634
rect 908 -4846 1040 -4761
rect 2806 -4846 2938 -4761
rect 53 -5153 119 -4874
rect 898 -4954 908 -4846
rect 1040 -4954 1050 -4846
rect 2796 -4954 2806 -4846
rect 2938 -4954 2948 -4846
rect 4421 -4798 4552 -4750
rect 4629 -4798 4635 -4446
rect 4421 -4822 4635 -4798
rect 4669 -4822 4675 -4446
rect 4421 -4834 4675 -4822
rect 4747 -4446 4793 -4434
rect 4747 -4822 4753 -4446
rect 4787 -4822 4793 -4446
rect 4747 -4834 4793 -4822
rect 4865 -4446 4911 -4434
rect 4865 -4822 4871 -4446
rect 4905 -4822 4911 -4446
rect 4865 -4834 4911 -4822
rect 4421 -4838 4669 -4834
rect 5570 -4836 5663 -3662
rect 6393 -3924 6549 -3918
rect 6393 -4022 6405 -3924
rect 6537 -4022 6549 -3924
rect 6393 -4028 6549 -4022
rect 5078 -4838 5663 -4836
rect 4421 -4882 4495 -4838
rect 5033 -4866 5663 -4838
rect 4678 -4872 4744 -4866
rect 4313 -4892 4421 -4882
rect 4678 -4906 4694 -4872
rect 4728 -4906 4744 -4872
rect 4678 -5002 4744 -4906
rect 4796 -4872 5663 -4866
rect 4796 -4906 4812 -4872
rect 4846 -4906 5663 -4872
rect 6610 -4878 6677 -3495
rect 6758 -4066 6792 -3283
rect 7461 -3345 7495 -3283
rect 7164 -3383 7906 -3345
rect 7164 -3507 7198 -3383
rect 7400 -3507 7434 -3383
rect 7636 -3507 7670 -3383
rect 7872 -3507 7906 -3383
rect 7158 -3519 7204 -3507
rect 7158 -3895 7164 -3519
rect 7198 -3895 7204 -3519
rect 7158 -3907 7204 -3895
rect 7276 -3519 7322 -3507
rect 7276 -3895 7282 -3519
rect 7316 -3895 7322 -3519
rect 7276 -3907 7322 -3895
rect 7394 -3519 7440 -3507
rect 7394 -3895 7400 -3519
rect 7434 -3895 7440 -3519
rect 7394 -3907 7440 -3895
rect 7512 -3519 7558 -3507
rect 7512 -3895 7518 -3519
rect 7552 -3895 7558 -3519
rect 7512 -3907 7558 -3895
rect 7630 -3519 7676 -3507
rect 7630 -3895 7636 -3519
rect 7670 -3895 7676 -3519
rect 7630 -3907 7676 -3895
rect 7748 -3519 7794 -3507
rect 7748 -3895 7754 -3519
rect 7788 -3895 7794 -3519
rect 7748 -3907 7794 -3895
rect 7866 -3519 7912 -3507
rect 7866 -3895 7872 -3519
rect 7906 -3895 7912 -3519
rect 7866 -3907 7912 -3895
rect 6758 -4067 7065 -4066
rect 7111 -4067 7180 -4066
rect 8174 -4067 8208 -3283
rect 6758 -4071 7180 -4067
rect 6758 -4082 7247 -4071
rect 7892 -4072 8208 -4067
rect 6758 -4110 7196 -4082
rect 6758 -4111 7065 -4110
rect 6758 -4239 6792 -4111
rect 7180 -4116 7196 -4110
rect 7230 -4116 7247 -4082
rect 7180 -4122 7247 -4116
rect 7825 -4083 8208 -4072
rect 7825 -4117 7842 -4083
rect 7876 -4110 8208 -4083
rect 7876 -4117 7892 -4110
rect 7825 -4123 7892 -4117
rect 6898 -4151 6954 -4139
rect 8011 -4150 8067 -4138
rect 8011 -4151 8027 -4150
rect 6898 -4185 6904 -4151
rect 6938 -4166 7508 -4151
rect 6938 -4185 7458 -4166
rect 6898 -4200 7458 -4185
rect 7492 -4200 7508 -4166
rect 6898 -4201 6954 -4200
rect 7441 -4210 7508 -4200
rect 7560 -4167 8027 -4151
rect 7560 -4201 7576 -4167
rect 7610 -4184 8027 -4167
rect 8061 -4184 8067 -4150
rect 7610 -4200 8067 -4184
rect 7610 -4201 7626 -4200
rect 7560 -4208 7626 -4201
rect 8174 -4239 8208 -4110
rect 8656 -4066 8690 -3283
rect 9359 -3345 9393 -3283
rect 9062 -3383 9804 -3345
rect 8723 -3490 8733 -3424
rect 8796 -3490 8806 -3424
rect 9062 -3507 9096 -3383
rect 9298 -3507 9332 -3383
rect 9534 -3507 9568 -3383
rect 9770 -3507 9804 -3383
rect 9056 -3519 9102 -3507
rect 9056 -3895 9062 -3519
rect 9096 -3895 9102 -3519
rect 9056 -3907 9102 -3895
rect 9174 -3519 9220 -3507
rect 9174 -3895 9180 -3519
rect 9214 -3895 9220 -3519
rect 9174 -3907 9220 -3895
rect 9292 -3519 9338 -3507
rect 9292 -3895 9298 -3519
rect 9332 -3895 9338 -3519
rect 9292 -3907 9338 -3895
rect 9410 -3519 9456 -3507
rect 9410 -3895 9416 -3519
rect 9450 -3895 9456 -3519
rect 9410 -3907 9456 -3895
rect 9528 -3519 9574 -3507
rect 9528 -3895 9534 -3519
rect 9568 -3895 9574 -3519
rect 9528 -3907 9574 -3895
rect 9646 -3519 9692 -3507
rect 9646 -3895 9652 -3519
rect 9686 -3895 9692 -3519
rect 9646 -3907 9692 -3895
rect 9764 -3519 9810 -3507
rect 9764 -3895 9770 -3519
rect 9804 -3895 9810 -3519
rect 9764 -3907 9810 -3895
rect 8656 -4067 8963 -4066
rect 10072 -4067 10106 -3283
rect 10866 -3292 10974 -3282
rect 11231 -3306 11247 -3272
rect 11281 -3306 11297 -3272
rect 11231 -3402 11297 -3306
rect 11349 -3272 11601 -3266
rect 11349 -3306 11365 -3272
rect 11399 -3306 11601 -3272
rect 11349 -3322 11601 -3306
rect 11586 -3324 11601 -3322
rect 11719 -3324 11729 -3206
rect 11586 -3338 11686 -3324
rect 11586 -3381 11686 -3380
rect 11960 -3381 12065 -2204
rect 11586 -3402 12065 -3381
rect 11231 -3450 12065 -3402
rect 11586 -3479 12065 -3450
rect 11586 -3480 11686 -3479
rect 11960 -3481 12065 -3479
rect 12128 -3587 12221 -1693
rect 12361 -1694 12650 -1693
rect 12344 -2104 12633 -1942
rect 12344 -2117 12384 -2104
rect 12342 -2210 12384 -2117
rect 12496 -2210 12633 -2104
rect 12342 -2221 12633 -2210
rect 12344 -2222 12633 -2221
rect 12962 -3051 13062 -1311
rect 13959 -1449 13993 -1303
rect 14143 -1318 14240 -1303
rect 14713 -1306 14748 -1214
rect 14183 -1385 14240 -1318
rect 14521 -1342 14748 -1306
rect 14521 -1376 14587 -1342
rect 14077 -1421 14346 -1385
rect 14521 -1410 14537 -1376
rect 14571 -1410 14587 -1376
rect 14521 -1416 14587 -1410
rect 14077 -1449 14110 -1421
rect 14313 -1449 14346 -1421
rect 14713 -1449 14748 -1342
rect 13953 -1461 13999 -1449
rect 13953 -1637 13959 -1461
rect 13993 -1637 13999 -1461
rect 13953 -1649 13999 -1637
rect 14071 -1461 14117 -1449
rect 14071 -1637 14077 -1461
rect 14111 -1637 14117 -1461
rect 14071 -1649 14117 -1637
rect 14189 -1461 14235 -1449
rect 14189 -1637 14195 -1461
rect 14229 -1637 14235 -1461
rect 14189 -1649 14235 -1637
rect 14307 -1461 14353 -1449
rect 14307 -1637 14313 -1461
rect 14347 -1516 14353 -1461
rect 14472 -1461 14518 -1449
rect 14472 -1516 14478 -1461
rect 14347 -1604 14478 -1516
rect 14347 -1637 14353 -1604
rect 14307 -1649 14353 -1637
rect 14472 -1637 14478 -1604
rect 14512 -1637 14518 -1461
rect 14472 -1649 14518 -1637
rect 14590 -1461 14636 -1449
rect 14590 -1637 14596 -1461
rect 14630 -1637 14636 -1461
rect 14590 -1649 14636 -1637
rect 14708 -1461 14754 -1449
rect 14708 -1637 14714 -1461
rect 14748 -1637 14754 -1461
rect 14708 -1649 14754 -1637
rect 14826 -1461 14872 -1449
rect 14826 -1637 14832 -1461
rect 14866 -1637 14872 -1461
rect 14826 -1649 14872 -1637
rect 13960 -1687 13993 -1649
rect 14196 -1687 14229 -1649
rect 13960 -1723 14229 -1687
rect 14596 -1688 14630 -1649
rect 14832 -1688 14866 -1649
rect 14596 -1724 14866 -1688
rect 14700 -1725 14866 -1724
rect 14700 -1804 14832 -1725
rect 14690 -1912 14700 -1804
rect 14832 -1912 14842 -1804
rect 14972 -2241 15034 -670
rect 15170 -682 15216 -670
rect 15170 -1058 15176 -682
rect 15210 -1058 15216 -682
rect 15170 -1070 15216 -1058
rect 15288 -682 15334 -670
rect 15288 -1058 15294 -682
rect 15328 -1058 15334 -682
rect 15288 -1070 15334 -1058
rect 15406 -682 15452 -670
rect 15406 -1058 15412 -682
rect 15446 -1058 15452 -682
rect 15406 -1070 15452 -1058
rect 15524 -682 15570 -670
rect 15524 -1058 15530 -682
rect 15564 -1058 15570 -682
rect 15524 -1070 15570 -1058
rect 15642 -682 15688 -670
rect 15642 -1058 15648 -682
rect 15682 -1058 15688 -682
rect 15642 -1070 15688 -1058
rect 15760 -682 15806 -670
rect 15760 -1058 15766 -682
rect 15800 -1058 15806 -682
rect 15760 -1070 15806 -1058
rect 15878 -682 15924 -670
rect 15973 -674 15983 -608
rect 16049 -674 16059 -608
rect 15878 -1058 15884 -682
rect 15918 -1058 15924 -682
rect 15878 -1070 15924 -1058
rect 15176 -1253 15210 -1070
rect 15294 -1111 15328 -1070
rect 15530 -1111 15564 -1070
rect 15294 -1140 15564 -1111
rect 15648 -1112 15682 -1070
rect 15884 -1112 15918 -1070
rect 15648 -1140 15918 -1112
rect 15884 -1188 15918 -1140
rect 15855 -1218 15918 -1188
rect 16908 -1147 16975 -557
rect 17626 -564 17670 -456
rect 17802 -564 17846 -456
rect 20544 -462 20554 -399
rect 20542 -473 20554 -462
rect 17626 -606 17846 -564
rect 20541 -507 20554 -473
rect 20686 -507 20696 -399
rect 21691 -462 21701 -399
rect 21689 -473 21701 -462
rect 21376 -483 21432 -481
rect 20541 -545 20686 -507
rect 20541 -573 20582 -545
rect 21366 -549 21376 -483
rect 21432 -549 21442 -483
rect 21688 -507 21701 -473
rect 21833 -507 21843 -399
rect 24139 -453 24359 -433
rect 22506 -495 22562 -487
rect 22506 -503 23488 -495
rect 21688 -545 21833 -507
rect 22506 -537 22512 -503
rect 22546 -537 23488 -503
rect 20541 -601 20817 -573
rect 17265 -636 18242 -606
rect 17265 -742 17299 -636
rect 17502 -742 17534 -636
rect 17738 -742 17770 -636
rect 17974 -742 18006 -636
rect 18210 -742 18242 -636
rect 20541 -663 20581 -601
rect 20783 -663 20817 -601
rect 20901 -601 21171 -573
rect 21688 -577 21729 -545
rect 22506 -553 23488 -537
rect 22509 -554 23488 -553
rect 20901 -663 20935 -601
rect 21137 -663 21171 -601
rect 21376 -617 21547 -601
rect 21376 -651 21382 -617
rect 21416 -651 21547 -617
rect 20541 -675 20587 -663
rect 17141 -754 17187 -742
rect 17141 -930 17147 -754
rect 17181 -930 17187 -754
rect 17141 -942 17187 -930
rect 17259 -754 17305 -742
rect 17259 -930 17265 -754
rect 17299 -930 17305 -754
rect 17259 -942 17305 -930
rect 17377 -754 17423 -742
rect 17377 -930 17383 -754
rect 17417 -930 17423 -754
rect 17377 -942 17423 -930
rect 17495 -754 17541 -742
rect 17495 -930 17501 -754
rect 17535 -930 17541 -754
rect 17495 -942 17541 -930
rect 17613 -754 17659 -742
rect 17613 -930 17619 -754
rect 17653 -930 17659 -754
rect 17613 -942 17659 -930
rect 17731 -754 17777 -742
rect 17731 -930 17737 -754
rect 17771 -930 17777 -754
rect 17731 -942 17777 -930
rect 17849 -754 17895 -742
rect 17849 -930 17855 -754
rect 17889 -930 17895 -754
rect 17849 -942 17895 -930
rect 17967 -754 18013 -742
rect 17967 -930 17973 -754
rect 18007 -930 18013 -754
rect 17967 -942 18013 -930
rect 18085 -754 18131 -742
rect 18085 -930 18091 -754
rect 18125 -930 18131 -754
rect 18085 -942 18131 -930
rect 18203 -754 18249 -742
rect 18203 -930 18209 -754
rect 18243 -930 18249 -754
rect 18203 -942 18249 -930
rect 17147 -1147 17182 -942
rect 17426 -990 17492 -983
rect 17426 -1024 17442 -990
rect 17476 -1024 17492 -990
rect 17426 -1035 17492 -1024
rect 17618 -1035 17654 -942
rect 17426 -1036 17654 -1035
rect 17854 -1036 17890 -942
rect 18090 -1036 18126 -942
rect 17426 -1065 18126 -1036
rect 20541 -1051 20547 -675
rect 20581 -1051 20587 -675
rect 20541 -1063 20587 -1051
rect 20659 -675 20705 -663
rect 20659 -1051 20665 -675
rect 20699 -1051 20705 -675
rect 20659 -1063 20705 -1051
rect 20777 -675 20823 -663
rect 20777 -1051 20783 -675
rect 20817 -1051 20823 -675
rect 20777 -1063 20823 -1051
rect 20895 -675 20941 -663
rect 20895 -1051 20901 -675
rect 20935 -1051 20941 -675
rect 20895 -1063 20941 -1051
rect 21013 -675 21059 -663
rect 21013 -1051 21019 -675
rect 21053 -1051 21059 -675
rect 21013 -1063 21059 -1051
rect 21131 -675 21177 -663
rect 21131 -1051 21137 -675
rect 21171 -1051 21177 -675
rect 21131 -1063 21177 -1051
rect 21249 -675 21295 -663
rect 21376 -667 21547 -651
rect 21688 -605 21959 -577
rect 21688 -667 21723 -605
rect 21925 -667 21959 -605
rect 22043 -605 22313 -577
rect 22043 -667 22077 -605
rect 22279 -667 22313 -605
rect 21249 -1051 21255 -675
rect 21289 -1051 21295 -675
rect 21249 -1063 21295 -1051
rect 16908 -1175 17182 -1147
rect 17544 -1066 18126 -1065
rect 17544 -1107 17610 -1066
rect 17544 -1141 17560 -1107
rect 17594 -1141 17610 -1107
rect 17544 -1148 17610 -1141
rect 16908 -1179 17536 -1175
rect 17972 -1179 18006 -1066
rect 16908 -1191 17541 -1179
rect 16908 -1204 17501 -1191
rect 15101 -1307 15210 -1253
rect 15101 -1453 15135 -1307
rect 15274 -1321 15284 -1224
rect 15383 -1321 15393 -1224
rect 15855 -1310 15890 -1218
rect 15285 -1322 15382 -1321
rect 15325 -1389 15382 -1322
rect 15663 -1346 15890 -1310
rect 15663 -1380 15729 -1346
rect 15219 -1425 15488 -1389
rect 15663 -1414 15679 -1380
rect 15713 -1414 15729 -1380
rect 15663 -1420 15729 -1414
rect 15219 -1453 15252 -1425
rect 15455 -1453 15488 -1425
rect 15855 -1453 15890 -1346
rect 17495 -1367 17501 -1204
rect 17535 -1367 17541 -1191
rect 17495 -1379 17541 -1367
rect 17613 -1191 17659 -1179
rect 17613 -1367 17619 -1191
rect 17653 -1367 17659 -1191
rect 17613 -1379 17659 -1367
rect 17730 -1191 17776 -1179
rect 15095 -1465 15141 -1453
rect 15095 -1641 15101 -1465
rect 15135 -1641 15141 -1465
rect 15095 -1653 15141 -1641
rect 15213 -1465 15259 -1453
rect 15213 -1641 15219 -1465
rect 15253 -1641 15259 -1465
rect 15213 -1653 15259 -1641
rect 15331 -1465 15377 -1453
rect 15331 -1641 15337 -1465
rect 15371 -1641 15377 -1465
rect 15331 -1653 15377 -1641
rect 15449 -1465 15495 -1453
rect 15449 -1641 15455 -1465
rect 15489 -1520 15495 -1465
rect 15614 -1465 15660 -1453
rect 15614 -1520 15620 -1465
rect 15489 -1608 15620 -1520
rect 15489 -1641 15495 -1608
rect 15449 -1653 15495 -1641
rect 15614 -1641 15620 -1608
rect 15654 -1641 15660 -1465
rect 15614 -1653 15660 -1641
rect 15732 -1465 15778 -1453
rect 15732 -1641 15738 -1465
rect 15772 -1641 15778 -1465
rect 15732 -1653 15778 -1641
rect 15850 -1465 15896 -1453
rect 15850 -1641 15856 -1465
rect 15890 -1641 15896 -1465
rect 15850 -1653 15896 -1641
rect 15968 -1465 16014 -1453
rect 15968 -1641 15974 -1465
rect 16008 -1641 16014 -1465
rect 17414 -1495 17522 -1485
rect 17618 -1495 17653 -1379
rect 17522 -1543 17653 -1495
rect 17730 -1543 17736 -1191
rect 17522 -1567 17736 -1543
rect 17770 -1567 17776 -1191
rect 17522 -1579 17776 -1567
rect 17848 -1191 17894 -1179
rect 17848 -1567 17854 -1191
rect 17888 -1567 17894 -1191
rect 17848 -1579 17894 -1567
rect 17966 -1191 18012 -1179
rect 17966 -1567 17972 -1191
rect 18006 -1567 18012 -1191
rect 19477 -1307 19577 -1232
rect 19645 -1307 19655 -1232
rect 20547 -1246 20581 -1063
rect 20665 -1104 20699 -1063
rect 20901 -1104 20935 -1063
rect 20665 -1133 20935 -1104
rect 21019 -1105 21053 -1063
rect 21255 -1105 21289 -1063
rect 21019 -1133 21289 -1105
rect 21255 -1181 21289 -1133
rect 21226 -1211 21289 -1181
rect 20472 -1300 20581 -1246
rect 20654 -1241 20754 -1220
rect 20654 -1295 20675 -1241
rect 20740 -1295 20754 -1241
rect 20654 -1300 20754 -1295
rect 19477 -1308 19628 -1307
rect 17966 -1579 18012 -1567
rect 17522 -1583 17770 -1579
rect 17522 -1627 17596 -1583
rect 18895 -1584 19184 -1409
rect 18134 -1611 19184 -1584
rect 17779 -1617 17845 -1611
rect 17414 -1637 17522 -1627
rect 15968 -1653 16014 -1641
rect 17779 -1651 17795 -1617
rect 17829 -1651 17845 -1617
rect 15102 -1691 15135 -1653
rect 15338 -1691 15371 -1653
rect 15102 -1727 15371 -1691
rect 15738 -1692 15772 -1653
rect 15974 -1692 16008 -1653
rect 15738 -1727 16008 -1692
rect 15738 -1728 15974 -1727
rect 15842 -1802 15974 -1728
rect 17779 -1747 17845 -1651
rect 17897 -1617 19184 -1611
rect 17897 -1651 17913 -1617
rect 17947 -1651 19184 -1617
rect 17897 -1667 19184 -1651
rect 18134 -1683 19184 -1667
rect 18197 -1684 19184 -1683
rect 18662 -1688 19184 -1684
rect 18133 -1747 18599 -1725
rect 17779 -1795 18599 -1747
rect 15832 -1910 15842 -1802
rect 15974 -1910 15984 -1802
rect 18133 -1826 18599 -1795
rect 18494 -2082 18599 -1826
rect 14971 -2258 15034 -2241
rect 17612 -2106 17832 -2086
rect 17612 -2214 17656 -2106
rect 17788 -2214 17832 -2106
rect 18414 -2188 18424 -2082
rect 18536 -2188 18599 -2082
rect 18450 -2199 18599 -2188
rect 17612 -2256 17832 -2214
rect 14971 -2262 15109 -2258
rect 14971 -2296 16941 -2262
rect 17251 -2286 18228 -2256
rect 14971 -2325 16943 -2296
rect 14971 -2327 15109 -2325
rect 16897 -2341 16943 -2325
rect 13935 -2557 13945 -2449
rect 14077 -2557 14087 -2449
rect 15833 -2557 15843 -2449
rect 15975 -2557 15985 -2449
rect 13945 -2597 14077 -2557
rect 15843 -2597 15975 -2557
rect 13945 -2663 14078 -2597
rect 15843 -2663 15976 -2597
rect 13276 -2706 14749 -2663
rect 13276 -3009 13310 -2706
rect 13641 -2809 13675 -2706
rect 13877 -2809 13911 -2706
rect 14113 -2809 14147 -2706
rect 14349 -2809 14383 -2706
rect 13635 -2821 13681 -2809
rect 12377 -3054 13062 -3051
rect 12345 -3152 13062 -3054
rect 13152 -3021 13198 -3009
rect 12345 -3153 12820 -3152
rect 12345 -3216 12633 -3153
rect 13152 -3197 13158 -3021
rect 13192 -3197 13198 -3021
rect 13152 -3209 13198 -3197
rect 13270 -3021 13316 -3009
rect 13270 -3197 13276 -3021
rect 13310 -3197 13316 -3021
rect 13270 -3209 13316 -3197
rect 13388 -3021 13434 -3009
rect 13388 -3197 13394 -3021
rect 13428 -3197 13434 -3021
rect 13388 -3209 13434 -3197
rect 13506 -3021 13552 -3009
rect 13635 -3021 13641 -2821
rect 13506 -3197 13512 -3021
rect 13546 -3197 13641 -3021
rect 13675 -3197 13681 -2821
rect 13506 -3209 13552 -3197
rect 13635 -3209 13681 -3197
rect 13753 -2821 13799 -2809
rect 13753 -3197 13759 -2821
rect 13793 -3197 13799 -2821
rect 13753 -3209 13799 -3197
rect 13871 -2821 13917 -2809
rect 13871 -3197 13877 -2821
rect 13911 -3197 13917 -2821
rect 13871 -3209 13917 -3197
rect 13989 -2821 14035 -2809
rect 13989 -3197 13995 -2821
rect 14029 -3197 14035 -2821
rect 13989 -3209 14035 -3197
rect 14107 -2821 14153 -2809
rect 14107 -3197 14113 -2821
rect 14147 -3197 14153 -2821
rect 14107 -3209 14153 -3197
rect 14225 -2821 14271 -2809
rect 14225 -3197 14231 -2821
rect 14265 -3197 14271 -2821
rect 14225 -3209 14271 -3197
rect 14343 -2821 14389 -2809
rect 14343 -3197 14349 -2821
rect 14383 -3021 14389 -2821
rect 14715 -3009 14749 -2706
rect 15174 -2706 16647 -2663
rect 15174 -3009 15208 -2706
rect 15539 -2809 15573 -2706
rect 15775 -2809 15809 -2706
rect 16011 -2809 16045 -2706
rect 16247 -2809 16281 -2706
rect 15533 -2821 15579 -2809
rect 14473 -3021 14519 -3009
rect 14383 -3197 14479 -3021
rect 14513 -3197 14519 -3021
rect 14343 -3209 14389 -3197
rect 14473 -3209 14519 -3197
rect 14591 -3021 14637 -3009
rect 14591 -3197 14597 -3021
rect 14631 -3197 14637 -3021
rect 14591 -3209 14637 -3197
rect 14709 -3021 14755 -3009
rect 14709 -3197 14715 -3021
rect 14749 -3197 14755 -3021
rect 14709 -3209 14755 -3197
rect 14827 -3021 14873 -3009
rect 14827 -3197 14833 -3021
rect 14867 -3197 14873 -3021
rect 14827 -3209 14873 -3197
rect 15050 -3021 15096 -3009
rect 15050 -3197 15056 -3021
rect 15090 -3197 15096 -3021
rect 15050 -3209 15096 -3197
rect 15168 -3021 15214 -3009
rect 15168 -3197 15174 -3021
rect 15208 -3197 15214 -3021
rect 15168 -3209 15214 -3197
rect 15286 -3021 15332 -3009
rect 15286 -3197 15292 -3021
rect 15326 -3197 15332 -3021
rect 15286 -3209 15332 -3197
rect 15404 -3021 15450 -3009
rect 15533 -3021 15539 -2821
rect 15404 -3197 15410 -3021
rect 15444 -3197 15539 -3021
rect 15573 -3197 15579 -2821
rect 15404 -3209 15450 -3197
rect 15533 -3209 15579 -3197
rect 15651 -2821 15697 -2809
rect 15651 -3197 15657 -2821
rect 15691 -3197 15697 -2821
rect 15651 -3209 15697 -3197
rect 15769 -2821 15815 -2809
rect 15769 -3197 15775 -2821
rect 15809 -3197 15815 -2821
rect 15769 -3209 15815 -3197
rect 15887 -2821 15933 -2809
rect 15887 -3197 15893 -2821
rect 15927 -3197 15933 -2821
rect 15887 -3209 15933 -3197
rect 16005 -2821 16051 -2809
rect 16005 -3197 16011 -2821
rect 16045 -3197 16051 -2821
rect 16005 -3209 16051 -3197
rect 16123 -2821 16169 -2809
rect 16123 -3197 16129 -2821
rect 16163 -3197 16169 -2821
rect 16123 -3209 16169 -3197
rect 16241 -2821 16287 -2809
rect 16241 -3197 16247 -2821
rect 16281 -3021 16287 -2821
rect 16613 -3009 16647 -2706
rect 16897 -2793 16944 -2341
rect 17251 -2392 17285 -2286
rect 17488 -2392 17520 -2286
rect 17724 -2392 17756 -2286
rect 17960 -2392 17992 -2286
rect 18196 -2392 18228 -2286
rect 17127 -2404 17173 -2392
rect 17127 -2580 17133 -2404
rect 17167 -2580 17173 -2404
rect 17127 -2592 17173 -2580
rect 17245 -2404 17291 -2392
rect 17245 -2580 17251 -2404
rect 17285 -2580 17291 -2404
rect 17245 -2592 17291 -2580
rect 17363 -2404 17409 -2392
rect 17363 -2580 17369 -2404
rect 17403 -2580 17409 -2404
rect 17363 -2592 17409 -2580
rect 17481 -2404 17527 -2392
rect 17481 -2580 17487 -2404
rect 17521 -2580 17527 -2404
rect 17481 -2592 17527 -2580
rect 17599 -2404 17645 -2392
rect 17599 -2580 17605 -2404
rect 17639 -2580 17645 -2404
rect 17599 -2592 17645 -2580
rect 17717 -2404 17763 -2392
rect 17717 -2580 17723 -2404
rect 17757 -2580 17763 -2404
rect 17717 -2592 17763 -2580
rect 17835 -2404 17881 -2392
rect 17835 -2580 17841 -2404
rect 17875 -2580 17881 -2404
rect 17835 -2592 17881 -2580
rect 17953 -2404 17999 -2392
rect 17953 -2580 17959 -2404
rect 17993 -2580 17999 -2404
rect 17953 -2592 17999 -2580
rect 18071 -2404 18117 -2392
rect 18071 -2580 18077 -2404
rect 18111 -2580 18117 -2404
rect 18071 -2592 18117 -2580
rect 18189 -2404 18235 -2392
rect 18189 -2580 18195 -2404
rect 18229 -2580 18235 -2404
rect 18189 -2592 18235 -2580
rect 16898 -2809 16944 -2793
rect 16898 -2810 16979 -2809
rect 17133 -2810 17168 -2592
rect 17412 -2640 17478 -2633
rect 17412 -2674 17428 -2640
rect 17462 -2674 17478 -2640
rect 17412 -2685 17478 -2674
rect 17604 -2685 17640 -2592
rect 17412 -2686 17640 -2685
rect 17840 -2686 17876 -2592
rect 18076 -2686 18112 -2592
rect 17412 -2715 18112 -2686
rect 17530 -2716 18112 -2715
rect 17530 -2757 17596 -2716
rect 17530 -2791 17546 -2757
rect 17580 -2791 17596 -2757
rect 17530 -2798 17596 -2791
rect 16898 -2825 17168 -2810
rect 16898 -2829 17522 -2825
rect 17958 -2829 17992 -2716
rect 16898 -2841 17527 -2829
rect 16898 -2853 17487 -2841
rect 16898 -2855 16979 -2853
rect 17245 -2854 17487 -2853
rect 16371 -3021 16417 -3009
rect 16281 -3197 16377 -3021
rect 16411 -3197 16417 -3021
rect 16241 -3209 16287 -3197
rect 16371 -3209 16417 -3197
rect 16489 -3021 16535 -3009
rect 16489 -3197 16495 -3021
rect 16529 -3197 16535 -3021
rect 16489 -3209 16535 -3197
rect 16607 -3021 16653 -3009
rect 16607 -3197 16613 -3021
rect 16647 -3197 16653 -3021
rect 16607 -3209 16653 -3197
rect 16725 -3021 16771 -3009
rect 16725 -3197 16731 -3021
rect 16765 -3197 16771 -3021
rect 17481 -3017 17487 -2854
rect 17521 -3017 17527 -2841
rect 17481 -3029 17527 -3017
rect 17599 -2841 17645 -2829
rect 17599 -3017 17605 -2841
rect 17639 -3017 17645 -2841
rect 17599 -3029 17645 -3017
rect 17716 -2841 17762 -2829
rect 16725 -3209 16771 -3197
rect 17400 -3145 17508 -3135
rect 17604 -3145 17639 -3029
rect 12345 -3218 12385 -3216
rect 12345 -3229 12379 -3218
rect 12344 -3324 12379 -3229
rect 12497 -3322 12633 -3216
rect 13158 -3243 13192 -3209
rect 13394 -3243 13428 -3209
rect 13158 -3278 13428 -3243
rect 13995 -3243 14029 -3209
rect 14231 -3243 14265 -3209
rect 14833 -3243 14867 -3209
rect 13995 -3278 14265 -3243
rect 14708 -3278 14867 -3243
rect 15056 -3243 15090 -3209
rect 15292 -3243 15326 -3209
rect 15056 -3278 15326 -3243
rect 15893 -3243 15927 -3209
rect 16129 -3243 16163 -3209
rect 16731 -3243 16765 -3209
rect 15893 -3278 16163 -3243
rect 16606 -3278 16765 -3243
rect 17508 -3193 17639 -3145
rect 17716 -3193 17722 -2841
rect 17508 -3217 17722 -3193
rect 17756 -3217 17762 -2841
rect 17508 -3229 17762 -3217
rect 17834 -2841 17880 -2829
rect 17834 -3217 17840 -2841
rect 17874 -3217 17880 -2841
rect 17834 -3229 17880 -3217
rect 17952 -2841 17998 -2829
rect 17952 -3217 17958 -2841
rect 17992 -3217 17998 -2841
rect 17952 -3229 17998 -3217
rect 17508 -3233 17756 -3229
rect 18125 -3233 18135 -3201
rect 17508 -3277 17582 -3233
rect 18120 -3261 18135 -3233
rect 17765 -3267 17831 -3261
rect 12491 -3324 12633 -3322
rect 12344 -3333 12633 -3324
rect 12345 -3334 12633 -3333
rect 12377 -3335 12633 -3334
rect 13144 -3456 13211 -3432
rect 13144 -3490 13160 -3456
rect 13194 -3490 13211 -3456
rect 12119 -3666 12129 -3587
rect 12222 -3666 12232 -3587
rect 11083 -3715 11303 -3695
rect 11083 -3823 11127 -3715
rect 11259 -3823 11303 -3715
rect 11083 -3865 11303 -3823
rect 10722 -3895 11699 -3865
rect 10722 -4001 10756 -3895
rect 10959 -4001 10991 -3895
rect 11195 -4001 11227 -3895
rect 11431 -4001 11463 -3895
rect 11667 -4001 11699 -3895
rect 8656 -4072 9076 -4067
rect 9790 -4072 10106 -4067
rect 8656 -4083 9143 -4072
rect 8656 -4110 9092 -4083
rect 8656 -4111 8963 -4110
rect 8656 -4239 8690 -4111
rect 9076 -4117 9092 -4110
rect 9126 -4117 9143 -4083
rect 9076 -4123 9143 -4117
rect 9723 -4083 10106 -4072
rect 9723 -4117 9740 -4083
rect 9774 -4110 10106 -4083
rect 9774 -4117 9790 -4110
rect 9723 -4123 9790 -4117
rect 8796 -4151 8852 -4139
rect 9909 -4150 9965 -4138
rect 9909 -4151 9925 -4150
rect 8796 -4185 8802 -4151
rect 8836 -4166 9406 -4151
rect 8836 -4185 9356 -4166
rect 8796 -4200 9356 -4185
rect 9390 -4200 9406 -4166
rect 8796 -4201 8852 -4200
rect 9339 -4210 9406 -4200
rect 9458 -4167 9925 -4151
rect 9458 -4201 9474 -4167
rect 9508 -4184 9925 -4167
rect 9959 -4184 9965 -4150
rect 9508 -4200 9965 -4184
rect 9508 -4201 9524 -4200
rect 9458 -4208 9524 -4201
rect 10072 -4239 10106 -4110
rect 10598 -4013 10644 -4001
rect 10598 -4189 10604 -4013
rect 10638 -4189 10644 -4013
rect 10598 -4201 10644 -4189
rect 10716 -4013 10762 -4001
rect 10716 -4189 10722 -4013
rect 10756 -4189 10762 -4013
rect 10716 -4201 10762 -4189
rect 10834 -4013 10880 -4001
rect 10834 -4189 10840 -4013
rect 10874 -4189 10880 -4013
rect 10834 -4201 10880 -4189
rect 10952 -4013 10998 -4001
rect 10952 -4189 10958 -4013
rect 10992 -4189 10998 -4013
rect 10952 -4201 10998 -4189
rect 11070 -4013 11116 -4001
rect 11070 -4189 11076 -4013
rect 11110 -4189 11116 -4013
rect 11070 -4201 11116 -4189
rect 11188 -4013 11234 -4001
rect 11188 -4189 11194 -4013
rect 11228 -4189 11234 -4013
rect 11188 -4201 11234 -4189
rect 11306 -4013 11352 -4001
rect 11306 -4189 11312 -4013
rect 11346 -4189 11352 -4013
rect 11306 -4201 11352 -4189
rect 11424 -4013 11470 -4001
rect 11424 -4189 11430 -4013
rect 11464 -4189 11470 -4013
rect 11424 -4201 11470 -4189
rect 11542 -4013 11588 -4001
rect 11542 -4189 11548 -4013
rect 11582 -4189 11588 -4013
rect 11542 -4201 11588 -4189
rect 11660 -4013 11706 -4001
rect 11660 -4189 11666 -4013
rect 11700 -4189 11706 -4013
rect 11660 -4201 11706 -4189
rect 6752 -4251 6798 -4239
rect 6752 -4427 6758 -4251
rect 6792 -4427 6798 -4251
rect 6752 -4439 6798 -4427
rect 6870 -4251 6916 -4239
rect 6870 -4427 6876 -4251
rect 6910 -4427 6916 -4251
rect 6870 -4439 6916 -4427
rect 7276 -4251 7322 -4239
rect 6877 -4733 6910 -4439
rect 7276 -4627 7282 -4251
rect 7316 -4627 7322 -4251
rect 7276 -4639 7322 -4627
rect 7394 -4251 7440 -4239
rect 7394 -4627 7400 -4251
rect 7434 -4627 7440 -4251
rect 7394 -4639 7440 -4627
rect 7512 -4251 7558 -4239
rect 7512 -4627 7518 -4251
rect 7552 -4627 7558 -4251
rect 7512 -4639 7558 -4627
rect 7630 -4251 7676 -4239
rect 7630 -4627 7636 -4251
rect 7670 -4627 7676 -4251
rect 7630 -4639 7676 -4627
rect 7748 -4251 7794 -4239
rect 7748 -4627 7754 -4251
rect 7788 -4627 7794 -4251
rect 8050 -4251 8096 -4239
rect 8050 -4427 8056 -4251
rect 8090 -4427 8096 -4251
rect 8050 -4439 8096 -4427
rect 8168 -4251 8214 -4239
rect 8168 -4427 8174 -4251
rect 8208 -4427 8214 -4251
rect 8168 -4439 8214 -4427
rect 8650 -4251 8696 -4239
rect 8650 -4427 8656 -4251
rect 8690 -4427 8696 -4251
rect 8650 -4439 8696 -4427
rect 8768 -4251 8814 -4239
rect 8768 -4427 8774 -4251
rect 8808 -4427 8814 -4251
rect 8768 -4439 8814 -4427
rect 9174 -4251 9220 -4239
rect 7748 -4639 7794 -4627
rect 7400 -4733 7434 -4639
rect 8057 -4733 8091 -4439
rect 6877 -4765 8091 -4733
rect 8775 -4733 8808 -4439
rect 9174 -4627 9180 -4251
rect 9214 -4627 9220 -4251
rect 9174 -4639 9220 -4627
rect 9292 -4251 9338 -4239
rect 9292 -4627 9298 -4251
rect 9332 -4627 9338 -4251
rect 9292 -4639 9338 -4627
rect 9410 -4251 9456 -4239
rect 9410 -4627 9416 -4251
rect 9450 -4627 9456 -4251
rect 9410 -4639 9456 -4627
rect 9528 -4251 9574 -4239
rect 9528 -4627 9534 -4251
rect 9568 -4627 9574 -4251
rect 9528 -4639 9574 -4627
rect 9646 -4251 9692 -4239
rect 9646 -4627 9652 -4251
rect 9686 -4627 9692 -4251
rect 9948 -4251 9994 -4239
rect 9948 -4427 9954 -4251
rect 9988 -4427 9994 -4251
rect 9948 -4439 9994 -4427
rect 10066 -4251 10112 -4239
rect 10066 -4427 10072 -4251
rect 10106 -4427 10112 -4251
rect 10066 -4439 10112 -4427
rect 10604 -4434 10639 -4201
rect 10883 -4249 10949 -4242
rect 10883 -4283 10899 -4249
rect 10933 -4283 10949 -4249
rect 10883 -4294 10949 -4283
rect 11075 -4294 11111 -4201
rect 10883 -4295 11111 -4294
rect 11311 -4295 11347 -4201
rect 11547 -4295 11583 -4201
rect 10883 -4324 11583 -4295
rect 11001 -4325 11583 -4324
rect 11001 -4366 11067 -4325
rect 11001 -4400 11017 -4366
rect 11051 -4400 11067 -4366
rect 11001 -4407 11067 -4400
rect 10604 -4438 10993 -4434
rect 11429 -4438 11463 -4325
rect 9646 -4639 9692 -4627
rect 9298 -4733 9332 -4639
rect 9955 -4733 9989 -4439
rect 10604 -4450 10998 -4438
rect 10604 -4463 10958 -4450
rect 10604 -4466 10682 -4463
rect 10599 -4518 10609 -4466
rect 10672 -4518 10682 -4466
rect 10604 -4524 10677 -4518
rect 10952 -4626 10958 -4463
rect 10992 -4626 10998 -4450
rect 10952 -4638 10998 -4626
rect 11070 -4450 11116 -4438
rect 11070 -4626 11076 -4450
rect 11110 -4626 11116 -4450
rect 11070 -4638 11116 -4626
rect 11187 -4450 11233 -4438
rect 8775 -4765 9989 -4733
rect 10871 -4754 10979 -4744
rect 11075 -4754 11110 -4638
rect 7466 -4850 7598 -4765
rect 9364 -4850 9496 -4765
rect 4796 -4922 5663 -4906
rect 5033 -4938 5663 -4922
rect 5078 -4942 5663 -4938
rect 5562 -4943 5663 -4942
rect 5033 -4991 5133 -4980
rect 5033 -5002 5047 -4991
rect 4678 -5050 5047 -5002
rect 4679 -5153 4745 -5050
rect 5033 -5080 5047 -5050
rect 5037 -5097 5047 -5080
rect 5159 -5097 5169 -4991
rect 53 -5233 4747 -5153
rect 6611 -5157 6677 -4878
rect 7456 -4958 7466 -4850
rect 7598 -4958 7608 -4850
rect 9354 -4958 9364 -4850
rect 9496 -4958 9506 -4850
rect 10979 -4802 11110 -4754
rect 11187 -4802 11193 -4450
rect 10979 -4826 11193 -4802
rect 11227 -4826 11233 -4450
rect 10979 -4838 11233 -4826
rect 11305 -4450 11351 -4438
rect 11305 -4826 11311 -4450
rect 11345 -4826 11351 -4450
rect 11305 -4838 11351 -4826
rect 11423 -4450 11469 -4438
rect 11423 -4826 11429 -4450
rect 11463 -4826 11469 -4450
rect 11423 -4838 11469 -4826
rect 10979 -4842 11227 -4838
rect 12128 -4840 12221 -3666
rect 12927 -3919 13083 -3913
rect 12927 -4017 12939 -3919
rect 13071 -4017 13083 -3919
rect 12927 -4023 13083 -4017
rect 11636 -4842 12221 -4840
rect 10979 -4886 11053 -4842
rect 11591 -4870 12221 -4842
rect 11236 -4876 11302 -4870
rect 10871 -4896 10979 -4886
rect 11236 -4910 11252 -4876
rect 11286 -4910 11302 -4876
rect 11236 -5006 11302 -4910
rect 11354 -4876 12221 -4870
rect 13144 -4873 13211 -3490
rect 13292 -4061 13326 -3278
rect 13995 -3340 14029 -3278
rect 13698 -3378 14440 -3340
rect 13698 -3502 13732 -3378
rect 13934 -3502 13968 -3378
rect 14170 -3502 14204 -3378
rect 14406 -3502 14440 -3378
rect 13692 -3514 13738 -3502
rect 13692 -3890 13698 -3514
rect 13732 -3890 13738 -3514
rect 13692 -3902 13738 -3890
rect 13810 -3514 13856 -3502
rect 13810 -3890 13816 -3514
rect 13850 -3890 13856 -3514
rect 13810 -3902 13856 -3890
rect 13928 -3514 13974 -3502
rect 13928 -3890 13934 -3514
rect 13968 -3890 13974 -3514
rect 13928 -3902 13974 -3890
rect 14046 -3514 14092 -3502
rect 14046 -3890 14052 -3514
rect 14086 -3890 14092 -3514
rect 14046 -3902 14092 -3890
rect 14164 -3514 14210 -3502
rect 14164 -3890 14170 -3514
rect 14204 -3890 14210 -3514
rect 14164 -3902 14210 -3890
rect 14282 -3514 14328 -3502
rect 14282 -3890 14288 -3514
rect 14322 -3890 14328 -3514
rect 14282 -3902 14328 -3890
rect 14400 -3514 14446 -3502
rect 14400 -3890 14406 -3514
rect 14440 -3890 14446 -3514
rect 14400 -3902 14446 -3890
rect 13292 -4062 13599 -4061
rect 13645 -4062 13714 -4061
rect 14708 -4062 14742 -3278
rect 13292 -4066 13714 -4062
rect 13292 -4077 13781 -4066
rect 14426 -4067 14742 -4062
rect 13292 -4105 13730 -4077
rect 13292 -4106 13599 -4105
rect 13292 -4234 13326 -4106
rect 13714 -4111 13730 -4105
rect 13764 -4111 13781 -4077
rect 13714 -4117 13781 -4111
rect 14359 -4078 14742 -4067
rect 14359 -4112 14376 -4078
rect 14410 -4105 14742 -4078
rect 14410 -4112 14426 -4105
rect 14359 -4118 14426 -4112
rect 13432 -4146 13488 -4134
rect 14545 -4145 14601 -4133
rect 14545 -4146 14561 -4145
rect 13432 -4180 13438 -4146
rect 13472 -4161 14042 -4146
rect 13472 -4180 13992 -4161
rect 13432 -4195 13992 -4180
rect 14026 -4195 14042 -4161
rect 13432 -4196 13488 -4195
rect 13975 -4205 14042 -4195
rect 14094 -4162 14561 -4146
rect 14094 -4196 14110 -4162
rect 14144 -4179 14561 -4162
rect 14595 -4179 14601 -4145
rect 14144 -4195 14601 -4179
rect 14144 -4196 14160 -4195
rect 14094 -4203 14160 -4196
rect 14708 -4234 14742 -4105
rect 15190 -4061 15224 -3278
rect 15893 -3340 15927 -3278
rect 15596 -3378 16338 -3340
rect 15257 -3485 15267 -3419
rect 15330 -3485 15340 -3419
rect 15596 -3502 15630 -3378
rect 15832 -3502 15866 -3378
rect 16068 -3502 16102 -3378
rect 16304 -3502 16338 -3378
rect 15590 -3514 15636 -3502
rect 15590 -3890 15596 -3514
rect 15630 -3890 15636 -3514
rect 15590 -3902 15636 -3890
rect 15708 -3514 15754 -3502
rect 15708 -3890 15714 -3514
rect 15748 -3890 15754 -3514
rect 15708 -3902 15754 -3890
rect 15826 -3514 15872 -3502
rect 15826 -3890 15832 -3514
rect 15866 -3890 15872 -3514
rect 15826 -3902 15872 -3890
rect 15944 -3514 15990 -3502
rect 15944 -3890 15950 -3514
rect 15984 -3890 15990 -3514
rect 15944 -3902 15990 -3890
rect 16062 -3514 16108 -3502
rect 16062 -3890 16068 -3514
rect 16102 -3890 16108 -3514
rect 16062 -3902 16108 -3890
rect 16180 -3514 16226 -3502
rect 16180 -3890 16186 -3514
rect 16220 -3890 16226 -3514
rect 16180 -3902 16226 -3890
rect 16298 -3514 16344 -3502
rect 16298 -3890 16304 -3514
rect 16338 -3890 16344 -3514
rect 16298 -3902 16344 -3890
rect 15190 -4062 15497 -4061
rect 16606 -4062 16640 -3278
rect 17400 -3287 17508 -3277
rect 17765 -3301 17781 -3267
rect 17815 -3301 17831 -3267
rect 17765 -3397 17831 -3301
rect 17883 -3267 18135 -3261
rect 17883 -3301 17899 -3267
rect 17933 -3301 18135 -3267
rect 17883 -3317 18135 -3301
rect 18120 -3319 18135 -3317
rect 18253 -3319 18263 -3201
rect 18120 -3333 18220 -3319
rect 18120 -3376 18220 -3375
rect 18494 -3376 18599 -2199
rect 18120 -3397 18599 -3376
rect 17765 -3445 18599 -3397
rect 18120 -3474 18599 -3445
rect 18120 -3475 18220 -3474
rect 18494 -3476 18599 -3474
rect 18662 -3582 18755 -1688
rect 18895 -1689 19184 -1688
rect 18878 -2099 19167 -1937
rect 18878 -2112 18918 -2099
rect 18876 -2205 18918 -2112
rect 19030 -2205 19167 -2099
rect 18876 -2216 19167 -2205
rect 18878 -2217 19167 -2216
rect 19477 -3049 19578 -1308
rect 20472 -1446 20506 -1300
rect 20656 -1315 20753 -1300
rect 21226 -1303 21261 -1211
rect 20696 -1382 20753 -1315
rect 21034 -1339 21261 -1303
rect 21034 -1373 21100 -1339
rect 20590 -1418 20859 -1382
rect 21034 -1407 21050 -1373
rect 21084 -1407 21100 -1373
rect 21034 -1413 21100 -1407
rect 20590 -1446 20623 -1418
rect 20826 -1446 20859 -1418
rect 21226 -1446 21261 -1339
rect 20466 -1458 20512 -1446
rect 20466 -1634 20472 -1458
rect 20506 -1634 20512 -1458
rect 20466 -1646 20512 -1634
rect 20584 -1458 20630 -1446
rect 20584 -1634 20590 -1458
rect 20624 -1634 20630 -1458
rect 20584 -1646 20630 -1634
rect 20702 -1458 20748 -1446
rect 20702 -1634 20708 -1458
rect 20742 -1634 20748 -1458
rect 20702 -1646 20748 -1634
rect 20820 -1458 20866 -1446
rect 20820 -1634 20826 -1458
rect 20860 -1513 20866 -1458
rect 20985 -1458 21031 -1446
rect 20985 -1513 20991 -1458
rect 20860 -1601 20991 -1513
rect 20860 -1634 20866 -1601
rect 20820 -1646 20866 -1634
rect 20985 -1634 20991 -1601
rect 21025 -1634 21031 -1458
rect 20985 -1646 21031 -1634
rect 21103 -1458 21149 -1446
rect 21103 -1634 21109 -1458
rect 21143 -1634 21149 -1458
rect 21103 -1646 21149 -1634
rect 21221 -1458 21267 -1446
rect 21221 -1634 21227 -1458
rect 21261 -1634 21267 -1458
rect 21221 -1646 21267 -1634
rect 21339 -1458 21385 -1446
rect 21339 -1634 21345 -1458
rect 21379 -1634 21385 -1458
rect 21339 -1646 21385 -1634
rect 20473 -1684 20506 -1646
rect 20709 -1684 20742 -1646
rect 20473 -1720 20742 -1684
rect 21109 -1685 21143 -1646
rect 21345 -1685 21379 -1646
rect 21109 -1721 21379 -1685
rect 21213 -1722 21379 -1721
rect 21213 -1801 21345 -1722
rect 21203 -1909 21213 -1801
rect 21345 -1909 21355 -1801
rect 21485 -2238 21547 -667
rect 21683 -679 21729 -667
rect 21683 -1055 21689 -679
rect 21723 -1055 21729 -679
rect 21683 -1067 21729 -1055
rect 21801 -679 21847 -667
rect 21801 -1055 21807 -679
rect 21841 -1055 21847 -679
rect 21801 -1067 21847 -1055
rect 21919 -679 21965 -667
rect 21919 -1055 21925 -679
rect 21959 -1055 21965 -679
rect 21919 -1067 21965 -1055
rect 22037 -679 22083 -667
rect 22037 -1055 22043 -679
rect 22077 -1055 22083 -679
rect 22037 -1067 22083 -1055
rect 22155 -679 22201 -667
rect 22155 -1055 22161 -679
rect 22195 -1055 22201 -679
rect 22155 -1067 22201 -1055
rect 22273 -679 22319 -667
rect 22273 -1055 22279 -679
rect 22313 -1055 22319 -679
rect 22273 -1067 22319 -1055
rect 22391 -679 22437 -667
rect 22486 -671 22496 -605
rect 22562 -671 22572 -605
rect 22391 -1055 22397 -679
rect 22431 -1055 22437 -679
rect 22391 -1067 22437 -1055
rect 21689 -1250 21723 -1067
rect 21807 -1108 21841 -1067
rect 22043 -1108 22077 -1067
rect 21807 -1137 22077 -1108
rect 22161 -1109 22195 -1067
rect 22397 -1109 22431 -1067
rect 22161 -1137 22431 -1109
rect 22397 -1185 22431 -1137
rect 22368 -1215 22431 -1185
rect 23421 -1144 23488 -554
rect 24139 -561 24183 -453
rect 24315 -561 24359 -453
rect 24139 -603 24359 -561
rect 23778 -633 24755 -603
rect 23778 -739 23812 -633
rect 24015 -739 24047 -633
rect 24251 -739 24283 -633
rect 24487 -739 24519 -633
rect 24723 -739 24755 -633
rect 23654 -751 23700 -739
rect 23654 -927 23660 -751
rect 23694 -927 23700 -751
rect 23654 -939 23700 -927
rect 23772 -751 23818 -739
rect 23772 -927 23778 -751
rect 23812 -927 23818 -751
rect 23772 -939 23818 -927
rect 23890 -751 23936 -739
rect 23890 -927 23896 -751
rect 23930 -927 23936 -751
rect 23890 -939 23936 -927
rect 24008 -751 24054 -739
rect 24008 -927 24014 -751
rect 24048 -927 24054 -751
rect 24008 -939 24054 -927
rect 24126 -751 24172 -739
rect 24126 -927 24132 -751
rect 24166 -927 24172 -751
rect 24126 -939 24172 -927
rect 24244 -751 24290 -739
rect 24244 -927 24250 -751
rect 24284 -927 24290 -751
rect 24244 -939 24290 -927
rect 24362 -751 24408 -739
rect 24362 -927 24368 -751
rect 24402 -927 24408 -751
rect 24362 -939 24408 -927
rect 24480 -751 24526 -739
rect 24480 -927 24486 -751
rect 24520 -927 24526 -751
rect 24480 -939 24526 -927
rect 24598 -751 24644 -739
rect 24598 -927 24604 -751
rect 24638 -927 24644 -751
rect 24598 -939 24644 -927
rect 24716 -751 24762 -739
rect 24716 -927 24722 -751
rect 24756 -927 24762 -751
rect 24716 -939 24762 -927
rect 23660 -1144 23695 -939
rect 23939 -987 24005 -980
rect 23939 -1021 23955 -987
rect 23989 -1021 24005 -987
rect 23939 -1032 24005 -1021
rect 24131 -1032 24167 -939
rect 23939 -1033 24167 -1032
rect 24367 -1033 24403 -939
rect 24603 -1033 24639 -939
rect 23939 -1062 24639 -1033
rect 23421 -1172 23695 -1144
rect 24057 -1063 24639 -1062
rect 24057 -1104 24123 -1063
rect 24057 -1138 24073 -1104
rect 24107 -1138 24123 -1104
rect 24057 -1145 24123 -1138
rect 23421 -1176 24049 -1172
rect 24485 -1176 24519 -1063
rect 23421 -1188 24054 -1176
rect 23421 -1201 24014 -1188
rect 21614 -1304 21723 -1250
rect 21614 -1450 21648 -1304
rect 21787 -1318 21797 -1221
rect 21896 -1318 21906 -1221
rect 22368 -1307 22403 -1215
rect 21798 -1319 21895 -1318
rect 21838 -1386 21895 -1319
rect 22176 -1343 22403 -1307
rect 22176 -1377 22242 -1343
rect 21732 -1422 22001 -1386
rect 22176 -1411 22192 -1377
rect 22226 -1411 22242 -1377
rect 22176 -1417 22242 -1411
rect 21732 -1450 21765 -1422
rect 21968 -1450 22001 -1422
rect 22368 -1450 22403 -1343
rect 24008 -1364 24014 -1201
rect 24048 -1364 24054 -1188
rect 24008 -1376 24054 -1364
rect 24126 -1188 24172 -1176
rect 24126 -1364 24132 -1188
rect 24166 -1364 24172 -1188
rect 24126 -1376 24172 -1364
rect 24243 -1188 24289 -1176
rect 21608 -1462 21654 -1450
rect 21608 -1638 21614 -1462
rect 21648 -1638 21654 -1462
rect 21608 -1650 21654 -1638
rect 21726 -1462 21772 -1450
rect 21726 -1638 21732 -1462
rect 21766 -1638 21772 -1462
rect 21726 -1650 21772 -1638
rect 21844 -1462 21890 -1450
rect 21844 -1638 21850 -1462
rect 21884 -1638 21890 -1462
rect 21844 -1650 21890 -1638
rect 21962 -1462 22008 -1450
rect 21962 -1638 21968 -1462
rect 22002 -1517 22008 -1462
rect 22127 -1462 22173 -1450
rect 22127 -1517 22133 -1462
rect 22002 -1605 22133 -1517
rect 22002 -1638 22008 -1605
rect 21962 -1650 22008 -1638
rect 22127 -1638 22133 -1605
rect 22167 -1638 22173 -1462
rect 22127 -1650 22173 -1638
rect 22245 -1462 22291 -1450
rect 22245 -1638 22251 -1462
rect 22285 -1638 22291 -1462
rect 22245 -1650 22291 -1638
rect 22363 -1462 22409 -1450
rect 22363 -1638 22369 -1462
rect 22403 -1638 22409 -1462
rect 22363 -1650 22409 -1638
rect 22481 -1462 22527 -1450
rect 22481 -1638 22487 -1462
rect 22521 -1638 22527 -1462
rect 23927 -1492 24035 -1482
rect 24131 -1492 24166 -1376
rect 24035 -1540 24166 -1492
rect 24243 -1540 24249 -1188
rect 24035 -1564 24249 -1540
rect 24283 -1564 24289 -1188
rect 24035 -1576 24289 -1564
rect 24361 -1188 24407 -1176
rect 24361 -1564 24367 -1188
rect 24401 -1564 24407 -1188
rect 24361 -1576 24407 -1564
rect 24479 -1188 24525 -1176
rect 24479 -1564 24485 -1188
rect 24519 -1564 24525 -1188
rect 24479 -1576 24525 -1564
rect 24035 -1580 24283 -1576
rect 24035 -1624 24109 -1580
rect 25408 -1581 25697 -1406
rect 24647 -1608 25697 -1581
rect 24292 -1614 24358 -1608
rect 23927 -1634 24035 -1624
rect 22481 -1650 22527 -1638
rect 24292 -1648 24308 -1614
rect 24342 -1648 24358 -1614
rect 21615 -1688 21648 -1650
rect 21851 -1688 21884 -1650
rect 21615 -1724 21884 -1688
rect 22251 -1689 22285 -1650
rect 22487 -1689 22521 -1650
rect 22251 -1724 22521 -1689
rect 22251 -1725 22487 -1724
rect 22355 -1799 22487 -1725
rect 24292 -1744 24358 -1648
rect 24410 -1614 25697 -1608
rect 24410 -1648 24426 -1614
rect 24460 -1648 25697 -1614
rect 24410 -1664 25697 -1648
rect 24647 -1680 25697 -1664
rect 24710 -1681 25697 -1680
rect 25175 -1685 25697 -1681
rect 24646 -1744 25112 -1722
rect 24292 -1792 25112 -1744
rect 22345 -1907 22355 -1799
rect 22487 -1907 22497 -1799
rect 24646 -1823 25112 -1792
rect 25007 -2079 25112 -1823
rect 21484 -2255 21547 -2238
rect 24125 -2103 24345 -2083
rect 24125 -2211 24169 -2103
rect 24301 -2211 24345 -2103
rect 24927 -2185 24937 -2079
rect 25049 -2185 25112 -2079
rect 24963 -2196 25112 -2185
rect 24125 -2253 24345 -2211
rect 21484 -2259 21622 -2255
rect 21484 -2293 23454 -2259
rect 23764 -2283 24741 -2253
rect 21484 -2322 23456 -2293
rect 21484 -2324 21622 -2322
rect 23410 -2338 23456 -2322
rect 20448 -2554 20458 -2446
rect 20590 -2554 20600 -2446
rect 22346 -2554 22356 -2446
rect 22488 -2554 22498 -2446
rect 20458 -2594 20590 -2554
rect 22356 -2594 22488 -2554
rect 20458 -2660 20591 -2594
rect 22356 -2660 22489 -2594
rect 19789 -2703 21262 -2660
rect 19789 -3006 19823 -2703
rect 20154 -2806 20188 -2703
rect 20390 -2806 20424 -2703
rect 20626 -2806 20660 -2703
rect 20862 -2806 20896 -2703
rect 20148 -2818 20194 -2806
rect 18879 -3151 19578 -3049
rect 19665 -3018 19711 -3006
rect 18879 -3211 19167 -3151
rect 19665 -3194 19671 -3018
rect 19705 -3194 19711 -3018
rect 19665 -3206 19711 -3194
rect 19783 -3018 19829 -3006
rect 19783 -3194 19789 -3018
rect 19823 -3194 19829 -3018
rect 19783 -3206 19829 -3194
rect 19901 -3018 19947 -3006
rect 19901 -3194 19907 -3018
rect 19941 -3194 19947 -3018
rect 19901 -3206 19947 -3194
rect 20019 -3018 20065 -3006
rect 20148 -3018 20154 -2818
rect 20019 -3194 20025 -3018
rect 20059 -3194 20154 -3018
rect 20188 -3194 20194 -2818
rect 20019 -3206 20065 -3194
rect 20148 -3206 20194 -3194
rect 20266 -2818 20312 -2806
rect 20266 -3194 20272 -2818
rect 20306 -3194 20312 -2818
rect 20266 -3206 20312 -3194
rect 20384 -2818 20430 -2806
rect 20384 -3194 20390 -2818
rect 20424 -3194 20430 -2818
rect 20384 -3206 20430 -3194
rect 20502 -2818 20548 -2806
rect 20502 -3194 20508 -2818
rect 20542 -3194 20548 -2818
rect 20502 -3206 20548 -3194
rect 20620 -2818 20666 -2806
rect 20620 -3194 20626 -2818
rect 20660 -3194 20666 -2818
rect 20620 -3206 20666 -3194
rect 20738 -2818 20784 -2806
rect 20738 -3194 20744 -2818
rect 20778 -3194 20784 -2818
rect 20738 -3206 20784 -3194
rect 20856 -2818 20902 -2806
rect 20856 -3194 20862 -2818
rect 20896 -3018 20902 -2818
rect 21228 -3006 21262 -2703
rect 21687 -2703 23160 -2660
rect 21687 -3006 21721 -2703
rect 22052 -2806 22086 -2703
rect 22288 -2806 22322 -2703
rect 22524 -2806 22558 -2703
rect 22760 -2806 22794 -2703
rect 22046 -2818 22092 -2806
rect 20986 -3018 21032 -3006
rect 20896 -3194 20992 -3018
rect 21026 -3194 21032 -3018
rect 20856 -3206 20902 -3194
rect 20986 -3206 21032 -3194
rect 21104 -3018 21150 -3006
rect 21104 -3194 21110 -3018
rect 21144 -3194 21150 -3018
rect 21104 -3206 21150 -3194
rect 21222 -3018 21268 -3006
rect 21222 -3194 21228 -3018
rect 21262 -3194 21268 -3018
rect 21222 -3206 21268 -3194
rect 21340 -3018 21386 -3006
rect 21340 -3194 21346 -3018
rect 21380 -3194 21386 -3018
rect 21340 -3206 21386 -3194
rect 21563 -3018 21609 -3006
rect 21563 -3194 21569 -3018
rect 21603 -3194 21609 -3018
rect 21563 -3206 21609 -3194
rect 21681 -3018 21727 -3006
rect 21681 -3194 21687 -3018
rect 21721 -3194 21727 -3018
rect 21681 -3206 21727 -3194
rect 21799 -3018 21845 -3006
rect 21799 -3194 21805 -3018
rect 21839 -3194 21845 -3018
rect 21799 -3206 21845 -3194
rect 21917 -3018 21963 -3006
rect 22046 -3018 22052 -2818
rect 21917 -3194 21923 -3018
rect 21957 -3194 22052 -3018
rect 22086 -3194 22092 -2818
rect 21917 -3206 21963 -3194
rect 22046 -3206 22092 -3194
rect 22164 -2818 22210 -2806
rect 22164 -3194 22170 -2818
rect 22204 -3194 22210 -2818
rect 22164 -3206 22210 -3194
rect 22282 -2818 22328 -2806
rect 22282 -3194 22288 -2818
rect 22322 -3194 22328 -2818
rect 22282 -3206 22328 -3194
rect 22400 -2818 22446 -2806
rect 22400 -3194 22406 -2818
rect 22440 -3194 22446 -2818
rect 22400 -3206 22446 -3194
rect 22518 -2818 22564 -2806
rect 22518 -3194 22524 -2818
rect 22558 -3194 22564 -2818
rect 22518 -3206 22564 -3194
rect 22636 -2818 22682 -2806
rect 22636 -3194 22642 -2818
rect 22676 -3194 22682 -2818
rect 22636 -3206 22682 -3194
rect 22754 -2818 22800 -2806
rect 22754 -3194 22760 -2818
rect 22794 -3018 22800 -2818
rect 23126 -3006 23160 -2703
rect 23410 -2790 23457 -2338
rect 23764 -2389 23798 -2283
rect 24001 -2389 24033 -2283
rect 24237 -2389 24269 -2283
rect 24473 -2389 24505 -2283
rect 24709 -2389 24741 -2283
rect 23640 -2401 23686 -2389
rect 23640 -2577 23646 -2401
rect 23680 -2577 23686 -2401
rect 23640 -2589 23686 -2577
rect 23758 -2401 23804 -2389
rect 23758 -2577 23764 -2401
rect 23798 -2577 23804 -2401
rect 23758 -2589 23804 -2577
rect 23876 -2401 23922 -2389
rect 23876 -2577 23882 -2401
rect 23916 -2577 23922 -2401
rect 23876 -2589 23922 -2577
rect 23994 -2401 24040 -2389
rect 23994 -2577 24000 -2401
rect 24034 -2577 24040 -2401
rect 23994 -2589 24040 -2577
rect 24112 -2401 24158 -2389
rect 24112 -2577 24118 -2401
rect 24152 -2577 24158 -2401
rect 24112 -2589 24158 -2577
rect 24230 -2401 24276 -2389
rect 24230 -2577 24236 -2401
rect 24270 -2577 24276 -2401
rect 24230 -2589 24276 -2577
rect 24348 -2401 24394 -2389
rect 24348 -2577 24354 -2401
rect 24388 -2577 24394 -2401
rect 24348 -2589 24394 -2577
rect 24466 -2401 24512 -2389
rect 24466 -2577 24472 -2401
rect 24506 -2577 24512 -2401
rect 24466 -2589 24512 -2577
rect 24584 -2401 24630 -2389
rect 24584 -2577 24590 -2401
rect 24624 -2577 24630 -2401
rect 24584 -2589 24630 -2577
rect 24702 -2401 24748 -2389
rect 24702 -2577 24708 -2401
rect 24742 -2577 24748 -2401
rect 24702 -2589 24748 -2577
rect 23411 -2806 23457 -2790
rect 23411 -2807 23492 -2806
rect 23646 -2807 23681 -2589
rect 23925 -2637 23991 -2630
rect 23925 -2671 23941 -2637
rect 23975 -2671 23991 -2637
rect 23925 -2682 23991 -2671
rect 24117 -2682 24153 -2589
rect 23925 -2683 24153 -2682
rect 24353 -2683 24389 -2589
rect 24589 -2683 24625 -2589
rect 23925 -2712 24625 -2683
rect 24043 -2713 24625 -2712
rect 24043 -2754 24109 -2713
rect 24043 -2788 24059 -2754
rect 24093 -2788 24109 -2754
rect 24043 -2795 24109 -2788
rect 23411 -2822 23681 -2807
rect 23411 -2826 24035 -2822
rect 24471 -2826 24505 -2713
rect 23411 -2838 24040 -2826
rect 23411 -2850 24000 -2838
rect 23411 -2852 23492 -2850
rect 23758 -2851 24000 -2850
rect 22884 -3018 22930 -3006
rect 22794 -3194 22890 -3018
rect 22924 -3194 22930 -3018
rect 22754 -3206 22800 -3194
rect 22884 -3206 22930 -3194
rect 23002 -3018 23048 -3006
rect 23002 -3194 23008 -3018
rect 23042 -3194 23048 -3018
rect 23002 -3206 23048 -3194
rect 23120 -3018 23166 -3006
rect 23120 -3194 23126 -3018
rect 23160 -3194 23166 -3018
rect 23120 -3206 23166 -3194
rect 23238 -3018 23284 -3006
rect 23238 -3194 23244 -3018
rect 23278 -3194 23284 -3018
rect 23994 -3014 24000 -2851
rect 24034 -3014 24040 -2838
rect 23994 -3026 24040 -3014
rect 24112 -2838 24158 -2826
rect 24112 -3014 24118 -2838
rect 24152 -3014 24158 -2838
rect 24112 -3026 24158 -3014
rect 24229 -2838 24275 -2826
rect 23238 -3206 23284 -3194
rect 23913 -3142 24021 -3132
rect 24117 -3142 24152 -3026
rect 18879 -3213 18919 -3211
rect 18879 -3224 18913 -3213
rect 18878 -3319 18913 -3224
rect 19031 -3317 19167 -3211
rect 19671 -3240 19705 -3206
rect 19907 -3240 19941 -3206
rect 19671 -3275 19941 -3240
rect 20508 -3240 20542 -3206
rect 20744 -3240 20778 -3206
rect 21346 -3240 21380 -3206
rect 20508 -3275 20778 -3240
rect 21221 -3275 21380 -3240
rect 21569 -3240 21603 -3206
rect 21805 -3240 21839 -3206
rect 21569 -3275 21839 -3240
rect 22406 -3240 22440 -3206
rect 22642 -3240 22676 -3206
rect 23244 -3240 23278 -3206
rect 22406 -3275 22676 -3240
rect 23119 -3275 23278 -3240
rect 24021 -3190 24152 -3142
rect 24229 -3190 24235 -2838
rect 24021 -3214 24235 -3190
rect 24269 -3214 24275 -2838
rect 24021 -3226 24275 -3214
rect 24347 -2838 24393 -2826
rect 24347 -3214 24353 -2838
rect 24387 -3214 24393 -2838
rect 24347 -3226 24393 -3214
rect 24465 -2838 24511 -2826
rect 24465 -3214 24471 -2838
rect 24505 -3214 24511 -2838
rect 24465 -3226 24511 -3214
rect 24021 -3230 24269 -3226
rect 24638 -3230 24648 -3198
rect 24021 -3274 24095 -3230
rect 24633 -3258 24648 -3230
rect 24278 -3264 24344 -3258
rect 19025 -3319 19167 -3317
rect 18878 -3328 19167 -3319
rect 18879 -3329 19167 -3328
rect 18911 -3330 19167 -3329
rect 19657 -3453 19724 -3429
rect 19657 -3487 19673 -3453
rect 19707 -3487 19724 -3453
rect 18653 -3661 18663 -3582
rect 18756 -3661 18766 -3582
rect 17617 -3710 17837 -3690
rect 17617 -3818 17661 -3710
rect 17793 -3818 17837 -3710
rect 17617 -3860 17837 -3818
rect 17256 -3890 18233 -3860
rect 17256 -3996 17290 -3890
rect 17493 -3996 17525 -3890
rect 17729 -3996 17761 -3890
rect 17965 -3996 17997 -3890
rect 18201 -3996 18233 -3890
rect 15190 -4067 15610 -4062
rect 16324 -4067 16640 -4062
rect 15190 -4078 15677 -4067
rect 15190 -4105 15626 -4078
rect 15190 -4106 15497 -4105
rect 15190 -4234 15224 -4106
rect 15610 -4112 15626 -4105
rect 15660 -4112 15677 -4078
rect 15610 -4118 15677 -4112
rect 16257 -4078 16640 -4067
rect 16257 -4112 16274 -4078
rect 16308 -4105 16640 -4078
rect 16308 -4112 16324 -4105
rect 16257 -4118 16324 -4112
rect 15330 -4146 15386 -4134
rect 16443 -4145 16499 -4133
rect 16443 -4146 16459 -4145
rect 15330 -4180 15336 -4146
rect 15370 -4161 15940 -4146
rect 15370 -4180 15890 -4161
rect 15330 -4195 15890 -4180
rect 15924 -4195 15940 -4161
rect 15330 -4196 15386 -4195
rect 15873 -4205 15940 -4195
rect 15992 -4162 16459 -4146
rect 15992 -4196 16008 -4162
rect 16042 -4179 16459 -4162
rect 16493 -4179 16499 -4145
rect 16042 -4195 16499 -4179
rect 16042 -4196 16058 -4195
rect 15992 -4203 16058 -4196
rect 16606 -4234 16640 -4105
rect 17132 -4008 17178 -3996
rect 17132 -4184 17138 -4008
rect 17172 -4184 17178 -4008
rect 17132 -4196 17178 -4184
rect 17250 -4008 17296 -3996
rect 17250 -4184 17256 -4008
rect 17290 -4184 17296 -4008
rect 17250 -4196 17296 -4184
rect 17368 -4008 17414 -3996
rect 17368 -4184 17374 -4008
rect 17408 -4184 17414 -4008
rect 17368 -4196 17414 -4184
rect 17486 -4008 17532 -3996
rect 17486 -4184 17492 -4008
rect 17526 -4184 17532 -4008
rect 17486 -4196 17532 -4184
rect 17604 -4008 17650 -3996
rect 17604 -4184 17610 -4008
rect 17644 -4184 17650 -4008
rect 17604 -4196 17650 -4184
rect 17722 -4008 17768 -3996
rect 17722 -4184 17728 -4008
rect 17762 -4184 17768 -4008
rect 17722 -4196 17768 -4184
rect 17840 -4008 17886 -3996
rect 17840 -4184 17846 -4008
rect 17880 -4184 17886 -4008
rect 17840 -4196 17886 -4184
rect 17958 -4008 18004 -3996
rect 17958 -4184 17964 -4008
rect 17998 -4184 18004 -4008
rect 17958 -4196 18004 -4184
rect 18076 -4008 18122 -3996
rect 18076 -4184 18082 -4008
rect 18116 -4184 18122 -4008
rect 18076 -4196 18122 -4184
rect 18194 -4008 18240 -3996
rect 18194 -4184 18200 -4008
rect 18234 -4184 18240 -4008
rect 18194 -4196 18240 -4184
rect 13286 -4246 13332 -4234
rect 13286 -4422 13292 -4246
rect 13326 -4422 13332 -4246
rect 13286 -4434 13332 -4422
rect 13404 -4246 13450 -4234
rect 13404 -4422 13410 -4246
rect 13444 -4422 13450 -4246
rect 13404 -4434 13450 -4422
rect 13810 -4246 13856 -4234
rect 13411 -4728 13444 -4434
rect 13810 -4622 13816 -4246
rect 13850 -4622 13856 -4246
rect 13810 -4634 13856 -4622
rect 13928 -4246 13974 -4234
rect 13928 -4622 13934 -4246
rect 13968 -4622 13974 -4246
rect 13928 -4634 13974 -4622
rect 14046 -4246 14092 -4234
rect 14046 -4622 14052 -4246
rect 14086 -4622 14092 -4246
rect 14046 -4634 14092 -4622
rect 14164 -4246 14210 -4234
rect 14164 -4622 14170 -4246
rect 14204 -4622 14210 -4246
rect 14164 -4634 14210 -4622
rect 14282 -4246 14328 -4234
rect 14282 -4622 14288 -4246
rect 14322 -4622 14328 -4246
rect 14584 -4246 14630 -4234
rect 14584 -4422 14590 -4246
rect 14624 -4422 14630 -4246
rect 14584 -4434 14630 -4422
rect 14702 -4246 14748 -4234
rect 14702 -4422 14708 -4246
rect 14742 -4422 14748 -4246
rect 14702 -4434 14748 -4422
rect 15184 -4246 15230 -4234
rect 15184 -4422 15190 -4246
rect 15224 -4422 15230 -4246
rect 15184 -4434 15230 -4422
rect 15302 -4246 15348 -4234
rect 15302 -4422 15308 -4246
rect 15342 -4422 15348 -4246
rect 15302 -4434 15348 -4422
rect 15708 -4246 15754 -4234
rect 14282 -4634 14328 -4622
rect 13934 -4728 13968 -4634
rect 14591 -4728 14625 -4434
rect 13411 -4760 14625 -4728
rect 15309 -4728 15342 -4434
rect 15708 -4622 15714 -4246
rect 15748 -4622 15754 -4246
rect 15708 -4634 15754 -4622
rect 15826 -4246 15872 -4234
rect 15826 -4622 15832 -4246
rect 15866 -4622 15872 -4246
rect 15826 -4634 15872 -4622
rect 15944 -4246 15990 -4234
rect 15944 -4622 15950 -4246
rect 15984 -4622 15990 -4246
rect 15944 -4634 15990 -4622
rect 16062 -4246 16108 -4234
rect 16062 -4622 16068 -4246
rect 16102 -4622 16108 -4246
rect 16062 -4634 16108 -4622
rect 16180 -4246 16226 -4234
rect 16180 -4622 16186 -4246
rect 16220 -4622 16226 -4246
rect 16482 -4246 16528 -4234
rect 16482 -4422 16488 -4246
rect 16522 -4422 16528 -4246
rect 16482 -4434 16528 -4422
rect 16600 -4246 16646 -4234
rect 16600 -4422 16606 -4246
rect 16640 -4422 16646 -4246
rect 16600 -4434 16646 -4422
rect 17138 -4429 17173 -4196
rect 17417 -4244 17483 -4237
rect 17417 -4278 17433 -4244
rect 17467 -4278 17483 -4244
rect 17417 -4289 17483 -4278
rect 17609 -4289 17645 -4196
rect 17417 -4290 17645 -4289
rect 17845 -4290 17881 -4196
rect 18081 -4290 18117 -4196
rect 17417 -4319 18117 -4290
rect 17535 -4320 18117 -4319
rect 17535 -4361 17601 -4320
rect 17535 -4395 17551 -4361
rect 17585 -4395 17601 -4361
rect 17535 -4402 17601 -4395
rect 17138 -4433 17527 -4429
rect 17963 -4433 17997 -4320
rect 16180 -4634 16226 -4622
rect 15832 -4728 15866 -4634
rect 16489 -4728 16523 -4434
rect 17138 -4445 17532 -4433
rect 17138 -4458 17492 -4445
rect 17138 -4461 17216 -4458
rect 17133 -4513 17143 -4461
rect 17206 -4513 17216 -4461
rect 17138 -4519 17211 -4513
rect 17486 -4621 17492 -4458
rect 17526 -4621 17532 -4445
rect 17486 -4633 17532 -4621
rect 17604 -4445 17650 -4433
rect 17604 -4621 17610 -4445
rect 17644 -4621 17650 -4445
rect 17604 -4633 17650 -4621
rect 17721 -4445 17767 -4433
rect 15309 -4760 16523 -4728
rect 17405 -4749 17513 -4739
rect 17609 -4749 17644 -4633
rect 14000 -4845 14132 -4760
rect 15898 -4845 16030 -4760
rect 11354 -4910 11370 -4876
rect 11404 -4910 12221 -4876
rect 11354 -4926 12221 -4910
rect 11591 -4942 12221 -4926
rect 11636 -4946 12221 -4942
rect 12120 -4947 12221 -4946
rect 11591 -4995 11691 -4984
rect 11591 -5006 11605 -4995
rect 11236 -5054 11605 -5006
rect 11237 -5157 11303 -5054
rect 11591 -5084 11605 -5054
rect 11595 -5101 11605 -5084
rect 11717 -5101 11727 -4995
rect 13145 -5152 13211 -4873
rect 13990 -4953 14000 -4845
rect 14132 -4953 14142 -4845
rect 15888 -4953 15898 -4845
rect 16030 -4953 16040 -4845
rect 17513 -4797 17644 -4749
rect 17721 -4797 17727 -4445
rect 17513 -4821 17727 -4797
rect 17761 -4821 17767 -4445
rect 17513 -4833 17767 -4821
rect 17839 -4445 17885 -4433
rect 17839 -4821 17845 -4445
rect 17879 -4821 17885 -4445
rect 17839 -4833 17885 -4821
rect 17957 -4445 18003 -4433
rect 17957 -4821 17963 -4445
rect 17997 -4821 18003 -4445
rect 17957 -4833 18003 -4821
rect 17513 -4837 17761 -4833
rect 18662 -4835 18755 -3661
rect 19440 -3916 19596 -3910
rect 19440 -4014 19452 -3916
rect 19584 -4014 19596 -3916
rect 19440 -4020 19596 -4014
rect 18170 -4837 18755 -4835
rect 17513 -4881 17587 -4837
rect 18125 -4865 18755 -4837
rect 17770 -4871 17836 -4865
rect 17405 -4891 17513 -4881
rect 17770 -4905 17786 -4871
rect 17820 -4905 17836 -4871
rect 17770 -5001 17836 -4905
rect 17888 -4871 18755 -4865
rect 19657 -4870 19724 -3487
rect 19805 -4058 19839 -3275
rect 20508 -3337 20542 -3275
rect 20211 -3375 20953 -3337
rect 20211 -3499 20245 -3375
rect 20447 -3499 20481 -3375
rect 20683 -3499 20717 -3375
rect 20919 -3499 20953 -3375
rect 20205 -3511 20251 -3499
rect 20205 -3887 20211 -3511
rect 20245 -3887 20251 -3511
rect 20205 -3899 20251 -3887
rect 20323 -3511 20369 -3499
rect 20323 -3887 20329 -3511
rect 20363 -3887 20369 -3511
rect 20323 -3899 20369 -3887
rect 20441 -3511 20487 -3499
rect 20441 -3887 20447 -3511
rect 20481 -3887 20487 -3511
rect 20441 -3899 20487 -3887
rect 20559 -3511 20605 -3499
rect 20559 -3887 20565 -3511
rect 20599 -3887 20605 -3511
rect 20559 -3899 20605 -3887
rect 20677 -3511 20723 -3499
rect 20677 -3887 20683 -3511
rect 20717 -3887 20723 -3511
rect 20677 -3899 20723 -3887
rect 20795 -3511 20841 -3499
rect 20795 -3887 20801 -3511
rect 20835 -3887 20841 -3511
rect 20795 -3899 20841 -3887
rect 20913 -3511 20959 -3499
rect 20913 -3887 20919 -3511
rect 20953 -3887 20959 -3511
rect 20913 -3899 20959 -3887
rect 19805 -4059 20112 -4058
rect 20158 -4059 20227 -4058
rect 21221 -4059 21255 -3275
rect 19805 -4063 20227 -4059
rect 19805 -4074 20294 -4063
rect 20939 -4064 21255 -4059
rect 19805 -4102 20243 -4074
rect 19805 -4103 20112 -4102
rect 19805 -4231 19839 -4103
rect 20227 -4108 20243 -4102
rect 20277 -4108 20294 -4074
rect 20227 -4114 20294 -4108
rect 20872 -4075 21255 -4064
rect 20872 -4109 20889 -4075
rect 20923 -4102 21255 -4075
rect 20923 -4109 20939 -4102
rect 20872 -4115 20939 -4109
rect 19945 -4143 20001 -4131
rect 21058 -4142 21114 -4130
rect 21058 -4143 21074 -4142
rect 19945 -4177 19951 -4143
rect 19985 -4158 20555 -4143
rect 19985 -4177 20505 -4158
rect 19945 -4192 20505 -4177
rect 20539 -4192 20555 -4158
rect 19945 -4193 20001 -4192
rect 20488 -4202 20555 -4192
rect 20607 -4159 21074 -4143
rect 20607 -4193 20623 -4159
rect 20657 -4176 21074 -4159
rect 21108 -4176 21114 -4142
rect 20657 -4192 21114 -4176
rect 20657 -4193 20673 -4192
rect 20607 -4200 20673 -4193
rect 21221 -4231 21255 -4102
rect 21703 -4058 21737 -3275
rect 22406 -3337 22440 -3275
rect 22109 -3375 22851 -3337
rect 21770 -3482 21780 -3416
rect 21843 -3482 21853 -3416
rect 22109 -3499 22143 -3375
rect 22345 -3499 22379 -3375
rect 22581 -3499 22615 -3375
rect 22817 -3499 22851 -3375
rect 22103 -3511 22149 -3499
rect 22103 -3887 22109 -3511
rect 22143 -3887 22149 -3511
rect 22103 -3899 22149 -3887
rect 22221 -3511 22267 -3499
rect 22221 -3887 22227 -3511
rect 22261 -3887 22267 -3511
rect 22221 -3899 22267 -3887
rect 22339 -3511 22385 -3499
rect 22339 -3887 22345 -3511
rect 22379 -3887 22385 -3511
rect 22339 -3899 22385 -3887
rect 22457 -3511 22503 -3499
rect 22457 -3887 22463 -3511
rect 22497 -3887 22503 -3511
rect 22457 -3899 22503 -3887
rect 22575 -3511 22621 -3499
rect 22575 -3887 22581 -3511
rect 22615 -3887 22621 -3511
rect 22575 -3899 22621 -3887
rect 22693 -3511 22739 -3499
rect 22693 -3887 22699 -3511
rect 22733 -3887 22739 -3511
rect 22693 -3899 22739 -3887
rect 22811 -3511 22857 -3499
rect 22811 -3887 22817 -3511
rect 22851 -3887 22857 -3511
rect 22811 -3899 22857 -3887
rect 21703 -4059 22010 -4058
rect 23119 -4059 23153 -3275
rect 23913 -3284 24021 -3274
rect 24278 -3298 24294 -3264
rect 24328 -3298 24344 -3264
rect 24278 -3394 24344 -3298
rect 24396 -3264 24648 -3258
rect 24396 -3298 24412 -3264
rect 24446 -3298 24648 -3264
rect 24396 -3314 24648 -3298
rect 24633 -3316 24648 -3314
rect 24766 -3316 24776 -3198
rect 24633 -3330 24733 -3316
rect 24633 -3373 24733 -3372
rect 25007 -3373 25112 -2196
rect 24633 -3394 25112 -3373
rect 24278 -3442 25112 -3394
rect 24633 -3471 25112 -3442
rect 24633 -3472 24733 -3471
rect 25007 -3473 25112 -3471
rect 25175 -3579 25268 -1685
rect 25408 -1686 25697 -1685
rect 25391 -2096 25680 -1934
rect 25391 -2109 25431 -2096
rect 25389 -2202 25431 -2109
rect 25543 -2202 25680 -2096
rect 25389 -2213 25680 -2202
rect 25391 -2214 25680 -2213
rect 25984 -3044 26111 3263
rect 25603 -3046 26111 -3044
rect 25392 -3200 26111 -3046
rect 25392 -3208 25680 -3200
rect 25392 -3210 25432 -3208
rect 25392 -3221 25426 -3210
rect 25391 -3316 25426 -3221
rect 25544 -3314 25680 -3208
rect 25538 -3316 25680 -3314
rect 25391 -3325 25680 -3316
rect 25392 -3326 25680 -3325
rect 25424 -3327 25680 -3326
rect 25166 -3658 25176 -3579
rect 25269 -3658 25279 -3579
rect 24130 -3707 24350 -3687
rect 24130 -3815 24174 -3707
rect 24306 -3815 24350 -3707
rect 24130 -3857 24350 -3815
rect 23769 -3887 24746 -3857
rect 23769 -3993 23803 -3887
rect 24006 -3993 24038 -3887
rect 24242 -3993 24274 -3887
rect 24478 -3993 24510 -3887
rect 24714 -3993 24746 -3887
rect 21703 -4064 22123 -4059
rect 22837 -4064 23153 -4059
rect 21703 -4075 22190 -4064
rect 21703 -4102 22139 -4075
rect 21703 -4103 22010 -4102
rect 21703 -4231 21737 -4103
rect 22123 -4109 22139 -4102
rect 22173 -4109 22190 -4075
rect 22123 -4115 22190 -4109
rect 22770 -4075 23153 -4064
rect 22770 -4109 22787 -4075
rect 22821 -4102 23153 -4075
rect 22821 -4109 22837 -4102
rect 22770 -4115 22837 -4109
rect 21843 -4143 21899 -4131
rect 22956 -4142 23012 -4130
rect 22956 -4143 22972 -4142
rect 21843 -4177 21849 -4143
rect 21883 -4158 22453 -4143
rect 21883 -4177 22403 -4158
rect 21843 -4192 22403 -4177
rect 22437 -4192 22453 -4158
rect 21843 -4193 21899 -4192
rect 22386 -4202 22453 -4192
rect 22505 -4159 22972 -4143
rect 22505 -4193 22521 -4159
rect 22555 -4176 22972 -4159
rect 23006 -4176 23012 -4142
rect 22555 -4192 23012 -4176
rect 22555 -4193 22571 -4192
rect 22505 -4200 22571 -4193
rect 23119 -4231 23153 -4102
rect 23645 -4005 23691 -3993
rect 23645 -4181 23651 -4005
rect 23685 -4181 23691 -4005
rect 23645 -4193 23691 -4181
rect 23763 -4005 23809 -3993
rect 23763 -4181 23769 -4005
rect 23803 -4181 23809 -4005
rect 23763 -4193 23809 -4181
rect 23881 -4005 23927 -3993
rect 23881 -4181 23887 -4005
rect 23921 -4181 23927 -4005
rect 23881 -4193 23927 -4181
rect 23999 -4005 24045 -3993
rect 23999 -4181 24005 -4005
rect 24039 -4181 24045 -4005
rect 23999 -4193 24045 -4181
rect 24117 -4005 24163 -3993
rect 24117 -4181 24123 -4005
rect 24157 -4181 24163 -4005
rect 24117 -4193 24163 -4181
rect 24235 -4005 24281 -3993
rect 24235 -4181 24241 -4005
rect 24275 -4181 24281 -4005
rect 24235 -4193 24281 -4181
rect 24353 -4005 24399 -3993
rect 24353 -4181 24359 -4005
rect 24393 -4181 24399 -4005
rect 24353 -4193 24399 -4181
rect 24471 -4005 24517 -3993
rect 24471 -4181 24477 -4005
rect 24511 -4181 24517 -4005
rect 24471 -4193 24517 -4181
rect 24589 -4005 24635 -3993
rect 24589 -4181 24595 -4005
rect 24629 -4181 24635 -4005
rect 24589 -4193 24635 -4181
rect 24707 -4005 24753 -3993
rect 24707 -4181 24713 -4005
rect 24747 -4181 24753 -4005
rect 24707 -4193 24753 -4181
rect 19799 -4243 19845 -4231
rect 19799 -4419 19805 -4243
rect 19839 -4419 19845 -4243
rect 19799 -4431 19845 -4419
rect 19917 -4243 19963 -4231
rect 19917 -4419 19923 -4243
rect 19957 -4419 19963 -4243
rect 19917 -4431 19963 -4419
rect 20323 -4243 20369 -4231
rect 19924 -4725 19957 -4431
rect 20323 -4619 20329 -4243
rect 20363 -4619 20369 -4243
rect 20323 -4631 20369 -4619
rect 20441 -4243 20487 -4231
rect 20441 -4619 20447 -4243
rect 20481 -4619 20487 -4243
rect 20441 -4631 20487 -4619
rect 20559 -4243 20605 -4231
rect 20559 -4619 20565 -4243
rect 20599 -4619 20605 -4243
rect 20559 -4631 20605 -4619
rect 20677 -4243 20723 -4231
rect 20677 -4619 20683 -4243
rect 20717 -4619 20723 -4243
rect 20677 -4631 20723 -4619
rect 20795 -4243 20841 -4231
rect 20795 -4619 20801 -4243
rect 20835 -4619 20841 -4243
rect 21097 -4243 21143 -4231
rect 21097 -4419 21103 -4243
rect 21137 -4419 21143 -4243
rect 21097 -4431 21143 -4419
rect 21215 -4243 21261 -4231
rect 21215 -4419 21221 -4243
rect 21255 -4419 21261 -4243
rect 21215 -4431 21261 -4419
rect 21697 -4243 21743 -4231
rect 21697 -4419 21703 -4243
rect 21737 -4419 21743 -4243
rect 21697 -4431 21743 -4419
rect 21815 -4243 21861 -4231
rect 21815 -4419 21821 -4243
rect 21855 -4419 21861 -4243
rect 21815 -4431 21861 -4419
rect 22221 -4243 22267 -4231
rect 20795 -4631 20841 -4619
rect 20447 -4725 20481 -4631
rect 21104 -4725 21138 -4431
rect 19924 -4757 21138 -4725
rect 21822 -4725 21855 -4431
rect 22221 -4619 22227 -4243
rect 22261 -4619 22267 -4243
rect 22221 -4631 22267 -4619
rect 22339 -4243 22385 -4231
rect 22339 -4619 22345 -4243
rect 22379 -4619 22385 -4243
rect 22339 -4631 22385 -4619
rect 22457 -4243 22503 -4231
rect 22457 -4619 22463 -4243
rect 22497 -4619 22503 -4243
rect 22457 -4631 22503 -4619
rect 22575 -4243 22621 -4231
rect 22575 -4619 22581 -4243
rect 22615 -4619 22621 -4243
rect 22575 -4631 22621 -4619
rect 22693 -4243 22739 -4231
rect 22693 -4619 22699 -4243
rect 22733 -4619 22739 -4243
rect 22995 -4243 23041 -4231
rect 22995 -4419 23001 -4243
rect 23035 -4419 23041 -4243
rect 22995 -4431 23041 -4419
rect 23113 -4243 23159 -4231
rect 23113 -4419 23119 -4243
rect 23153 -4419 23159 -4243
rect 23113 -4431 23159 -4419
rect 23651 -4426 23686 -4193
rect 23930 -4241 23996 -4234
rect 23930 -4275 23946 -4241
rect 23980 -4275 23996 -4241
rect 23930 -4286 23996 -4275
rect 24122 -4286 24158 -4193
rect 23930 -4287 24158 -4286
rect 24358 -4287 24394 -4193
rect 24594 -4287 24630 -4193
rect 23930 -4316 24630 -4287
rect 24048 -4317 24630 -4316
rect 24048 -4358 24114 -4317
rect 24048 -4392 24064 -4358
rect 24098 -4392 24114 -4358
rect 24048 -4399 24114 -4392
rect 23651 -4430 24040 -4426
rect 24476 -4430 24510 -4317
rect 22693 -4631 22739 -4619
rect 22345 -4725 22379 -4631
rect 23002 -4725 23036 -4431
rect 23651 -4442 24045 -4430
rect 23651 -4455 24005 -4442
rect 23651 -4458 23729 -4455
rect 23646 -4510 23656 -4458
rect 23719 -4510 23729 -4458
rect 23651 -4516 23724 -4510
rect 23999 -4618 24005 -4455
rect 24039 -4618 24045 -4442
rect 23999 -4630 24045 -4618
rect 24117 -4442 24163 -4430
rect 24117 -4618 24123 -4442
rect 24157 -4618 24163 -4442
rect 24117 -4630 24163 -4618
rect 24234 -4442 24280 -4430
rect 21822 -4757 23036 -4725
rect 23918 -4746 24026 -4736
rect 24122 -4746 24157 -4630
rect 20513 -4842 20645 -4757
rect 22411 -4842 22543 -4757
rect 17888 -4905 17904 -4871
rect 17938 -4905 18755 -4871
rect 17888 -4921 18755 -4905
rect 18125 -4937 18755 -4921
rect 18170 -4941 18755 -4937
rect 18654 -4942 18755 -4941
rect 18125 -4990 18225 -4979
rect 18125 -5001 18139 -4990
rect 17770 -5049 18139 -5001
rect 17771 -5152 17837 -5049
rect 18125 -5079 18139 -5049
rect 18129 -5096 18139 -5079
rect 18251 -5096 18261 -4990
rect 19658 -5149 19724 -4870
rect 20503 -4950 20513 -4842
rect 20645 -4950 20655 -4842
rect 22401 -4950 22411 -4842
rect 22543 -4950 22553 -4842
rect 24026 -4794 24157 -4746
rect 24234 -4794 24240 -4442
rect 24026 -4818 24240 -4794
rect 24274 -4818 24280 -4442
rect 24026 -4830 24280 -4818
rect 24352 -4442 24398 -4430
rect 24352 -4818 24358 -4442
rect 24392 -4818 24398 -4442
rect 24352 -4830 24398 -4818
rect 24470 -4442 24516 -4430
rect 24470 -4818 24476 -4442
rect 24510 -4818 24516 -4442
rect 24470 -4830 24516 -4818
rect 24026 -4834 24274 -4830
rect 25175 -4832 25268 -3658
rect 24683 -4834 25268 -4832
rect 24026 -4878 24100 -4834
rect 24638 -4862 25268 -4834
rect 24283 -4868 24349 -4862
rect 23918 -4888 24026 -4878
rect 24283 -4902 24299 -4868
rect 24333 -4902 24349 -4868
rect 24283 -4998 24349 -4902
rect 24401 -4868 25268 -4862
rect 24401 -4902 24417 -4868
rect 24451 -4902 25268 -4868
rect 24401 -4918 25268 -4902
rect 24638 -4934 25268 -4918
rect 24683 -4938 25268 -4934
rect 25167 -4939 25268 -4938
rect 24638 -4987 24738 -4976
rect 24638 -4998 24652 -4987
rect 24283 -5046 24652 -4998
rect 24284 -5149 24350 -5046
rect 24638 -5076 24652 -5046
rect 24642 -5093 24652 -5076
rect 24764 -5093 24774 -4987
rect 6611 -5237 11305 -5157
rect 13145 -5232 17839 -5152
rect 19658 -5229 24352 -5149
<< via1 >>
rect 1372 5043 1504 5151
rect 3854 5097 3986 5205
rect 4255 5107 4311 5121
rect 4255 5073 4271 5107
rect 4271 5073 4305 5107
rect 4305 5073 4311 5107
rect 4255 5055 4311 5073
rect 5001 5097 5133 5205
rect 3125 4983 3191 4999
rect 3125 4949 3141 4983
rect 3141 4949 3175 4983
rect 3175 4949 3191 4983
rect 3125 4933 3191 4949
rect 7885 5040 8017 5148
rect 10367 5094 10499 5202
rect 3791 4286 3890 4383
rect 1652 3980 1760 4112
rect 144 3402 256 3508
rect 143 2394 255 2396
rect 143 2290 261 2394
rect 149 2288 261 2290
rect 3200 3697 3332 3805
rect 638 3419 750 3525
rect 1386 3393 1518 3501
rect 4947 4309 5012 4363
rect 10768 5104 10824 5118
rect 10768 5070 10784 5104
rect 10784 5070 10818 5104
rect 10818 5070 10824 5104
rect 10768 5052 10824 5070
rect 11514 5094 11646 5202
rect 9638 4980 9704 4996
rect 9638 4946 9654 4980
rect 9654 4946 9688 4980
rect 9688 4946 9704 4980
rect 9638 4930 9704 4946
rect 14419 5035 14551 5143
rect 16901 5089 17033 5197
rect 6042 4297 6110 4372
rect 4342 3695 4474 3803
rect 3199 3050 3331 3158
rect 5097 3050 5229 3158
rect 921 2288 1039 2406
rect 1666 2330 1774 2462
rect 10304 4283 10403 4380
rect 8165 3977 8273 4109
rect 6657 3399 6769 3505
rect 418 1946 511 2025
rect 1381 1789 1513 1897
rect 3844 2172 3907 2188
rect 3844 2138 3873 2172
rect 3873 2138 3907 2172
rect 3844 2122 3907 2138
rect 6656 2391 6768 2393
rect 6656 2287 6774 2391
rect 6662 2285 6774 2287
rect 1968 1094 2031 1146
rect 1661 726 1769 858
rect 923 511 1035 617
rect 3144 654 3276 762
rect 5042 654 5174 762
rect 9713 3694 9845 3802
rect 7151 3416 7263 3522
rect 7899 3390 8031 3498
rect 11460 4306 11525 4360
rect 17302 5099 17358 5113
rect 17302 5065 17318 5099
rect 17318 5065 17352 5099
rect 17352 5065 17358 5099
rect 17302 5047 17358 5065
rect 18048 5089 18180 5197
rect 16172 4975 16238 4991
rect 16172 4941 16188 4975
rect 16188 4941 16222 4975
rect 16222 4941 16238 4975
rect 16172 4925 16238 4941
rect 20977 5039 21109 5147
rect 23459 5093 23591 5201
rect 12555 4294 12623 4369
rect 10855 3692 10987 3800
rect 9712 3047 9844 3155
rect 11610 3047 11742 3155
rect 7434 2285 7552 2403
rect 8179 2327 8287 2459
rect 16838 4278 16937 4375
rect 14699 3972 14807 4104
rect 13191 3394 13303 3500
rect 6931 1943 7024 2022
rect 7894 1786 8026 1894
rect 10357 2169 10420 2185
rect 10357 2135 10386 2169
rect 10386 2135 10420 2169
rect 10357 2119 10420 2135
rect 13190 2386 13302 2388
rect 13190 2282 13308 2386
rect 13196 2280 13308 2282
rect 8481 1091 8544 1143
rect 8174 723 8282 855
rect 7436 508 7548 614
rect 9657 651 9789 759
rect 11555 651 11687 759
rect 16247 3689 16379 3797
rect 13685 3411 13797 3517
rect 14433 3385 14565 3493
rect 17994 4301 18059 4355
rect 23860 5103 23916 5117
rect 23860 5069 23876 5103
rect 23876 5069 23910 5103
rect 23910 5069 23916 5103
rect 23860 5051 23916 5069
rect 24606 5093 24738 5201
rect 22730 4979 22796 4995
rect 22730 4945 22746 4979
rect 22746 4945 22780 4979
rect 22780 4945 22796 4979
rect 22730 4929 22796 4945
rect 19089 4289 19157 4364
rect 17389 3687 17521 3795
rect 16246 3042 16378 3150
rect 18144 3042 18276 3150
rect 13968 2280 14086 2398
rect 14713 2322 14821 2454
rect 23396 4282 23495 4379
rect 21257 3976 21365 4108
rect 19749 3398 19861 3504
rect 13465 1938 13558 2017
rect 14428 1781 14560 1889
rect 16891 2164 16954 2180
rect 16891 2130 16920 2164
rect 16920 2130 16954 2164
rect 16891 2114 16954 2130
rect 19748 2390 19860 2392
rect 19748 2286 19866 2390
rect 19754 2284 19866 2286
rect 15015 1086 15078 1138
rect 14708 718 14816 850
rect 13970 503 14082 609
rect 16191 646 16323 754
rect 18089 646 18221 754
rect 22805 3693 22937 3801
rect 20243 3415 20355 3521
rect 20991 3389 21123 3497
rect 24552 4305 24617 4359
rect 25647 4293 25715 4368
rect 23947 3691 24079 3799
rect 22804 3046 22936 3154
rect 24702 3046 24834 3154
rect 20526 2284 20644 2402
rect 21271 2326 21379 2458
rect 20023 1942 20116 2021
rect 20986 1785 21118 1893
rect 23449 2168 23512 2184
rect 23449 2134 23478 2168
rect 23478 2134 23512 2168
rect 23449 2118 23512 2134
rect 21573 1090 21636 1142
rect 21266 722 21374 854
rect 20528 507 20640 613
rect 22749 650 22881 758
rect 24647 650 24779 758
rect 949 -511 1081 -403
rect 1771 -501 1827 -487
rect 1771 -535 1777 -501
rect 1777 -535 1811 -501
rect 1811 -535 1827 -501
rect 1771 -553 1827 -535
rect 2096 -511 2228 -403
rect -28 -1311 40 -1236
rect 1070 -1299 1135 -1245
rect 1608 -1913 1740 -1805
rect 2891 -625 2957 -609
rect 2891 -659 2907 -625
rect 2907 -659 2941 -625
rect 2941 -659 2957 -625
rect 2891 -675 2957 -659
rect 4578 -565 4710 -457
rect 7507 -515 7639 -407
rect 8329 -505 8385 -491
rect 8329 -539 8335 -505
rect 8335 -539 8369 -505
rect 8369 -539 8385 -505
rect 8329 -557 8385 -539
rect 8654 -515 8786 -407
rect 2192 -1322 2291 -1225
rect 4322 -1628 4430 -1496
rect 6530 -1315 6598 -1240
rect 7628 -1303 7693 -1249
rect 2750 -1911 2882 -1803
rect 4564 -2215 4696 -2107
rect 5332 -2189 5444 -2083
rect 853 -2558 985 -2450
rect 2751 -2558 2883 -2450
rect 4308 -3278 4416 -3146
rect 2175 -3436 2238 -3420
rect 2175 -3470 2209 -3436
rect 2209 -3470 2238 -3436
rect 2175 -3486 2238 -3470
rect 5043 -3320 5161 -3202
rect 5826 -2206 5938 -2100
rect 8166 -1917 8298 -1809
rect 9449 -629 9515 -613
rect 9449 -663 9465 -629
rect 9465 -663 9499 -629
rect 9499 -663 9515 -629
rect 9449 -679 9515 -663
rect 11136 -569 11268 -461
rect 14041 -510 14173 -402
rect 14863 -500 14919 -486
rect 14863 -534 14869 -500
rect 14869 -534 14903 -500
rect 14903 -534 14919 -500
rect 14863 -552 14919 -534
rect 15188 -510 15320 -402
rect 8750 -1326 8849 -1229
rect 10880 -1632 10988 -1500
rect 13064 -1310 13132 -1235
rect 14162 -1298 14227 -1244
rect 9308 -1915 9440 -1807
rect 11122 -2219 11254 -2111
rect 11890 -2193 12002 -2087
rect 7411 -2562 7543 -2454
rect 9309 -2562 9441 -2454
rect 5827 -3214 5939 -3212
rect 5821 -3318 5939 -3214
rect 10866 -3282 10974 -3150
rect 5821 -3320 5933 -3318
rect 5571 -3662 5664 -3583
rect 4569 -3819 4701 -3711
rect 4051 -4514 4114 -4462
rect 908 -4954 1040 -4846
rect 2806 -4954 2938 -4846
rect 4313 -4882 4421 -4750
rect 8733 -3440 8796 -3424
rect 8733 -3474 8767 -3440
rect 8767 -3474 8796 -3440
rect 8733 -3490 8796 -3474
rect 11601 -3324 11719 -3206
rect 12384 -2210 12496 -2104
rect 14700 -1912 14832 -1804
rect 15983 -624 16049 -608
rect 15983 -658 15999 -624
rect 15999 -658 16033 -624
rect 16033 -658 16049 -624
rect 15983 -674 16049 -658
rect 17670 -564 17802 -456
rect 20554 -507 20686 -399
rect 21376 -497 21432 -483
rect 21376 -531 21382 -497
rect 21382 -531 21416 -497
rect 21416 -531 21432 -497
rect 21376 -549 21432 -531
rect 21701 -507 21833 -399
rect 15284 -1321 15383 -1224
rect 17414 -1627 17522 -1495
rect 19577 -1307 19645 -1232
rect 20675 -1295 20740 -1241
rect 15842 -1910 15974 -1802
rect 17656 -2214 17788 -2106
rect 18424 -2188 18536 -2082
rect 13945 -2557 14077 -2449
rect 15843 -2557 15975 -2449
rect 12385 -3218 12497 -3216
rect 12379 -3322 12497 -3218
rect 17400 -3277 17508 -3145
rect 12379 -3324 12491 -3322
rect 12129 -3666 12222 -3587
rect 11127 -3823 11259 -3715
rect 10609 -4518 10672 -4466
rect 5047 -5097 5159 -4991
rect 7466 -4958 7598 -4850
rect 9364 -4958 9496 -4850
rect 10871 -4886 10979 -4754
rect 15267 -3435 15330 -3419
rect 15267 -3469 15301 -3435
rect 15301 -3469 15330 -3435
rect 15267 -3485 15330 -3469
rect 18135 -3319 18253 -3201
rect 18918 -2205 19030 -2099
rect 21213 -1909 21345 -1801
rect 22496 -621 22562 -605
rect 22496 -655 22512 -621
rect 22512 -655 22546 -621
rect 22546 -655 22562 -621
rect 22496 -671 22562 -655
rect 24183 -561 24315 -453
rect 21797 -1318 21896 -1221
rect 23927 -1624 24035 -1492
rect 22355 -1907 22487 -1799
rect 24169 -2211 24301 -2103
rect 24937 -2185 25049 -2079
rect 20458 -2554 20590 -2446
rect 22356 -2554 22488 -2446
rect 18919 -3213 19031 -3211
rect 18913 -3317 19031 -3213
rect 23913 -3274 24021 -3142
rect 18913 -3319 19025 -3317
rect 18663 -3661 18756 -3582
rect 17661 -3818 17793 -3710
rect 17143 -4513 17206 -4461
rect 11605 -5101 11717 -4995
rect 14000 -4953 14132 -4845
rect 15898 -4953 16030 -4845
rect 17405 -4881 17513 -4749
rect 21780 -3432 21843 -3416
rect 21780 -3466 21814 -3432
rect 21814 -3466 21843 -3432
rect 21780 -3482 21843 -3466
rect 24648 -3316 24766 -3198
rect 25431 -2202 25543 -2096
rect 25432 -3210 25544 -3208
rect 25426 -3314 25544 -3210
rect 25426 -3316 25538 -3314
rect 25176 -3658 25269 -3579
rect 24174 -3815 24306 -3707
rect 23656 -4510 23719 -4458
rect 18139 -5096 18251 -4990
rect 20513 -4950 20645 -4842
rect 22411 -4950 22543 -4842
rect 23918 -4878 24026 -4746
rect 24652 -5093 24764 -4987
<< metal2 >>
rect 3843 5216 3996 5226
rect 1361 5162 1514 5172
rect 4990 5216 5143 5226
rect 4255 5121 4311 5131
rect 3843 5077 3996 5087
rect 1361 5023 1514 5033
rect 4130 5055 4255 5117
rect 4311 5055 4312 5117
rect 10356 5213 10509 5223
rect 4990 5077 5143 5087
rect 7874 5159 8027 5169
rect 3125 5006 3191 5009
rect 2199 4999 3191 5006
rect 2199 4933 3125 4999
rect 1632 3970 1642 4123
rect 1771 3970 1781 4123
rect 132 3535 299 3536
rect 639 3535 755 3536
rect 132 3525 755 3535
rect 132 3508 638 3525
rect 132 3402 144 3508
rect 256 3419 638 3508
rect 750 3419 755 3525
rect 256 3402 755 3419
rect 132 3393 755 3402
rect 1375 3512 1528 3522
rect 1375 3373 1528 3383
rect 131 2414 296 2424
rect 131 2413 299 2414
rect 921 2413 1039 2416
rect 131 2406 1039 2413
rect 131 2396 921 2406
rect 131 2290 143 2396
rect 255 2394 921 2396
rect 131 2288 149 2290
rect 261 2288 921 2394
rect 1646 2320 1656 2473
rect 1785 2320 1795 2473
rect 131 2281 1039 2288
rect 137 2279 1039 2281
rect 174 2278 1039 2279
rect 408 2034 523 2044
rect 408 1927 523 1937
rect 918 627 1034 2278
rect 1370 1908 1523 1918
rect 1370 1769 1523 1779
rect 1968 1150 2031 1156
rect 2199 1150 2267 4933
rect 3125 4923 3191 4933
rect 4130 4394 4190 5055
rect 4255 5045 4311 5055
rect 11503 5213 11656 5223
rect 10768 5118 10824 5128
rect 10356 5074 10509 5084
rect 7874 5020 8027 5030
rect 10643 5052 10768 5114
rect 10824 5052 10825 5114
rect 16890 5208 17043 5218
rect 11503 5074 11656 5084
rect 14408 5154 14561 5164
rect 9638 5003 9704 5006
rect 4052 4393 4190 4394
rect 3790 4383 4190 4393
rect 3790 4286 3791 4383
rect 3890 4286 4190 4383
rect 8712 4996 9704 5003
rect 8712 4930 9638 4996
rect 4947 4372 5012 4373
rect 6042 4372 6110 4382
rect 4946 4363 6042 4372
rect 4946 4309 4947 4363
rect 5012 4309 6042 4363
rect 4946 4298 6042 4309
rect 6042 4287 6110 4297
rect 3790 4278 4190 4286
rect 3790 4274 4099 4278
rect 8145 3967 8155 4120
rect 8284 3967 8294 4120
rect 3190 3815 3343 3825
rect 3190 3676 3343 3686
rect 4332 3813 4485 3823
rect 4332 3674 4485 3684
rect 6645 3532 6812 3533
rect 7152 3532 7268 3533
rect 6645 3522 7268 3532
rect 6645 3505 7151 3522
rect 6645 3399 6657 3505
rect 6769 3416 7151 3505
rect 7263 3416 7268 3522
rect 6769 3399 7268 3416
rect 6645 3390 7268 3399
rect 7888 3509 8041 3519
rect 7888 3370 8041 3380
rect 3188 3169 3341 3179
rect 3188 3030 3341 3040
rect 5086 3169 5239 3179
rect 5086 3030 5239 3040
rect 6644 2411 6809 2421
rect 6644 2410 6812 2411
rect 7434 2410 7552 2413
rect 6644 2403 7552 2410
rect 6644 2393 7434 2403
rect 6644 2287 6656 2393
rect 6768 2391 7434 2393
rect 6644 2285 6662 2287
rect 6774 2285 7434 2391
rect 8159 2317 8169 2470
rect 8298 2317 8308 2470
rect 6644 2278 7552 2285
rect 6650 2276 7552 2278
rect 6687 2275 7552 2276
rect 3829 2198 3907 2208
rect 3829 2102 3907 2112
rect 6921 2031 7036 2041
rect 6921 1924 7036 1934
rect 1963 1146 2267 1150
rect 1963 1094 1968 1146
rect 2031 1094 2267 1146
rect 1963 1088 2267 1094
rect 1968 1084 2031 1088
rect 1641 716 1651 869
rect 1780 716 1790 869
rect 3134 772 3287 782
rect 3134 633 3287 643
rect 5032 772 5185 782
rect 5032 633 5185 643
rect 918 617 1035 627
rect 918 511 923 617
rect 918 501 1035 511
rect 7431 624 7547 2275
rect 7883 1905 8036 1915
rect 7883 1766 8036 1776
rect 8481 1147 8544 1153
rect 8712 1147 8780 4930
rect 9638 4920 9704 4930
rect 10643 4391 10703 5052
rect 10768 5042 10824 5052
rect 18037 5208 18190 5218
rect 17302 5113 17358 5123
rect 16890 5069 17043 5079
rect 14408 5015 14561 5025
rect 17177 5047 17302 5109
rect 17358 5047 17359 5109
rect 23448 5212 23601 5222
rect 18037 5069 18190 5079
rect 20966 5158 21119 5168
rect 16172 4998 16238 5001
rect 10565 4390 10703 4391
rect 10303 4380 10703 4390
rect 10303 4283 10304 4380
rect 10403 4283 10703 4380
rect 15246 4991 16238 4998
rect 15246 4925 16172 4991
rect 11460 4369 11525 4370
rect 12555 4369 12623 4379
rect 11459 4360 12555 4369
rect 11459 4306 11460 4360
rect 11525 4306 12555 4360
rect 11459 4295 12555 4306
rect 12555 4284 12623 4294
rect 10303 4275 10703 4283
rect 10303 4271 10612 4275
rect 14679 3962 14689 4115
rect 14818 3962 14828 4115
rect 9703 3812 9856 3822
rect 9703 3673 9856 3683
rect 10845 3810 10998 3820
rect 10845 3671 10998 3681
rect 13179 3527 13346 3528
rect 13686 3527 13802 3528
rect 13179 3517 13802 3527
rect 13179 3500 13685 3517
rect 13179 3394 13191 3500
rect 13303 3411 13685 3500
rect 13797 3411 13802 3517
rect 13303 3394 13802 3411
rect 13179 3385 13802 3394
rect 14422 3504 14575 3514
rect 14422 3365 14575 3375
rect 9701 3166 9854 3176
rect 9701 3027 9854 3037
rect 11599 3166 11752 3176
rect 11599 3027 11752 3037
rect 13178 2406 13343 2416
rect 13178 2405 13346 2406
rect 13968 2405 14086 2408
rect 13178 2398 14086 2405
rect 13178 2388 13968 2398
rect 13178 2282 13190 2388
rect 13302 2386 13968 2388
rect 13178 2280 13196 2282
rect 13308 2280 13968 2386
rect 14693 2312 14703 2465
rect 14832 2312 14842 2465
rect 13178 2273 14086 2280
rect 13184 2271 14086 2273
rect 13221 2270 14086 2271
rect 10342 2195 10420 2205
rect 10342 2099 10420 2109
rect 13455 2026 13570 2036
rect 13455 1919 13570 1929
rect 8476 1143 8780 1147
rect 8476 1091 8481 1143
rect 8544 1091 8780 1143
rect 8476 1085 8780 1091
rect 8481 1081 8544 1085
rect 8154 713 8164 866
rect 8293 713 8303 866
rect 9647 769 9800 779
rect 9647 630 9800 640
rect 11545 769 11698 779
rect 11545 630 11698 640
rect 7431 614 7548 624
rect 7431 508 7436 614
rect 918 500 1034 501
rect 7431 498 7548 508
rect 13965 619 14081 2270
rect 14417 1900 14570 1910
rect 14417 1761 14570 1771
rect 15015 1142 15078 1148
rect 15246 1142 15314 4925
rect 16172 4915 16238 4925
rect 17177 4386 17237 5047
rect 17302 5037 17358 5047
rect 24595 5212 24748 5222
rect 23860 5117 23916 5127
rect 23448 5073 23601 5083
rect 20966 5019 21119 5029
rect 23735 5051 23860 5113
rect 23916 5051 23917 5113
rect 24595 5073 24748 5083
rect 22730 5002 22796 5005
rect 17099 4385 17237 4386
rect 16837 4375 17237 4385
rect 16837 4278 16838 4375
rect 16937 4278 17237 4375
rect 21804 4995 22796 5002
rect 21804 4929 22730 4995
rect 17994 4364 18059 4365
rect 19089 4364 19157 4374
rect 17993 4355 19089 4364
rect 17993 4301 17994 4355
rect 18059 4301 19089 4355
rect 17993 4290 19089 4301
rect 19089 4279 19157 4289
rect 16837 4270 17237 4278
rect 16837 4266 17146 4270
rect 21237 3966 21247 4119
rect 21376 3966 21386 4119
rect 16237 3807 16390 3817
rect 16237 3668 16390 3678
rect 17379 3805 17532 3815
rect 17379 3666 17532 3676
rect 19737 3531 19904 3532
rect 20244 3531 20360 3532
rect 19737 3521 20360 3531
rect 19737 3504 20243 3521
rect 19737 3398 19749 3504
rect 19861 3415 20243 3504
rect 20355 3415 20360 3521
rect 19861 3398 20360 3415
rect 19737 3389 20360 3398
rect 20980 3508 21133 3518
rect 20980 3369 21133 3379
rect 16235 3161 16388 3171
rect 16235 3022 16388 3032
rect 18133 3161 18286 3171
rect 18133 3022 18286 3032
rect 19736 2410 19901 2420
rect 19736 2409 19904 2410
rect 20526 2409 20644 2412
rect 19736 2402 20644 2409
rect 19736 2392 20526 2402
rect 19736 2286 19748 2392
rect 19860 2390 20526 2392
rect 19736 2284 19754 2286
rect 19866 2284 20526 2390
rect 21251 2316 21261 2469
rect 21390 2316 21400 2469
rect 19736 2277 20644 2284
rect 19742 2275 20644 2277
rect 19779 2274 20644 2275
rect 16876 2190 16954 2200
rect 16876 2094 16954 2104
rect 20013 2030 20128 2040
rect 20013 1923 20128 1933
rect 15010 1138 15314 1142
rect 15010 1086 15015 1138
rect 15078 1086 15314 1138
rect 15010 1080 15314 1086
rect 15015 1076 15078 1080
rect 14688 708 14698 861
rect 14827 708 14837 861
rect 16181 764 16334 774
rect 16181 625 16334 635
rect 18079 764 18232 774
rect 18079 625 18232 635
rect 20523 623 20639 2274
rect 20975 1904 21128 1914
rect 20975 1765 21128 1775
rect 21573 1146 21636 1152
rect 21804 1146 21872 4929
rect 22730 4919 22796 4929
rect 23735 4390 23795 5051
rect 23860 5041 23916 5051
rect 23657 4389 23795 4390
rect 23395 4379 23795 4389
rect 23395 4282 23396 4379
rect 23495 4282 23795 4379
rect 24552 4368 24617 4369
rect 25647 4368 25715 4378
rect 24551 4359 25647 4368
rect 24551 4305 24552 4359
rect 24617 4305 25647 4359
rect 24551 4294 25647 4305
rect 25647 4283 25715 4293
rect 23395 4274 23795 4282
rect 23395 4270 23704 4274
rect 22795 3811 22948 3821
rect 22795 3672 22948 3682
rect 23937 3809 24090 3819
rect 23937 3670 24090 3680
rect 22793 3165 22946 3175
rect 22793 3026 22946 3036
rect 24691 3165 24844 3175
rect 24691 3026 24844 3036
rect 23434 2194 23512 2204
rect 23434 2098 23512 2108
rect 21568 1142 21872 1146
rect 21568 1090 21573 1142
rect 21636 1090 21872 1142
rect 21568 1084 21872 1090
rect 21573 1080 21636 1084
rect 21246 712 21256 865
rect 21385 712 21395 865
rect 22739 768 22892 778
rect 22739 629 22892 639
rect 24637 768 24790 778
rect 24637 629 24790 639
rect 13965 609 14082 619
rect 13965 503 13970 609
rect 7431 497 7547 498
rect 13965 493 14082 503
rect 20523 613 20640 623
rect 20523 507 20528 613
rect 20523 497 20640 507
rect 20523 496 20639 497
rect 13965 492 14081 493
rect 939 -392 1092 -382
rect 2086 -392 2239 -382
rect 1771 -487 1827 -477
rect 939 -531 1092 -521
rect 1770 -553 1771 -491
rect 1827 -553 1952 -491
rect 7497 -396 7650 -386
rect 2086 -531 2239 -521
rect 4568 -446 4721 -436
rect 1771 -563 1827 -553
rect 1892 -1214 1952 -553
rect 8644 -396 8797 -386
rect 8329 -491 8385 -481
rect 7497 -535 7650 -525
rect 8328 -557 8329 -495
rect 8385 -557 8510 -495
rect 14031 -391 14184 -381
rect 8644 -535 8797 -525
rect 11126 -450 11279 -440
rect 8329 -567 8385 -557
rect 4568 -585 4721 -575
rect 2891 -602 2957 -599
rect 2891 -609 3883 -602
rect 2957 -675 3883 -609
rect 2891 -685 2957 -675
rect 1892 -1215 2030 -1214
rect 1892 -1225 2292 -1215
rect -28 -1236 40 -1226
rect 1070 -1236 1135 -1235
rect 40 -1245 1136 -1236
rect 40 -1299 1070 -1245
rect 1135 -1299 1136 -1245
rect 40 -1310 1136 -1299
rect -28 -1321 40 -1311
rect 1892 -1322 2192 -1225
rect 2291 -1322 2292 -1225
rect 1892 -1330 2292 -1322
rect 1983 -1334 2292 -1330
rect 1597 -1795 1750 -1785
rect 1597 -1934 1750 -1924
rect 2739 -1793 2892 -1783
rect 2739 -1932 2892 -1922
rect 843 -2439 996 -2429
rect 843 -2578 996 -2568
rect 2741 -2439 2894 -2429
rect 2741 -2578 2894 -2568
rect 2175 -3410 2253 -3400
rect 2175 -3506 2253 -3496
rect 3815 -4458 3883 -675
rect 8450 -1218 8510 -557
rect 15178 -391 15331 -381
rect 14863 -486 14919 -476
rect 14031 -530 14184 -520
rect 14862 -552 14863 -490
rect 14919 -552 15044 -490
rect 20544 -388 20697 -378
rect 15178 -530 15331 -520
rect 17660 -445 17813 -435
rect 14863 -562 14919 -552
rect 11126 -589 11279 -579
rect 9449 -606 9515 -603
rect 9449 -613 10441 -606
rect 9515 -679 10441 -613
rect 9449 -689 9515 -679
rect 8450 -1219 8588 -1218
rect 8450 -1229 8850 -1219
rect 6530 -1240 6598 -1230
rect 7628 -1240 7693 -1239
rect 6598 -1249 7694 -1240
rect 6598 -1303 7628 -1249
rect 7693 -1303 7694 -1249
rect 6598 -1314 7694 -1303
rect 6530 -1325 6598 -1315
rect 8450 -1326 8750 -1229
rect 8849 -1326 8850 -1229
rect 8450 -1334 8850 -1326
rect 8541 -1338 8850 -1334
rect 4301 -1638 4311 -1485
rect 4440 -1638 4450 -1485
rect 8155 -1799 8308 -1789
rect 8155 -1938 8308 -1928
rect 9297 -1797 9450 -1787
rect 9297 -1936 9450 -1926
rect 5327 -2073 5443 -2072
rect 5783 -2073 5950 -2072
rect 5327 -2083 5950 -2073
rect 4554 -2096 4707 -2086
rect 5327 -2189 5332 -2083
rect 5444 -2100 5950 -2083
rect 5444 -2189 5826 -2100
rect 5327 -2206 5826 -2189
rect 5938 -2206 5950 -2100
rect 5327 -2215 5950 -2206
rect 4554 -2235 4707 -2225
rect 7401 -2443 7554 -2433
rect 7401 -2582 7554 -2572
rect 9299 -2443 9452 -2433
rect 9299 -2582 9452 -2572
rect 4287 -3288 4297 -3135
rect 4426 -3288 4436 -3135
rect 5043 -3195 5161 -3192
rect 5786 -3194 5951 -3184
rect 5783 -3195 5951 -3194
rect 5043 -3202 5951 -3195
rect 5161 -3212 5951 -3202
rect 5161 -3214 5827 -3212
rect 5161 -3320 5821 -3214
rect 5939 -3318 5951 -3212
rect 5933 -3320 5951 -3318
rect 5043 -3327 5951 -3320
rect 5043 -3329 5945 -3327
rect 5043 -3330 5908 -3329
rect 4559 -3700 4712 -3690
rect 4559 -3839 4712 -3829
rect 4051 -4458 4114 -4452
rect 3815 -4462 4119 -4458
rect 3815 -4514 4051 -4462
rect 4114 -4514 4119 -4462
rect 3815 -4520 4119 -4514
rect 4051 -4524 4114 -4520
rect 897 -4836 1050 -4826
rect 897 -4975 1050 -4965
rect 2795 -4836 2948 -4826
rect 4292 -4892 4302 -4739
rect 4431 -4892 4441 -4739
rect 2795 -4975 2948 -4965
rect 5048 -4981 5164 -3330
rect 8733 -3414 8811 -3404
rect 8733 -3510 8811 -3500
rect 5559 -3574 5674 -3564
rect 5559 -3681 5674 -3671
rect 10373 -4462 10441 -679
rect 14984 -1213 15044 -552
rect 21691 -388 21844 -378
rect 21376 -483 21432 -473
rect 20544 -527 20697 -517
rect 21375 -549 21376 -487
rect 21432 -549 21557 -487
rect 21691 -527 21844 -517
rect 24173 -442 24326 -432
rect 21376 -559 21432 -549
rect 17660 -584 17813 -574
rect 15983 -601 16049 -598
rect 15983 -608 16975 -601
rect 16049 -674 16975 -608
rect 15983 -684 16049 -674
rect 14984 -1214 15122 -1213
rect 14984 -1224 15384 -1214
rect 13064 -1235 13132 -1225
rect 14162 -1235 14227 -1234
rect 13132 -1244 14228 -1235
rect 13132 -1298 14162 -1244
rect 14227 -1298 14228 -1244
rect 13132 -1309 14228 -1298
rect 13064 -1320 13132 -1310
rect 14984 -1321 15284 -1224
rect 15383 -1321 15384 -1224
rect 14984 -1329 15384 -1321
rect 15075 -1333 15384 -1329
rect 10859 -1642 10869 -1489
rect 10998 -1642 11008 -1489
rect 14689 -1794 14842 -1784
rect 14689 -1933 14842 -1923
rect 15831 -1792 15984 -1782
rect 15831 -1931 15984 -1921
rect 11885 -2077 12001 -2076
rect 12341 -2077 12508 -2076
rect 11885 -2087 12508 -2077
rect 11112 -2100 11265 -2090
rect 11885 -2193 11890 -2087
rect 12002 -2104 12508 -2087
rect 12002 -2193 12384 -2104
rect 11885 -2210 12384 -2193
rect 12496 -2210 12508 -2104
rect 11885 -2219 12508 -2210
rect 11112 -2239 11265 -2229
rect 13935 -2438 14088 -2428
rect 13935 -2577 14088 -2567
rect 15833 -2438 15986 -2428
rect 15833 -2577 15986 -2567
rect 10845 -3292 10855 -3139
rect 10984 -3292 10994 -3139
rect 11601 -3199 11719 -3196
rect 12344 -3198 12509 -3188
rect 12341 -3199 12509 -3198
rect 11601 -3206 12509 -3199
rect 11719 -3216 12509 -3206
rect 11719 -3218 12385 -3216
rect 11719 -3324 12379 -3218
rect 12497 -3322 12509 -3216
rect 12491 -3324 12509 -3322
rect 11601 -3331 12509 -3324
rect 11601 -3333 12503 -3331
rect 11601 -3334 12466 -3333
rect 11117 -3704 11270 -3694
rect 11117 -3843 11270 -3833
rect 10609 -4462 10672 -4456
rect 10373 -4466 10677 -4462
rect 10373 -4518 10609 -4466
rect 10672 -4518 10677 -4466
rect 10373 -4524 10677 -4518
rect 10609 -4528 10672 -4524
rect 7455 -4840 7608 -4830
rect 7455 -4979 7608 -4969
rect 9353 -4840 9506 -4830
rect 10850 -4896 10860 -4743
rect 10989 -4896 10999 -4743
rect 9353 -4979 9506 -4969
rect 5047 -4991 5164 -4981
rect 11606 -4985 11722 -3334
rect 15267 -3409 15345 -3399
rect 15267 -3505 15345 -3495
rect 12117 -3578 12232 -3568
rect 12117 -3685 12232 -3675
rect 16907 -4457 16975 -674
rect 21497 -1210 21557 -549
rect 24173 -581 24326 -571
rect 22496 -598 22562 -595
rect 22496 -605 23488 -598
rect 22562 -671 23488 -605
rect 22496 -681 22562 -671
rect 21497 -1211 21635 -1210
rect 21497 -1221 21897 -1211
rect 19577 -1232 19645 -1222
rect 20675 -1232 20740 -1231
rect 19645 -1241 20741 -1232
rect 19645 -1295 20675 -1241
rect 20740 -1295 20741 -1241
rect 19645 -1306 20741 -1295
rect 19577 -1317 19645 -1307
rect 21497 -1318 21797 -1221
rect 21896 -1318 21897 -1221
rect 21497 -1326 21897 -1318
rect 21588 -1330 21897 -1326
rect 17393 -1637 17403 -1484
rect 17532 -1637 17542 -1484
rect 21202 -1791 21355 -1781
rect 21202 -1930 21355 -1920
rect 22344 -1789 22497 -1779
rect 22344 -1928 22497 -1918
rect 18419 -2072 18535 -2071
rect 18875 -2072 19042 -2071
rect 18419 -2082 19042 -2072
rect 17646 -2095 17799 -2085
rect 18419 -2188 18424 -2082
rect 18536 -2099 19042 -2082
rect 18536 -2188 18918 -2099
rect 18419 -2205 18918 -2188
rect 19030 -2205 19042 -2099
rect 18419 -2214 19042 -2205
rect 17646 -2234 17799 -2224
rect 20448 -2435 20601 -2425
rect 20448 -2574 20601 -2564
rect 22346 -2435 22499 -2425
rect 22346 -2574 22499 -2564
rect 17379 -3287 17389 -3134
rect 17518 -3287 17528 -3134
rect 18135 -3194 18253 -3191
rect 18878 -3193 19043 -3183
rect 18875 -3194 19043 -3193
rect 18135 -3201 19043 -3194
rect 18253 -3211 19043 -3201
rect 18253 -3213 18919 -3211
rect 18253 -3319 18913 -3213
rect 19031 -3317 19043 -3211
rect 19025 -3319 19043 -3317
rect 18135 -3326 19043 -3319
rect 18135 -3328 19037 -3326
rect 18135 -3329 19000 -3328
rect 17651 -3699 17804 -3689
rect 17651 -3838 17804 -3828
rect 17143 -4457 17206 -4451
rect 16907 -4461 17211 -4457
rect 16907 -4513 17143 -4461
rect 17206 -4513 17211 -4461
rect 16907 -4519 17211 -4513
rect 17143 -4523 17206 -4519
rect 13989 -4835 14142 -4825
rect 13989 -4974 14142 -4964
rect 15887 -4835 16040 -4825
rect 17384 -4891 17394 -4738
rect 17523 -4891 17533 -4738
rect 15887 -4974 16040 -4964
rect 18140 -4980 18256 -3329
rect 21780 -3406 21858 -3396
rect 21780 -3502 21858 -3492
rect 18651 -3573 18766 -3563
rect 18651 -3680 18766 -3670
rect 23420 -4454 23488 -671
rect 23906 -1634 23916 -1481
rect 24045 -1634 24055 -1481
rect 24932 -2069 25048 -2068
rect 25388 -2069 25555 -2068
rect 24932 -2079 25555 -2069
rect 24159 -2092 24312 -2082
rect 24932 -2185 24937 -2079
rect 25049 -2096 25555 -2079
rect 25049 -2185 25431 -2096
rect 24932 -2202 25431 -2185
rect 25543 -2202 25555 -2096
rect 24932 -2211 25555 -2202
rect 24159 -2231 24312 -2221
rect 23892 -3284 23902 -3131
rect 24031 -3284 24041 -3131
rect 24648 -3191 24766 -3188
rect 25391 -3190 25556 -3180
rect 25388 -3191 25556 -3190
rect 24648 -3198 25556 -3191
rect 24766 -3208 25556 -3198
rect 24766 -3210 25432 -3208
rect 24766 -3316 25426 -3210
rect 25544 -3314 25556 -3208
rect 25538 -3316 25556 -3314
rect 24648 -3323 25556 -3316
rect 24648 -3325 25550 -3323
rect 24648 -3326 25513 -3325
rect 24164 -3696 24317 -3686
rect 24164 -3835 24317 -3825
rect 23656 -4454 23719 -4448
rect 23420 -4458 23724 -4454
rect 23420 -4510 23656 -4458
rect 23719 -4510 23724 -4458
rect 23420 -4516 23724 -4510
rect 23656 -4520 23719 -4516
rect 20502 -4832 20655 -4822
rect 20502 -4971 20655 -4961
rect 22400 -4832 22553 -4822
rect 23897 -4888 23907 -4735
rect 24036 -4888 24046 -4735
rect 22400 -4971 22553 -4961
rect 24653 -4977 24769 -3326
rect 25164 -3570 25279 -3560
rect 25164 -3677 25279 -3667
rect 5159 -5097 5164 -4991
rect 5047 -5107 5164 -5097
rect 5048 -5108 5164 -5107
rect 11605 -4995 11722 -4985
rect 11717 -5101 11722 -4995
rect 11605 -5111 11722 -5101
rect 18139 -4990 18256 -4980
rect 18251 -5096 18256 -4990
rect 18139 -5106 18256 -5096
rect 24652 -4987 24769 -4977
rect 24764 -5093 24769 -4987
rect 24652 -5103 24769 -5093
rect 24653 -5104 24769 -5103
rect 18140 -5107 18256 -5106
rect 11606 -5112 11722 -5111
<< via2 >>
rect 3843 5205 3996 5216
rect 1361 5151 1514 5162
rect 1361 5043 1372 5151
rect 1372 5043 1504 5151
rect 1504 5043 1514 5151
rect 3843 5097 3854 5205
rect 3854 5097 3986 5205
rect 3986 5097 3996 5205
rect 4990 5205 5143 5216
rect 3843 5087 3996 5097
rect 1361 5033 1514 5043
rect 4990 5097 5001 5205
rect 5001 5097 5133 5205
rect 5133 5097 5143 5205
rect 10356 5202 10509 5213
rect 4990 5087 5143 5097
rect 7874 5148 8027 5159
rect 1642 4112 1771 4123
rect 1642 3980 1652 4112
rect 1652 3980 1760 4112
rect 1760 3980 1771 4112
rect 1642 3970 1771 3980
rect 1375 3501 1528 3512
rect 1375 3393 1386 3501
rect 1386 3393 1518 3501
rect 1518 3393 1528 3501
rect 1375 3383 1528 3393
rect 1656 2462 1785 2473
rect 1656 2330 1666 2462
rect 1666 2330 1774 2462
rect 1774 2330 1785 2462
rect 1656 2320 1785 2330
rect 408 2025 523 2034
rect 408 1946 418 2025
rect 418 1946 511 2025
rect 511 1946 523 2025
rect 408 1937 523 1946
rect 1370 1897 1523 1908
rect 1370 1789 1381 1897
rect 1381 1789 1513 1897
rect 1513 1789 1523 1897
rect 1370 1779 1523 1789
rect 7874 5040 7885 5148
rect 7885 5040 8017 5148
rect 8017 5040 8027 5148
rect 10356 5094 10367 5202
rect 10367 5094 10499 5202
rect 10499 5094 10509 5202
rect 11503 5202 11656 5213
rect 10356 5084 10509 5094
rect 7874 5030 8027 5040
rect 11503 5094 11514 5202
rect 11514 5094 11646 5202
rect 11646 5094 11656 5202
rect 16890 5197 17043 5208
rect 11503 5084 11656 5094
rect 14408 5143 14561 5154
rect 8155 4109 8284 4120
rect 8155 3977 8165 4109
rect 8165 3977 8273 4109
rect 8273 3977 8284 4109
rect 8155 3967 8284 3977
rect 3190 3805 3343 3815
rect 3190 3697 3200 3805
rect 3200 3697 3332 3805
rect 3332 3697 3343 3805
rect 3190 3686 3343 3697
rect 4332 3803 4485 3813
rect 4332 3695 4342 3803
rect 4342 3695 4474 3803
rect 4474 3695 4485 3803
rect 4332 3684 4485 3695
rect 7888 3498 8041 3509
rect 7888 3390 7899 3498
rect 7899 3390 8031 3498
rect 8031 3390 8041 3498
rect 7888 3380 8041 3390
rect 3188 3158 3341 3169
rect 3188 3050 3199 3158
rect 3199 3050 3331 3158
rect 3331 3050 3341 3158
rect 3188 3040 3341 3050
rect 5086 3158 5239 3169
rect 5086 3050 5097 3158
rect 5097 3050 5229 3158
rect 5229 3050 5239 3158
rect 5086 3040 5239 3050
rect 8169 2459 8298 2470
rect 8169 2327 8179 2459
rect 8179 2327 8287 2459
rect 8287 2327 8298 2459
rect 8169 2317 8298 2327
rect 3829 2188 3907 2198
rect 3829 2122 3844 2188
rect 3844 2122 3907 2188
rect 3829 2112 3907 2122
rect 6921 2022 7036 2031
rect 6921 1943 6931 2022
rect 6931 1943 7024 2022
rect 7024 1943 7036 2022
rect 6921 1934 7036 1943
rect 1651 858 1780 869
rect 1651 726 1661 858
rect 1661 726 1769 858
rect 1769 726 1780 858
rect 1651 716 1780 726
rect 3134 762 3287 772
rect 3134 654 3144 762
rect 3144 654 3276 762
rect 3276 654 3287 762
rect 3134 643 3287 654
rect 5032 762 5185 772
rect 5032 654 5042 762
rect 5042 654 5174 762
rect 5174 654 5185 762
rect 5032 643 5185 654
rect 7883 1894 8036 1905
rect 7883 1786 7894 1894
rect 7894 1786 8026 1894
rect 8026 1786 8036 1894
rect 7883 1776 8036 1786
rect 14408 5035 14419 5143
rect 14419 5035 14551 5143
rect 14551 5035 14561 5143
rect 16890 5089 16901 5197
rect 16901 5089 17033 5197
rect 17033 5089 17043 5197
rect 18037 5197 18190 5208
rect 16890 5079 17043 5089
rect 14408 5025 14561 5035
rect 18037 5089 18048 5197
rect 18048 5089 18180 5197
rect 18180 5089 18190 5197
rect 23448 5201 23601 5212
rect 18037 5079 18190 5089
rect 20966 5147 21119 5158
rect 14689 4104 14818 4115
rect 14689 3972 14699 4104
rect 14699 3972 14807 4104
rect 14807 3972 14818 4104
rect 14689 3962 14818 3972
rect 9703 3802 9856 3812
rect 9703 3694 9713 3802
rect 9713 3694 9845 3802
rect 9845 3694 9856 3802
rect 9703 3683 9856 3694
rect 10845 3800 10998 3810
rect 10845 3692 10855 3800
rect 10855 3692 10987 3800
rect 10987 3692 10998 3800
rect 10845 3681 10998 3692
rect 14422 3493 14575 3504
rect 14422 3385 14433 3493
rect 14433 3385 14565 3493
rect 14565 3385 14575 3493
rect 14422 3375 14575 3385
rect 9701 3155 9854 3166
rect 9701 3047 9712 3155
rect 9712 3047 9844 3155
rect 9844 3047 9854 3155
rect 9701 3037 9854 3047
rect 11599 3155 11752 3166
rect 11599 3047 11610 3155
rect 11610 3047 11742 3155
rect 11742 3047 11752 3155
rect 11599 3037 11752 3047
rect 14703 2454 14832 2465
rect 14703 2322 14713 2454
rect 14713 2322 14821 2454
rect 14821 2322 14832 2454
rect 14703 2312 14832 2322
rect 10342 2185 10420 2195
rect 10342 2119 10357 2185
rect 10357 2119 10420 2185
rect 10342 2109 10420 2119
rect 13455 2017 13570 2026
rect 13455 1938 13465 2017
rect 13465 1938 13558 2017
rect 13558 1938 13570 2017
rect 13455 1929 13570 1938
rect 8164 855 8293 866
rect 8164 723 8174 855
rect 8174 723 8282 855
rect 8282 723 8293 855
rect 8164 713 8293 723
rect 9647 759 9800 769
rect 9647 651 9657 759
rect 9657 651 9789 759
rect 9789 651 9800 759
rect 9647 640 9800 651
rect 11545 759 11698 769
rect 11545 651 11555 759
rect 11555 651 11687 759
rect 11687 651 11698 759
rect 11545 640 11698 651
rect 14417 1889 14570 1900
rect 14417 1781 14428 1889
rect 14428 1781 14560 1889
rect 14560 1781 14570 1889
rect 14417 1771 14570 1781
rect 20966 5039 20977 5147
rect 20977 5039 21109 5147
rect 21109 5039 21119 5147
rect 23448 5093 23459 5201
rect 23459 5093 23591 5201
rect 23591 5093 23601 5201
rect 24595 5201 24748 5212
rect 23448 5083 23601 5093
rect 20966 5029 21119 5039
rect 24595 5093 24606 5201
rect 24606 5093 24738 5201
rect 24738 5093 24748 5201
rect 24595 5083 24748 5093
rect 21247 4108 21376 4119
rect 21247 3976 21257 4108
rect 21257 3976 21365 4108
rect 21365 3976 21376 4108
rect 21247 3966 21376 3976
rect 16237 3797 16390 3807
rect 16237 3689 16247 3797
rect 16247 3689 16379 3797
rect 16379 3689 16390 3797
rect 16237 3678 16390 3689
rect 17379 3795 17532 3805
rect 17379 3687 17389 3795
rect 17389 3687 17521 3795
rect 17521 3687 17532 3795
rect 17379 3676 17532 3687
rect 20980 3497 21133 3508
rect 20980 3389 20991 3497
rect 20991 3389 21123 3497
rect 21123 3389 21133 3497
rect 20980 3379 21133 3389
rect 16235 3150 16388 3161
rect 16235 3042 16246 3150
rect 16246 3042 16378 3150
rect 16378 3042 16388 3150
rect 16235 3032 16388 3042
rect 18133 3150 18286 3161
rect 18133 3042 18144 3150
rect 18144 3042 18276 3150
rect 18276 3042 18286 3150
rect 18133 3032 18286 3042
rect 21261 2458 21390 2469
rect 21261 2326 21271 2458
rect 21271 2326 21379 2458
rect 21379 2326 21390 2458
rect 21261 2316 21390 2326
rect 16876 2180 16954 2190
rect 16876 2114 16891 2180
rect 16891 2114 16954 2180
rect 16876 2104 16954 2114
rect 20013 2021 20128 2030
rect 20013 1942 20023 2021
rect 20023 1942 20116 2021
rect 20116 1942 20128 2021
rect 20013 1933 20128 1942
rect 14698 850 14827 861
rect 14698 718 14708 850
rect 14708 718 14816 850
rect 14816 718 14827 850
rect 14698 708 14827 718
rect 16181 754 16334 764
rect 16181 646 16191 754
rect 16191 646 16323 754
rect 16323 646 16334 754
rect 16181 635 16334 646
rect 18079 754 18232 764
rect 18079 646 18089 754
rect 18089 646 18221 754
rect 18221 646 18232 754
rect 18079 635 18232 646
rect 20975 1893 21128 1904
rect 20975 1785 20986 1893
rect 20986 1785 21118 1893
rect 21118 1785 21128 1893
rect 20975 1775 21128 1785
rect 22795 3801 22948 3811
rect 22795 3693 22805 3801
rect 22805 3693 22937 3801
rect 22937 3693 22948 3801
rect 22795 3682 22948 3693
rect 23937 3799 24090 3809
rect 23937 3691 23947 3799
rect 23947 3691 24079 3799
rect 24079 3691 24090 3799
rect 23937 3680 24090 3691
rect 22793 3154 22946 3165
rect 22793 3046 22804 3154
rect 22804 3046 22936 3154
rect 22936 3046 22946 3154
rect 22793 3036 22946 3046
rect 24691 3154 24844 3165
rect 24691 3046 24702 3154
rect 24702 3046 24834 3154
rect 24834 3046 24844 3154
rect 24691 3036 24844 3046
rect 23434 2184 23512 2194
rect 23434 2118 23449 2184
rect 23449 2118 23512 2184
rect 23434 2108 23512 2118
rect 21256 854 21385 865
rect 21256 722 21266 854
rect 21266 722 21374 854
rect 21374 722 21385 854
rect 21256 712 21385 722
rect 22739 758 22892 768
rect 22739 650 22749 758
rect 22749 650 22881 758
rect 22881 650 22892 758
rect 22739 639 22892 650
rect 24637 758 24790 768
rect 24637 650 24647 758
rect 24647 650 24779 758
rect 24779 650 24790 758
rect 24637 639 24790 650
rect 939 -403 1092 -392
rect 939 -511 949 -403
rect 949 -511 1081 -403
rect 1081 -511 1092 -403
rect 2086 -403 2239 -392
rect 939 -521 1092 -511
rect 2086 -511 2096 -403
rect 2096 -511 2228 -403
rect 2228 -511 2239 -403
rect 7497 -407 7650 -396
rect 2086 -521 2239 -511
rect 4568 -457 4721 -446
rect 4568 -565 4578 -457
rect 4578 -565 4710 -457
rect 4710 -565 4721 -457
rect 7497 -515 7507 -407
rect 7507 -515 7639 -407
rect 7639 -515 7650 -407
rect 8644 -407 8797 -396
rect 7497 -525 7650 -515
rect 8644 -515 8654 -407
rect 8654 -515 8786 -407
rect 8786 -515 8797 -407
rect 14031 -402 14184 -391
rect 8644 -525 8797 -515
rect 11126 -461 11279 -450
rect 4568 -575 4721 -565
rect 1597 -1805 1750 -1795
rect 1597 -1913 1608 -1805
rect 1608 -1913 1740 -1805
rect 1740 -1913 1750 -1805
rect 1597 -1924 1750 -1913
rect 2739 -1803 2892 -1793
rect 2739 -1911 2750 -1803
rect 2750 -1911 2882 -1803
rect 2882 -1911 2892 -1803
rect 2739 -1922 2892 -1911
rect 843 -2450 996 -2439
rect 843 -2558 853 -2450
rect 853 -2558 985 -2450
rect 985 -2558 996 -2450
rect 843 -2568 996 -2558
rect 2741 -2450 2894 -2439
rect 2741 -2558 2751 -2450
rect 2751 -2558 2883 -2450
rect 2883 -2558 2894 -2450
rect 2741 -2568 2894 -2558
rect 2175 -3420 2253 -3410
rect 2175 -3486 2238 -3420
rect 2238 -3486 2253 -3420
rect 2175 -3496 2253 -3486
rect 11126 -569 11136 -461
rect 11136 -569 11268 -461
rect 11268 -569 11279 -461
rect 14031 -510 14041 -402
rect 14041 -510 14173 -402
rect 14173 -510 14184 -402
rect 15178 -402 15331 -391
rect 14031 -520 14184 -510
rect 15178 -510 15188 -402
rect 15188 -510 15320 -402
rect 15320 -510 15331 -402
rect 20544 -399 20697 -388
rect 15178 -520 15331 -510
rect 17660 -456 17813 -445
rect 11126 -579 11279 -569
rect 4311 -1496 4440 -1485
rect 4311 -1628 4322 -1496
rect 4322 -1628 4430 -1496
rect 4430 -1628 4440 -1496
rect 4311 -1638 4440 -1628
rect 8155 -1809 8308 -1799
rect 8155 -1917 8166 -1809
rect 8166 -1917 8298 -1809
rect 8298 -1917 8308 -1809
rect 8155 -1928 8308 -1917
rect 9297 -1807 9450 -1797
rect 9297 -1915 9308 -1807
rect 9308 -1915 9440 -1807
rect 9440 -1915 9450 -1807
rect 9297 -1926 9450 -1915
rect 4554 -2107 4707 -2096
rect 4554 -2215 4564 -2107
rect 4564 -2215 4696 -2107
rect 4696 -2215 4707 -2107
rect 4554 -2225 4707 -2215
rect 7401 -2454 7554 -2443
rect 7401 -2562 7411 -2454
rect 7411 -2562 7543 -2454
rect 7543 -2562 7554 -2454
rect 7401 -2572 7554 -2562
rect 9299 -2454 9452 -2443
rect 9299 -2562 9309 -2454
rect 9309 -2562 9441 -2454
rect 9441 -2562 9452 -2454
rect 9299 -2572 9452 -2562
rect 4297 -3146 4426 -3135
rect 4297 -3278 4308 -3146
rect 4308 -3278 4416 -3146
rect 4416 -3278 4426 -3146
rect 4297 -3288 4426 -3278
rect 4559 -3711 4712 -3700
rect 4559 -3819 4569 -3711
rect 4569 -3819 4701 -3711
rect 4701 -3819 4712 -3711
rect 4559 -3829 4712 -3819
rect 897 -4846 1050 -4836
rect 897 -4954 908 -4846
rect 908 -4954 1040 -4846
rect 1040 -4954 1050 -4846
rect 897 -4965 1050 -4954
rect 2795 -4846 2948 -4836
rect 2795 -4954 2806 -4846
rect 2806 -4954 2938 -4846
rect 2938 -4954 2948 -4846
rect 4302 -4750 4431 -4739
rect 4302 -4882 4313 -4750
rect 4313 -4882 4421 -4750
rect 4421 -4882 4431 -4750
rect 4302 -4892 4431 -4882
rect 2795 -4965 2948 -4954
rect 8733 -3424 8811 -3414
rect 8733 -3490 8796 -3424
rect 8796 -3490 8811 -3424
rect 8733 -3500 8811 -3490
rect 5559 -3583 5674 -3574
rect 5559 -3662 5571 -3583
rect 5571 -3662 5664 -3583
rect 5664 -3662 5674 -3583
rect 5559 -3671 5674 -3662
rect 17660 -564 17670 -456
rect 17670 -564 17802 -456
rect 17802 -564 17813 -456
rect 20544 -507 20554 -399
rect 20554 -507 20686 -399
rect 20686 -507 20697 -399
rect 21691 -399 21844 -388
rect 20544 -517 20697 -507
rect 21691 -507 21701 -399
rect 21701 -507 21833 -399
rect 21833 -507 21844 -399
rect 21691 -517 21844 -507
rect 24173 -453 24326 -442
rect 17660 -574 17813 -564
rect 10869 -1500 10998 -1489
rect 10869 -1632 10880 -1500
rect 10880 -1632 10988 -1500
rect 10988 -1632 10998 -1500
rect 10869 -1642 10998 -1632
rect 14689 -1804 14842 -1794
rect 14689 -1912 14700 -1804
rect 14700 -1912 14832 -1804
rect 14832 -1912 14842 -1804
rect 14689 -1923 14842 -1912
rect 15831 -1802 15984 -1792
rect 15831 -1910 15842 -1802
rect 15842 -1910 15974 -1802
rect 15974 -1910 15984 -1802
rect 15831 -1921 15984 -1910
rect 11112 -2111 11265 -2100
rect 11112 -2219 11122 -2111
rect 11122 -2219 11254 -2111
rect 11254 -2219 11265 -2111
rect 11112 -2229 11265 -2219
rect 13935 -2449 14088 -2438
rect 13935 -2557 13945 -2449
rect 13945 -2557 14077 -2449
rect 14077 -2557 14088 -2449
rect 13935 -2567 14088 -2557
rect 15833 -2449 15986 -2438
rect 15833 -2557 15843 -2449
rect 15843 -2557 15975 -2449
rect 15975 -2557 15986 -2449
rect 15833 -2567 15986 -2557
rect 10855 -3150 10984 -3139
rect 10855 -3282 10866 -3150
rect 10866 -3282 10974 -3150
rect 10974 -3282 10984 -3150
rect 10855 -3292 10984 -3282
rect 11117 -3715 11270 -3704
rect 11117 -3823 11127 -3715
rect 11127 -3823 11259 -3715
rect 11259 -3823 11270 -3715
rect 11117 -3833 11270 -3823
rect 7455 -4850 7608 -4840
rect 7455 -4958 7466 -4850
rect 7466 -4958 7598 -4850
rect 7598 -4958 7608 -4850
rect 7455 -4969 7608 -4958
rect 9353 -4850 9506 -4840
rect 9353 -4958 9364 -4850
rect 9364 -4958 9496 -4850
rect 9496 -4958 9506 -4850
rect 10860 -4754 10989 -4743
rect 10860 -4886 10871 -4754
rect 10871 -4886 10979 -4754
rect 10979 -4886 10989 -4754
rect 10860 -4896 10989 -4886
rect 9353 -4969 9506 -4958
rect 15267 -3419 15345 -3409
rect 15267 -3485 15330 -3419
rect 15330 -3485 15345 -3419
rect 15267 -3495 15345 -3485
rect 12117 -3587 12232 -3578
rect 12117 -3666 12129 -3587
rect 12129 -3666 12222 -3587
rect 12222 -3666 12232 -3587
rect 12117 -3675 12232 -3666
rect 24173 -561 24183 -453
rect 24183 -561 24315 -453
rect 24315 -561 24326 -453
rect 24173 -571 24326 -561
rect 17403 -1495 17532 -1484
rect 17403 -1627 17414 -1495
rect 17414 -1627 17522 -1495
rect 17522 -1627 17532 -1495
rect 17403 -1637 17532 -1627
rect 21202 -1801 21355 -1791
rect 21202 -1909 21213 -1801
rect 21213 -1909 21345 -1801
rect 21345 -1909 21355 -1801
rect 21202 -1920 21355 -1909
rect 22344 -1799 22497 -1789
rect 22344 -1907 22355 -1799
rect 22355 -1907 22487 -1799
rect 22487 -1907 22497 -1799
rect 22344 -1918 22497 -1907
rect 17646 -2106 17799 -2095
rect 17646 -2214 17656 -2106
rect 17656 -2214 17788 -2106
rect 17788 -2214 17799 -2106
rect 17646 -2224 17799 -2214
rect 20448 -2446 20601 -2435
rect 20448 -2554 20458 -2446
rect 20458 -2554 20590 -2446
rect 20590 -2554 20601 -2446
rect 20448 -2564 20601 -2554
rect 22346 -2446 22499 -2435
rect 22346 -2554 22356 -2446
rect 22356 -2554 22488 -2446
rect 22488 -2554 22499 -2446
rect 22346 -2564 22499 -2554
rect 17389 -3145 17518 -3134
rect 17389 -3277 17400 -3145
rect 17400 -3277 17508 -3145
rect 17508 -3277 17518 -3145
rect 17389 -3287 17518 -3277
rect 17651 -3710 17804 -3699
rect 17651 -3818 17661 -3710
rect 17661 -3818 17793 -3710
rect 17793 -3818 17804 -3710
rect 17651 -3828 17804 -3818
rect 13989 -4845 14142 -4835
rect 13989 -4953 14000 -4845
rect 14000 -4953 14132 -4845
rect 14132 -4953 14142 -4845
rect 13989 -4964 14142 -4953
rect 15887 -4845 16040 -4835
rect 15887 -4953 15898 -4845
rect 15898 -4953 16030 -4845
rect 16030 -4953 16040 -4845
rect 17394 -4749 17523 -4738
rect 17394 -4881 17405 -4749
rect 17405 -4881 17513 -4749
rect 17513 -4881 17523 -4749
rect 17394 -4891 17523 -4881
rect 15887 -4964 16040 -4953
rect 21780 -3416 21858 -3406
rect 21780 -3482 21843 -3416
rect 21843 -3482 21858 -3416
rect 21780 -3492 21858 -3482
rect 18651 -3582 18766 -3573
rect 18651 -3661 18663 -3582
rect 18663 -3661 18756 -3582
rect 18756 -3661 18766 -3582
rect 18651 -3670 18766 -3661
rect 23916 -1492 24045 -1481
rect 23916 -1624 23927 -1492
rect 23927 -1624 24035 -1492
rect 24035 -1624 24045 -1492
rect 23916 -1634 24045 -1624
rect 24159 -2103 24312 -2092
rect 24159 -2211 24169 -2103
rect 24169 -2211 24301 -2103
rect 24301 -2211 24312 -2103
rect 24159 -2221 24312 -2211
rect 23902 -3142 24031 -3131
rect 23902 -3274 23913 -3142
rect 23913 -3274 24021 -3142
rect 24021 -3274 24031 -3142
rect 23902 -3284 24031 -3274
rect 24164 -3707 24317 -3696
rect 24164 -3815 24174 -3707
rect 24174 -3815 24306 -3707
rect 24306 -3815 24317 -3707
rect 24164 -3825 24317 -3815
rect 20502 -4842 20655 -4832
rect 20502 -4950 20513 -4842
rect 20513 -4950 20645 -4842
rect 20645 -4950 20655 -4842
rect 20502 -4961 20655 -4950
rect 22400 -4842 22553 -4832
rect 22400 -4950 22411 -4842
rect 22411 -4950 22543 -4842
rect 22543 -4950 22553 -4842
rect 23907 -4746 24036 -4735
rect 23907 -4878 23918 -4746
rect 23918 -4878 24026 -4746
rect 24026 -4878 24036 -4746
rect 23907 -4888 24036 -4878
rect 22400 -4961 22553 -4950
rect 25164 -3579 25279 -3570
rect 25164 -3658 25176 -3579
rect 25176 -3658 25269 -3579
rect 25269 -3658 25279 -3579
rect 25164 -3667 25279 -3658
<< metal3 >>
rect 1329 5014 1339 5193
rect 1538 5014 1548 5193
rect 3811 5068 3821 5247
rect 4020 5068 4030 5247
rect 4958 5068 4968 5247
rect 5167 5068 5177 5247
rect 7842 5011 7852 5190
rect 8051 5011 8061 5190
rect 10324 5065 10334 5244
rect 10533 5065 10543 5244
rect 11471 5065 11481 5244
rect 11680 5065 11690 5244
rect 14376 5006 14386 5185
rect 14585 5006 14595 5185
rect 16858 5060 16868 5239
rect 17067 5060 17077 5239
rect 18005 5060 18015 5239
rect 18214 5060 18224 5239
rect 20934 5010 20944 5189
rect 21143 5010 21153 5189
rect 23416 5064 23426 5243
rect 23625 5064 23635 5243
rect 24563 5064 24573 5243
rect 24772 5064 24782 5243
rect 1623 4145 1802 4155
rect 1623 3937 1802 3946
rect 8136 4142 8315 4152
rect 8136 3934 8315 3943
rect 14670 4137 14849 4147
rect 14670 3929 14849 3938
rect 21228 4141 21407 4151
rect 21228 3933 21407 3942
rect 3157 3655 3166 3834
rect 3365 3655 3375 3834
rect 4299 3653 4308 3832
rect 4507 3653 4517 3832
rect 9670 3652 9679 3831
rect 9878 3652 9888 3831
rect 10812 3650 10821 3829
rect 11020 3650 11030 3829
rect 16204 3647 16213 3826
rect 16412 3647 16422 3826
rect 17346 3645 17355 3824
rect 17554 3645 17564 3824
rect 22762 3651 22771 3830
rect 22970 3651 22980 3830
rect 23904 3649 23913 3828
rect 24112 3649 24122 3828
rect 1343 3364 1353 3543
rect 1552 3364 1562 3543
rect 7856 3361 7866 3540
rect 8065 3361 8075 3540
rect 14390 3356 14400 3535
rect 14599 3356 14609 3535
rect 20948 3360 20958 3539
rect 21157 3360 21167 3539
rect 3156 3021 3166 3200
rect 3365 3021 3375 3200
rect 5054 3021 5064 3200
rect 5263 3021 5273 3200
rect 9669 3018 9679 3197
rect 9878 3018 9888 3197
rect 11567 3018 11577 3197
rect 11776 3018 11786 3197
rect 16203 3013 16213 3192
rect 16412 3013 16422 3192
rect 18101 3013 18111 3192
rect 18310 3013 18320 3192
rect 22761 3017 22771 3196
rect 22970 3017 22980 3196
rect 24659 3017 24669 3196
rect 24868 3017 24878 3196
rect 1637 2495 1816 2505
rect 1637 2287 1816 2296
rect 8150 2492 8329 2502
rect 8150 2284 8329 2293
rect 14684 2487 14863 2497
rect 14684 2279 14863 2288
rect 21242 2491 21421 2501
rect 21242 2283 21421 2292
rect 419 2202 511 2203
rect 3817 2202 3921 2204
rect 419 2198 3921 2202
rect 419 2112 3829 2198
rect 3907 2112 3921 2198
rect 419 2099 3921 2112
rect 6932 2199 7024 2200
rect 10330 2199 10434 2201
rect 6932 2195 10434 2199
rect 20024 2198 20116 2199
rect 23422 2198 23526 2200
rect 6932 2109 10342 2195
rect 10420 2109 10434 2195
rect 419 2039 511 2099
rect 6932 2096 10434 2109
rect 13466 2194 13558 2195
rect 16864 2194 16968 2196
rect 13466 2190 16968 2194
rect 13466 2104 16876 2190
rect 16954 2104 16968 2190
rect 398 2034 533 2039
rect 6932 2036 7024 2096
rect 13466 2091 16968 2104
rect 20024 2194 23526 2198
rect 20024 2108 23434 2194
rect 23512 2108 23526 2194
rect 20024 2095 23526 2108
rect 398 1937 408 2034
rect 523 1937 533 2034
rect 6911 2031 7046 2036
rect 13466 2031 13558 2091
rect 20024 2035 20116 2095
rect 398 1932 533 1937
rect 1338 1760 1348 1939
rect 1547 1760 1557 1939
rect 6911 1934 6921 2031
rect 7036 1934 7046 2031
rect 13445 2026 13580 2031
rect 6911 1929 7046 1934
rect 7851 1757 7861 1936
rect 8060 1757 8070 1936
rect 13445 1929 13455 2026
rect 13570 1929 13580 2026
rect 20003 2030 20138 2035
rect 20003 1933 20013 2030
rect 20128 1933 20138 2030
rect 13445 1924 13580 1929
rect 14385 1752 14395 1931
rect 14594 1752 14604 1931
rect 20003 1928 20138 1933
rect 20943 1756 20953 1935
rect 21152 1756 21162 1935
rect 1632 891 1811 901
rect 8145 888 8324 898
rect 1632 683 1811 692
rect 3100 612 3110 791
rect 3309 612 3319 791
rect 4998 612 5008 791
rect 5207 612 5217 791
rect 14679 883 14858 893
rect 8145 680 8324 689
rect 9613 609 9623 788
rect 9822 609 9832 788
rect 11511 609 11521 788
rect 11720 609 11730 788
rect 21237 887 21416 897
rect 14679 675 14858 684
rect 16147 604 16157 783
rect 16356 604 16366 783
rect 18045 604 18055 783
rect 18254 604 18264 783
rect 21237 679 21416 688
rect 22705 608 22715 787
rect 22914 608 22924 787
rect 24603 608 24613 787
rect 24812 608 24822 787
rect 905 -540 915 -361
rect 1114 -540 1124 -361
rect 2052 -540 2062 -361
rect 2261 -540 2271 -361
rect 4534 -594 4544 -415
rect 4743 -594 4753 -415
rect 7463 -544 7473 -365
rect 7672 -544 7682 -365
rect 8610 -544 8620 -365
rect 8819 -544 8829 -365
rect 11092 -598 11102 -419
rect 11301 -598 11311 -419
rect 13997 -539 14007 -360
rect 14206 -539 14216 -360
rect 15144 -539 15154 -360
rect 15353 -539 15363 -360
rect 17626 -593 17636 -414
rect 17835 -593 17845 -414
rect 20510 -536 20520 -357
rect 20719 -536 20729 -357
rect 21657 -536 21667 -357
rect 21866 -536 21876 -357
rect 24139 -590 24149 -411
rect 24348 -590 24358 -411
rect 4280 -1463 4459 -1453
rect 4280 -1671 4459 -1662
rect 10838 -1467 11017 -1457
rect 10838 -1675 11017 -1666
rect 17372 -1462 17551 -1452
rect 17372 -1670 17551 -1661
rect 23885 -1459 24064 -1449
rect 23885 -1667 24064 -1658
rect 1565 -1955 1575 -1776
rect 1774 -1955 1783 -1776
rect 2707 -1953 2717 -1774
rect 2916 -1953 2925 -1774
rect 8123 -1959 8133 -1780
rect 8332 -1959 8341 -1780
rect 9265 -1957 9275 -1778
rect 9474 -1957 9483 -1778
rect 14657 -1954 14667 -1775
rect 14866 -1954 14875 -1775
rect 15799 -1952 15809 -1773
rect 16008 -1952 16017 -1773
rect 21170 -1951 21180 -1772
rect 21379 -1951 21388 -1772
rect 22312 -1949 22322 -1770
rect 22521 -1949 22530 -1770
rect 4520 -2244 4530 -2065
rect 4729 -2244 4739 -2065
rect 11078 -2248 11088 -2069
rect 11287 -2248 11297 -2069
rect 17612 -2243 17622 -2064
rect 17821 -2243 17831 -2064
rect 24125 -2240 24135 -2061
rect 24334 -2240 24344 -2061
rect 809 -2587 819 -2408
rect 1018 -2587 1028 -2408
rect 2707 -2587 2717 -2408
rect 2916 -2587 2926 -2408
rect 7367 -2591 7377 -2412
rect 7576 -2591 7586 -2412
rect 9265 -2591 9275 -2412
rect 9474 -2591 9484 -2412
rect 13901 -2586 13911 -2407
rect 14110 -2586 14120 -2407
rect 15799 -2586 15809 -2407
rect 16008 -2586 16018 -2407
rect 20414 -2583 20424 -2404
rect 20623 -2583 20633 -2404
rect 22312 -2583 22322 -2404
rect 22521 -2583 22531 -2404
rect 4266 -3113 4445 -3103
rect 4266 -3321 4445 -3312
rect 10824 -3117 11003 -3107
rect 10824 -3325 11003 -3316
rect 17358 -3112 17537 -3102
rect 17358 -3320 17537 -3311
rect 23871 -3109 24050 -3099
rect 23871 -3317 24050 -3308
rect 21766 -3402 21870 -3400
rect 25176 -3402 25268 -3401
rect 2161 -3406 2265 -3404
rect 15253 -3405 15357 -3403
rect 18663 -3405 18755 -3404
rect 5571 -3406 5663 -3405
rect 2161 -3410 5663 -3406
rect 2161 -3496 2175 -3410
rect 2253 -3496 5663 -3410
rect 2161 -3509 5663 -3496
rect 5571 -3569 5663 -3509
rect 8719 -3410 8823 -3408
rect 15253 -3409 18755 -3405
rect 12129 -3410 12221 -3409
rect 8719 -3414 12221 -3410
rect 8719 -3500 8733 -3414
rect 8811 -3500 12221 -3414
rect 8719 -3513 12221 -3500
rect 15253 -3495 15267 -3409
rect 15345 -3495 18755 -3409
rect 15253 -3508 18755 -3495
rect 21766 -3406 25268 -3402
rect 21766 -3492 21780 -3406
rect 21858 -3492 25268 -3406
rect 21766 -3505 25268 -3492
rect 5549 -3574 5684 -3569
rect 12129 -3573 12221 -3513
rect 18663 -3568 18755 -3508
rect 25176 -3565 25268 -3505
rect 18641 -3573 18776 -3568
rect 4525 -3848 4535 -3669
rect 4734 -3848 4744 -3669
rect 5549 -3671 5559 -3574
rect 5674 -3671 5684 -3574
rect 5549 -3676 5684 -3671
rect 12107 -3578 12242 -3573
rect 11083 -3852 11093 -3673
rect 11292 -3852 11302 -3673
rect 12107 -3675 12117 -3578
rect 12232 -3675 12242 -3578
rect 12107 -3680 12242 -3675
rect 17617 -3847 17627 -3668
rect 17826 -3847 17836 -3668
rect 18641 -3670 18651 -3573
rect 18766 -3670 18776 -3573
rect 25154 -3570 25289 -3565
rect 18641 -3675 18776 -3670
rect 24130 -3844 24140 -3665
rect 24339 -3844 24349 -3665
rect 25154 -3667 25164 -3570
rect 25279 -3667 25289 -3570
rect 25154 -3672 25289 -3667
rect 4271 -4717 4450 -4707
rect 865 -4996 875 -4817
rect 1074 -4996 1084 -4817
rect 2763 -4996 2773 -4817
rect 2972 -4996 2982 -4817
rect 10829 -4721 11008 -4711
rect 4271 -4925 4450 -4916
rect 7423 -5000 7433 -4821
rect 7632 -5000 7642 -4821
rect 9321 -5000 9331 -4821
rect 9530 -5000 9540 -4821
rect 17363 -4716 17542 -4706
rect 10829 -4929 11008 -4920
rect 13957 -4995 13967 -4816
rect 14166 -4995 14176 -4816
rect 15855 -4995 15865 -4816
rect 16064 -4995 16074 -4816
rect 23876 -4713 24055 -4703
rect 17363 -4924 17542 -4915
rect 20470 -4992 20480 -4813
rect 20679 -4992 20689 -4813
rect 22368 -4992 22378 -4813
rect 22577 -4992 22587 -4813
rect 23876 -4921 24055 -4912
<< via3 >>
rect 1339 5162 1538 5193
rect 1339 5033 1361 5162
rect 1361 5033 1514 5162
rect 1514 5033 1538 5162
rect 1339 5014 1538 5033
rect 3821 5216 4020 5247
rect 3821 5087 3843 5216
rect 3843 5087 3996 5216
rect 3996 5087 4020 5216
rect 3821 5068 4020 5087
rect 4968 5216 5167 5247
rect 4968 5087 4990 5216
rect 4990 5087 5143 5216
rect 5143 5087 5167 5216
rect 4968 5068 5167 5087
rect 7852 5159 8051 5190
rect 7852 5030 7874 5159
rect 7874 5030 8027 5159
rect 8027 5030 8051 5159
rect 7852 5011 8051 5030
rect 10334 5213 10533 5244
rect 10334 5084 10356 5213
rect 10356 5084 10509 5213
rect 10509 5084 10533 5213
rect 10334 5065 10533 5084
rect 11481 5213 11680 5244
rect 11481 5084 11503 5213
rect 11503 5084 11656 5213
rect 11656 5084 11680 5213
rect 11481 5065 11680 5084
rect 14386 5154 14585 5185
rect 14386 5025 14408 5154
rect 14408 5025 14561 5154
rect 14561 5025 14585 5154
rect 14386 5006 14585 5025
rect 16868 5208 17067 5239
rect 16868 5079 16890 5208
rect 16890 5079 17043 5208
rect 17043 5079 17067 5208
rect 16868 5060 17067 5079
rect 18015 5208 18214 5239
rect 18015 5079 18037 5208
rect 18037 5079 18190 5208
rect 18190 5079 18214 5208
rect 18015 5060 18214 5079
rect 20944 5158 21143 5189
rect 20944 5029 20966 5158
rect 20966 5029 21119 5158
rect 21119 5029 21143 5158
rect 20944 5010 21143 5029
rect 23426 5212 23625 5243
rect 23426 5083 23448 5212
rect 23448 5083 23601 5212
rect 23601 5083 23625 5212
rect 23426 5064 23625 5083
rect 24573 5212 24772 5243
rect 24573 5083 24595 5212
rect 24595 5083 24748 5212
rect 24748 5083 24772 5212
rect 24573 5064 24772 5083
rect 1623 4123 1802 4145
rect 1623 3970 1642 4123
rect 1642 3970 1771 4123
rect 1771 3970 1802 4123
rect 1623 3946 1802 3970
rect 8136 4120 8315 4142
rect 8136 3967 8155 4120
rect 8155 3967 8284 4120
rect 8284 3967 8315 4120
rect 8136 3943 8315 3967
rect 14670 4115 14849 4137
rect 14670 3962 14689 4115
rect 14689 3962 14818 4115
rect 14818 3962 14849 4115
rect 14670 3938 14849 3962
rect 21228 4119 21407 4141
rect 21228 3966 21247 4119
rect 21247 3966 21376 4119
rect 21376 3966 21407 4119
rect 21228 3942 21407 3966
rect 3166 3815 3365 3834
rect 3166 3686 3190 3815
rect 3190 3686 3343 3815
rect 3343 3686 3365 3815
rect 3166 3655 3365 3686
rect 4308 3813 4507 3832
rect 4308 3684 4332 3813
rect 4332 3684 4485 3813
rect 4485 3684 4507 3813
rect 4308 3653 4507 3684
rect 9679 3812 9878 3831
rect 9679 3683 9703 3812
rect 9703 3683 9856 3812
rect 9856 3683 9878 3812
rect 9679 3652 9878 3683
rect 10821 3810 11020 3829
rect 10821 3681 10845 3810
rect 10845 3681 10998 3810
rect 10998 3681 11020 3810
rect 10821 3650 11020 3681
rect 16213 3807 16412 3826
rect 16213 3678 16237 3807
rect 16237 3678 16390 3807
rect 16390 3678 16412 3807
rect 16213 3647 16412 3678
rect 17355 3805 17554 3824
rect 17355 3676 17379 3805
rect 17379 3676 17532 3805
rect 17532 3676 17554 3805
rect 17355 3645 17554 3676
rect 22771 3811 22970 3830
rect 22771 3682 22795 3811
rect 22795 3682 22948 3811
rect 22948 3682 22970 3811
rect 22771 3651 22970 3682
rect 23913 3809 24112 3828
rect 23913 3680 23937 3809
rect 23937 3680 24090 3809
rect 24090 3680 24112 3809
rect 23913 3649 24112 3680
rect 1353 3512 1552 3543
rect 1353 3383 1375 3512
rect 1375 3383 1528 3512
rect 1528 3383 1552 3512
rect 1353 3364 1552 3383
rect 7866 3509 8065 3540
rect 7866 3380 7888 3509
rect 7888 3380 8041 3509
rect 8041 3380 8065 3509
rect 7866 3361 8065 3380
rect 14400 3504 14599 3535
rect 14400 3375 14422 3504
rect 14422 3375 14575 3504
rect 14575 3375 14599 3504
rect 14400 3356 14599 3375
rect 20958 3508 21157 3539
rect 20958 3379 20980 3508
rect 20980 3379 21133 3508
rect 21133 3379 21157 3508
rect 20958 3360 21157 3379
rect 3166 3169 3365 3200
rect 3166 3040 3188 3169
rect 3188 3040 3341 3169
rect 3341 3040 3365 3169
rect 3166 3021 3365 3040
rect 5064 3169 5263 3200
rect 5064 3040 5086 3169
rect 5086 3040 5239 3169
rect 5239 3040 5263 3169
rect 5064 3021 5263 3040
rect 9679 3166 9878 3197
rect 9679 3037 9701 3166
rect 9701 3037 9854 3166
rect 9854 3037 9878 3166
rect 9679 3018 9878 3037
rect 11577 3166 11776 3197
rect 11577 3037 11599 3166
rect 11599 3037 11752 3166
rect 11752 3037 11776 3166
rect 11577 3018 11776 3037
rect 16213 3161 16412 3192
rect 16213 3032 16235 3161
rect 16235 3032 16388 3161
rect 16388 3032 16412 3161
rect 16213 3013 16412 3032
rect 18111 3161 18310 3192
rect 18111 3032 18133 3161
rect 18133 3032 18286 3161
rect 18286 3032 18310 3161
rect 18111 3013 18310 3032
rect 22771 3165 22970 3196
rect 22771 3036 22793 3165
rect 22793 3036 22946 3165
rect 22946 3036 22970 3165
rect 22771 3017 22970 3036
rect 24669 3165 24868 3196
rect 24669 3036 24691 3165
rect 24691 3036 24844 3165
rect 24844 3036 24868 3165
rect 24669 3017 24868 3036
rect 1637 2473 1816 2495
rect 1637 2320 1656 2473
rect 1656 2320 1785 2473
rect 1785 2320 1816 2473
rect 1637 2296 1816 2320
rect 8150 2470 8329 2492
rect 8150 2317 8169 2470
rect 8169 2317 8298 2470
rect 8298 2317 8329 2470
rect 8150 2293 8329 2317
rect 14684 2465 14863 2487
rect 14684 2312 14703 2465
rect 14703 2312 14832 2465
rect 14832 2312 14863 2465
rect 14684 2288 14863 2312
rect 21242 2469 21421 2491
rect 21242 2316 21261 2469
rect 21261 2316 21390 2469
rect 21390 2316 21421 2469
rect 21242 2292 21421 2316
rect 1348 1908 1547 1939
rect 1348 1779 1370 1908
rect 1370 1779 1523 1908
rect 1523 1779 1547 1908
rect 1348 1760 1547 1779
rect 7861 1905 8060 1936
rect 7861 1776 7883 1905
rect 7883 1776 8036 1905
rect 8036 1776 8060 1905
rect 7861 1757 8060 1776
rect 14395 1900 14594 1931
rect 14395 1771 14417 1900
rect 14417 1771 14570 1900
rect 14570 1771 14594 1900
rect 14395 1752 14594 1771
rect 20953 1904 21152 1935
rect 20953 1775 20975 1904
rect 20975 1775 21128 1904
rect 21128 1775 21152 1904
rect 20953 1756 21152 1775
rect 1632 869 1811 891
rect 1632 716 1651 869
rect 1651 716 1780 869
rect 1780 716 1811 869
rect 8145 866 8324 888
rect 1632 692 1811 716
rect 3110 772 3309 791
rect 3110 643 3134 772
rect 3134 643 3287 772
rect 3287 643 3309 772
rect 3110 612 3309 643
rect 5008 772 5207 791
rect 5008 643 5032 772
rect 5032 643 5185 772
rect 5185 643 5207 772
rect 5008 612 5207 643
rect 8145 713 8164 866
rect 8164 713 8293 866
rect 8293 713 8324 866
rect 14679 861 14858 883
rect 8145 689 8324 713
rect 9623 769 9822 788
rect 9623 640 9647 769
rect 9647 640 9800 769
rect 9800 640 9822 769
rect 9623 609 9822 640
rect 11521 769 11720 788
rect 11521 640 11545 769
rect 11545 640 11698 769
rect 11698 640 11720 769
rect 11521 609 11720 640
rect 14679 708 14698 861
rect 14698 708 14827 861
rect 14827 708 14858 861
rect 21237 865 21416 887
rect 14679 684 14858 708
rect 16157 764 16356 783
rect 16157 635 16181 764
rect 16181 635 16334 764
rect 16334 635 16356 764
rect 16157 604 16356 635
rect 18055 764 18254 783
rect 18055 635 18079 764
rect 18079 635 18232 764
rect 18232 635 18254 764
rect 18055 604 18254 635
rect 21237 712 21256 865
rect 21256 712 21385 865
rect 21385 712 21416 865
rect 21237 688 21416 712
rect 22715 768 22914 787
rect 22715 639 22739 768
rect 22739 639 22892 768
rect 22892 639 22914 768
rect 22715 608 22914 639
rect 24613 768 24812 787
rect 24613 639 24637 768
rect 24637 639 24790 768
rect 24790 639 24812 768
rect 24613 608 24812 639
rect 915 -392 1114 -361
rect 915 -521 939 -392
rect 939 -521 1092 -392
rect 1092 -521 1114 -392
rect 915 -540 1114 -521
rect 2062 -392 2261 -361
rect 2062 -521 2086 -392
rect 2086 -521 2239 -392
rect 2239 -521 2261 -392
rect 2062 -540 2261 -521
rect 4544 -446 4743 -415
rect 4544 -575 4568 -446
rect 4568 -575 4721 -446
rect 4721 -575 4743 -446
rect 4544 -594 4743 -575
rect 7473 -396 7672 -365
rect 7473 -525 7497 -396
rect 7497 -525 7650 -396
rect 7650 -525 7672 -396
rect 7473 -544 7672 -525
rect 8620 -396 8819 -365
rect 8620 -525 8644 -396
rect 8644 -525 8797 -396
rect 8797 -525 8819 -396
rect 8620 -544 8819 -525
rect 11102 -450 11301 -419
rect 11102 -579 11126 -450
rect 11126 -579 11279 -450
rect 11279 -579 11301 -450
rect 11102 -598 11301 -579
rect 14007 -391 14206 -360
rect 14007 -520 14031 -391
rect 14031 -520 14184 -391
rect 14184 -520 14206 -391
rect 14007 -539 14206 -520
rect 15154 -391 15353 -360
rect 15154 -520 15178 -391
rect 15178 -520 15331 -391
rect 15331 -520 15353 -391
rect 15154 -539 15353 -520
rect 17636 -445 17835 -414
rect 17636 -574 17660 -445
rect 17660 -574 17813 -445
rect 17813 -574 17835 -445
rect 17636 -593 17835 -574
rect 20520 -388 20719 -357
rect 20520 -517 20544 -388
rect 20544 -517 20697 -388
rect 20697 -517 20719 -388
rect 20520 -536 20719 -517
rect 21667 -388 21866 -357
rect 21667 -517 21691 -388
rect 21691 -517 21844 -388
rect 21844 -517 21866 -388
rect 21667 -536 21866 -517
rect 24149 -442 24348 -411
rect 24149 -571 24173 -442
rect 24173 -571 24326 -442
rect 24326 -571 24348 -442
rect 24149 -590 24348 -571
rect 4280 -1485 4459 -1463
rect 4280 -1638 4311 -1485
rect 4311 -1638 4440 -1485
rect 4440 -1638 4459 -1485
rect 4280 -1662 4459 -1638
rect 10838 -1489 11017 -1467
rect 10838 -1642 10869 -1489
rect 10869 -1642 10998 -1489
rect 10998 -1642 11017 -1489
rect 10838 -1666 11017 -1642
rect 17372 -1484 17551 -1462
rect 17372 -1637 17403 -1484
rect 17403 -1637 17532 -1484
rect 17532 -1637 17551 -1484
rect 17372 -1661 17551 -1637
rect 23885 -1481 24064 -1459
rect 23885 -1634 23916 -1481
rect 23916 -1634 24045 -1481
rect 24045 -1634 24064 -1481
rect 23885 -1658 24064 -1634
rect 1575 -1795 1774 -1776
rect 1575 -1924 1597 -1795
rect 1597 -1924 1750 -1795
rect 1750 -1924 1774 -1795
rect 1575 -1955 1774 -1924
rect 2717 -1793 2916 -1774
rect 2717 -1922 2739 -1793
rect 2739 -1922 2892 -1793
rect 2892 -1922 2916 -1793
rect 2717 -1953 2916 -1922
rect 8133 -1799 8332 -1780
rect 8133 -1928 8155 -1799
rect 8155 -1928 8308 -1799
rect 8308 -1928 8332 -1799
rect 8133 -1959 8332 -1928
rect 9275 -1797 9474 -1778
rect 9275 -1926 9297 -1797
rect 9297 -1926 9450 -1797
rect 9450 -1926 9474 -1797
rect 9275 -1957 9474 -1926
rect 14667 -1794 14866 -1775
rect 14667 -1923 14689 -1794
rect 14689 -1923 14842 -1794
rect 14842 -1923 14866 -1794
rect 14667 -1954 14866 -1923
rect 15809 -1792 16008 -1773
rect 15809 -1921 15831 -1792
rect 15831 -1921 15984 -1792
rect 15984 -1921 16008 -1792
rect 15809 -1952 16008 -1921
rect 21180 -1791 21379 -1772
rect 21180 -1920 21202 -1791
rect 21202 -1920 21355 -1791
rect 21355 -1920 21379 -1791
rect 21180 -1951 21379 -1920
rect 22322 -1789 22521 -1770
rect 22322 -1918 22344 -1789
rect 22344 -1918 22497 -1789
rect 22497 -1918 22521 -1789
rect 22322 -1949 22521 -1918
rect 4530 -2096 4729 -2065
rect 4530 -2225 4554 -2096
rect 4554 -2225 4707 -2096
rect 4707 -2225 4729 -2096
rect 4530 -2244 4729 -2225
rect 11088 -2100 11287 -2069
rect 11088 -2229 11112 -2100
rect 11112 -2229 11265 -2100
rect 11265 -2229 11287 -2100
rect 11088 -2248 11287 -2229
rect 17622 -2095 17821 -2064
rect 17622 -2224 17646 -2095
rect 17646 -2224 17799 -2095
rect 17799 -2224 17821 -2095
rect 17622 -2243 17821 -2224
rect 24135 -2092 24334 -2061
rect 24135 -2221 24159 -2092
rect 24159 -2221 24312 -2092
rect 24312 -2221 24334 -2092
rect 24135 -2240 24334 -2221
rect 819 -2439 1018 -2408
rect 819 -2568 843 -2439
rect 843 -2568 996 -2439
rect 996 -2568 1018 -2439
rect 819 -2587 1018 -2568
rect 2717 -2439 2916 -2408
rect 2717 -2568 2741 -2439
rect 2741 -2568 2894 -2439
rect 2894 -2568 2916 -2439
rect 2717 -2587 2916 -2568
rect 7377 -2443 7576 -2412
rect 7377 -2572 7401 -2443
rect 7401 -2572 7554 -2443
rect 7554 -2572 7576 -2443
rect 7377 -2591 7576 -2572
rect 9275 -2443 9474 -2412
rect 9275 -2572 9299 -2443
rect 9299 -2572 9452 -2443
rect 9452 -2572 9474 -2443
rect 9275 -2591 9474 -2572
rect 13911 -2438 14110 -2407
rect 13911 -2567 13935 -2438
rect 13935 -2567 14088 -2438
rect 14088 -2567 14110 -2438
rect 13911 -2586 14110 -2567
rect 15809 -2438 16008 -2407
rect 15809 -2567 15833 -2438
rect 15833 -2567 15986 -2438
rect 15986 -2567 16008 -2438
rect 15809 -2586 16008 -2567
rect 20424 -2435 20623 -2404
rect 20424 -2564 20448 -2435
rect 20448 -2564 20601 -2435
rect 20601 -2564 20623 -2435
rect 20424 -2583 20623 -2564
rect 22322 -2435 22521 -2404
rect 22322 -2564 22346 -2435
rect 22346 -2564 22499 -2435
rect 22499 -2564 22521 -2435
rect 22322 -2583 22521 -2564
rect 4266 -3135 4445 -3113
rect 4266 -3288 4297 -3135
rect 4297 -3288 4426 -3135
rect 4426 -3288 4445 -3135
rect 4266 -3312 4445 -3288
rect 10824 -3139 11003 -3117
rect 10824 -3292 10855 -3139
rect 10855 -3292 10984 -3139
rect 10984 -3292 11003 -3139
rect 10824 -3316 11003 -3292
rect 17358 -3134 17537 -3112
rect 17358 -3287 17389 -3134
rect 17389 -3287 17518 -3134
rect 17518 -3287 17537 -3134
rect 17358 -3311 17537 -3287
rect 23871 -3131 24050 -3109
rect 23871 -3284 23902 -3131
rect 23902 -3284 24031 -3131
rect 24031 -3284 24050 -3131
rect 23871 -3308 24050 -3284
rect 4535 -3700 4734 -3669
rect 4535 -3829 4559 -3700
rect 4559 -3829 4712 -3700
rect 4712 -3829 4734 -3700
rect 4535 -3848 4734 -3829
rect 11093 -3704 11292 -3673
rect 11093 -3833 11117 -3704
rect 11117 -3833 11270 -3704
rect 11270 -3833 11292 -3704
rect 11093 -3852 11292 -3833
rect 17627 -3699 17826 -3668
rect 17627 -3828 17651 -3699
rect 17651 -3828 17804 -3699
rect 17804 -3828 17826 -3699
rect 17627 -3847 17826 -3828
rect 24140 -3696 24339 -3665
rect 24140 -3825 24164 -3696
rect 24164 -3825 24317 -3696
rect 24317 -3825 24339 -3696
rect 24140 -3844 24339 -3825
rect 4271 -4739 4450 -4717
rect 875 -4836 1074 -4817
rect 875 -4965 897 -4836
rect 897 -4965 1050 -4836
rect 1050 -4965 1074 -4836
rect 875 -4996 1074 -4965
rect 2773 -4836 2972 -4817
rect 2773 -4965 2795 -4836
rect 2795 -4965 2948 -4836
rect 2948 -4965 2972 -4836
rect 2773 -4996 2972 -4965
rect 4271 -4892 4302 -4739
rect 4302 -4892 4431 -4739
rect 4431 -4892 4450 -4739
rect 10829 -4743 11008 -4721
rect 4271 -4916 4450 -4892
rect 7433 -4840 7632 -4821
rect 7433 -4969 7455 -4840
rect 7455 -4969 7608 -4840
rect 7608 -4969 7632 -4840
rect 7433 -5000 7632 -4969
rect 9331 -4840 9530 -4821
rect 9331 -4969 9353 -4840
rect 9353 -4969 9506 -4840
rect 9506 -4969 9530 -4840
rect 9331 -5000 9530 -4969
rect 10829 -4896 10860 -4743
rect 10860 -4896 10989 -4743
rect 10989 -4896 11008 -4743
rect 17363 -4738 17542 -4716
rect 10829 -4920 11008 -4896
rect 13967 -4835 14166 -4816
rect 13967 -4964 13989 -4835
rect 13989 -4964 14142 -4835
rect 14142 -4964 14166 -4835
rect 13967 -4995 14166 -4964
rect 15865 -4835 16064 -4816
rect 15865 -4964 15887 -4835
rect 15887 -4964 16040 -4835
rect 16040 -4964 16064 -4835
rect 15865 -4995 16064 -4964
rect 17363 -4891 17394 -4738
rect 17394 -4891 17523 -4738
rect 17523 -4891 17542 -4738
rect 23876 -4735 24055 -4713
rect 17363 -4915 17542 -4891
rect 20480 -4832 20679 -4813
rect 20480 -4961 20502 -4832
rect 20502 -4961 20655 -4832
rect 20655 -4961 20679 -4832
rect 20480 -4992 20679 -4961
rect 22378 -4832 22577 -4813
rect 22378 -4961 22400 -4832
rect 22400 -4961 22553 -4832
rect 22553 -4961 22577 -4832
rect 22378 -4992 22577 -4961
rect 23876 -4888 23907 -4735
rect 23907 -4888 24036 -4735
rect 24036 -4888 24055 -4735
rect 23876 -4912 24055 -4888
<< metal4 >>
rect 473 5544 1325 5555
rect 473 5514 22173 5544
rect 473 5349 25355 5514
rect 473 5247 25351 5349
rect 473 5193 3821 5247
rect 473 5014 1339 5193
rect 1538 5068 3821 5193
rect 4020 5068 4968 5247
rect 5167 5244 25351 5247
rect 5167 5190 10334 5244
rect 5167 5068 7852 5190
rect 1538 5014 7852 5068
rect 473 5011 7852 5014
rect 8051 5065 10334 5190
rect 10533 5065 11481 5244
rect 11680 5243 25351 5244
rect 11680 5239 23426 5243
rect 11680 5185 16868 5239
rect 11680 5065 14386 5185
rect 8051 5011 14386 5065
rect 473 5006 14386 5011
rect 14585 5060 16868 5185
rect 17067 5060 18015 5239
rect 18214 5189 23426 5239
rect 18214 5060 20944 5189
rect 14585 5010 20944 5060
rect 21143 5064 23426 5189
rect 23625 5064 24573 5243
rect 24772 5064 25351 5243
rect 21143 5010 25351 5064
rect 14585 5006 25351 5010
rect 473 4804 25351 5006
rect 473 3757 1325 4804
rect 473 3543 1693 3757
rect 473 3364 1353 3543
rect 1552 3375 1693 3543
rect 1552 3370 2038 3375
rect 3916 3370 4263 3373
rect 5130 3370 5746 4804
rect 1552 3364 5746 3370
rect 473 3200 5746 3364
rect 473 3021 3166 3200
rect 3365 3021 5064 3200
rect 5263 3021 5746 3200
rect 473 2865 5746 3021
rect 473 2135 1325 2865
rect 5130 2860 5746 2865
rect 7311 3540 8206 3754
rect 7311 3361 7866 3540
rect 8065 3372 8206 3540
rect 8065 3367 8551 3372
rect 10429 3367 10776 3370
rect 11643 3367 12259 4804
rect 14365 4800 18793 4804
rect 8065 3361 12259 3367
rect 7311 3197 12259 3361
rect 7311 3018 9679 3197
rect 9878 3018 11577 3197
rect 11776 3018 12259 3197
rect 7311 2862 12259 3018
rect 473 1939 2066 2135
rect 473 1760 1348 1939
rect 1547 1760 2066 1939
rect 473 1491 2066 1760
rect 7311 2132 7481 2862
rect 11643 2857 12259 2862
rect 13845 3535 14740 3749
rect 13845 3356 14400 3535
rect 14599 3367 14740 3535
rect 14599 3362 15085 3367
rect 16963 3362 17310 3365
rect 18177 3362 18793 4800
rect 14599 3356 18793 3362
rect 13845 3192 18793 3356
rect 13845 3013 16213 3192
rect 16412 3013 18111 3192
rect 18310 3013 18793 3192
rect 13845 2857 18793 3013
rect 7311 1936 8579 2132
rect 7311 1757 7861 1936
rect 8060 1757 8579 1936
rect 473 204 1325 1491
rect 7311 1488 8579 1757
rect 13845 2127 14015 2857
rect 18177 2852 18793 2857
rect 20403 3539 21298 3753
rect 20403 3360 20958 3539
rect 21157 3371 21298 3539
rect 21157 3366 21643 3371
rect 23521 3366 23868 3369
rect 24735 3366 25351 4804
rect 21157 3360 25351 3366
rect 20403 3196 25351 3360
rect 20403 3017 22771 3196
rect 22970 3017 24669 3196
rect 24868 3017 25351 3196
rect 20403 2861 25351 3017
rect 20403 2131 20573 2861
rect 24735 2856 25351 2861
rect 13845 1931 15113 2127
rect 13845 1752 14395 1931
rect 14594 1752 15113 1931
rect 13845 1483 15113 1752
rect 20403 1935 21671 2131
rect 20403 1756 20953 1935
rect 21152 1756 21671 1935
rect 20403 1487 21671 1756
rect 3086 791 3331 794
rect 3086 773 3110 791
rect 3309 773 3331 791
rect 4984 791 5229 794
rect 4984 773 5008 791
rect 5207 773 5229 791
rect 2982 469 3006 706
rect 3516 469 4852 655
rect 9599 788 9844 791
rect 9599 770 9623 788
rect 9822 770 9844 788
rect 11497 788 11742 791
rect 11497 770 11521 788
rect 11720 770 11742 788
rect 2982 464 5349 469
rect 9495 466 9519 703
rect 10029 466 11365 652
rect 16133 783 16378 786
rect 16133 765 16157 783
rect 16356 765 16378 783
rect 18031 783 18276 786
rect 18031 765 18055 783
rect 18254 765 18276 783
rect 3370 462 5041 464
rect 9495 461 11862 466
rect 16029 461 16053 698
rect 16563 461 17899 647
rect 22691 787 22936 790
rect 22691 769 22715 787
rect 22914 769 22936 787
rect 24589 787 24834 790
rect 24589 769 24613 787
rect 24812 769 24834 787
rect 22587 465 22611 702
rect 23121 465 24457 651
rect 9883 459 11554 461
rect 16029 456 18396 461
rect 22587 460 24954 465
rect 22975 458 24646 460
rect 16417 454 18088 456
rect 469 -90 1326 204
rect 24362 -72 25214 -60
rect 3526 -90 25214 -72
rect 465 -357 25214 -90
rect 465 -360 20520 -357
rect 465 -361 14007 -360
rect 465 -540 915 -361
rect 1114 -540 2062 -361
rect 2261 -365 14007 -361
rect 2261 -415 7473 -365
rect 2261 -540 4544 -415
rect 465 -594 4544 -540
rect 4743 -544 7473 -415
rect 7672 -544 8620 -365
rect 8819 -419 14007 -365
rect 8819 -544 11102 -419
rect 4743 -594 11102 -544
rect 465 -598 11102 -594
rect 11301 -539 14007 -419
rect 14206 -539 15154 -360
rect 15353 -414 20520 -360
rect 15353 -539 17636 -414
rect 11301 -593 17636 -539
rect 17835 -536 20520 -414
rect 20719 -536 21667 -357
rect 21866 -411 25214 -357
rect 21866 -536 24149 -411
rect 17835 -590 24149 -536
rect 24348 -590 25214 -411
rect 17835 -593 25214 -590
rect 11301 -598 25214 -593
rect 465 -800 25214 -598
rect 465 -2238 952 -800
rect 3526 -812 25214 -800
rect 4389 -2065 5284 -1851
rect 4389 -2233 4530 -2065
rect 1819 -2238 2166 -2235
rect 4044 -2238 4530 -2233
rect 465 -2244 4530 -2238
rect 4729 -2244 5284 -2065
rect 465 -2408 5284 -2244
rect 465 -2587 819 -2408
rect 1018 -2587 2717 -2408
rect 2916 -2587 5284 -2408
rect 465 -2743 5284 -2587
rect 465 -2748 952 -2743
rect 5114 -3473 5284 -2743
rect 6894 -2242 7510 -812
rect 10947 -2069 11842 -1855
rect 10947 -2237 11088 -2069
rect 8377 -2242 8724 -2239
rect 10602 -2242 11088 -2237
rect 6894 -2248 11088 -2242
rect 11287 -2248 11842 -2069
rect 6894 -2412 11842 -2248
rect 6894 -2591 7377 -2412
rect 7576 -2591 9275 -2412
rect 9474 -2591 11842 -2412
rect 6894 -2747 11842 -2591
rect 13428 -2237 14044 -812
rect 17481 -2064 18376 -1850
rect 17481 -2232 17622 -2064
rect 14911 -2237 15258 -2234
rect 17136 -2237 17622 -2232
rect 13428 -2243 17622 -2237
rect 17821 -2243 18376 -2064
rect 13428 -2407 18376 -2243
rect 13428 -2586 13911 -2407
rect 14110 -2586 15809 -2407
rect 16008 -2586 18376 -2407
rect 13428 -2742 18376 -2586
rect 13428 -2747 14044 -2742
rect 6894 -2752 7510 -2747
rect 4016 -3669 5284 -3473
rect 11672 -3477 11842 -2747
rect 18206 -3472 18376 -2742
rect 19941 -2234 20557 -812
rect 24362 -845 25214 -812
rect 23994 -2061 24889 -1847
rect 23994 -2229 24135 -2061
rect 21424 -2234 21771 -2231
rect 23649 -2234 24135 -2229
rect 19941 -2240 24135 -2234
rect 24334 -2240 24889 -2061
rect 19941 -2404 24889 -2240
rect 19941 -2583 20424 -2404
rect 20623 -2583 22322 -2404
rect 22521 -2583 24889 -2404
rect 19941 -2739 24889 -2583
rect 19941 -2744 20557 -2739
rect 24719 -3469 24889 -2739
rect 4016 -3848 4535 -3669
rect 4734 -3848 5284 -3669
rect 4016 -4117 5284 -3848
rect 10574 -3673 11842 -3477
rect 10574 -3852 11093 -3673
rect 11292 -3852 11842 -3673
rect 10574 -4121 11842 -3852
rect 17108 -3668 18376 -3472
rect 17108 -3847 17627 -3668
rect 17826 -3847 18376 -3668
rect 17108 -4116 18376 -3847
rect 23621 -3665 24889 -3469
rect 23621 -3844 24140 -3665
rect 24339 -3844 24889 -3665
rect 23621 -4113 24889 -3844
rect 853 -4817 1098 -4814
rect 853 -4835 875 -4817
rect 1074 -4835 1098 -4817
rect 2751 -4817 2996 -4814
rect 2751 -4835 2773 -4817
rect 2972 -4835 2996 -4817
rect 1230 -5139 2566 -4953
rect 3076 -5139 3100 -4902
rect 7411 -4821 7656 -4818
rect 7411 -4839 7433 -4821
rect 7632 -4839 7656 -4821
rect 9309 -4821 9554 -4818
rect 9309 -4839 9331 -4821
rect 9530 -4839 9554 -4821
rect 733 -5144 3100 -5139
rect 7788 -5143 9124 -4957
rect 9634 -5143 9658 -4906
rect 13945 -4816 14190 -4813
rect 13945 -4834 13967 -4816
rect 14166 -4834 14190 -4816
rect 15843 -4816 16088 -4813
rect 15843 -4834 15865 -4816
rect 16064 -4834 16088 -4816
rect 14322 -5138 15658 -4952
rect 16168 -5138 16192 -4901
rect 20458 -4813 20703 -4810
rect 20458 -4831 20480 -4813
rect 20679 -4831 20703 -4813
rect 22356 -4813 22601 -4810
rect 22356 -4831 22378 -4813
rect 22577 -4831 22601 -4813
rect 20835 -5135 22171 -4949
rect 22681 -5135 22705 -4898
rect 13825 -5143 16192 -5138
rect 20338 -5140 22705 -5135
rect 20646 -5142 22317 -5140
rect 1041 -5146 2712 -5144
rect 7291 -5148 9658 -5143
rect 14133 -5145 15804 -5143
rect 7599 -5150 9270 -5148
<< via4 >>
rect 1564 4145 2074 4223
rect 1564 3946 1623 4145
rect 1623 3946 1802 4145
rect 1802 3946 2074 4145
rect 1564 3919 2074 3946
rect 3132 3834 3436 3985
rect 3132 3655 3166 3834
rect 3166 3655 3365 3834
rect 3365 3655 3436 3834
rect 3132 3475 3436 3655
rect 4266 3832 4570 3995
rect 4266 3653 4308 3832
rect 4308 3653 4507 3832
rect 4507 3653 4570 3832
rect 4266 3485 4570 3653
rect 8077 4142 8587 4220
rect 8077 3943 8136 4142
rect 8136 3943 8315 4142
rect 8315 3943 8587 4142
rect 8077 3916 8587 3943
rect 9645 3831 9949 3982
rect 9645 3652 9679 3831
rect 9679 3652 9878 3831
rect 9878 3652 9949 3831
rect 9645 3472 9949 3652
rect 10779 3829 11083 3992
rect 10779 3650 10821 3829
rect 10821 3650 11020 3829
rect 11020 3650 11083 3829
rect 10779 3482 11083 3650
rect 14611 4137 15121 4215
rect 14611 3938 14670 4137
rect 14670 3938 14849 4137
rect 14849 3938 15121 4137
rect 14611 3911 15121 3938
rect 16179 3826 16483 3977
rect 1558 2495 2068 2563
rect 1558 2296 1637 2495
rect 1637 2296 1816 2495
rect 1816 2296 2068 2495
rect 1558 2259 2068 2296
rect 16179 3647 16213 3826
rect 16213 3647 16412 3826
rect 16412 3647 16483 3826
rect 16179 3467 16483 3647
rect 17313 3824 17617 3987
rect 17313 3645 17355 3824
rect 17355 3645 17554 3824
rect 17554 3645 17617 3824
rect 17313 3477 17617 3645
rect 21169 4141 21679 4219
rect 21169 3942 21228 4141
rect 21228 3942 21407 4141
rect 21407 3942 21679 4141
rect 21169 3915 21679 3942
rect 22737 3830 23041 3981
rect 8071 2492 8581 2560
rect 8071 2293 8150 2492
rect 8150 2293 8329 2492
rect 8329 2293 8581 2492
rect 8071 2256 8581 2293
rect 22737 3651 22771 3830
rect 22771 3651 22970 3830
rect 22970 3651 23041 3830
rect 22737 3471 23041 3651
rect 23871 3828 24175 3991
rect 23871 3649 23913 3828
rect 23913 3649 24112 3828
rect 24112 3649 24175 3828
rect 23871 3481 24175 3649
rect 14605 2487 15115 2555
rect 14605 2288 14684 2487
rect 14684 2288 14863 2487
rect 14863 2288 15115 2487
rect 14605 2251 15115 2288
rect 21163 2491 21673 2559
rect 21163 2292 21242 2491
rect 21242 2292 21421 2491
rect 21421 2292 21673 2491
rect 21163 2255 21673 2292
rect 1557 891 2067 958
rect 1557 692 1632 891
rect 1632 692 1811 891
rect 1811 692 2067 891
rect 8070 888 8580 955
rect 1557 654 2067 692
rect 3006 612 3110 773
rect 3110 612 3309 773
rect 3309 612 3516 773
rect 3006 469 3516 612
rect 4852 612 5008 773
rect 5008 612 5207 773
rect 5207 612 5362 773
rect 8070 689 8145 888
rect 8145 689 8324 888
rect 8324 689 8580 888
rect 14604 883 15114 950
rect 8070 651 8580 689
rect 4852 469 5362 612
rect 9519 609 9623 770
rect 9623 609 9822 770
rect 9822 609 10029 770
rect 9519 466 10029 609
rect 11365 609 11521 770
rect 11521 609 11720 770
rect 11720 609 11875 770
rect 14604 684 14679 883
rect 14679 684 14858 883
rect 14858 684 15114 883
rect 21162 887 21672 954
rect 14604 646 15114 684
rect 11365 466 11875 609
rect 16053 604 16157 765
rect 16157 604 16356 765
rect 16356 604 16563 765
rect 16053 461 16563 604
rect 17899 604 18055 765
rect 18055 604 18254 765
rect 18254 604 18409 765
rect 21162 688 21237 887
rect 21237 688 21416 887
rect 21416 688 21672 887
rect 21162 650 21672 688
rect 17899 461 18409 604
rect 22611 608 22715 769
rect 22715 608 22914 769
rect 22914 608 23121 769
rect 22611 465 23121 608
rect 24457 608 24613 769
rect 24613 608 24812 769
rect 24812 608 24967 769
rect 24457 465 24967 608
rect 4008 -1463 4518 -1385
rect 1512 -1776 1816 -1613
rect 1512 -1955 1575 -1776
rect 1575 -1955 1774 -1776
rect 1774 -1955 1816 -1776
rect 1512 -2123 1816 -1955
rect 2646 -1774 2950 -1623
rect 4008 -1662 4280 -1463
rect 4280 -1662 4459 -1463
rect 4459 -1662 4518 -1463
rect 4008 -1689 4518 -1662
rect 2646 -1953 2717 -1774
rect 2717 -1953 2916 -1774
rect 2916 -1953 2950 -1774
rect 2646 -2133 2950 -1953
rect 4014 -3113 4524 -3045
rect 4014 -3312 4266 -3113
rect 4266 -3312 4445 -3113
rect 4445 -3312 4524 -3113
rect 4014 -3349 4524 -3312
rect 10566 -1467 11076 -1389
rect 8070 -1780 8374 -1617
rect 8070 -1959 8133 -1780
rect 8133 -1959 8332 -1780
rect 8332 -1959 8374 -1780
rect 8070 -2127 8374 -1959
rect 9204 -1778 9508 -1627
rect 10566 -1666 10838 -1467
rect 10838 -1666 11017 -1467
rect 11017 -1666 11076 -1467
rect 10566 -1693 11076 -1666
rect 9204 -1957 9275 -1778
rect 9275 -1957 9474 -1778
rect 9474 -1957 9508 -1778
rect 9204 -2137 9508 -1957
rect 17100 -1462 17610 -1384
rect 14604 -1775 14908 -1612
rect 14604 -1954 14667 -1775
rect 14667 -1954 14866 -1775
rect 14866 -1954 14908 -1775
rect 14604 -2122 14908 -1954
rect 15738 -1773 16042 -1622
rect 17100 -1661 17372 -1462
rect 17372 -1661 17551 -1462
rect 17551 -1661 17610 -1462
rect 17100 -1688 17610 -1661
rect 15738 -1952 15809 -1773
rect 15809 -1952 16008 -1773
rect 16008 -1952 16042 -1773
rect 15738 -2132 16042 -1952
rect 10572 -3117 11082 -3049
rect 10572 -3316 10824 -3117
rect 10824 -3316 11003 -3117
rect 11003 -3316 11082 -3117
rect 10572 -3353 11082 -3316
rect 17106 -3112 17616 -3044
rect 17106 -3311 17358 -3112
rect 17358 -3311 17537 -3112
rect 17537 -3311 17616 -3112
rect 17106 -3348 17616 -3311
rect 23613 -1459 24123 -1381
rect 21117 -1772 21421 -1609
rect 21117 -1951 21180 -1772
rect 21180 -1951 21379 -1772
rect 21379 -1951 21421 -1772
rect 21117 -2119 21421 -1951
rect 22251 -1770 22555 -1619
rect 23613 -1658 23885 -1459
rect 23885 -1658 24064 -1459
rect 24064 -1658 24123 -1459
rect 23613 -1685 24123 -1658
rect 22251 -1949 22322 -1770
rect 22322 -1949 22521 -1770
rect 22521 -1949 22555 -1770
rect 22251 -2129 22555 -1949
rect 23619 -3109 24129 -3041
rect 23619 -3308 23871 -3109
rect 23871 -3308 24050 -3109
rect 24050 -3308 24129 -3109
rect 23619 -3345 24129 -3308
rect 4015 -4717 4525 -4650
rect 720 -4996 875 -4835
rect 875 -4996 1074 -4835
rect 1074 -4996 1230 -4835
rect 720 -5139 1230 -4996
rect 2566 -4996 2773 -4835
rect 2773 -4996 2972 -4835
rect 2972 -4996 3076 -4835
rect 2566 -5139 3076 -4996
rect 4015 -4916 4271 -4717
rect 4271 -4916 4450 -4717
rect 4450 -4916 4525 -4717
rect 10573 -4721 11083 -4654
rect 4015 -4954 4525 -4916
rect 7278 -5000 7433 -4839
rect 7433 -5000 7632 -4839
rect 7632 -5000 7788 -4839
rect 7278 -5143 7788 -5000
rect 9124 -5000 9331 -4839
rect 9331 -5000 9530 -4839
rect 9530 -5000 9634 -4839
rect 9124 -5143 9634 -5000
rect 10573 -4920 10829 -4721
rect 10829 -4920 11008 -4721
rect 11008 -4920 11083 -4721
rect 17107 -4716 17617 -4649
rect 10573 -4958 11083 -4920
rect 13812 -4995 13967 -4834
rect 13967 -4995 14166 -4834
rect 14166 -4995 14322 -4834
rect 13812 -5138 14322 -4995
rect 15658 -4995 15865 -4834
rect 15865 -4995 16064 -4834
rect 16064 -4995 16168 -4834
rect 15658 -5138 16168 -4995
rect 17107 -4915 17363 -4716
rect 17363 -4915 17542 -4716
rect 17542 -4915 17617 -4716
rect 23620 -4713 24130 -4646
rect 17107 -4953 17617 -4915
rect 20325 -4992 20480 -4831
rect 20480 -4992 20679 -4831
rect 20679 -4992 20835 -4831
rect 20325 -5135 20835 -4992
rect 22171 -4992 22378 -4831
rect 22378 -4992 22577 -4831
rect 22577 -4992 22681 -4831
rect 22171 -5135 22681 -4992
rect 23620 -4912 23876 -4713
rect 23876 -4912 24055 -4713
rect 24055 -4912 24130 -4713
rect 23620 -4950 24130 -4912
<< metal5 >>
rect 1413 4223 5387 4387
rect 1413 3919 1564 4223
rect 2074 3995 5387 4223
rect 2074 3985 4266 3995
rect 2074 3919 3132 3985
rect 1413 3475 3132 3919
rect 3436 3485 4266 3985
rect 4570 3485 5387 3995
rect 3436 3475 5387 3485
rect 1413 3262 5387 3475
rect 7926 4220 11900 4384
rect 7926 3916 8077 4220
rect 8587 3992 11900 4220
rect 8587 3982 10779 3992
rect 8587 3916 9645 3982
rect 7926 3472 9645 3916
rect 9949 3482 10779 3982
rect 11083 3482 11900 3992
rect 9949 3472 11900 3482
rect 7926 3262 11900 3472
rect 14460 4215 18434 4379
rect 14460 3911 14611 4215
rect 15121 3987 18434 4215
rect 15121 3977 17313 3987
rect 15121 3911 16179 3977
rect 14460 3467 16179 3911
rect 16483 3477 17313 3977
rect 17617 3477 18434 3987
rect 16483 3467 18434 3477
rect 14460 3262 18434 3467
rect 21018 4219 24992 4383
rect 21018 3915 21169 4219
rect 21679 3991 24992 4219
rect 21679 3981 23871 3991
rect 21679 3915 22737 3981
rect 21018 3471 22737 3915
rect 23041 3481 23871 3981
rect 24175 3481 24992 3991
rect 23041 3471 24992 3481
rect 21018 3262 24992 3471
rect 25634 3262 26647 3263
rect 1401 2716 26647 3262
rect 1413 2563 5387 2716
rect 1413 2259 1558 2563
rect 2068 2259 5387 2563
rect 1413 958 5387 2259
rect 1413 654 1557 958
rect 2067 773 5387 958
rect 2067 654 3006 773
rect 1413 469 3006 654
rect 3516 469 4852 773
rect 5362 469 5387 773
rect 1413 455 5387 469
rect 7926 2560 11900 2716
rect 7926 2256 8071 2560
rect 8581 2256 11900 2560
rect 7926 955 11900 2256
rect 7926 651 8070 955
rect 8580 770 11900 955
rect 8580 651 9519 770
rect 7926 466 9519 651
rect 10029 466 11365 770
rect 11875 466 11900 770
rect 7926 455 11900 466
rect 14460 2555 18434 2716
rect 14460 2251 14605 2555
rect 15115 2251 18434 2555
rect 14460 950 18434 2251
rect 14460 646 14604 950
rect 15114 765 18434 950
rect 15114 646 16053 765
rect 14460 461 16053 646
rect 16563 461 17899 765
rect 18409 461 18434 765
rect 14460 455 18434 461
rect 21018 2559 24992 2716
rect 21018 2255 21163 2559
rect 21673 2255 24992 2559
rect 21018 954 24992 2255
rect 21018 650 21162 954
rect 21672 769 24992 954
rect 21672 650 22611 769
rect 21018 465 22611 650
rect 23121 465 24457 769
rect 24967 465 24992 769
rect 25890 623 26647 2716
rect 21018 455 24992 465
rect 25889 455 26650 623
rect 1413 0 26650 455
rect 5065 -24 26650 0
rect 695 -1385 4669 -1221
rect 695 -1613 4008 -1385
rect 695 -2123 1512 -1613
rect 1816 -1623 4008 -1613
rect 1816 -2123 2646 -1623
rect 695 -2133 2646 -2123
rect 2950 -1689 4008 -1623
rect 4518 -1689 4669 -1385
rect 2950 -2133 4669 -1689
rect 695 -2362 4669 -2133
rect 7253 -1389 11227 -1225
rect 7253 -1617 10566 -1389
rect 7253 -2127 8070 -1617
rect 8374 -1627 10566 -1617
rect 8374 -2127 9204 -1627
rect 7253 -2137 9204 -2127
rect 9508 -1693 10566 -1627
rect 11076 -1693 11227 -1389
rect 9508 -2137 11227 -1693
rect 7253 -2362 11227 -2137
rect 13787 -1384 17761 -1220
rect 13787 -1612 17100 -1384
rect 13787 -2122 14604 -1612
rect 14908 -1622 17100 -1612
rect 14908 -2122 15738 -1622
rect 13787 -2132 15738 -2122
rect 16042 -1688 17100 -1622
rect 17610 -1688 17761 -1384
rect 16042 -2132 17761 -1688
rect 13787 -2362 17761 -2132
rect 20300 -1381 24274 -1217
rect 20300 -1609 23613 -1381
rect 20300 -2119 21117 -1609
rect 21421 -1619 23613 -1609
rect 21421 -2119 22251 -1619
rect 20300 -2129 22251 -2119
rect 22555 -1685 23613 -1619
rect 24123 -1685 24274 -1381
rect 22555 -2129 24274 -1685
rect 20300 -2359 24274 -2129
rect 25889 -2359 26650 -24
rect 18587 -2362 26650 -2359
rect 465 -2908 26650 -2362
rect 695 -3045 4669 -2908
rect 695 -3349 4014 -3045
rect 4524 -3349 4669 -3045
rect 695 -4650 4669 -3349
rect 695 -4835 4015 -4650
rect 695 -5135 720 -4835
rect 465 -5139 720 -5135
rect 1230 -5139 2566 -4835
rect 3076 -4954 4015 -4835
rect 4525 -4954 4669 -4650
rect 3076 -5135 4669 -4954
rect 7253 -3049 11227 -2908
rect 7253 -3353 10572 -3049
rect 11082 -3353 11227 -3049
rect 7253 -4654 11227 -3353
rect 7253 -4839 10573 -4654
rect 7253 -5135 7278 -4839
rect 3076 -5139 7278 -5135
rect 465 -5143 7278 -5139
rect 7788 -5143 9124 -4839
rect 9634 -4958 10573 -4839
rect 11083 -4958 11227 -4654
rect 9634 -5135 11227 -4958
rect 13787 -3044 17761 -2908
rect 18587 -2922 26650 -2908
rect 13787 -3348 17106 -3044
rect 17616 -3348 17761 -3044
rect 13787 -4649 17761 -3348
rect 13787 -4834 17107 -4649
rect 13787 -5135 13812 -4834
rect 9634 -5138 13812 -5135
rect 14322 -5138 15658 -4834
rect 16168 -4953 17107 -4834
rect 17617 -4953 17761 -4649
rect 16168 -5135 17761 -4953
rect 20300 -3041 24274 -2922
rect 20300 -3345 23619 -3041
rect 24129 -3345 24274 -3041
rect 20300 -4646 24274 -3345
rect 20300 -4831 23620 -4646
rect 20300 -5135 20325 -4831
rect 20835 -5135 22171 -4831
rect 22681 -4950 23620 -4831
rect 24130 -4950 24274 -4646
rect 22681 -5129 24274 -4950
rect 25889 -5129 26650 -2922
rect 22681 -5135 26650 -5129
rect 16168 -5138 26650 -5135
rect 9634 -5143 26650 -5138
rect 465 -5625 26650 -5143
rect 23224 -5634 26650 -5625
rect 23224 -5646 26648 -5634
<< labels >>
flabel metal1 16 3956 246 4163 1 FreeSans 400 0 0 0 A[0]
port 1 n
flabel metal1 29 3425 259 3632 1 FreeSans 400 0 0 0 B[0]
port 2 n
flabel metal1 29 2306 259 2513 1 FreeSans 400 0 0 0 carry_in
port 3 n
flabel viali 6103 1591 6235 1688 1 FreeSans 400 0 0 0 Y[0]
port 4 n
flabel metal1 6522 3944 6771 4155 1 FreeSans 400 0 0 0 A[1]
port 5 n
flabel metal1 6536 3424 6785 3635 1 FreeSans 400 0 0 0 B[1]
port 6 n
flabel metal1 13058 3941 13307 4152 1 FreeSans 400 0 0 0 A[2]
port 7 n
flabel metal1 13075 3415 13324 3626 1 FreeSans 400 0 0 0 B[2]
port 8 n
flabel metal1 19616 3946 19865 4154 1 FreeSans 400 0 0 0 A[3]
port 9 n
flabel metal1 19634 3409 19883 3617 1 FreeSans 400 0 0 0 B[3]
port 10 n
flabel metal1 12616 1587 12750 1686 1 FreeSans 400 0 0 0 Y[1]
port 11 n
flabel metal1 19150 1582 19284 1681 1 FreeSans 400 0 0 0 Y[2]
port 12 n
flabel metal1 25707 1586 25841 1685 1 FreeSans 400 0 0 0 Y[3]
port 13 n
flabel metal1 25425 -1653 25677 -1445 1 FreeSans 400 0 0 0 A[4]
port 14 n
flabel metal1 25413 -2182 25665 -1974 1 FreeSans 400 0 0 0 B[4]
port 15 n
flabel metal1 18913 -1654 19165 -1446 1 FreeSans 400 0 0 0 A[5]
port 16 n
flabel metal1 18896 -2180 19148 -1972 1 FreeSans 400 0 0 0 B[5]
port 17 n
flabel metal1 12363 -2180 12615 -1972 1 FreeSans 400 0 0 0 B[6]
port 18 n
flabel metal1 12380 -1658 12632 -1450 1 FreeSans 400 0 0 0 A[6]
port 19 n
flabel metal1 5821 -1658 6073 -1450 1 FreeSans 400 0 0 0 A[7]
port 20 n
flabel metal1 5804 -2182 6056 -1974 1 FreeSans 400 0 0 0 B[7]
port 21 n
flabel metal1 19452 -4014 19586 -3913 1 FreeSans 400 0 0 0 Y[4]
port 22 n
flabel metal1 12938 -4017 13072 -3916 1 FreeSans 400 0 0 0 Y[5]
port 23 n
flabel metal1 6405 -4023 6539 -3922 1 FreeSans 400 0 0 0 Y[6]
port 24 n
flabel metal1 -154 -4019 -20 -3918 1 FreeSans 400 0 0 0 Y[7]
port 25 n
flabel metal5 11869 -5605 13554 -5281 1 FreeSans 1600 0 0 0 VSS
port 27 n
flabel metal4 11874 5051 13559 5375 1 FreeSans 1600 0 0 0 VDD
port 28 n
flabel metal1 -120 -1302 42 -1246 1 FreeSans 480 0 0 0 carry_out
port 29 n
<< end >>
