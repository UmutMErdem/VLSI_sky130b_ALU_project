* NGSPICE file created from array_multiplier_pex.ext - technology: sky130B

.subckt array_multiplier A[0],A[1],A[2],A[3] B[0],B[1],B[2],B[3] VDD VSS Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7]
X0 a_16803_n2942.t3 a_16213_n2505.t7 VSS.t95 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1 VDD.t641 a_6818_316.t8 a_32246_4888.t2 VDD.t640 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2 a_13367_404.t4 a_12822_1097.t4 a_13249_404.t1 VDD.t397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3 VDD.t262 a_16227_42.t7 a_16817_n395.t3 VDD.t261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4 a_7112_290.t3 a_2969_1600.t4 VDD.t399 VDD.t398 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 a_13367_404.t1 a_12822_1097.t5 a_13367_n328.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X6 a_24630_404.t7 a_19826_n3212.t4 VDD.t202 VDD.t201 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 a_10918_n4773.t3 a_7414_n7824.t4 VDD.t1570 VDD.t1569 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8 a_18425_3168.t3 a_16817_n395.t4 a_18543_3168.t2 VDD.t1611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X9 a_3619_1189.t3 a_3029_1626.t7 VDD.t350 VDD.t349 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10 Y[3].t6 a_30337_n7043.t4 a_30882_n8468.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 a_12035_2653.t3 a_11771_3236.t5 VDD.t510 VDD.t509 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X12 VDD.t1467 a_25042_n2632.t5 a_25306_n3215.t3 VDD.t1466 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X13 VDD.t485 a_11463_n5466.t8 a_12816_n4773.t3 VDD.t484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X14 VDD.t1414 A[0].t0 a_28645_5296.t3 VDD.t1413 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X15 a_26302_n2628.t2 a_25306_n3215.t4 VDD.t823 VDD.t822 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X16 a_25160_n2632.t4 a_23425_n2941.t4 VDD.t1213 VDD.t1212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 VDD.t1598 a_18689_2585.t4 a_19685_3172.t3 VDD.t1597 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 VDD.t601 a_13367_404.t8 a_16232_1646.t5 VDD.t600 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X19 a_28640_n308.t3 A[1].t0 VDD.t855 VDD.t854 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X20 VDD.t901 B[1].t0 a_125_3543.t6 VDD.t900 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X21 a_19903_336.t9 a_18123_336.t8 VDD.t952 VDD.t951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X22 a_16822_1209.t3 a_16232_1646.t7 VDD.t833 VDD.t832 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X23 a_9573_110.t4 a_7379_5006.t4 VDD.t1282 VDD.t1281 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X24 a_23072_n3141.t0 a_20016_n5465.t8 a_22835_n2504.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X25 a_6692_n5464.t4 a_2961_n4180.t4 VDD.t1310 VDD.t1309 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X26 VDD.t245 a_19562_n2629.t5 a_19826_n3212.t0 VDD.t244 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X27 a_22789_n4180.t0 a_32248_n2698.t7 VSS.t28 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 a_31176_n7762.t0 a_13361_n5466.t8 VSS.t69 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X29 a_26520_n5464.t4 a_24740_n5464.t8 VDD.t1491 VDD.t1490 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X30 a_715_3106.t3 a_125_3543.t7 VDD.t909 VDD.t908 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X31 a_16822_1209.t0 a_16232_1646.t8 VSS.t109 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X32 a_30764_107.t2 a_29301_n2665.t4 VDD.t257 VDD.t256 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X33 VDD.t689 a_29305_n8580.t4 a_32248_n7046.t2 VDD.t688 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X34 VDD.t467 a_22844_n5758.t7 a_23434_n6195.t3 VDD.t466 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X35 a_715_3106.t0 a_125_3543.t8 VSS.t149 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X36 VDD.t825 a_25306_n3215.t5 a_26302_n2628.t1 VDD.t824 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X37 VDD.t259 a_16172_1620.t4 a_19903_336.t2 VDD.t258 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X38 VDD.t1209 a_23425_n2941.t5 a_25160_n2632.t3 VDD.t1208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 a_16222_n5759.t3 a_13177_2657.t4 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X40 a_3605_2839.t3 a_3015_3276.t7 VDD.t1447 VDD.t1446 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X41 a_6700_316.t2 a_4920_316.t8 VDD.t538 VDD.t537 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X42 VDD.t149 a_3024_22.t7 a_3614_n415.t3 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X43 VSS.t142 a_707_521.t4 a_4375_1009.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X44 a_10163_n327.t3 a_9573_110.t7 VDD.t1249 VDD.t1248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X45 a_6824_n8261.t5 B[2].t0 VDD.t548 VDD.t547 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X46 a_32248_797.t2 a_29301_n2665.t5 VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X47 Y[1].t5 a_31176_81.t4 a_30764_107.t7 VDD.t877 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X48 a_24976_n6196.t1 a_20617_n7831.t4 a_24740_n5464.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X49 VDD.t603 a_13367_404.t9 a_16218_3296.t6 VDD.t602 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X50 VDD.t1106 a_11469_404.t8 a_12822_1097.t0 VDD.t1105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X51 VSS.t91 a_20617_n7831.t5 a_23072_n3141.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X52 VDD.t1312 a_2961_n4180.t5 a_6692_n5464.t3 VDD.t1311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X53 a_19826_n3212.t1 a_19562_n2629.t6 VDD.t247 VDD.t246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X54 a_26932_n5490.t0 a_22789_n4180.t4 VSS.t105 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X55 a_26520_n5464.t8 a_26932_n5490.t4 Y[5].t2 VDD.t686 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X56 VDD.t1493 a_24740_n5464.t9 a_26520_n5464.t3 VDD.t1492 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X57 a_9512_n4182.t0 a_32246_4888.t7 VSS.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X58 VSS.t79 a_13367_404.t10 a_16469_1009.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X59 a_23447_1277.t3 a_22857_1714.t7 VDD.t1062 VDD.t1061 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X60 a_24203_1097.t3 a_19826_n3212.t5 VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X61 a_12907_n2630.t0 a_10162_n4593.t4 VSS.t37 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X62 a_16172_1620.t3 a_32248_n7046.t7 VDD.t74 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 a_18000_n5465.t4 a_13968_n7819.t4 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X64 VDD.t550 B[2].t1 a_6824_n8261.t4 VDD.t549 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X65 a_22844_n5758.t3 a_20016_n5465.t9 VDD.t1241 VDD.t1240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X66 VDD.t368 a_704_n5517.t4 a_4794_n5464.t9 VDD.t367 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X67 VDD.t1058 a_22849_n4154.t7 a_23439_n4591.t3 VDD.t1057 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X68 a_13928_5005.t3 a_13338_5442.t7 VDD.t685 VDD.t684 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X69 a_12913_3240.t3 a_10168_1277.t4 a_13031_3240.t1 VDD.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X70 a_22852_110.t2 a_20582_5026.t4 VDD.t301 VDD.t300 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X71 Y[6].t6 a_26940_378.t4 a_26528_404.t4 VDD.t610 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X72 VDD.t249 a_19562_n2629.t7 a_19826_n3212.t2 VDD.t248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X73 a_13968_n7819.t0 a_13378_n8256.t7 VDD.t516 VDD.t515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X74 a_26520_n5464.t2 a_24740_n5464.t10 VDD.t1495 VDD.t1494 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X75 a_13177_2657.t0 a_12913_3240.t5 VDD.t348 VDD.t347 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X76 a_29230_2288.t3 a_28640_2725.t7 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X77 a_20582_5026.t0 a_19992_5463.t7 VDD.t293 VDD.t292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X78 VSS.t148 a_12029_n3217.t4 a_12907_n2630.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X79 a_29301_n2665.t0 a_28711_n2228.t7 VDD.t1422 VDD.t1421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X80 a_20582_5026.t1 a_19992_5463.t8 VSS.t34 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X81 a_11351_404.t2 a_11763_378.t4 a_11469_404.t5 VDD.t1394 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X82 a_31176_81.t1 a_29230_n745.t4 VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X83 a_30762_4198.t2 a_6818_316.t9 VDD.t639 VDD.t638 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X84 VDD.t637 a_6818_316.t10 a_32246_4888.t4 VDD.t636 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X85 a_29230_n745.t0 a_28640_n308.t7 VSS.t26 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X86 a_18412_n5491.t0 a_13177_2657.t5 VSS.t13 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X87 VDD.t15 a_13968_n7819.t5 a_18000_n5465.t3 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 VDD.t378 a_9512_n4182.t4 a_9567_n5760.t6 VDD.t377 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X89 a_30762_4198.t11 a_31174_4172.t4 Y[2].t7 VDD.t1187 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X90 a_7112_290.t2 a_2969_1600.t5 VDD.t1479 VDD.t1478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X91 a_6789_5443.t6 A[3].t0 VDD.t372 VDD.t371 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X92 VDD.t1323 a_16808_2859.t4 a_18543_3168.t5 VDD.t1322 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X93 a_23433_2927.t3 a_22843_3364.t7 VDD.t1359 VDD.t1358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X94 a_26528_404.t9 a_22797_1688.t4 VDD.t1347 VDD.t1346 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X95 a_4794_n5464.t8 a_704_n5517.t5 VDD.t370 VDD.t369 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X96 a_23439_n4591.t2 a_22849_n4154.t8 VDD.t1060 VDD.t1059 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X97 a_6273_1009.t3 a_4920_316.t9 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X98 a_18359_n396.t1 a_13367_404.t11 a_18123_336.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X99 VSS.t116 a_13968_n7819.t6 a_16450_n3142.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X100 a_20016_n6197.t1 a_20310_n5491.t4 VSS.t58 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X101 a_12035_2653.t0 a_11771_3236.t6 VSS.t119 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X102 a_19903_336.t5 a_20315_310.t4 a_20021_336.t4 VDD.t453 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X103 a_31176_n7762.t3 a_13361_n5466.t9 VDD.t552 VDD.t551 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X104 VDD.t518 a_13378_n8256.t8 a_13968_n7819.t1 VDD.t517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X105 a_7054_n416.t0 a_4920_316.t10 a_6818_316.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X106 VDD.t303 a_20582_5026.t5 a_24630_404.t3 VDD.t302 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X107 a_11765_n2634.t1 a_10157_n6197.t4 VSS.t36 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X108 VDD.t402 a_7414_n7824.t5 a_10918_n4773.t2 VDD.t401 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X109 a_3619_1189.t2 a_3029_1626.t8 VDD.t426 VDD.t425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X110 VDD.t1430 a_28711_n2228.t8 a_29301_n2665.t1 VDD.t1429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X111 a_22849_n4154.t2 a_22789_n4180.t5 VDD.t800 VDD.t799 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X112 VDD.t1424 a_28645_5296.t7 Y[0].t3 VDD.t1423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X113 VDD.t807 a_715_3106.t4 a_5214_290.t3 VDD.t806 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X114 a_11705_n328.t1 a_6620_n3211.t4 a_11469_404.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X115 a_13361_n5466.t2 a_12816_n4773.t4 a_13361_n6198.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X116 a_16167_n4181.t3 a_19567_3172.t5 VDD.t458 VDD.t457 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X117 VSS.t39 a_20617_n7831.t6 a_24195_n4771.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X118 a_18000_n5465.t2 a_13968_n7819.t7 VDD.t917 VDD.t916 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X119 a_6810_n5464.t5 a_6265_n4771.t4 a_6810_n6196.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X120 VDD.t1110 a_707_521.t5 a_4375_1009.t3 VDD.t1109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X121 VDD.t323 a_12907_n2630.t5 a_9518_1688.t3 VDD.t322 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X122 a_3015_3276.t3 a_715_3106.t5 VDD.t809 VDD.t808 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X123 VDD.t1537 a_688_n2757.t4 a_4794_n5464.t5 VDD.t1536 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X124 a_6818_316.t4 a_6273_1009.t4 a_6700_316.t3 VDD.t240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X125 a_19476_1029.t3 a_18123_336.t9 VDD.t954 VDD.t953 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X126 a_6474_n2628.t2 a_3611_n4591.t4 a_6356_n2628.t3 VDD.t1107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X127 a_5332_n2632.t2 a_3606_n6195.t4 a_5214_n2632.t1 VDD.t437 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X128 a_24622_n5464.t2 a_25034_n5490.t4 a_24740_n5464.t0 VDD.t589 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X129 a_11771_3236.t1 a_10163_n327.t4 a_11889_3236.t2 VDD.t704 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X130 VDD.t554 a_13361_n5466.t10 a_31176_n7762.t2 VDD.t553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X131 a_13968_n7819.t2 a_13378_n8256.t9 VDD.t520 VDD.t519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X132 a_28708_n5298.t2 A[1].t1 VDD.t857 VDD.t856 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X133 a_26932_n5490.t3 a_22789_n4180.t6 VDD.t802 VDD.t801 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X134 VDD.t811 a_715_3106.t6 a_3015_3276.t2 VDD.t810 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X135 VSS.t66 a_10148_n2943.t4 a_11765_n2634.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X136 a_29301_n2665.t2 a_28711_n2228.t9 VDD.t1432 VDD.t1431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X137 a_13597_n6198.t0 a_11463_n5466.t9 a_13361_n5466.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X138 a_11889_3236.t1 a_10163_n327.t5 a_11771_3236.t2 VDD.t995 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X139 a_7046_n6196.t1 a_4912_n5464.t8 a_6810_n5464.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X140 a_13338_5442.t0 A[2].t0 VDD.t214 VDD.t213 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X141 VDD.t1481 a_2969_1600.t6 a_6700_316.t11 VDD.t1480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X142 a_19680_n2629.t5 a_16817_n4592.t4 a_19562_n2629.t3 VDD.t1070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X143 VDD.t1314 a_2961_n4180.t6 a_3016_n5758.t6 VDD.t1313 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X144 a_4794_n5464.t6 a_688_n2757.t5 VDD.t1539 VDD.t1538 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X145 a_5222_3148.t1 a_3614_n415.t4 VSS.t24 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X146 a_6356_n2628.t0 a_3611_n4591.t5 a_6474_n2628.t1 VDD.t1108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X147 a_19898_n5465.t4 a_18118_n5465.t8 VDD.t1525 VDD.t1524 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X148 a_5214_n2632.t3 a_3606_n6195.t5 a_5332_n2632.t1 VDD.t438 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X149 a_24740_n5464.t1 a_25034_n5490.t5 a_24622_n5464.t1 VDD.t590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X150 a_31174_4172.t3 a_29230_2288.t4 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X151 a_30764_107.t3 a_31176_81.t5 Y[1].t4 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X152 a_31176_n7762.t1 a_13361_n5466.t11 VDD.t717 VDD.t716 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X153 VDD.t222 A[1].t2 a_28708_n5298.t1 VDD.t221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X154 VDD.t804 a_22789_n4180.t7 a_26932_n5490.t2 VDD.t803 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X155 a_30335_4891.t3 a_6818_316.t11 VDD.t635 VDD.t634 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X156 VDD.t663 a_18684_n3216.t4 a_19680_n2629.t1 VDD.t662 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X157 a_30764_n3388.t11 a_29298_n5735.t4 VDD.t691 VDD.t690 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X158 Y[3].t5 a_30337_n7043.t5 a_30764_n7736.t11 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X159 VSS.t45 a_9512_n4182.t5 a_13597_n6198.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X160 a_4802_316.t2 a_707_521.t6 VDD.t1112 VDD.t1111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X161 a_9558_n2506.t3 a_6810_n5464.t8 VDD.t1434 VDD.t1433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X162 a_16808_2859.t3 a_16218_3296.t7 VDD.t1080 VDD.t1079 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X163 a_3024_22.t2 a_715_3106.t7 VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X164 a_32485_160.t1 a_29230_n745.t5 a_32248_797.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X165 VDD.t27 a_11765_n2634.t5 a_12029_n3217.t0 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X166 a_23425_n2941.t0 a_22835_n2504.t7 VDD.t1286 VDD.t1285 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X167 VDD.t1436 a_6810_n5464.t9 a_11345_n5466.t2 VDD.t1435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X168 a_13025_n2630.t5 a_10162_n4593.t5 a_12907_n2630.t3 VDD.t309 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X169 a_6474_n2628.t0 a_3611_n4591.t6 a_6356_n2628.t1 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X170 a_24622_n5464.t0 a_25034_n5490.t6 a_24740_n5464.t5 VDD.t786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X171 VDD.t1527 a_18118_n5465.t9 a_19898_n5465.t3 VDD.t1526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X172 Y[7].t3 a_26192_3240.t5 VDD.t879 VDD.t878 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X173 a_3029_1626.t6 a_2969_1600.t7 VDD.t1483 VDD.t1482 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X174 a_28708_n5298.t0 A[1].t3 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X175 a_20582_5026.t2 a_19992_5463.t9 VDD.t835 VDD.t834 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X176 VDD.t1451 a_12035_2653.t4 a_13031_3240.t5 VDD.t1450 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X177 a_24748_404.t2 a_24203_1097.t4 a_24630_404.t8 VDD.t680 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X178 VDD.t380 a_9512_n4182.t6 a_13243_n5466.t11 VDD.t379 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X179 a_4794_n5464.t7 a_704_n5517.t6 VDD.t352 VDD.t351 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X180 a_16227_n4155.t6 a_16167_n4181.t4 VDD.t1170 VDD.t1169 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X181 a_4802_316.t8 a_5214_290.t4 a_4920_316.t7 VDD.t1533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X182 a_23094_1077.t0 a_22797_1688.t5 a_22857_1714.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X183 VDD.t693 a_29298_n5735.t5 a_30764_n3388.t10 VDD.t692 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X184 a_29230_2288.t2 a_28640_2725.t8 VDD.t905 VDD.t904 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X185 VDD.t354 a_704_n5517.t7 a_3021_n4154.t6 VDD.t353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X186 VDD.t374 A[3].t1 a_13378_n8256.t0 VDD.t373 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X187 VDD.t1485 a_2969_1600.t8 a_3029_1626.t5 VDD.t1484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X188 a_13249_404.t3 a_12822_1097.t6 a_13367_404.t3 VDD.t1609 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X189 a_30764_n7736.t10 a_30337_n7043.t6 Y[3].t4 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X190 a_23086_n4791.t0 a_22789_n4180.t8 a_22849_n4154.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X191 a_13361_n6198.t1 a_13655_n5492.t4 VSS.t112 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X192 a_7379_5006.t2 a_6789_5443.t7 VDD.t1034 VDD.t1033 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X193 VDD.t1134 a_20021_336.t8 a_32248_n2698.t5 VDD.t1133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X194 a_31118_n8468.t0 a_29305_n8580.t5 Y[3].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X195 VDD.t83 a_13177_2657.t6 a_18412_n5491.t3 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X196 VDD.t446 a_25050_3236.t5 a_25314_2653.t3 VDD.t445 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X197 a_12029_n3217.t1 a_11765_n2634.t6 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X198 a_7379_5006.t3 a_6789_5443.t8 VSS.t128 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X199 a_29298_n5735.t0 a_28708_n5298.t7 VSS.t75 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X200 a_11351_404.t4 a_6620_n3211.t5 VDD.t669 VDD.t668 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X201 VSS.t170 a_22797_1688.t6 a_26882_n328.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X202 VSS.t32 a_29230_n745.t6 a_31118_n625.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X203 a_10154_2927.t3 a_9564_3364.t7 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X204 a_20617_n7831.t2 a_20027_n8268.t7 VSS.t200 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X205 VDD.t118 a_29230_2288.t5 a_30762_4198.t5 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X206 a_9512_n4182.t3 a_32246_4888.t8 VDD.t619 VDD.t618 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X207 a_9815_1077.t0 a_9518_1688.t4 a_9578_1714.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X208 a_18123_n396.t0 a_18417_310.t4 VSS.t143 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X209 a_22835_n2504.t6 a_20016_n5465.t10 VDD.t1243 VDD.t1242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X210 a_5206_n5490.t0 a_688_n2757.t6 VSS.t57 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X211 VDD.t919 a_13968_n7819.t8 a_16227_n4155.t2 VDD.t918 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X212 a_125_3543.t3 A[1].t4 VDD.t226 VDD.t225 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X213 a_23081_n6395.t0 a_20016_n5465.t11 a_22844_n5758.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X214 VDD.t1284 a_7379_5006.t5 a_9564_3364.t3 VDD.t1283 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X215 VDD.t186 a_16172_1620.t5 a_16232_1646.t0 VDD.t185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X216 VDD.t305 a_20582_5026.t6 a_24630_404.t4 VDD.t304 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X217 a_3021_n4154.t5 a_704_n5517.t8 VDD.t356 VDD.t355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X218 a_6482_3152.t3 a_3619_1189.t4 a_6364_3152.t4 VDD.t1504 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X219 VDD.t1114 a_707_521.t7 a_4375_1009.t2 VDD.t1113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X220 a_28640_n308.t2 A[1].t5 VDD.t228 VDD.t227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X221 VSS.t40 a_20617_n7831.t7 a_23086_n4791.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X222 a_16817_n4592.t0 a_16227_n4155.t7 VSS.t68 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X223 a_32248_n2698.t6 a_20021_336.t9 VDD.t1203 VDD.t1202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X224 VSS.t94 a_13361_n5466.t12 a_31118_n8468.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X225 a_3606_n6195.t3 a_3016_n5758.t7 VSS.t43 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X226 VDD.t775 A[1].t6 a_125_3543.t2 VDD.t774 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X227 VSS.t144 a_11469_404.t9 a_12822_1097.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X228 VDD.t176 a_29301_n2665.t6 a_30764_107.t1 VDD.t175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X229 VSS.t101 a_707_521.t8 a_3252_2639.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X230 a_18417_310.t3 a_13928_5005.t4 VDD.t342 VDD.t341 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X231 a_30337_n7043.t0 a_29305_n8580.t6 VDD.t767 VDD.t766 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X232 VDD.t96 a_24740_n5464.t11 a_26093_n4771.t3 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X233 a_18000_n5465.t9 a_18412_n5491.t4 a_18118_n5465.t7 VDD.t963 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X234 a_6364_3152.t2 a_3619_1189.t5 VSS.t190 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X235 a_16822_1209.t2 a_16232_1646.t9 VDD.t218 VDD.t217 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X236 a_3614_n415.t0 a_3024_22.t8 VSS.t23 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X237 VDD.t168 a_28640_n308.t8 a_29230_n745.t3 VDD.t167 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X238 a_13575_4805.t0 A[2].t1 a_13338_5442.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X239 VDD.t344 a_13928_5005.t5 a_18417_310.t2 VDD.t343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X240 a_24740_n5464.t6 a_24195_n4771.t4 a_24622_n5464.t8 VDD.t1065 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X241 VDD.t404 a_7414_n7824.t6 a_9572_n4156.t2 VDD.t403 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X242 a_16812_n6196.t0 a_16222_n5759.t7 VSS.t22 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X243 a_351_n5717.t0 B[0].t0 a_114_n5080.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X244 a_11469_404.t6 a_11763_378.t5 a_11351_404.t1 VDD.t1395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X245 VDD.t921 a_13367_404.t12 a_17578_1029.t3 VDD.t920 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X246 VDD.t739 a_704_n5517.t9 a_3021_n4154.t4 VDD.t738 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X247 a_11463_n5466.t2 a_10918_n4773.t4 a_11463_n6198.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X248 a_16218_3296.t1 a_13928_5005.t6 VDD.t346 VDD.t345 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X249 VDD.t1132 a_117_958.t7 a_707_521.t0 VDD.t1131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X250 VDD.t239 a_9518_1688.t5 a_9573_110.t0 VDD.t238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X251 a_23425_n2941.t1 a_22835_n2504.t8 VSS.t163 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X252 a_4912_n5464.t1 a_4367_n4771.t4 a_4912_n6196.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X253 VDD.t1173 a_5222_3148.t5 a_5486_2565.t3 VDD.t1172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X254 a_30880_3466.t1 a_31174_4172.t5 VSS.t96 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X255 a_23433_2927.t0 a_22843_3364.t8 VSS.t172 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X256 VDD.t881 a_29298_n5735.t6 a_32248_n2698.t3 VDD.t880 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X257 a_30882_n8468.t0 a_31176_n7762.t4 VSS.t150 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X258 VDD.t178 a_29301_n2665.t7 a_32248_797.t1 VDD.t177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X259 a_30764_107.t4 a_31176_81.t6 Y[1].t3 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X260 a_11889_3236.t3 a_10154_2927.t4 VDD.t682 VDD.t681 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X261 a_13338_5442.t2 A[2].t2 VDD.t273 VDD.t272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X262 VDD.t1191 a_11469_404.t10 a_12822_1097.t2 VDD.t1190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X263 VDD.t769 a_29305_n8580.t7 a_30337_n7043.t1 VDD.t768 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X264 VDD.t827 a_2969_1600.t9 a_6700_316.t10 VDD.t826 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X265 a_28711_n2228.t3 B[1].t1 VDD.t903 VDD.t902 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X266 VDD.t701 a_6810_n5464.t10 a_11345_n5466.t1 VDD.t700 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X267 a_11883_n2634.t2 a_10157_n6197.t5 a_11765_n2634.t0 VDD.t308 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X268 a_10168_1277.t3 a_9578_1714.t7 VDD.t1150 VDD.t1149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X269 a_4802_316.t5 a_715_3106.t8 VDD.t794 VDD.t793 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X270 a_10162_n4593.t0 a_9572_n4156.t7 VDD.t255 VDD.t254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X271 VSS.t72 a_19826_n3212.t6 a_23080_2727.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X272 VDD.t431 a_9518_1688.t6 a_9578_1714.t3 VDD.t430 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X273 a_32248_n2698.t4 a_29298_n5735.t7 VDD.t883 VDD.t882 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X274 a_20027_n8268.t2 A[2].t3 VDD.t275 VDD.t274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X275 VDD.t376 A[3].t2 a_19992_5463.t0 VDD.t375 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X276 a_10924_1097.t3 a_6620_n3211.t6 VDD.t659 VDD.t658 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X277 a_24748_404.t1 a_24203_1097.t5 a_24630_404.t0 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X278 a_5222_3148.t3 a_3614_n415.t5 a_5340_3148.t5 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X279 VDD.t923 a_13367_404.t13 a_18005_336.t8 VDD.t922 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X280 VDD.t382 a_18118_n5465.t10 a_19471_n4772.t3 VDD.t381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X281 a_32246_4888.t5 a_29230_2288.t6 VDD.t1088 VDD.t1087 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X282 VDD.t33 a_13968_n7819.t9 a_16213_n2505.t0 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X283 a_20027_n8268.t4 B[3].t0 VDD.t975 VDD.t974 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X284 a_11345_n5466.t0 a_6810_n5464.t11 VDD.t703 VDD.t702 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X285 a_9578_1714.t6 a_6620_n3211.t7 VDD.t661 VDD.t660 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X286 a_11765_n2634.t3 a_10157_n6197.t6 a_11883_n2634.t1 VDD.t724 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X287 a_5206_n5490.t3 a_688_n2757.t7 VDD.t450 VDD.t449 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X288 VDD.t568 a_19826_n3212.t7 a_22843_3364.t6 VDD.t567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X289 VSS.t76 a_16167_n4181.t5 a_16459_n6396.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X290 a_20016_n5465.t2 a_20310_n5491.t5 a_19898_n5465.t11 VDD.t451 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X291 VDD.t433 a_9518_1688.t7 a_13249_404.t4 VDD.t432 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X292 a_18005_336.t5 a_13928_5005.t7 VDD.t1040 VDD.t1039 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X293 VDD.t184 a_24748_404.t8 a_26528_404.t0 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X294 VDD.t289 a_29230_n745.t7 a_31176_81.t0 VDD.t288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X295 a_3007_n2504.t6 a_704_n5517.t10 VDD.t741 VDD.t740 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X296 VDD.t1471 B[0].t1 a_28645_5296.t6 VDD.t1470 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X297 a_30764_n3388.t1 a_31176_n3414.t4 Y[4].t6 VDD.t1218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X298 a_7414_n7824.t0 a_6824_n8261.t7 VSS.t174 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X299 VSS.t82 a_6620_n3211.t8 a_9801_2727.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X300 a_3619_1189.t0 a_3029_1626.t9 VSS.t53 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X301 a_9810_n527.t1 a_7379_5006.t6 a_9573_110.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X302 a_18420_n2633.t3 a_16812_n6196.t4 VSS.t131 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X303 VDD.t719 a_13361_n5466.t13 a_30764_n7736.t8 VDD.t718 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X304 VDD.t1592 A[2].t4 a_20027_n8268.t1 VDD.t1591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X305 VDD.t788 a_707_521.t9 a_3029_1626.t2 VDD.t787 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X306 a_20016_n5465.t6 a_19471_n4772.t4 a_19898_n5465.t8 VDD.t1223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X307 a_19471_n4772.t2 a_18118_n5465.t11 VDD.t384 VDD.t383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X308 a_10154_2927.t2 a_9564_3364.t8 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X309 a_23433_2927.t2 a_22843_3364.t9 VDD.t1351 VDD.t1350 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X310 VSS.t92 B[2].t2 a_28877_2088.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X311 VDD.t362 A[3].t3 a_114_n5080.t6 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X312 a_20021_336.t3 a_20315_310.t5 a_19903_336.t6 VDD.t454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X313 a_13243_n5466.t4 a_12816_n4773.t5 a_13361_n5466.t3 VDD.t1419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X314 a_18412_n5491.t2 a_13177_2657.t7 VDD.t277 VDD.t276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X315 VDD.t1090 a_29230_2288.t7 a_30762_4198.t4 VDD.t1089 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X316 a_25314_2653.t0 a_25050_3236.t6 VSS.t56 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X317 a_24748_404.t3 a_24203_1097.t6 a_24748_n328.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X318 a_6692_n5464.t11 a_6265_n4771.t5 a_6810_n5464.t4 VDD.t1519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X319 VDD.t1625 a_6810_n5464.t12 a_11757_n5492.t3 VDD.t1624 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X320 VDD.t43 a_4912_n5464.t9 a_6265_n4771.t0 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X321 a_31176_n3414.t0 a_20021_336.t10 VSS.t152 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X322 a_11351_404.t3 a_6620_n3211.t9 VDD.t609 VDD.t608 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X323 a_16213_n2505.t1 a_13968_n7819.t10 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X324 VSS.t113 B[1].t2 a_362_2906.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X325 VDD.t540 a_6620_n3211.t10 a_9564_3364.t6 VDD.t539 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X326 VDD.t813 a_688_n2757.t8 a_5206_n5490.t2 VDD.t812 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X327 a_20310_n5491.t0 a_16167_n4181.t6 VSS.t77 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X328 a_19898_n5465.t10 a_20310_n5491.t6 a_20016_n5465.t3 VDD.t957 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X329 a_6482_3152.t2 a_3619_1189.t6 a_6364_3152.t3 VDD.t1505 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X330 VDD.t743 a_704_n5517.t11 a_3007_n2504.t5 VDD.t742 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X331 VSS.t27 a_24748_404.t9 a_26101_1097.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X332 a_20617_n7831.t0 a_20027_n8268.t8 VDD.t235 VDD.t234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X333 a_6700_316.t4 a_6273_1009.t5 a_6818_316.t5 VDD.t241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X334 VDD.t621 a_18118_n5465.t12 a_19471_n4772.t1 VDD.t620 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X335 a_2961_n4180.t1 a_6364_3152.t5 VSS.t192 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X336 a_7414_n7824.t1 a_6824_n8261.t8 VDD.t1361 VDD.t1360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X337 a_114_n5080.t5 A[3].t4 VDD.t364 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X338 VSS.t103 a_715_3106.t9 a_5156_n416.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X339 a_98_n2320.t2 A[2].t5 VDD.t1594 VDD.t1593 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X340 a_13361_n5466.t5 a_12816_n4773.t6 a_13243_n5466.t3 VDD.t1420 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X341 a_6356_n2628.t2 a_3611_n4591.t7 VSS.t15 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X342 a_6810_n5464.t3 a_6265_n4771.t6 a_6692_n5464.t9 VDD.t1155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X343 a_11757_n5492.t2 a_6810_n5464.t13 VDD.t1627 VDD.t1626 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X344 a_25050_3236.t2 a_23442_n327.t4 a_25168_3236.t2 VDD.t1378 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X345 VDD.t37 a_13968_n7819.t11 a_16213_n2505.t2 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X346 a_10148_n2943.t2 a_9558_n2506.t7 VDD.t1168 VDD.t1167 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X347 a_5206_n5490.t1 a_688_n2757.t9 VDD.t815 VDD.t814 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X348 VDD.t790 a_707_521.t10 a_3015_3276.t5 VDD.t789 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X349 Y[4].t3 a_30337_n2695.t4 a_30882_n4120.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X350 a_19685_3172.t4 a_16822_1209.t4 a_19567_3172.t4 VDD.t1246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X351 a_3597_n2941.t3 a_3007_n2504.t7 VDD.t243 VDD.t242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X352 VSS.t7 a_3605_2839.t4 a_5222_3148.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X353 VSS.t63 a_11463_n5466.t10 a_12816_n4773.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X354 a_25168_3236.t5 a_23433_2927.t4 VDD.t1355 VDD.t1354 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X355 a_18005_336.t2 a_18417_310.t5 a_18123_336.t4 VDD.t1102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X356 VDD.t237 a_20027_n8268.t9 a_20617_n7831.t1 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X357 a_16167_n4181.t0 a_19567_3172.t6 VSS.t60 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X358 VDD.t1158 a_24748_404.t10 a_26101_1097.t3 VDD.t1157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X359 a_18417_310.t0 a_13928_5005.t8 VSS.t129 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X360 a_19562_n2629.t4 a_16817_n4592.t5 VSS.t132 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X361 VDD.t366 A[3].t5 a_114_n5080.t4 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X362 VSS.t106 B[3].t1 a_20229_4826.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X363 VDD.t76 a_32248_n7046.t8 a_16172_1620.t2 VDD.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X364 a_13243_n5466.t8 a_13655_n5492.t5 a_13361_n5466.t7 VDD.t886 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X365 a_7112_290.t0 a_2969_1600.t10 VSS.t108 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X366 VSS.t156 a_5478_n3215.t4 a_6356_n2628.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X367 a_16803_n2942.t2 a_16213_n2505.t8 VDD.t737 VDD.t736 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X368 VDD.t1582 a_29298_n5735.t8 a_30337_n2695.t3 VDD.t1581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X369 VDD.t1222 a_26184_n2628.t5 a_22797_1688.t3 VDD.t1221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X370 a_23434_n6195.t2 a_22844_n5758.t8 VDD.t469 VDD.t468 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X371 VDD.t544 a_9558_n2506.t8 a_10148_n2943.t0 VDD.t543 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X372 a_11763_378.t0 a_7379_5006.t7 VSS.t162 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X373 a_6824_n8261.t3 B[2].t3 VDD.t707 VDD.t706 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X374 VSS.t167 a_16808_2859.t5 a_18425_3168.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X375 VDD.t412 a_18425_3168.t5 a_18689_2585.t3 VDD.t411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X376 a_28640_2725.t2 A[0].t1 VDD.t1416 VDD.t1415 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X377 VDD.t753 a_3007_n2504.t8 a_3597_n2941.t2 VDD.t752 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X378 a_28948_n2865.t0 B[1].t3 a_28711_n2228.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X379 VDD.t821 B[3].t2 a_19992_5463.t3 VDD.t820 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X380 a_30762_4198.t9 a_30335_4891.t4 Y[2].t3 VDD.t1159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X381 a_6789_5443.t3 B[1].t4 VDD.t781 VDD.t780 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X382 a_13031_3240.t0 a_10168_1277.t5 a_12913_3240.t2 VDD.t605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X383 a_704_n5517.t1 a_114_n5080.t7 VDD.t986 VDD.t985 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X384 Y[2].t4 a_30335_4891.t5 a_30762_4198.t10 VDD.t1160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X385 VDD.t188 a_16172_1620.t6 a_20315_310.t3 VDD.t187 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X386 a_9518_1688.t0 a_12907_n2630.t6 VSS.t38 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X387 a_16172_1620.t1 a_32248_n7046.t9 VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X388 a_13361_n5466.t0 a_13655_n5492.t6 a_13243_n5466.t0 VDD.t470 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X389 VDD.t1562 a_704_n5517.t12 a_4367_n4771.t3 VDD.t1561 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X390 VDD.t296 a_3605_2839.t5 a_5340_3148.t2 VDD.t295 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X391 a_12913_3240.t0 a_10168_1277.t6 VSS.t80 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X392 a_4920_316.t5 a_5214_290.t5 a_4802_316.t7 VDD.t1528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X393 a_24630_404.t1 a_24203_1097.t7 a_24748_404.t0 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X394 a_688_n2757.t2 a_98_n2320.t7 VSS.t175 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X395 a_6620_n3211.t3 a_6356_n2628.t5 VSS.t214 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X396 Y[3].t7 a_30337_n7043.t7 a_30764_n7736.t9 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X397 VDD.t504 a_25314_2653.t4 a_26310_3240.t5 VDD.t503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X398 VDD.t1343 a_22797_1688.t7 a_26528_404.t8 VDD.t1342 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X399 a_32246_4888.t6 a_29230_2288.t8 VDD.t1092 VDD.t1091 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X400 a_10148_n2943.t1 a_9558_n2506.t9 VDD.t546 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X401 Y[5].t4 a_26093_n4771.t4 a_26638_n6196.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X402 VDD.t1418 A[0].t2 a_28645_5296.t2 VDD.t1417 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X403 a_20315_310.t2 a_16172_1620.t7 VDD.t190 VDD.t189 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X404 a_20310_n5491.t3 a_16167_n4181.t7 VDD.t945 VDD.t944 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X405 VSS.t208 a_6818_316.t12 a_32483_4251.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X406 a_13367_404.t2 a_12822_1097.t7 a_13249_404.t2 VDD.t1610 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X407 a_3597_n2941.t1 a_3007_n2504.t9 VDD.t456 VDD.t455 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X408 VDD.t1 a_707_521.t11 a_3029_1626.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X409 a_20021_336.t0 a_19476_1029.t4 a_19903_336.t0 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X410 a_32248_n7046.t6 a_13361_n5466.t14 VDD.t721 VDD.t720 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X411 a_22844_n5758.t2 a_20016_n5465.t12 VDD.t1258 VDD.t1257 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X412 VDD.t1260 a_20016_n5465.t13 a_24622_n5464.t5 VDD.t1259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X413 a_19992_5463.t6 A[3].t6 VDD.t1457 VDD.t1456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X414 a_26302_n2628.t3 a_23439_n4591.t4 a_26184_n2628.t4 VDD.t884 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X415 a_28645_5296.t1 A[0].t3 VDD.t1406 VDD.t1405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X416 VDD.t931 a_11771_3236.t7 a_12035_2653.t2 VDD.t930 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X417 a_98_n2320.t6 B[1].t5 VDD.t783 VDD.t782 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X418 VDD.t462 a_13968_n7819.t12 a_17573_n4772.t3 VDD.t461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X419 a_11463_n5466.t1 a_10918_n4773.t5 a_11345_n5466.t5 VDD.t748 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X420 VSS.t140 a_9518_1688.t8 a_13603_n328.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X421 a_4912_n5464.t2 a_4367_n4771.t5 a_4794_n5464.t1 VDD.t705 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X422 VDD.t1516 a_114_n5080.t8 a_704_n5517.t2 VDD.t1515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X423 a_16232_1646.t1 a_16172_1620.t8 VDD.t1531 VDD.t1530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X424 a_11351_404.t7 a_7379_5006.t8 VDD.t1274 VDD.t1273 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X425 a_24630_404.t6 a_19826_n3212.t8 VDD.t570 VDD.t569 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X426 VSS.t155 a_3597_n2941.t4 a_5214_n2632.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X427 VDD.t960 a_22789_n4180.t9 a_26520_n5464.t7 VDD.t959 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X428 a_13243_n5466.t1 a_13655_n5492.t7 a_13361_n5466.t1 VDD.t471 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X429 a_4367_n4771.t2 a_704_n5517.t13 VDD.t1564 VDD.t1563 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X430 a_30764_n7736.t5 a_31176_n7762.t5 Y[3].t1 VDD.t948 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X431 VDD.t829 a_2969_1600.t11 a_3024_22.t6 VDD.t828 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X432 VDD.t1408 A[0].t4 a_28715_n8143.t6 VDD.t1407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X433 a_28952_n8780.t0 B[3].t3 a_28715_n8143.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X434 VDD.t1276 a_7379_5006.t9 a_11351_404.t6 VDD.t1275 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X435 a_22852_110.t1 a_20582_5026.t7 VDD.t479 VDD.t478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X436 VDD.t925 a_13367_404.t14 a_16232_1646.t4 VDD.t924 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X437 a_30764_107.t0 a_29301_n2665.t8 VDD.t1473 VDD.t1472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X438 a_26184_n2628.t3 a_23439_n4591.t5 a_26302_n2628.t4 VDD.t1073 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X439 VDD.t785 B[1].t6 a_125_3543.t5 VDD.t784 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X440 a_23442_n327.t3 a_22852_110.t7 VDD.t317 VDD.t316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X441 a_18118_n5465.t2 a_17573_n4772.t4 a_18118_n6197.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X442 a_11345_n5466.t4 a_10918_n4773.t6 a_11463_n5466.t0 VDD.t749 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X443 VDD.t406 a_7414_n7824.t7 a_10918_n4773.t1 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X444 a_4794_n5464.t2 a_4367_n4771.t6 a_4912_n5464.t3 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X445 a_19903_336.t8 a_18123_336.t10 VDD.t956 VDD.t955 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X446 VDD.t1076 B[0].t2 a_28640_n308.t4 VDD.t1075 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X447 a_5148_n6196.t1 a_704_n5517.t14 a_4912_n5464.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X448 VDD.t1084 a_704_n5517.t15 a_4367_n4771.t1 VDD.t1083 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X449 VDD.t998 a_5486_2565.t4 a_6482_3152.t4 VDD.t997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X450 Y[3].t2 a_31176_n7762.t6 a_30764_n7736.t4 VDD.t949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X451 a_22849_n4154.t1 a_22789_n4180.t10 VDD.t962 VDD.t961 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X452 a_16227_42.t1 a_13928_5005.t9 VDD.t1042 VDD.t1041 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X453 a_28715_n8143.t5 A[0].t5 VDD.t1410 VDD.t1409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X454 a_26940_378.t3 a_22797_1688.t8 VDD.t1345 VDD.t1344 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X455 a_31176_81.t2 a_29230_n745.t8 VSS.t178 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X456 VSS.t166 a_2961_n4180.t7 a_7046_n6196.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X457 a_11351_404.t0 a_11763_378.t6 a_11469_404.t7 VDD.t1396 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X458 a_707_521.t2 a_117_958.t8 VDD.t1546 VDD.t1545 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X459 a_9795_n3143.t0 a_6810_n5464.t14 a_9558_n2506.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X460 VDD.t279 a_13177_2657.t8 a_18000_n5465.t7 VDD.t278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X461 Y[1].t7 a_30337_800.t4 a_30764_107.t11 VDD.t1617 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X462 a_18538_n2633.t2 a_16812_n6196.t5 a_18420_n2633.t2 VDD.t1048 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X463 a_10154_2927.t0 a_9564_3364.t9 VSS.t9 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X464 a_32248_797.t6 a_29230_n745.t9 VDD.t1389 VDD.t1388 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X465 a_16469_1009.t0 a_16172_1620.t9 a_16232_1646.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X466 a_18354_n6197.t0 a_13968_n7819.t13 a_18118_n5465.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X467 a_24622_n5464.t11 a_20617_n7831.t8 VDD.t340 VDD.t339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X468 a_707_521.t3 a_117_958.t9 VDD.t1548 VDD.t1547 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X469 VDD.t481 a_20582_5026.t8 a_25042_378.t3 VDD.t480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X470 VDD.t1082 a_16218_3296.t8 a_16808_2859.t2 VDD.t1081 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X471 a_25042_378.t0 a_20582_5026.t9 VSS.t62 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X472 a_12029_n3217.t2 a_11765_n2634.t7 VSS.t130 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X473 VDD.t1412 A[0].t6 a_28715_n8143.t4 VDD.t1411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X474 VDD.t327 a_20617_n7831.t9 a_22849_n4154.t6 VDD.t326 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X475 a_16817_n395.t2 a_16227_42.t8 VDD.t194 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X476 a_23447_1277.t2 a_22857_1714.t8 VDD.t1064 VDD.t1063 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X477 a_6810_n6196.t1 a_7104_n5490.t4 VSS.t199 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X478 VDD.t23 a_13338_5442.t8 a_13928_5005.t2 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X479 a_9573_110.t6 a_9518_1688.t9 VDD.t1095 VDD.t1094 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X480 VSS.t48 a_7414_n7824.t8 a_9795_n3143.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X481 a_23439_n4591.t0 a_22849_n4154.t9 VSS.t52 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X482 VDD.t947 a_16167_n4181.t8 a_16222_n5759.t6 VDD.t946 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X483 a_18000_n5465.t6 a_13177_2657.t9 VDD.t281 VDD.t280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X484 a_18420_n2633.t1 a_16812_n6196.t6 a_18538_n2633.t1 VDD.t496 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X485 a_19562_n2629.t1 a_16817_n4592.t6 a_19680_n2629.t4 VDD.t1067 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X486 a_4920_316.t1 a_4375_1009.t4 a_4802_316.t11 VDD.t597 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X487 a_11883_n2634.t0 a_10157_n6197.t7 a_11765_n2634.t2 VDD.t725 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X488 VDD.t1186 B[3].t4 a_28708_n5298.t5 VDD.t1185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X489 a_3016_n5758.t5 a_2961_n4180.t8 VDD.t1306 VDD.t1305 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X490 VDD.t1116 a_688_n2757.t10 a_4794_n5464.t4 VDD.t1115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X491 VDD.t1184 B[3].t5 a_19992_5463.t4 VDD.t1183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X492 a_22843_3364.t2 a_20582_5026.t10 VDD.t849 VDD.t848 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X493 a_25034_n5490.t0 a_20016_n5465.t14 VSS.t159 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X494 VDD.t329 a_20617_n7831.t10 a_24622_n5464.t10 VDD.t328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X495 a_30764_n3388.t9 a_29298_n5735.t9 VDD.t1584 VDD.t1583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X496 a_32246_4888.t3 a_6818_316.t13 VDD.t633 VDD.t632 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X497 a_29305_n8580.t2 a_28715_n8143.t7 VDD.t584 VDD.t583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X498 a_22849_n4154.t5 a_20617_n7831.t11 VDD.t331 VDD.t330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X499 VDD.t1353 a_22843_3364.t10 a_23433_2927.t1 VDD.t1352 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X500 a_31176_81.t3 a_29230_n745.t10 VDD.t1391 VDD.t1390 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X501 a_23434_n6195.t0 a_22844_n5758.t9 VSS.t201 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X502 a_18543_3168.t1 a_16817_n395.t5 a_18425_3168.t2 VDD.t1612 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X503 VDD.t1193 a_11469_404.t11 a_13249_404.t11 VDD.t1192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X504 a_20315_310.t0 a_16172_1620.t10 VSS.t195 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X505 a_16222_n5759.t4 a_16167_n4181.t9 VDD.t859 VDD.t858 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X506 VSS.t89 a_10154_2927.t5 a_11771_3236.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X507 a_19680_n2629.t3 a_16817_n4592.t7 a_19562_n2629.t2 VDD.t1068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X508 a_2969_1600.t1 a_32248_797.t7 VDD.t1371 VDD.t1370 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X509 a_9572_n4156.t6 a_9512_n4182.t7 VDD.t971 VDD.t970 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X510 a_6818_316.t6 a_6273_1009.t6 a_6818_n416.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X511 a_16817_n395.t0 a_16227_42.t9 VSS.t29 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X512 VDD.t508 a_10148_n2943.t5 a_11883_n2634.t5 VDD.t507 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X513 VDD.t1138 a_12029_n3217.t5 a_13025_n2630.t2 VDD.t1137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X514 a_28708_n5298.t4 B[3].t6 VDD.t613 VDD.t612 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X515 VDD.t1308 a_2961_n4180.t9 a_3016_n5758.t4 VDD.t1307 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X516 a_19903_336.t4 a_20315_310.t6 a_20021_336.t2 VDD.t452 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X517 VDD.t1266 a_5478_n3215.t5 a_6474_n2628.t5 VDD.t1265 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X518 VDD.t1262 a_20016_n5465.t15 a_22844_n5758.t1 VDD.t1261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X519 a_24622_n5464.t9 a_20617_n7831.t12 VDD.t333 VDD.t332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X520 a_19898_n5465.t2 a_18118_n5465.t13 VDD.t623 VDD.t622 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X521 a_5214_290.t2 a_715_3106.t10 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X522 a_11469_404.t0 a_10924_1097.t4 a_11469_n328.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X523 VDD.t1205 a_20021_336.t11 a_30764_n3388.t7 VDD.t1204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X524 VDD.t512 a_19567_3172.t7 a_16167_n4181.t2 VDD.t511 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X525 VDD.t891 a_28715_n8143.t8 a_29305_n8580.t3 VDD.t890 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X526 a_20016_n5465.t5 a_19471_n4772.t5 a_20016_n6197.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X527 VDD.t220 a_16232_1646.t10 a_16822_1209.t1 VDD.t219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X528 VDD.t871 a_18123_336.t11 a_19476_1029.t2 VDD.t870 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X529 a_11469_n328.t0 a_11763_378.t7 VSS.t33 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X530 VDD.t1047 a_11765_n2634.t8 a_12029_n3217.t3 VDD.t1046 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X531 VDD.t861 a_16167_n4181.t10 a_16222_n5759.t5 VDD.t860 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X532 a_18412_n5491.t1 a_13177_2657.t10 VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X533 a_24630_404.t11 a_25042_378.t4 a_24748_404.t7 VDD.t1045 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X534 VDD.t665 a_18684_n3216.t5 a_19680_n2629.t2 VDD.t664 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X535 a_10157_n6197.t3 a_9567_n5760.t7 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X536 a_11889_3236.t0 a_10163_n327.t6 a_11771_3236.t3 VDD.t996 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X537 VDD.t1542 a_6364_3152.t6 a_2961_n4180.t2 VDD.t1541 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X538 a_117_958.t6 B[0].t3 VDD.t1078 VDD.t1077 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X539 a_6818_316.t7 a_6273_1009.t7 a_6700_316.t8 VDD.t1093 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X540 VDD.t973 a_9512_n4182.t8 a_9572_n4156.t5 VDD.t972 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X541 VDD.t851 a_20582_5026.t11 a_22852_110.t0 VDD.t850 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X542 a_26528_404.t6 a_26940_378.t5 Y[6].t5 VDD.t611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X543 a_11883_n2634.t4 a_10148_n2943.t6 VDD.t1497 VDD.t1496 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X544 a_13025_n2630.t1 a_12029_n3217.t6 VDD.t1140 VDD.t1139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X545 VDD.t522 a_6356_n2628.t6 a_6620_n3211.t1 VDD.t521 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X546 a_3606_n6195.t0 a_3016_n5758.t8 VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X547 a_6474_n2628.t3 a_5478_n3215.t6 VDD.t1245 VDD.t1244 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X548 VDD.t105 a_16167_n4181.t11 a_19898_n5465.t7 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X549 a_31118_n4120.t1 a_29298_n5735.t10 Y[4].t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X550 VDD.t335 a_20617_n7831.t13 a_22835_n2504.t0 VDD.t334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X551 a_30764_n3388.t6 a_20021_336.t12 VDD.t671 VDD.t670 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X552 a_16227_n4155.t1 a_13968_n7819.t14 VDD.t464 VDD.t463 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X553 a_22857_1714.t5 a_22797_1688.t9 VDD.t1337 VDD.t1336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X554 a_32248_797.t4 a_29230_n745.t11 VDD.t965 VDD.t964 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X555 VSS.t121 a_22789_n4180.t11 a_23081_n6395.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X556 a_20252_n6197.t0 a_18118_n5465.t14 a_20016_n5465.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X557 a_12822_1097.t3 a_11469_404.t12 VDD.t1195 VDD.t1194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X558 a_13243_n5466.t7 a_11463_n5466.t11 VDD.t528 VDD.t527 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X559 VDD.t1014 a_22789_n4180.t12 a_22849_n4154.t0 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X560 a_13661_378.t3 a_9518_1688.t10 VDD.t500 VDD.t499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X561 a_3244_n3141.t0 a_688_n2757.t11 a_3007_n2504.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X562 a_16812_n6196.t3 a_16222_n5759.t8 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X563 a_18123_336.t2 a_18417_310.t6 a_18005_336.t1 VDD.t642 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X564 VDD.t128 a_9567_n5760.t8 a_10157_n6197.t2 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X565 VDD.t1086 a_29230_2288.t9 a_31174_4172.t2 VDD.t1085 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X566 a_4802_316.t1 a_707_521.t12 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X567 a_9518_1688.t2 a_12907_n2630.t7 VDD.t325 VDD.t324 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X568 a_13378_n8256.t5 B[2].t4 VDD.t709 VDD.t708 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X569 Y[5].t5 a_26093_n4771.t5 a_26520_n5464.t9 VDD.t984 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X570 a_26093_n4771.t2 a_24740_n5464.t12 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X571 a_10168_1277.t1 a_9578_1714.t8 VSS.t85 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X572 VDD.t937 a_12029_n3217.t7 a_13025_n2630.t0 VDD.t936 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X573 a_6620_n3211.t2 a_6356_n2628.t7 VDD.t524 VDD.t523 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X574 VDD.t60 a_3016_n5758.t9 a_3606_n6195.t1 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X575 a_25034_n5490.t3 a_20016_n5465.t16 VDD.t1233 VDD.t1232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X576 a_19898_n5465.t6 a_16167_n4181.t12 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X577 VSS.t86 a_20021_336.t13 a_31118_n4120.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X578 VSS.t206 a_16172_1620.t11 a_16464_n595.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X579 VDD.t5 a_707_521.t13 a_4802_316.t0 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X580 VDD.t542 a_6620_n3211.t11 a_10924_1097.t2 VDD.t541 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X581 a_22835_n2504.t1 a_20617_n7831.t14 VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X582 VSS.t98 a_29305_n8580.t8 a_30337_n7043.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X583 VDD.t64 a_13968_n7819.t15 a_16227_n4155.t0 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X584 a_16450_n3142.t1 a_13177_2657.t11 a_16213_n2505.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X585 a_3611_n4591.t1 a_3021_n4154.t7 VDD.t1586 VDD.t1585 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X586 a_11699_n6198.t1 a_7414_n7824.t9 a_11463_n5466.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X587 a_28640_2725.t1 A[0].t7 VDD.t1404 VDD.t1403 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X588 a_13655_n5492.t0 a_9512_n4182.t9 VSS.t122 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X589 VDD.t530 a_11463_n5466.t12 a_13243_n5466.t6 VDD.t529 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X590 VDD.t408 a_26192_3240.t6 Y[7].t2 VDD.t407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X591 a_13031_3240.t2 a_10168_1277.t7 a_12913_3240.t1 VDD.t606 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X592 a_26310_3240.t2 a_23447_1277.t4 a_26192_3240.t3 VDD.t306 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X593 a_16227_42.t6 a_16172_1620.t12 VDD.t1588 VDD.t1587 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X594 a_16803_n2942.t1 a_16213_n2505.t9 VDD.t735 VDD.t734 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X595 a_10157_n6197.t1 a_9567_n5760.t9 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X596 VDD.t837 a_19992_5463.t10 a_20582_5026.t3 VDD.t836 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X597 VDD.t1507 a_5214_n2632.t5 a_5478_n3215.t3 VDD.t1506 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X598 VDD.t695 a_12907_n2630.t8 a_9518_1688.t1 VDD.t694 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X599 VDD.t727 B[2].t5 a_13378_n8256.t4 VDD.t726 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X600 a_26520_n5464.t10 a_26093_n4771.t6 Y[5].t6 VDD.t987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X601 VDD.t100 a_24740_n5464.t13 a_26093_n4771.t1 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X602 VDD.t907 a_28640_2725.t9 a_29230_2288.t1 VDD.t906 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X603 VDD.t939 B[1].t7 a_28711_n2228.t2 VDD.t938 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X604 VDD.t1235 a_20016_n5465.t17 a_25034_n5490.t2 VDD.t1234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X605 a_30882_n4120.t1 a_31176_n3414.t5 VSS.t176 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X606 a_4802_316.t6 a_5214_290.t6 a_4920_316.t6 VDD.t1529 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X607 a_13177_2657.t1 a_12913_3240.t6 VSS.t41 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X608 a_26192_3240.t0 a_23447_1277.t5 VSS.t35 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X609 VDD.t388 a_20617_n7831.t15 a_22835_n2504.t2 VDD.t387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X610 a_16817_n4592.t1 a_16227_n4155.t8 VDD.t1054 VDD.t1053 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X611 VDD.t1459 A[3].t7 a_6789_5443.t5 VDD.t1458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X612 VDD.t1453 a_12035_2653.t5 a_13031_3240.t4 VDD.t1452 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X613 VDD.t1146 a_9572_n4156.t8 a_10162_n4593.t2 VDD.t1145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X614 a_18118_n5465.t1 a_17573_n4772.t5 a_18000_n5465.t8 VDD.t489 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X615 VDD.t1614 a_3021_n4154.t8 a_3611_n4591.t2 VDD.t1613 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X616 VSS.t146 a_6810_n5464.t15 a_11699_n6198.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X617 a_19903_336.t1 a_19476_1029.t5 a_20021_336.t1 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X618 a_26882_n328.t1 a_24748_404.t11 Y[6].t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X619 a_31118_n625.t0 a_29301_n2665.t9 Y[1].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X620 a_13243_n5466.t5 a_11463_n5466.t13 VDD.t532 VDD.t531 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X621 a_31174_4172.t0 a_29230_2288.t10 VSS.t138 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X622 VDD.t416 a_29298_n5735.t11 a_32248_n2698.t2 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X623 VDD.t1606 a_6810_n5464.t16 a_9558_n2506.t2 VDD.t1605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X624 a_7379_5006.t0 a_6789_5443.t9 VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X625 a_30762_4198.t1 a_6818_316.t14 VDD.t631 VDD.t630 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X626 VDD.t617 a_32246_4888.t9 a_9512_n4182.t2 VDD.t616 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X627 VDD.t251 a_25050_3236.t7 a_25314_2653.t2 VDD.t250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X628 VSS.t50 a_13928_5005.t10 a_18359_n396.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X629 a_26184_n2628.t1 a_23439_n4591.t6 VSS.t134 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X630 a_13378_n8256.t3 B[2].t6 VDD.t729 VDD.t728 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X631 Y[0].t2 a_28645_5296.t8 VDD.t1426 VDD.t1425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X632 a_20310_n5491.t1 a_16167_n4181.t13 VDD.t893 VDD.t892 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X633 a_9564_3364.t2 a_7379_5006.t10 VDD.t1278 VDD.t1277 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X634 a_24630_404.t9 a_20582_5026.t12 VDD.t853 VDD.t852 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X635 a_28711_n2228.t1 B[1].t8 VDD.t941 VDD.t940 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X636 a_16232_1646.t6 a_16172_1620.t13 VDD.t1590 VDD.t1589 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X637 a_354_321.t1 B[0].t4 a_117_958.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X638 a_707_521.t1 a_117_958.t10 VSS.t191 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X639 a_32485_n7683.t1 a_13361_n5466.t15 a_32248_n7046.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X640 a_9809_n4793.t1 a_9512_n4182.t10 a_9572_n4156.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X641 a_23425_n2941.t2 a_22835_n2504.t9 VDD.t1288 VDD.t1287 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X642 VDD.t1056 a_16227_n4155.t9 a_16817_n4592.t2 VDD.t1055 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X643 a_29301_n2665.t3 a_28711_n2228.t10 VSS.t183 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X644 a_10162_n4593.t3 a_9572_n4156.t9 VDD.t1148 VDD.t1147 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X645 a_18000_n5465.t11 a_17573_n4772.t6 a_18118_n5465.t4 VDD.t1315 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X646 a_3024_22.t5 a_2969_1600.t12 VDD.t831 VDD.t830 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X647 a_11463_n6198.t1 a_11757_n5492.t4 VSS.t147 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X648 VSS.t74 a_4912_n5464.t10 a_6265_n4771.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X649 a_6818_n416.t0 a_7112_290.t4 VSS.t44 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X650 a_4912_n5464.t4 a_4367_n4771.t7 a_4794_n5464.t3 VDD.t888 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X651 VSS.t117 a_13367_404.t15 a_17578_1029.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X652 a_22789_n4180.t3 a_32248_n2698.t8 VDD.t192 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X653 VDD.t319 a_22852_110.t8 a_23442_n327.t2 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X654 VSS.t78 B[0].t5 a_28877_n945.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X655 a_9558_n2506.t1 a_6810_n5464.t17 VDD.t1608 VDD.t1607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X656 VSS.t107 a_25306_n3215.t6 a_26184_n2628.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X657 VDD.t1461 A[3].t8 a_13378_n8256.t6 VDD.t1460 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X658 a_6692_n5464.t5 a_7104_n5490.t5 a_6810_n5464.t6 VDD.t751 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X659 a_9804_n6397.t0 a_6810_n5464.t18 a_9567_n5760.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X660 a_16455_2659.t0 a_13928_5005.t11 a_16218_3296.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X661 a_13249_404.t5 a_13661_378.t4 a_13367_404.t5 VDD.t488 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X662 a_17578_1029.t2 a_13367_404.t16 VDD.t841 VDD.t840 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X663 VSS.t73 a_29305_n8580.t9 a_32485_n7683.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X664 VSS.t207 a_18118_n5465.t15 a_19471_n4772.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X665 VSS.t189 a_7414_n7824.t10 a_9809_n4793.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X666 a_5486_2565.t2 a_5222_3148.t6 VDD.t1443 VDD.t1442 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X667 VSS.t139 a_29230_2288.t11 a_31116_3466.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X668 a_18123_336.t0 a_17578_1029.t4 a_18005_336.t11 VDD.t494 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X669 a_18118_n5465.t3 a_17573_n4772.t7 a_18000_n5465.t10 VDD.t1252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X670 a_13661_378.t2 a_9518_1688.t11 VDD.t502 VDD.t501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X671 a_11469_404.t4 a_10924_1097.t5 a_11351_404.t10 VDD.t876 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X672 VDD.t420 a_13928_5005.t12 a_16227_42.t0 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X673 a_26940_378.t2 a_22797_1688.t10 VDD.t1339 VDD.t1338 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X674 a_20021_336.t5 a_19476_1029.t6 a_19903_336.t3 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X675 VDD.t386 A[2].t6 a_117_958.t2 VDD.t385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X676 a_13655_n5492.t3 a_9512_n4182.t11 VDD.t1189 VDD.t1188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X677 a_16218_3296.t0 a_13928_5005.t13 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X678 a_23447_1277.t0 a_22857_1714.t9 VSS.t51 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X679 VDD.t967 a_29230_n745.t12 a_32248_797.t5 VDD.t966 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X680 VDD.t629 a_6818_316.t15 a_30335_4891.t2 VDD.t628 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X681 a_20257_n396.t1 a_18123_336.t12 a_20021_336.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X682 VDD.t1487 a_7414_n7824.t11 a_9558_n2506.t6 VDD.t1486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X683 a_25042_n2632.t2 a_23434_n6195.t4 VSS.t111 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X684 VDD.t390 a_20617_n7831.t16 a_24195_n4771.t3 VDD.t389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X685 VDD.t1475 a_29301_n2665.t10 a_30337_800.t3 VDD.t1474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X686 a_13378_n8256.t1 A[3].t9 VDD.t745 VDD.t744 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X687 a_6810_n5464.t1 a_7104_n5490.t6 a_6692_n5464.t0 VDD.t400 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X688 VDD.t586 a_6620_n3211.t12 a_9578_1714.t5 VDD.t585 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X689 VDD.t572 a_19826_n3212.t9 a_22857_1714.t2 VDD.t571 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X690 VSS.t151 a_9512_n4182.t12 a_9804_n6397.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X691 a_13338_5442.t5 B[2].t7 VDD.t731 VDD.t730 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X692 VSS.t180 A[0].t8 a_28948_n2865.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X693 VDD.t1280 a_7379_5006.t11 a_11763_378.t3 VDD.t1279 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X694 a_9578_1714.t2 a_9518_1688.t12 VDD.t558 VDD.t557 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X695 VDD.t560 a_9518_1688.t13 a_9573_110.t1 VDD.t559 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X696 a_20264_n7831.t1 B[3].t7 a_20027_n8268.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X697 a_10168_1277.t2 a_9578_1714.t9 VDD.t667 VDD.t666 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X698 a_31176_n3414.t3 a_20021_336.t14 VDD.t673 VDD.t672 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X699 VDD.t1341 a_22797_1688.t11 a_22852_110.t6 VDD.t1340 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X700 a_11345_n5466.t9 a_7414_n7824.t12 VDD.t1489 VDD.t1488 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X701 a_26310_3240.t1 a_23447_1277.t6 a_26192_3240.t2 VDD.t307 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X702 VDD.t969 a_29230_n745.t13 a_30764_107.t8 VDD.t968 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X703 VSS.t30 a_18684_n3216.t6 a_19562_n2629.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X704 a_24740_n5464.t7 a_24195_n4771.t5 a_24622_n5464.t7 VDD.t1066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X705 a_3261_n615.t0 a_715_3106.t11 a_3024_22.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X706 a_24748_404.t4 a_25042_378.t5 a_24630_404.t2 VDD.t260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X707 a_9558_n2506.t5 a_7414_n7824.t13 VDD.t283 VDD.t282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X708 a_24195_n4771.t2 a_20617_n7831.t17 VDD.t392 VDD.t391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X709 VDD.t410 a_26192_3240.t7 Y[7].t1 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X710 VDD.t588 a_6620_n3211.t13 a_9578_1714.t4 VDD.t587 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X711 a_6692_n5464.t8 a_7104_n5490.t7 a_6810_n5464.t7 VDD.t1069 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X712 VSS.t181 A[0].t9 a_28882_4659.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X713 a_22843_3364.t1 a_20582_5026.t13 VDD.t313 VDD.t312 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X714 a_29230_2288.t0 a_28640_2725.t10 VSS.t114 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X715 Y[7].t0 a_26192_3240.t8 VSS.t65 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X716 VDD.t19 a_13928_5005.t14 a_18005_336.t4 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X717 a_26528_404.t10 a_24748_404.t12 VDD.t1521 VDD.t1520 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X718 VDD.t733 a_16213_n2505.t10 a_16803_n2942.t0 VDD.t732 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X719 VDD.t460 B[3].t8 a_20027_n8268.t3 VDD.t459 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X720 VDD.t9 a_715_3106.t12 a_3024_22.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X721 VDD.t777 A[1].t7 a_6824_n8261.t2 VDD.t776 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X722 VSS.t46 A[2].t7 a_20264_n7831.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X723 VDD.t85 a_19826_n3212.t10 a_22843_3364.t5 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X724 a_3029_1626.t4 a_2969_1600.t13 VDD.t264 VDD.t263 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X725 VDD.t1197 a_20021_336.t15 a_31176_n3414.t2 VDD.t1196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X726 a_18543_3168.t0 a_16817_n395.t6 a_18425_3168.t1 VDD.t1441 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X727 a_28877_2088.t0 A[0].t10 a_28640_2725.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X728 VDD.t1126 a_9518_1688.t14 a_13249_404.t7 VDD.t1125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X729 a_16213_n2505.t4 a_13177_2657.t12 VDD.t200 VDD.t199 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X730 VDD.t1373 a_32248_797.t8 a_2969_1600.t2 VDD.t1372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X731 a_30762_4198.t3 a_29230_2288.t12 VDD.t440 VDD.t439 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X732 VSS.t171 a_23433_2927.t5 a_25050_3236.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X733 a_19826_n3212.t3 a_19562_n2629.t8 VSS.t102 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X734 a_19898_n5465.t1 a_19471_n4772.t6 a_20016_n5465.t1 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X735 a_26520_n5464.t6 a_22789_n4180.t13 VDD.t1016 VDD.t1015 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X736 VDD.t110 a_688_n2757.t12 a_3007_n2504.t3 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X737 a_362_2906.t0 A[1].t8 a_125_3543.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X738 a_19685_3172.t2 a_18689_2585.t5 VDD.t1600 VDD.t1599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X739 VDD.t779 A[1].t9 a_28640_n308.t1 VDD.t778 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X740 VSS.t179 A[0].t11 a_28952_n8780.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X741 a_3258_n4791.t0 a_2961_n4180.t10 a_3021_n4154.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X742 a_6824_n8261.t1 A[1].t10 VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X743 VDD.t895 a_16167_n4181.t14 a_20310_n5491.t2 VDD.t894 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X744 VSS.t133 A[2].t8 a_354_321.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X745 a_31176_n3414.t1 a_20021_336.t16 VDD.t1199 VDD.t1198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X746 a_125_3543.t1 A[1].t11 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X747 VDD.t927 a_13177_2657.t13 a_16213_n2505.t6 VDD.t926 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X748 VDD.t1018 a_22789_n4180.t14 a_22844_n5758.t6 VDD.t1017 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X749 a_6482_3152.t5 a_5486_2565.t5 VDD.t1000 VDD.t999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X750 a_24748_n328.t1 a_25042_378.t6 VSS.t87 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X751 a_17573_n4772.t2 a_13968_n7819.t16 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X752 a_25168_3236.t1 a_23442_n327.t5 a_25050_3236.t3 VDD.t1379 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X753 VSS.t6 a_4920_316.t11 a_6273_1009.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X754 VDD.t943 B[1].t9 a_98_n2320.t5 VDD.t942 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X755 VSS.t203 a_16803_n2942.t4 a_18420_n2633.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X756 a_20016_n5465.t0 a_19471_n4772.t7 a_19898_n5465.t0 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X757 VDD.t1020 a_22789_n4180.t15 a_26520_n5464.t5 VDD.t1019 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X758 Y[6].t2 a_26101_1097.t4 a_26528_404.t3 VDD.t599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X759 a_3007_n2504.t2 a_688_n2757.t13 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X760 a_3015_3276.t6 a_707_521.t14 VDD.t1030 VDD.t1029 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X761 a_704_n5517.t3 a_114_n5080.t9 VDD.t1518 VDD.t1517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X762 a_19567_3172.t3 a_16822_1209.t5 a_19685_3172.t5 VDD.t1247 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X763 VSS.t84 a_6620_n3211.t14 a_10924_1097.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X764 a_5478_n3215.t0 a_5214_n2632.t6 VSS.t64 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X765 a_3253_n6395.t0 a_688_n2757.t14 a_3016_n5758.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X766 a_26638_n6196.t0 a_26932_n5490.t5 VSS.t90 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X767 a_3021_n4154.t2 a_2961_n4180.t11 VDD.t1298 VDD.t1297 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X768 VSS.t31 a_7414_n7824.t14 a_10918_n4773.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X769 VDD.t1602 a_10154_2927.t6 a_11889_3236.t4 VDD.t1601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X770 VDD.t1357 a_23433_2927.t6 a_25168_3236.t4 VDD.t1356 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X771 VDD.t147 A[1].t12 a_6824_n8261.t0 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X772 VSS.t136 a_704_n5517.t16 a_4367_n4771.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X773 VDD.t1152 B[0].t6 a_114_n5080.t3 VDD.t1151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X774 VDD.t1449 a_3015_3276.t8 a_3605_2839.t2 VDD.t1448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X775 VSS.t209 a_18689_2585.t6 a_19567_3172.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X776 a_26101_1097.t2 a_24748_404.t13 VDD.t1523 VDD.t1522 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X777 VDD.t1509 a_29301_n2665.t11 a_30337_800.t2 VDD.t1508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X778 VDD.t448 a_6356_n2628.t8 a_6620_n3211.t0 VDD.t447 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X779 a_20229_4826.t1 A[3].t10 a_19992_5463.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X780 a_18005_336.t0 a_18417_310.t7 a_18123_336.t3 VDD.t643 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X781 a_22844_n5758.t5 a_22789_n4180.t16 VDD.t911 VDD.t910 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X782 a_26302_n2628.t5 a_23439_n4591.t7 a_26184_n2628.t2 VDD.t1074 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X783 VDD.t68 a_13968_n7819.t17 a_17573_n4772.t1 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X784 Y[0].t0 a_28645_5296.t9 VSS.t182 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X785 VDD.t87 a_19826_n3212.t11 a_22857_1714.t1 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X786 a_688_n2757.t3 a_98_n2320.t8 VDD.t1621 VDD.t1620 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X787 a_18684_n3216.t1 a_18420_n2633.t5 VSS.t61 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X788 a_7061_n7824.t1 B[2].t8 a_6824_n8261.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X789 a_3614_n415.t2 a_3024_22.t9 VDD.t162 VDD.t161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X790 a_11463_n5466.t3 a_10918_n4773.t7 a_11345_n5466.t3 VDD.t750 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X791 a_13928_5005.t1 a_13338_5442.t9 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X792 a_16218_3296.t5 a_13367_404.t17 VDD.t843 VDD.t842 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X793 VSS.t127 a_707_521.t15 a_3266_989.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X794 a_20021_n396.t0 a_20315_310.t7 VSS.t59 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X795 a_10148_n2943.t3 a_9558_n2506.t10 VSS.t197 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X796 a_13928_5005.t0 a_13338_5442.t10 VSS.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X797 a_9567_n5760.t3 a_6810_n5464.t19 VDD.t711 VDD.t710 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X798 a_7026_4806.t0 B[1].t10 a_6789_5443.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X799 VDD.t657 a_6620_n3211.t15 a_10924_1097.t1 VDD.t656 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X800 VDD.t89 a_19826_n3212.t12 a_24203_1097.t2 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X801 VSS.t169 a_22797_1688.t12 a_23089_n527.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X802 a_19992_5463.t2 A[3].t11 VDD.t747 VDD.t746 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X803 VDD.t796 a_715_3106.t13 a_4802_316.t4 VDD.t795 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X804 a_7414_n7824.t2 a_6824_n8261.t9 VDD.t1363 VDD.t1362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X805 a_114_n5080.t2 B[0].t7 VDD.t1154 VDD.t1153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X806 a_20315_310.t1 a_16172_1620.t14 VDD.t1162 VDD.t1161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X807 VDD.t913 a_22789_n4180.t17 a_22844_n5758.t4 VDD.t912 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X808 VSS.t20 A[3].t12 a_7026_4806.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X809 VDD.t1207 a_25306_n3215.t7 a_26302_n2628.t0 VDD.t1206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X810 a_5340_3148.t4 a_3614_n415.t6 a_5222_3148.t2 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X811 a_6700_316.t7 a_7112_290.t5 a_6818_316.t1 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X812 a_23442_n327.t1 a_22852_110.t9 VDD.t321 VDD.t320 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X813 VDD.t1369 a_98_n2320.t9 a_688_n2757.t1 VDD.t1368 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X814 a_6789_5443.t2 B[1].t11 VDD.t865 VDD.t864 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X815 a_26310_3240.t4 a_25314_2653.t5 VDD.t506 VDD.t505 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X816 VDD.t1164 a_16172_1620.t15 a_16227_42.t2 VDD.t1163 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X817 a_26528_404.t11 a_24748_404.t14 VDD.t1566 VDD.t1565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X818 a_20617_n7831.t3 a_20027_n8268.t10 VDD.t1619 VDD.t1618 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X819 a_11345_n5466.t10 a_11757_n5492.t5 a_11463_n5466.t6 VDD.t805 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X820 VDD.t442 a_29230_2288.t13 a_32246_4888.t0 VDD.t441 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X821 VDD.t757 B[2].t9 a_28640_2725.t6 VDD.t756 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X822 a_32483_4251.t1 a_29230_2288.t14 a_32246_4888.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X823 VDD.t1050 a_12913_3240.t7 a_13177_2657.t2 VDD.t1049 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X824 VSS.t145 a_9518_1688.t15 a_9810_n527.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X825 a_18684_n3216.t2 a_18420_n2633.t6 VDD.t839 VDD.t838 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X826 VDD.t592 a_6810_n5464.t20 a_9567_n5760.t0 VDD.t591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X827 Y[2].t6 a_31174_4172.t6 a_30762_4198.t7 VDD.t754 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X828 VDD.t21 a_13928_5005.t15 a_18005_336.t3 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X829 Y[4].t1 a_30337_n2695.t5 a_30764_n3388.t3 VDD.t1317 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X830 VDD.t135 A[3].t13 a_6789_5443.t4 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X831 VDD.t298 a_3605_2839.t6 a_5340_3148.t1 VDD.t297 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X832 a_18005_336.t10 a_17578_1029.t5 a_18123_336.t1 VDD.t495 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X833 a_30337_n2695.t2 a_29298_n5735.t12 VDD.t1438 VDD.t1437 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X834 VDD.t1365 a_6824_n8261.t10 a_7414_n7824.t3 VDD.t1364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X835 a_30764_n7736.t2 a_29305_n8580.t10 VDD.t574 VDD.t573 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X836 a_16808_2859.t0 a_16218_3296.t9 VSS.t135 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X837 a_13603_n328.t1 a_11469_404.t13 a_13367_404.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X838 VDD.t91 a_19826_n3212.t13 a_24630_404.t5 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X839 VDD.t1220 a_26184_n2628.t6 a_22797_1688.t2 VDD.t1219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X840 a_23434_n6195.t1 a_22844_n5758.t10 VDD.t1554 VDD.t1553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X841 VDD.t266 a_2969_1600.t14 a_7112_290.t1 VDD.t265 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X842 a_16227_42.t3 a_13928_5005.t16 VDD.t1550 VDD.t1549 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X843 VDD.t428 a_3029_1626.t10 a_3619_1189.t1 VDD.t427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X844 a_688_n2757.t0 a_98_n2320.t10 VDD.t1367 VDD.t1366 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X845 a_25160_n2632.t5 a_23434_n6195.t5 a_25042_n2632.t3 VDD.t885 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X846 VDD.t933 a_11771_3236.t8 a_12035_2653.t1 VDD.t932 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X847 VDD.t761 a_4920_316.t12 a_6273_1009.t2 VDD.t760 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X848 a_18123_336.t5 a_17578_1029.t6 a_18123_n396.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X849 a_11463_n5466.t7 a_11757_n5492.t6 a_11345_n5466.t11 VDD.t1180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X850 Y[0].t1 a_28645_5296.t10 VDD.t1428 VDD.t1427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X851 a_3007_n2504.t1 a_688_n2757.t15 VDD.t1128 VDD.t1127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X852 VDD.t39 a_20617_n7831.t18 a_22849_n4154.t4 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X853 VDD.t1022 a_18420_n2633.t7 a_18684_n3216.t3 VDD.t1021 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X854 a_24740_n5464.t2 a_24195_n4771.t6 a_24740_n6196.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X855 a_9567_n5760.t1 a_6810_n5464.t21 VDD.t594 VDD.t593 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X856 a_16232_1646.t3 a_13367_404.t18 VDD.t845 VDD.t844 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X857 VDD.t1576 B[0].t8 a_28640_n308.t5 VDD.t1575 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X858 a_30764_n3388.t4 a_30337_n2695.t6 Y[4].t2 VDD.t1376 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X859 VDD.t1440 a_29298_n5735.t13 a_30337_n2695.t1 VDD.t1439 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X860 a_125_3543.t4 B[1].t12 VDD.t867 VDD.t866 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X861 Y[6].t1 a_26101_1097.t5 a_26528_404.t2 VDD.t555 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X862 a_26874_n6196.t0 a_24740_n5464.t14 Y[5].t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X863 VDD.t576 a_29305_n8580.t11 a_30764_n7736.t1 VDD.t575 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X864 VDD.t268 a_2969_1600.t15 a_3024_22.t4 VDD.t267 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X865 VDD.t873 a_18123_336.t13 a_19903_336.t7 VDD.t872 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X866 a_30764_107.t9 a_29230_n745.t14 VDD.t1572 VDD.t1571 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X867 a_28640_n308.t6 B[0].t9 VDD.t1578 VDD.t1577 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X868 VDD.t1264 a_5478_n3215.t7 a_6474_n2628.t4 VDD.t1263 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X869 VDD.t578 a_13361_n5466.t16 a_32248_n7046.t5 VDD.t577 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X870 VSS.t70 a_19826_n3212.t14 a_24203_1097.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X871 VDD.t1385 B[3].t9 a_28708_n5298.t6 VDD.t1384 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X872 VDD.t1177 a_125_3543.t9 a_715_3106.t2 VDD.t1176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X873 VDD.t1215 a_18689_2585.t7 a_19685_3172.t1 VDD.t1214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X874 a_11345_n5466.t6 a_11757_n5492.t7 a_11463_n5466.t4 VDD.t556 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X875 a_13367_404.t7 a_13661_378.t5 a_13249_404.t10 VDD.t1171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X876 a_23439_n4591.t1 a_22849_n4154.t10 VDD.t424 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X877 VDD.t1349 a_23433_2927.t7 a_25168_3236.t3 VDD.t1348 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X878 a_19903_336.t10 a_16172_1620.t16 VDD.t1166 VDD.t1165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X879 a_29305_n8580.t0 a_28715_n8143.t9 VDD.t396 VDD.t395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X880 VDD.t675 a_9512_n4182.t13 a_9567_n5760.t5 VDD.t674 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X881 VSS.t193 a_29298_n5735.t14 a_30337_n2695.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X882 VDD.t763 a_4920_316.t13 a_6700_316.t1 VDD.t762 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X883 a_3024_22.t0 a_715_3106.t14 VDD.t798 VDD.t797 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X884 a_11351_404.t8 a_10924_1097.t6 a_11469_404.t2 VDD.t714 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X885 a_117_958.t1 A[2].t9 VDD.t1072 VDD.t1071 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X886 VSS.t115 a_22789_n4180.t18 a_26874_n6196.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X887 a_28945_n5935.t1 A[1].t13 a_28708_n5298.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X888 a_6700_316.t0 a_4920_316.t14 VDD.t765 VDD.t764 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X889 a_9572_n4156.t4 a_9512_n4182.t14 VDD.t677 VDD.t676 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X890 a_32248_n7046.t4 a_13361_n5466.t17 VDD.t580 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X891 VDD.t627 a_6818_316.t16 a_30335_4891.t1 VDD.t626 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X892 a_16808_2859.t1 a_16218_3296.t10 VDD.t1104 VDD.t1103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X893 a_30337_800.t1 a_29301_n2665.t12 VDD.t1511 VDD.t1510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X894 a_29298_n5735.t3 a_28708_n5298.t8 VDD.t1099 VDD.t1098 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X895 a_18689_2585.t0 a_18425_3168.t6 VSS.t49 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X896 VDD.t422 a_22857_1714.t10 a_23447_1277.t1 VDD.t421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X897 VDD.t1201 a_20021_336.t17 a_30764_n3388.t5 VDD.t1200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X898 VDD.t564 a_19826_n3212.t15 a_24203_1097.t1 VDD.t563 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X899 a_30764_n7736.t3 a_31176_n7762.t7 Y[3].t3 VDD.t950 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X900 VSS.t18 a_688_n2757.t16 a_5148_n6196.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X901 a_9573_110.t3 a_7379_5006.t12 VDD.t1270 VDD.t1269 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X902 a_5214_290.t0 a_715_3106.t15 VSS.t104 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X903 a_22852_110.t5 a_22797_1688.t13 VDD.t1333 VDD.t1332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X904 a_6692_n5464.t1 a_4912_n5464.t11 VDD.t596 VDD.t595 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X905 VDD.t141 a_16222_n5759.t9 a_16812_n6196.t2 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X906 a_19992_5463.t5 B[3].t10 VDD.t1381 VDD.t1380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X907 VSS.t186 a_12035_2653.t6 a_12913_3240.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X908 a_24630_404.t10 a_25042_378.t7 a_24748_404.t6 VDD.t889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X909 VDD.t285 a_7414_n7824.t15 a_9572_n4156.t1 VDD.t284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X910 VDD.t1024 a_29305_n8580.t12 a_32248_n7046.t1 VDD.t1023 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X911 VDD.t534 a_11463_n5466.t14 a_12816_n4773.t2 VDD.t533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X912 VDD.t1101 a_28708_n5298.t9 a_29298_n5735.t2 VDD.t1100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X913 VDD.t1052 a_12913_3240.t8 a_13177_2657.t3 VDD.t1051 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X914 VSS.t118 a_13177_2657.t14 a_18354_n6197.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X915 a_16222_n5759.t2 a_13177_2657.t15 VDD.t929 VDD.t928 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X916 a_10163_n327.t2 a_9573_110.t8 VDD.t1251 VDD.t1250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X917 a_5332_n2632.t0 a_3606_n6195.t6 a_5214_n2632.t2 VDD.t435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X918 a_117_958.t5 B[0].t10 VDD.t180 VDD.t179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X919 a_13249_404.t8 a_11469_404.t14 VDD.t1142 VDD.t1141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X920 VSS.t88 a_24740_n5464.t15 a_26093_n4771.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X921 a_16172_1620.t0 a_32248_n7046.t10 VSS.t42 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X922 a_26932_n5490.t1 a_22789_n4180.t19 VDD.t915 VDD.t914 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X923 a_2969_1600.t3 a_32248_797.t9 VDD.t1375 VDD.t1374 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X924 a_4912_n6196.t1 a_5206_n5490.t4 VSS.t81 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X925 VDD.t122 a_688_n2757.t17 a_3016_n5758.t3 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X926 VDD.t625 a_6818_316.t17 a_30762_4198.t0 VDD.t624 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X927 a_9512_n4182.t1 a_32246_4888.t10 VDD.t615 VDD.t614 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X928 a_11771_3236.t4 a_10163_n327.t7 VSS.t125 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X929 Y[1].t6 a_30337_800.t5 a_30882_n625.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X930 VDD.t1300 a_2961_n4180.t12 a_6692_n5464.t2 VDD.t1299 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X931 VDD.t1006 a_6620_n3211.t16 a_9564_3364.t5 VDD.t1005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X932 a_13367_n328.t1 a_13661_378.t6 VSS.t157 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X933 a_335_n2957.t0 A[2].t10 a_98_n2320.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X934 VDD.t56 a_18420_n2633.t8 a_18684_n3216.t0 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X935 a_18543_3168.t3 a_16808_2859.t6 VDD.t1319 VDD.t1318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X936 VDD.t1335 a_22797_1688.t14 a_26528_404.t7 VDD.t1334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X937 a_30764_107.t6 a_30337_800.t6 Y[1].t2 VDD.t338 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X938 VDD.t473 a_13177_2657.t16 a_18000_n5465.t5 VDD.t472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X939 VDD.t536 a_4920_316.t15 a_6273_1009.t1 VDD.t535 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X940 a_5478_n3215.t2 a_5214_n2632.t7 VDD.t487 VDD.t486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X941 a_18538_n2633.t0 a_16812_n6196.t7 a_18420_n2633.t0 VDD.t497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X942 VDD.t1398 A[0].t12 a_28711_n2228.t6 VDD.t1397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X943 a_9572_n4156.t0 a_7414_n7824.t16 VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X944 a_32248_n7046.t0 a_29305_n8580.t13 VDD.t1026 VDD.t1025 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X945 a_12816_n4773.t1 a_11463_n5466.t15 VDD.t483 VDD.t482 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X946 a_29298_n5735.t1 a_28708_n5298.t10 VDD.t1175 VDD.t1174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X947 a_16817_n4592.t3 a_16227_n4155.t10 VDD.t1387 VDD.t1386 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X948 a_18118_n6197.t1 a_18412_n5491.t5 VSS.t8 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X949 VDD.t475 a_13177_2657.t17 a_16222_n5759.t1 VDD.t474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X950 VDD.t1321 a_16808_2859.t7 a_18543_3168.t4 VDD.t1320 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X951 VDD.t1229 a_3597_n2941.t5 a_5332_n2632.t5 VDD.t1228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X952 VSS.t161 a_7379_5006.t13 a_11705_n328.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X953 a_3016_n5758.t2 a_688_n2757.t18 VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X954 a_3252_2639.t1 a_715_3106.t16 a_3015_3276.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X955 VDD.t514 a_19567_3172.t8 a_16167_n4181.t1 VDD.t513 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X956 a_5214_290.t1 a_715_3106.t17 VDD.t817 VDD.t816 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X957 VDD.t649 a_32248_n2698.t9 a_22789_n4180.t2 VDD.t648 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X958 a_4375_1009.t1 a_707_521.t16 VDD.t1032 VDD.t1031 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X959 a_10163_n327.t0 a_9573_110.t9 VSS.t160 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X960 a_704_n5517.t0 a_114_n5080.t10 VSS.t10 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X961 VSS.t110 B[1].t13 a_335_n2957.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X962 a_16227_n4155.t5 a_16167_n4181.t15 VDD.t1002 VDD.t1001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X963 a_29230_n745.t2 a_28640_n308.t9 VDD.t170 VDD.t169 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X964 a_19680_n2629.t0 a_18684_n3216.t7 VDD.t216 VDD.t215 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X965 Y[5].t1 a_26932_n5490.t6 a_26520_n5464.t0 VDD.t393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X966 VDD.t875 a_18123_336.t14 a_19476_1029.t1 VDD.t874 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X967 VDD.t1302 a_2961_n4180.t13 a_3021_n4154.t1 VDD.t1301 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X968 a_6818_316.t2 a_7112_290.t6 a_6700_316.t6 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X969 a_26528_404.t1 a_26101_1097.t6 Y[6].t0 VDD.t434 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X970 VDD.t1596 a_5214_n2632.t8 a_5478_n3215.t1 VDD.t1595 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X971 VDD.t994 a_16803_n2942.t5 a_18538_n2633.t5 VDD.t993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X972 a_28711_n2228.t5 A[0].t13 VDD.t1400 VDD.t1399 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X973 a_3015_3276.t1 a_715_3106.t18 VDD.t819 VDD.t818 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X974 a_13968_n7819.t3 a_13378_n8256.t10 VSS.t120 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X975 a_5332_n2632.t4 a_3597_n2941.t6 VDD.t1227 VDD.t1226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X976 a_12907_n2630.t2 a_10162_n4593.t6 a_13025_n2630.t4 VDD.t310 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X977 VDD.t1604 a_10154_2927.t7 a_11889_3236.t5 VDD.t1603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X978 a_22789_n4180.t1 a_32248_n2698.t10 VDD.t651 VDD.t650 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X979 a_31174_4172.t1 a_29230_2288.t15 VDD.t444 VDD.t443 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X980 a_32485_n3335.t0 a_20021_336.t18 a_32248_n2698.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X981 VDD.t1535 A[2].t11 a_13338_5442.t6 VDD.t1534 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X982 a_6700_316.t9 a_2969_1600.t16 VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X983 VDD.t1004 a_16167_n4181.t16 a_16227_n4155.t4 VDD.t1003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X984 a_25042_378.t2 a_20582_5026.t14 VDD.t315 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X985 a_16464_n595.t0 a_13928_5005.t17 a_16227_42.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X986 a_22797_1688.t1 a_26184_n2628.t7 VSS.t154 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X987 a_3021_n4154.t0 a_2961_n4180.t14 VDD.t1304 VDD.t1303 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X988 a_6692_n5464.t6 a_4912_n5464.t12 VDD.t897 VDD.t896 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X989 a_18538_n2633.t4 a_16803_n2942.t6 VDD.t992 VDD.t991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X990 VDD.t1402 A[0].t14 a_28711_n2228.t4 VDD.t1401 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X991 a_3266_989.t1 a_2969_1600.t17 a_3029_1626.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X992 a_28715_n8143.t3 B[3].t11 VDD.t1631 VDD.t1630 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X993 VDD.t1499 a_10148_n2943.t7 a_11883_n2634.t3 VDD.t1498 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X994 a_32248_n2698.t1 a_20021_336.t19 VDD.t358 VDD.t357 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X995 a_29305_n8580.t1 a_28715_n8143.t10 VSS.t67 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X996 VDD.t1225 a_3597_n2941.t7 a_5332_n2632.t3 VDD.t1224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X997 VSS.t0 a_6818_316.t18 a_30335_4891.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X998 VDD.t1182 a_715_3106.t19 a_4802_316.t3 VDD.t1181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X999 VSS.t16 a_16167_n4181.t17 a_20252_n6197.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1000 VSS.t21 A[3].t14 a_351_n5717.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1001 VSS.t194 a_29298_n5735.t15 a_32485_n3335.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1002 a_23080_2727.t0 a_20582_5026.t15 a_22843_3364.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1003 a_4802_316.t10 a_4375_1009.t5 a_4920_316.t2 VDD.t598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1004 VSS.t137 a_704_n5517.t17 a_3244_n3141.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1005 VSS.t153 a_23425_n2941.t6 a_25042_n2632.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1006 a_7104_n5490.t0 a_2961_n4180.t15 VSS.t165 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1007 VDD.t899 a_4912_n5464.t13 a_6692_n5464.t7 VDD.t898 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1008 a_5340_3148.t3 a_3614_n415.t7 a_5222_3148.t4 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1009 VDD.t70 a_20582_5026.t16 a_22843_3364.t0 VDD.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1010 a_18005_336.t7 a_13367_404.t19 VDD.t847 VDD.t846 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1011 a_13031_3240.t3 a_12035_2653.t7 VDD.t1455 VDD.t1454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1012 VDD.t1383 B[3].t12 a_28715_n8143.t2 VDD.t1382 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1013 a_3606_n6195.t2 a_3016_n5758.t10 VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1014 a_28645_5296.t0 B[0].t11 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1015 VSS.t71 a_19826_n3212.t16 a_23094_1077.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1016 a_16817_n395.t1 a_16227_42.t10 VDD.t196 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1017 VDD.t114 a_16167_n4181.t18 a_19898_n5465.t5 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1018 a_13249_404.t0 a_13661_378.t7 a_13367_404.t0 VDD.t233 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1019 a_715_3106.t1 a_125_3543.t10 VDD.t1179 VDD.t1178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1020 Y[6].t3 a_26101_1097.t7 a_26646_n328.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1021 a_13615_n7819.t0 B[2].t10 a_13378_n8256.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1022 a_13249_404.t9 a_11469_404.t15 VDD.t1144 VDD.t1143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1023 a_18123_336.t6 a_17578_1029.t7 a_18005_336.t9 VDD.t1514 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1024 VDD.t1028 a_29305_n8580.t14 a_30337_n7043.t3 VDD.t1027 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1025 VDD.t158 a_6789_5443.t10 a_7379_5006.t1 VDD.t157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1026 a_11757_n5492.t0 a_6810_n5464.t22 VSS.t14 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1027 VDD.t208 a_7414_n7824.t17 a_11345_n5466.t8 VDD.t207 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1028 a_9801_2727.t0 a_7379_5006.t14 a_9564_3364.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1029 a_25314_2653.t1 a_25050_3236.t8 VDD.t253 VDD.t252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1030 VDD.t230 A[2].t12 a_117_958.t0 VDD.t229 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1031 a_3016_n5758.t1 a_688_n2757.t19 VDD.t493 VDD.t492 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1032 VSS.t5 a_18123_336.t15 a_19476_1029.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1033 a_30882_n625.t0 a_31176_81.t7 VSS.t11 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1034 a_24622_n5464.t6 a_24195_n4771.t7 a_24740_n5464.t3 VDD.t604 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1035 VDD.t41 a_20617_n7831.t19 a_24195_n4771.t1 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1036 VDD.t418 a_9564_3364.t10 a_10154_2927.t1 VDD.t417 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1037 VDD.t1008 a_6620_n3211.t17 a_11351_404.t11 VDD.t1007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1038 a_25306_n3215.t0 a_25042_n2632.t6 VSS.t187 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1039 VDD.t1556 a_16172_1620.t17 a_16227_42.t5 VDD.t1555 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1040 Y[4].t0 a_30337_n2695.t7 a_30764_n3388.t2 VDD.t1316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1041 Y[5].t7 a_26093_n4771.t7 a_26520_n5464.t11 VDD.t988 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1042 a_10157_n6197.t0 a_9567_n5760.t10 VSS.t19 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1043 VSS.t123 a_6620_n3211.t18 a_9815_1077.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1044 a_28715_n8143.t1 B[3].t13 VDD.t1629 VDD.t1628 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1045 a_4920_316.t3 a_4375_1009.t6 a_4920_n416.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1046 a_25034_n5490.t1 a_20016_n5465.t18 VDD.t1237 VDD.t1236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1047 VSS.t210 a_2969_1600.t18 a_7054_n416.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1048 a_9564_3364.t1 a_7379_5006.t15 VDD.t1272 VDD.t1271 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1049 VSS.t3 A[3].t15 a_13615_n7819.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1050 a_2961_n4180.t3 a_6364_3152.t7 VDD.t1544 VDD.t1543 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1051 a_23442_n327.t0 a_22852_110.t10 VSS.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1052 a_6364_3152.t1 a_3619_1189.t7 a_6482_3152.t1 VDD.t498 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1053 VDD.t1118 a_7379_5006.t16 a_9573_110.t2 VDD.t1117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1054 a_28877_n945.t0 A[1].t14 a_28640_n308.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1055 a_11345_n5466.t7 a_7414_n7824.t18 VDD.t210 VDD.t209 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1056 Y[2].t1 a_30335_4891.t6 a_30880_3466.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1057 a_5156_n416.t0 a_707_521.t17 a_4920_316.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1058 a_3611_n4591.t3 a_3021_n4154.t9 VDD.t1616 VDD.t1615 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1059 a_3614_n415.t1 a_3024_22.t10 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1060 VDD.t1574 a_29230_n745.t15 a_30764_107.t10 VDD.t1573 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1061 VDD.t679 a_9512_n4182.t15 a_13243_n5466.t10 VDD.t678 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1062 VSS.t93 a_5486_2565.t6 a_6364_3152.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1063 VDD.t1477 a_6364_3152.t8 a_2961_n4180.t0 VDD.t1476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1064 VDD.t771 a_13367_404.t20 a_17578_1029.t1 VDD.t770 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1065 VDD.t1558 a_16172_1620.t18 a_19903_336.t11 VDD.t1557 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1066 a_29230_n745.t1 a_28640_n308.t10 VDD.t172 VDD.t171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1067 a_30764_n3388.t0 a_31176_n3414.t6 Y[4].t5 VDD.t294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1068 a_26520_n5464.t1 a_26932_n5490.t7 Y[5].t0 VDD.t394 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1069 VDD.t1445 a_5222_3148.t7 a_5486_2565.t1 VDD.t1444 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1070 a_31116_3466.t0 a_6818_316.t19 Y[2].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1071 VSS.t83 B[2].t11 a_13575_4805.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1072 VDD.t120 a_9518_1688.t16 a_13661_378.t1 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1073 a_18417_310.t1 a_13928_5005.t18 VDD.t1552 VDD.t1551 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1074 VDD.t1327 a_22797_1688.t15 a_22857_1714.t3 VDD.t1326 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1075 VDD.t1290 a_22835_n2504.t10 a_23425_n2941.t3 VDD.t1289 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1076 VDD.t1136 a_13928_5005.t19 a_16218_3296.t3 VDD.t1135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1077 a_11469_404.t3 a_10924_1097.t7 a_11351_404.t9 VDD.t715 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1078 a_20021_336.t6 a_19476_1029.t7 a_20021_n396.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1079 a_16213_n2505.t5 a_13177_2657.t18 VDD.t477 VDD.t476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1080 a_22857_1714.t4 a_22797_1688.t16 VDD.t1329 VDD.t1328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1081 a_13661_378.t0 a_9518_1688.t17 VSS.t17 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1082 a_13025_n2630.t3 a_10162_n4593.t7 a_12907_n2630.t1 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1083 a_16459_n6396.t0 a_13177_2657.t19 a_16222_n5759.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1084 VDD.t653 B[2].t12 a_13338_5442.t4 VDD.t652 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1085 a_13243_n5466.t9 a_9512_n4182.t16 VDD.t979 VDD.t978 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1086 a_4794_n5464.t0 a_5206_n5490.t5 a_4912_n5464.t0 VDD.t607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1087 a_11763_378.t2 a_7379_5006.t17 VDD.t1120 VDD.t1119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1088 a_7104_n5490.t3 a_2961_n4180.t16 VDD.t1292 VDD.t1291 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1089 VDD.t414 a_18425_3168.t7 a_18689_2585.t2 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1090 a_2969_1600.t0 a_32248_797.t10 VSS.t173 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1091 Y[4].t4 a_31176_n3414.t7 a_30764_n3388.t8 VDD.t1540 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1092 VDD.t1393 A[0].t15 a_28640_2725.t0 VDD.t1392 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1093 VSS.t212 a_13968_n7819.t18 a_17573_n4772.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1094 a_18425_3168.t0 a_16817_n395.t7 VSS.t184 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1095 VDD.t31 a_9578_1714.t10 a_10168_1277.t0 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1096 a_26192_3240.t1 a_23447_1277.t7 a_26310_3240.t0 VDD.t299 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1097 a_18689_2585.t1 a_18425_3168.t8 VDD.t287 VDD.t286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1098 VDD.t1331 a_22797_1688.t17 a_22852_110.t4 VDD.t1330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1099 a_26528_404.t5 a_26940_378.t6 Y[6].t4 VDD.t1532 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1100 a_18000_n5465.t0 a_18412_n5491.t6 a_18118_n5465.t6 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1101 a_11757_n5492.t1 a_6810_n5464.t23 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1102 Y[2].t2 a_30335_4891.t7 a_30762_4198.t6 VDD.t687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1103 a_9578_1714.t1 a_9518_1688.t18 VDD.t697 VDD.t696 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1104 a_28882_4659.t1 B[0].t12 a_28645_5296.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1105 VSS.t141 a_25314_2653.t6 a_26192_3240.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1106 a_18005_336.t6 a_13367_404.t21 VDD.t773 VDD.t772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1107 VDD.t981 a_9512_n4182.t17 a_13655_n5492.t2 VDD.t980 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1108 VSS.t25 A[1].t15 a_7061_n7824.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1109 a_4912_n5464.t6 a_5206_n5490.t6 a_4794_n5464.t10 VDD.t1579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1110 a_22835_n2504.t5 a_20016_n5465.t19 VDD.t1239 VDD.t1238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1111 VDD.t1294 a_2961_n4180.t17 a_7104_n5490.t2 VDD.t1293 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1112 a_3605_2839.t0 a_3015_3276.t9 VSS.t185 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1113 VDD.t1268 a_9573_110.t10 a_10163_n327.t1 VDD.t1267 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1114 a_22843_3364.t4 a_19826_n3212.t17 VDD.t566 VDD.t565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1115 VDD.t723 B[0].t13 a_117_958.t4 VDD.t722 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1116 a_13249_404.t6 a_9518_1688.t19 VDD.t699 VDD.t698 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1117 VDD.t1513 a_29301_n2665.t13 a_32248_797.t0 VDD.t1512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1118 a_10162_n4593.t1 a_9572_n4156.t10 VSS.t124 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1119 a_28645_5296.t5 B[0].t14 VDD.t1010 VDD.t1009 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1120 a_25050_3236.t4 a_23442_n327.t6 VSS.t215 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1121 a_3611_n4591.t0 a_3021_n4154.t10 VSS.t47 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1122 a_26646_n328.t0 a_26940_378.t7 VSS.t196 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1123 a_18118_n5465.t5 a_18412_n5491.t7 a_18000_n5465.t1 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1124 a_3029_1626.t1 a_707_521.t18 VDD.t152 VDD.t151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1125 Y[1].t1 a_30337_800.t7 a_30764_107.t5 VDD.t271 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1126 VDD.t1130 a_7414_n7824.t19 a_9558_n2506.t4 VDD.t1129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1127 a_13655_n5492.t1 a_9512_n4182.t18 VDD.t983 VDD.t982 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1128 a_4794_n5464.t11 a_5206_n5490.t7 a_4912_n5464.t7 VDD.t1580 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1129 a_24984_n328.t1 a_19826_n3212.t18 a_24748_404.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1130 VDD.t1254 a_20016_n5465.t20 a_22835_n2504.t4 VDD.t1253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1131 a_7104_n5490.t1 a_2961_n4180.t18 VDD.t1296 VDD.t1295 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1132 VDD.t1122 a_7379_5006.t18 a_11351_404.t5 VDD.t1121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1133 a_9564_3364.t4 a_6620_n3211.t19 VDD.t977 VDD.t976 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1134 VDD.t232 A[2].t13 a_98_n2320.t1 VDD.t231 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1135 VDD.t713 a_5486_2565.t7 a_6482_3152.t0 VDD.t712 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1136 a_30764_n7736.t0 a_29305_n8580.t15 VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1137 a_20027_n8268.t6 B[3].t14 VDD.t1623 VDD.t1622 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1138 VSS.t12 a_20582_5026.t17 a_24984_n328.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1139 VSS.t204 a_29301_n2665.t14 a_30337_800.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1140 a_22797_1688.t0 a_26184_n2628.t8 VDD.t1217 VDD.t1216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1141 VDD.t154 a_707_521.t19 a_3015_3276.t0 VDD.t153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1142 a_24622_n5464.t4 a_20016_n5465.t21 VDD.t1256 VDD.t1255 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1143 a_19685_3172.t0 a_16822_1209.t6 a_19567_3172.t2 VDD.t436 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1144 a_4920_316.t4 a_4375_1009.t7 a_4802_316.t9 VDD.t683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1145 a_6700_316.t5 a_7112_290.t7 a_6818_316.t3 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1146 a_4920_n416.t0 a_5214_290.t7 VSS.t188 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1147 a_25042_n2632.t0 a_23434_n6195.t6 a_25160_n2632.t0 VDD.t359 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1148 VSS.t99 a_13367_404.t22 a_16455_2659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1149 VDD.t1325 a_22797_1688.t18 a_26940_378.t0 VDD.t1324 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1150 a_25168_3236.t0 a_23442_n327.t7 a_25050_3236.t1 VDD.t1377 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1151 VSS.t158 a_20016_n5465.t22 a_24976_n6196.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1152 a_16464_n4792.t1 a_16167_n4181.t19 a_16227_n4155.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1153 VDD.t1568 a_24748_404.t15 a_26101_1097.t1 VDD.t1567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1154 a_3605_2839.t1 a_3015_3276.t10 VDD.t1501 VDD.t1500 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1155 a_19567_3172.t1 a_16822_1209.t7 VSS.t55 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1156 a_98_n2320.t0 A[2].t14 VDD.t1463 VDD.t1462 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1157 VDD.t582 a_13361_n5466.t18 a_30764_n7736.t7 VDD.t581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1158 VDD.t1465 A[2].t15 a_20027_n8268.t0 VDD.t1464 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1159 VSS.t97 a_704_n5517.t18 a_3258_n4791.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1160 a_5486_2565.t0 a_5222_3148.t8 VSS.t198 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1161 VSS.t177 B[3].t15 a_28945_n5935.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1162 a_22857_1714.t0 a_19826_n3212.t19 VDD.t1044 VDD.t1043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1163 a_26940_378.t1 a_22797_1688.t19 VSS.t168 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1164 VDD.t990 a_16803_n2942.t7 a_18538_n2633.t3 VDD.t989 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1165 VDD.t1469 a_25042_n2632.t7 a_25306_n3215.t2 VDD.t1468 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1166 VDD.t655 B[2].t13 a_13338_5442.t3 VDD.t654 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1167 VDD.t1560 a_13367_404.t23 a_16218_3296.t4 VDD.t1559 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1168 VSS.t202 a_16172_1620.t19 a_20257_n396.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1169 VDD.t1231 a_20016_n5465.t23 a_24622_n5464.t3 VDD.t1230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1170 VDD.t1036 a_4912_n5464.t14 a_6265_n4771.t2 VDD.t1035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1171 a_11763_378.t1 a_7379_5006.t19 VDD.t1124 VDD.t1123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1172 a_25042_378.t1 a_20582_5026.t18 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1173 a_114_n5080.t1 B[0].t15 VDD.t1012 VDD.t1011 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1174 a_23089_n527.t1 a_20582_5026.t19 a_22852_110.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1175 a_25160_n2632.t1 a_23434_n6195.t7 a_25042_n2632.t1 VDD.t360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1176 VDD.t759 a_704_n5517.t19 a_3007_n2504.t4 VDD.t758 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1177 a_19898_n5465.t9 a_20310_n5491.t7 a_20016_n5465.t4 VDD.t958 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1178 a_24740_n6196.t0 a_25034_n5490.t7 VSS.t100 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1179 VSS.t213 a_13968_n7819.t19 a_16464_n4792.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1180 VSS.t164 a_2961_n4180.t19 a_3253_n6395.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1181 a_9567_n5760.t4 a_9512_n4182.t19 VDD.t526 VDD.t525 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1182 VSS.t205 a_29301_n2665.t15 a_32485_160.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1183 VDD.t869 B[1].t14 a_98_n2320.t4 VDD.t868 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1184 VDD.t645 B[2].t14 a_28640_2725.t5 VDD.t644 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1185 a_3597_n2941.t0 a_3007_n2504.t10 VSS.t126 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1186 a_30764_n7736.t6 a_13361_n5466.t19 VDD.t562 VDD.t561 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1187 a_16812_n6196.t1 a_16222_n5759.t10 VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1188 VSS.t211 a_2969_1600.t19 a_3261_n615.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1189 VDD.t1097 a_25314_2653.t7 a_26310_3240.t3 VDD.t1096 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1190 a_5214_n2632.t0 a_3606_n6195.t7 VSS.t54 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1191 a_13361_n5466.t4 a_12816_n4773.t7 a_13243_n5466.t2 VDD.t465 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1192 VDD.t863 B[1].t15 a_6789_5443.t1 VDD.t862 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1193 a_25306_n3215.t1 a_25042_n2632.t8 VDD.t1503 VDD.t1502 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1194 a_6810_n5464.t2 a_6265_n4771.t7 a_6692_n5464.t10 VDD.t1156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1195 a_6265_n4771.t3 a_4912_n5464.t15 VDD.t1038 VDD.t1037 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1196 a_28640_2725.t4 B[2].t15 VDD.t647 VDD.t646 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1197 VDD.t1211 a_23425_n2941.t7 a_25160_n2632.t2 VDD.t1210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1198 a_30762_4198.t8 a_31174_4172.t7 Y[2].t5 VDD.t755 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1199 a_5340_3148.t0 a_3605_2839.t7 VDD.t935 VDD.t934 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
R0 a_16213_n2505.n2 a_16213_n2505.t9 214.335
R1 a_16213_n2505.t8 a_16213_n2505.n2 214.335
R2 a_16213_n2505.n3 a_16213_n2505.t8 143.851
R3 a_16213_n2505.n3 a_16213_n2505.t7 135.658
R4 a_16213_n2505.n2 a_16213_n2505.t10 80.333
R5 a_16213_n2505.n4 a_16213_n2505.t2 28.565
R6 a_16213_n2505.n4 a_16213_n2505.t1 28.565
R7 a_16213_n2505.n0 a_16213_n2505.t6 28.565
R8 a_16213_n2505.n0 a_16213_n2505.t4 28.565
R9 a_16213_n2505.t0 a_16213_n2505.n7 28.565
R10 a_16213_n2505.n7 a_16213_n2505.t5 28.565
R11 a_16213_n2505.n1 a_16213_n2505.t3 9.714
R12 a_16213_n2505.n1 a_16213_n2505.n0 1.003
R13 a_16213_n2505.n6 a_16213_n2505.n5 0.833
R14 a_16213_n2505.n5 a_16213_n2505.n4 0.653
R15 a_16213_n2505.n7 a_16213_n2505.n6 0.653
R16 a_16213_n2505.n6 a_16213_n2505.n1 0.341
R17 a_16213_n2505.n5 a_16213_n2505.n3 0.032
R18 VSS.n77 VSS.t165 20.763
R19 VSS.n103 VSS.t57 20.763
R20 VSS.n148 VSS.t14 20.763
R21 VSS.n163 VSS.t122 20.763
R22 VSS.n194 VSS.t13 20.763
R23 VSS.n207 VSS.t77 20.763
R24 VSS.n234 VSS.t105 20.763
R25 VSS.n226 VSS.t159 20.763
R26 VSS.n318 VSS.t129 20.763
R27 VSS.n201 VSS.t195 20.763
R28 VSS.n153 VSS.t162 20.763
R29 VSS.n168 VSS.t17 20.763
R30 VSS.n74 VSS.t108 20.763
R31 VSS.n93 VSS.t104 20.763
R32 VSS.n260 VSS.t168 20.763
R33 VSS.n280 VSS.t62 20.763
R34 VSS.n78 VSS.t74 20.606
R35 VSS.n104 VSS.t136 20.606
R36 VSS.n149 VSS.t31 20.606
R37 VSS.n164 VSS.t63 20.606
R38 VSS.n195 VSS.t212 20.606
R39 VSS.n208 VSS.t207 20.606
R40 VSS.n235 VSS.t88 20.606
R41 VSS.n227 VSS.t39 20.606
R42 VSS.n319 VSS.t117 20.606
R43 VSS.n202 VSS.t5 20.606
R44 VSS.n154 VSS.t84 20.606
R45 VSS.n169 VSS.t144 20.606
R46 VSS.n75 VSS.t6 20.606
R47 VSS.n94 VSS.t142 20.606
R48 VSS.n261 VSS.t27 20.606
R49 VSS.n281 VSS.t70 20.606
R50 VSS.n243 VSS.t69 20.5
R51 VSS.n250 VSS.t152 20.5
R52 VSS.n248 VSS.t178 20.5
R53 VSS.n246 VSS.t138 20.5
R54 VSS.n244 VSS.t98 20.224
R55 VSS.n256 VSS.t193 20.223
R56 VSS.n256 VSS.t204 20.223
R57 VSS.n256 VSS.t0 20.223
R58 VSS.n57 VSS.t19 18.185
R59 VSS.n133 VSS.t43 18.185
R60 VSS.n284 VSS.t201 18.185
R61 VSS.n51 VSS.t124 18.185
R62 VSS.n224 VSS.t52 18.185
R63 VSS.n113 VSS.t47 18.185
R64 VSS.n69 VSS.t197 18.185
R65 VSS.n297 VSS.t163 18.185
R66 VSS.n122 VSS.t126 18.185
R67 VSS.n45 VSS.t160 18.185
R68 VSS.n107 VSS.t23 18.185
R69 VSS.n219 VSS.t1 18.185
R70 VSS.n117 VSS.t53 18.185
R71 VSS.n213 VSS.t51 18.185
R72 VSS.n39 VSS.t85 18.185
R73 VSS.n119 VSS.t185 18.185
R74 VSS.n292 VSS.t172 18.185
R75 VSS.n63 VSS.t9 18.185
R76 VSS.n10 VSS.t109 18.185
R77 VSS.n188 VSS.t29 18.185
R78 VSS.n181 VSS.t68 18.185
R79 VSS.n17 VSS.t22 18.185
R80 VSS.n174 VSS.t135 18.185
R81 VSS.n1 VSS.t95 18.185
R82 VSS.n170 VSS.t2 18.178
R83 VSS.n211 VSS.t34 18.178
R84 VSS.n257 VSS.t182 18.178
R85 VSS.n241 VSS.t67 18.178
R86 VSS.n251 VSS.t42 18.178
R87 VSS.n239 VSS.t75 18.178
R88 VSS.n129 VSS.t10 18.178
R89 VSS.n128 VSS.t175 18.178
R90 VSS.n252 VSS.t28 18.178
R91 VSS.n240 VSS.t183 18.178
R92 VSS.n238 VSS.t26 18.178
R93 VSS.n253 VSS.t173 18.178
R94 VSS.n127 VSS.t191 18.178
R95 VSS.n237 VSS.t114 18.178
R96 VSS.n126 VSS.t149 18.178
R97 VSS.n254 VSS.t4 18.178
R98 VSS.n144 VSS.t128 18.178
R99 VSS.n299 VSS.t200 18.176
R100 VSS.n171 VSS.t120 18.176
R101 VSS.n143 VSS.t174 18.176
R102 VSS.n87 VSS.t15 17.929
R103 VSS.n25 VSS.t37 17.929
R104 VSS.n307 VSS.t132 17.929
R105 VSS.n269 VSS.t134 17.929
R106 VSS.n30 VSS.t80 17.929
R107 VSS.n82 VSS.t190 17.929
R108 VSS.n302 VSS.t55 17.929
R109 VSS.n264 VSS.t35 17.929
R110 VSS.n197 VSS.t131 17.925
R111 VSS.n230 VSS.t111 17.925
R112 VSS.n101 VSS.t54 17.925
R113 VSS.n151 VSS.t36 17.925
R114 VSS.n34 VSS.t125 17.925
R115 VSS.n97 VSS.t24 17.925
R116 VSS.n313 VSS.t184 17.925
R117 VSS.n275 VSS.t215 17.925
R118 VSS.n86 VSS.t214 17.4
R119 VSS.n86 VSS.t156 17.4
R120 VSS.n24 VSS.t38 17.4
R121 VSS.n24 VSS.t148 17.4
R122 VSS.n196 VSS.t61 17.4
R123 VSS.n196 VSS.t203 17.4
R124 VSS.n229 VSS.t187 17.4
R125 VSS.n229 VSS.t153 17.4
R126 VSS.n306 VSS.t102 17.4
R127 VSS.n306 VSS.t30 17.4
R128 VSS.n100 VSS.t64 17.4
R129 VSS.n100 VSS.t155 17.4
R130 VSS.n150 VSS.t130 17.4
R131 VSS.n150 VSS.t66 17.4
R132 VSS.n268 VSS.t154 17.4
R133 VSS.n268 VSS.t107 17.4
R134 VSS.n33 VSS.t119 17.4
R135 VSS.n33 VSS.t89 17.4
R136 VSS.n29 VSS.t41 17.4
R137 VSS.n29 VSS.t186 17.4
R138 VSS.n96 VSS.t198 17.4
R139 VSS.n96 VSS.t7 17.4
R140 VSS.n81 VSS.t192 17.4
R141 VSS.n81 VSS.t93 17.4
R142 VSS.n312 VSS.t49 17.4
R143 VSS.n312 VSS.t167 17.4
R144 VSS.n301 VSS.t60 17.4
R145 VSS.n301 VSS.t209 17.4
R146 VSS.n274 VSS.t56 17.4
R147 VSS.n274 VSS.t171 17.4
R148 VSS.n263 VSS.t65 17.4
R149 VSS.n263 VSS.t141 17.4
R150 VSS.n57 VSS.t151 9.568
R151 VSS.n133 VSS.t164 9.568
R152 VSS.n284 VSS.t121 9.568
R153 VSS.n51 VSS.t189 9.568
R154 VSS.n224 VSS.t40 9.568
R155 VSS.n113 VSS.t97 9.568
R156 VSS.n69 VSS.t48 9.568
R157 VSS.n297 VSS.t91 9.568
R158 VSS.n122 VSS.t137 9.568
R159 VSS.n45 VSS.t145 9.568
R160 VSS.n107 VSS.t211 9.568
R161 VSS.n219 VSS.t169 9.568
R162 VSS.n117 VSS.t127 9.568
R163 VSS.n213 VSS.t71 9.568
R164 VSS.n39 VSS.t123 9.568
R165 VSS.n119 VSS.t101 9.568
R166 VSS.n292 VSS.t72 9.568
R167 VSS.n63 VSS.t82 9.568
R168 VSS.n10 VSS.t79 9.568
R169 VSS.n188 VSS.t206 9.568
R170 VSS.n181 VSS.t213 9.568
R171 VSS.n17 VSS.t76 9.568
R172 VSS.n174 VSS.t99 9.568
R173 VSS.n1 VSS.t116 9.568
R174 VSS.n170 VSS.t83 9.319
R175 VSS.n211 VSS.t106 9.319
R176 VSS.n257 VSS.t181 9.319
R177 VSS.n241 VSS.t179 9.319
R178 VSS.n251 VSS.t73 9.319
R179 VSS.n239 VSS.t177 9.319
R180 VSS.n129 VSS.t21 9.319
R181 VSS.n128 VSS.t110 9.319
R182 VSS.n252 VSS.t194 9.319
R183 VSS.n240 VSS.t180 9.319
R184 VSS.n238 VSS.t78 9.319
R185 VSS.n253 VSS.t205 9.319
R186 VSS.n127 VSS.t133 9.319
R187 VSS.n237 VSS.t92 9.319
R188 VSS.n126 VSS.t113 9.319
R189 VSS.n254 VSS.t208 9.319
R190 VSS.n144 VSS.t20 9.319
R191 VSS.n299 VSS.t46 9.317
R192 VSS.n171 VSS.t3 9.317
R193 VSS.n143 VSS.t25 9.317
R194 VSS.n137 VSS.n131 9.041
R195 VSS.n132 VSS.n131 9
R196 VSS.n242 VSS.t150 8.7
R197 VSS.n242 VSS.t94 8.7
R198 VSS.n76 VSS.t199 8.7
R199 VSS.n76 VSS.t166 8.7
R200 VSS.n102 VSS.t81 8.7
R201 VSS.n102 VSS.t18 8.7
R202 VSS.n147 VSS.t147 8.7
R203 VSS.n147 VSS.t146 8.7
R204 VSS.n162 VSS.t112 8.7
R205 VSS.n162 VSS.t45 8.7
R206 VSS.n193 VSS.t8 8.7
R207 VSS.n193 VSS.t118 8.7
R208 VSS.n206 VSS.t58 8.7
R209 VSS.n206 VSS.t16 8.7
R210 VSS.n233 VSS.t90 8.7
R211 VSS.n233 VSS.t115 8.7
R212 VSS.n225 VSS.t100 8.7
R213 VSS.n225 VSS.t158 8.7
R214 VSS.n249 VSS.t176 8.7
R215 VSS.n249 VSS.t86 8.7
R216 VSS.n317 VSS.t143 8.7
R217 VSS.n317 VSS.t50 8.7
R218 VSS.n200 VSS.t59 8.7
R219 VSS.n200 VSS.t202 8.7
R220 VSS.n152 VSS.t33 8.7
R221 VSS.n152 VSS.t161 8.7
R222 VSS.n167 VSS.t157 8.7
R223 VSS.n167 VSS.t140 8.7
R224 VSS.n73 VSS.t44 8.7
R225 VSS.n73 VSS.t210 8.7
R226 VSS.n92 VSS.t188 8.7
R227 VSS.n92 VSS.t103 8.7
R228 VSS.n247 VSS.t11 8.7
R229 VSS.n247 VSS.t32 8.7
R230 VSS.n259 VSS.t196 8.7
R231 VSS.n259 VSS.t170 8.7
R232 VSS.n279 VSS.t87 8.7
R233 VSS.n279 VSS.t12 8.7
R234 VSS.n245 VSS.t96 8.7
R235 VSS.n245 VSS.t139 8.7
R236 VSS.n166 VSS.n165 3.487
R237 VSS.n47 VSS.n43 3.483
R238 VSS.n109 VSS.n105 3.482
R239 VSS.n41 VSS.n37 3.481
R240 VSS.n53 VSS.n49 3.481
R241 VSS.n65 VSS.n61 3.48
R242 VSS.n115 VSS.n111 3.48
R243 VSS.n60 VSS.n59 3.466
R244 VSS.n125 VSS.n124 3.462
R245 VSS.n72 VSS.n71 3.458
R246 VSS.n132 VSS.n118 3.445
R247 VSS.n161 VSS.n160 3.435
R248 VSS.n35 VSS.n32 3.42
R249 VSS.n98 VSS.n95 3.42
R250 VSS.n159 VSS.n31 3.416
R251 VSS.n83 VSS.n80 3.416
R252 VSS.n146 VSS.n60 3.414
R253 VSS.n146 VSS.n72 3.414
R254 VSS.n138 VSS.n125 3.414
R255 VSS.n88 VSS.n85 3.41
R256 VSS.n27 VSS.n26 3.41
R257 VSS.n77 VSS.n76 0.948
R258 VSS.n103 VSS.n102 0.948
R259 VSS.n148 VSS.n147 0.948
R260 VSS.n163 VSS.n162 0.948
R261 VSS.n194 VSS.n193 0.948
R262 VSS.n207 VSS.n206 0.948
R263 VSS.n234 VSS.n233 0.948
R264 VSS.n226 VSS.n225 0.948
R265 VSS.n318 VSS.n317 0.948
R266 VSS.n201 VSS.n200 0.948
R267 VSS.n153 VSS.n152 0.948
R268 VSS.n168 VSS.n167 0.948
R269 VSS.n74 VSS.n73 0.948
R270 VSS.n93 VSS.n92 0.948
R271 VSS.n260 VSS.n259 0.948
R272 VSS.n280 VSS.n279 0.948
R273 VSS.n243 VSS.n242 0.889
R274 VSS.n250 VSS.n249 0.889
R275 VSS.n248 VSS.n247 0.889
R276 VSS.n246 VSS.n245 0.889
R277 VSS.n87 VSS.n86 0.72
R278 VSS.n25 VSS.n24 0.72
R279 VSS.n197 VSS.n196 0.72
R280 VSS.n230 VSS.n229 0.72
R281 VSS.n307 VSS.n306 0.72
R282 VSS.n101 VSS.n100 0.72
R283 VSS.n151 VSS.n150 0.72
R284 VSS.n269 VSS.n268 0.72
R285 VSS.n34 VSS.n33 0.72
R286 VSS.n30 VSS.n29 0.72
R287 VSS.n97 VSS.n96 0.72
R288 VSS.n82 VSS.n81 0.72
R289 VSS.n313 VSS.n312 0.72
R290 VSS.n302 VSS.n301 0.72
R291 VSS.n275 VSS.n274 0.72
R292 VSS.n264 VSS.n263 0.72
R293 VSS.n157 VSS.n156 0.439
R294 VSS.n156 VSS.n21 0.416
R295 VSS.n85 VSS.n79 0.395
R296 VSS.n172 VSS.n27 0.395
R297 VSS.n142 VSS.n141 0.393
R298 VSS.n141 VSS.n91 0.385
R299 VSS.n157 VSS.n22 0.38
R300 VSS.n139 VSS.n91 0.38
R301 VSS.n139 VSS.n79 0.375
R302 VSS.n172 VSS.n22 0.365
R303 VSS.n138 VSS.n137 0.357
R304 VSS.n146 VSS.n49 0.322
R305 VSS.n138 VSS.n111 0.322
R306 VSS.n146 VSS.n43 0.322
R307 VSS.n138 VSS.n105 0.322
R308 VSS.n146 VSS.n37 0.322
R309 VSS.n146 VSS.n61 0.322
R310 VSS.n300 VSS.n299 0.311
R311 VSS.n172 VSS.n171 0.311
R312 VSS.n145 VSS.n143 0.311
R313 VSS.n172 VSS.n170 0.309
R314 VSS.n300 VSS.n211 0.309
R315 VSS.n258 VSS.n257 0.309
R316 VSS.n258 VSS.n241 0.309
R317 VSS.n255 VSS.n251 0.309
R318 VSS.n258 VSS.n239 0.309
R319 VSS.n130 VSS.n129 0.309
R320 VSS.n130 VSS.n128 0.309
R321 VSS.n255 VSS.n252 0.309
R322 VSS.n258 VSS.n240 0.309
R323 VSS.n258 VSS.n238 0.309
R324 VSS.n255 VSS.n253 0.309
R325 VSS.n130 VSS.n127 0.309
R326 VSS.n258 VSS.n237 0.309
R327 VSS.n130 VSS.n126 0.309
R328 VSS.n255 VSS.n254 0.309
R329 VSS.n145 VSS.n144 0.309
R330 VSS.n172 VSS.n159 0.191
R331 VSS.n80 VSS.n79 0.191
R332 VSS.n236 VSS.n235 0.147
R333 VSS.n79 VSS.n78 0.146
R334 VSS.n165 VSS.n164 0.146
R335 VSS.n209 VSS.n208 0.146
R336 VSS.n300 VSS.n202 0.146
R337 VSS.n172 VSS.n169 0.146
R338 VSS.n145 VSS.n75 0.146
R339 VSS.n262 VSS.n261 0.146
R340 VSS.n140 VSS.n104 0.142
R341 VSS.n155 VSS.n149 0.142
R342 VSS.n321 VSS.n195 0.142
R343 VSS.n155 VSS.n154 0.142
R344 VSS.n282 VSS.n281 0.142
R345 VSS.n26 VSS.n25 0.141
R346 VSS.n321 VSS.n319 0.141
R347 VSS.n282 VSS.n227 0.14
R348 VSS.n140 VSS.n94 0.14
R349 VSS.n88 VSS.n87 0.138
R350 VSS.n265 VSS.n264 0.138
R351 VSS.n270 VSS.n269 0.137
R352 VSS.n31 VSS.n30 0.137
R353 VSS.n155 VSS.n151 0.136
R354 VSS.n83 VSS.n82 0.136
R355 VSS.n140 VSS.n101 0.135
R356 VSS.n276 VSS.n275 0.135
R357 VSS.n321 VSS.n197 0.134
R358 VSS.n282 VSS.n230 0.133
R359 VSS.n308 VSS.n307 0.133
R360 VSS.n98 VSS.n97 0.133
R361 VSS.n303 VSS.n302 0.133
R362 VSS.n314 VSS.n313 0.131
R363 VSS.n35 VSS.n34 0.129
R364 VSS.n78 VSS.n77 0.125
R365 VSS.n104 VSS.n103 0.125
R366 VSS.n149 VSS.n148 0.125
R367 VSS.n164 VSS.n163 0.125
R368 VSS.n195 VSS.n194 0.125
R369 VSS.n208 VSS.n207 0.125
R370 VSS.n235 VSS.n234 0.125
R371 VSS.n227 VSS.n226 0.125
R372 VSS.n319 VSS.n318 0.125
R373 VSS.n202 VSS.n201 0.125
R374 VSS.n154 VSS.n153 0.125
R375 VSS.n169 VSS.n168 0.125
R376 VSS.n75 VSS.n74 0.125
R377 VSS.n94 VSS.n93 0.125
R378 VSS.n261 VSS.n260 0.125
R379 VSS.n281 VSS.n280 0.125
R380 VSS.n298 VSS.n224 0.119
R381 VSS.n138 VSS.n117 0.119
R382 VSS.n18 VSS.n17 0.118
R383 VSS.n138 VSS.n119 0.118
R384 VSS.n298 VSS.n297 0.117
R385 VSS.n46 VSS.n45 0.116
R386 VSS.n108 VSS.n107 0.116
R387 VSS.n189 VSS.n188 0.116
R388 VSS.n2 VSS.n1 0.116
R389 VSS.n220 VSS.n219 0.115
R390 VSS.n40 VSS.n39 0.115
R391 VSS.n52 VSS.n51 0.114
R392 VSS.n293 VSS.n292 0.114
R393 VSS.n182 VSS.n181 0.114
R394 VSS.n134 VSS.n133 0.113
R395 VSS.n285 VSS.n284 0.113
R396 VSS.n70 VSS.n69 0.113
R397 VSS.n123 VSS.n122 0.113
R398 VSS.n64 VSS.n63 0.113
R399 VSS.n11 VSS.n10 0.112
R400 VSS.n58 VSS.n57 0.111
R401 VSS.n175 VSS.n174 0.111
R402 VSS.n114 VSS.n113 0.11
R403 VSS.n214 VSS.n213 0.11
R404 VSS.n256 VSS.n250 0.062
R405 VSS.n256 VSS.n248 0.062
R406 VSS.n256 VSS.n246 0.062
R407 VSS.n244 VSS.n243 0.061
R408 VSS.n134 VSS.n132 0.04
R409 VSS.n293 VSS.n291 0.04
R410 VSS.n172 VSS.n21 0.028
R411 VSS.n141 VSS.n140 0.023
R412 VSS.n321 VSS.n316 0.022
R413 VSS.n155 VSS.n22 0.022
R414 VSS.n282 VSS.n278 0.022
R415 VSS.n282 VSS.n228 0.022
R416 VSS.n140 VSS.n139 0.022
R417 VSS.n60 VSS.n56 0.018
R418 VSS.n287 VSS.n286 0.018
R419 VSS.n72 VSS.n68 0.018
R420 VSS.n125 VSS.n121 0.018
R421 VSS.n13 VSS.n12 0.018
R422 VSS.n191 VSS.n190 0.018
R423 VSS.n184 VSS.n183 0.018
R424 VSS.n16 VSS.n15 0.018
R425 VSS.n177 VSS.n176 0.018
R426 VSS.n4 VSS.n3 0.018
R427 VSS.n116 VSS.n115 0.014
R428 VSS.n59 VSS.n55 0.013
R429 VSS.n71 VSS.n67 0.012
R430 VSS.n124 VSS.n120 0.012
R431 VSS.n161 VSS.n21 0.012
R432 VSS.n204 VSS.n203 0.012
R433 VSS.n90 VSS.n85 0.011
R434 VSS.n158 VSS.n27 0.011
R435 VSS.n310 VSS.n305 0.011
R436 VSS.n272 VSS.n267 0.011
R437 VSS.n66 VSS.n65 0.011
R438 VSS.n287 VSS.n285 0.01
R439 VSS.n70 VSS.n68 0.01
R440 VSS.n54 VSS.n53 0.01
R441 VSS.n42 VSS.n41 0.009
R442 VSS.n110 VSS.n109 0.008
R443 VSS.n48 VSS.n47 0.008
R444 VSS.n222 VSS.n220 0.007
R445 VSS.n114 VSS.n112 0.006
R446 VSS.n123 VSS.n121 0.006
R447 VSS.n216 VSS.n214 0.006
R448 VSS.n272 VSS.n232 0.006
R449 VSS.n310 VSS.n199 0.006
R450 VSS.n90 VSS.n80 0.006
R451 VSS.n159 VSS.n158 0.006
R452 VSS.n20 VSS.n19 0.006
R453 VSS.n89 VSS.n88 0.005
R454 VSS.n26 VSS.n23 0.005
R455 VSS.n271 VSS.n270 0.005
R456 VSS.n309 VSS.n308 0.005
R457 VSS.n52 VSS.n50 0.005
R458 VSS.n40 VSS.n38 0.005
R459 VSS.n64 VSS.n62 0.005
R460 VSS.n13 VSS.n11 0.005
R461 VSS.n191 VSS.n189 0.005
R462 VSS.n300 VSS.n298 0.005
R463 VSS.n146 VSS.n145 0.005
R464 VSS.n138 VSS.n130 0.005
R465 VSS.n166 VSS.n161 0.004
R466 VSS.n108 VSS.n106 0.004
R467 VSS.n184 VSS.n182 0.004
R468 VSS.n177 VSS.n175 0.004
R469 VSS.n304 VSS.n303 0.004
R470 VSS.n99 VSS.n98 0.004
R471 VSS.n84 VSS.n83 0.004
R472 VSS.n266 VSS.n265 0.004
R473 VSS.n31 VSS.n28 0.004
R474 VSS.n36 VSS.n35 0.004
R475 VSS.n315 VSS.n314 0.004
R476 VSS.n277 VSS.n276 0.004
R477 VSS.n262 VSS.n236 0.003
R478 VSS.n205 VSS.n204 0.003
R479 VSS.n46 VSS.n44 0.003
R480 VSS.n4 VSS.n2 0.003
R481 VSS.n258 VSS.n256 0.003
R482 VSS.n262 VSS.n258 0.003
R483 VSS VSS.n172 0.003
R484 VSS.n140 VSS.n95 0.003
R485 VSS.n155 VSS.n32 0.003
R486 VSS.n50 VSS.n49 0.003
R487 VSS.n112 VSS.n111 0.003
R488 VSS.n44 VSS.n43 0.003
R489 VSS.n106 VSS.n105 0.003
R490 VSS.n222 VSS.n221 0.003
R491 VSS.n216 VSS.n215 0.003
R492 VSS.n38 VSS.n37 0.003
R493 VSS.n135 VSS.n134 0.003
R494 VSS.n142 VSS.n79 0.002
R495 VSS.n62 VSS.n61 0.002
R496 VSS.n58 VSS.n56 0.002
R497 VSS.n256 VSS.n255 0.002
R498 VSS.n298 VSS.n282 0.002
R499 VSS VSS.n321 0.002
R500 VSS.n155 VSS.n146 0.002
R501 VSS.n140 VSS.n138 0.002
R502 VSS.n294 VSS.n293 0.002
R503 VSS VSS.n8 0.002
R504 VSS VSS.n186 0.002
R505 VSS VSS.n179 0.002
R506 VSS.n146 VSS.n67 0.001
R507 VSS.n68 VSS.n67 0.001
R508 VSS.n138 VSS.n120 0.001
R509 VSS.n121 VSS.n120 0.001
R510 VSS.n321 VSS.n320 0.001
R511 VSS.n156 VSS.n155 0.001
R512 VSS.n256 VSS.n244 0.001
R513 VSS VSS.n5 0.001
R514 VSS.n273 VSS.n272 0.001
R515 VSS.n311 VSS.n310 0.001
R516 VSS.n158 VSS.n157 0.001
R517 VSS.n91 VSS.n90 0.001
R518 VSS.n136 VSS.n118 0.001
R519 VSS.n138 VSS.n118 0.001
R520 VSS.n146 VSS.n55 0.001
R521 VSS.n56 VSS.n55 0.001
R522 VSS.n298 VSS.n288 0.001
R523 VSS.n288 VSS.n287 0.001
R524 VSS.n157 VSS.n32 0.001
R525 VSS.n95 VSS.n91 0.001
R526 VSS.n311 VSS.n198 0.001
R527 VSS.n273 VSS.n231 0.001
R528 VSS VSS.n6 0.001
R529 VSS VSS.n7 0.001
R530 VSS.n145 VSS.n142 0.001
R531 VSS.n137 VSS.n136 0.001
R532 VSS.n295 VSS.n289 0.001
R533 VSS.n300 VSS.n205 0.001
R534 VSS.n115 VSS.n114 0.001
R535 VSS.n214 VSS.n212 0.001
R536 VSS.n59 VSS.n58 0.001
R537 VSS.n175 VSS.n173 0.001
R538 VSS.n11 VSS.n9 0.001
R539 VSS.n124 VSS.n123 0.001
R540 VSS.n65 VSS.n64 0.001
R541 VSS.n285 VSS.n283 0.001
R542 VSS.n71 VSS.n70 0.001
R543 VSS.n182 VSS.n180 0.001
R544 VSS.n53 VSS.n52 0.001
R545 VSS.n41 VSS.n40 0.001
R546 VSS.n220 VSS.n218 0.001
R547 VSS.n47 VSS.n46 0.001
R548 VSS.n2 VSS.n0 0.001
R549 VSS.n109 VSS.n108 0.001
R550 VSS.n189 VSS.n187 0.001
R551 VSS.n19 VSS.n18 0.001
R552 VSS.n172 VSS.n166 0.001
R553 VSS.n135 VSS.n131 0.001
R554 VSS.n136 VSS.n135 0.001
R555 VSS.n165 VSS.n160 0.001
R556 VSS.n172 VSS.n160 0.001
R557 VSS.n210 VSS.n209 0.001
R558 VSS.n300 VSS.n210 0.001
R559 VSS.n146 VSS.n54 0.001
R560 VSS.n138 VSS.n116 0.001
R561 VSS.n89 VSS.n79 0.001
R562 VSS.n172 VSS.n23 0.001
R563 VSS.n146 VSS.n48 0.001
R564 VSS.n138 VSS.n110 0.001
R565 VSS.n298 VSS.n223 0.001
R566 VSS.n298 VSS.n217 0.001
R567 VSS.n146 VSS.n42 0.001
R568 VSS.n157 VSS.n36 0.001
R569 VSS.n172 VSS.n28 0.001
R570 VSS.n99 VSS.n91 0.001
R571 VSS.n84 VSS.n79 0.001
R572 VSS.n315 VSS.n311 0.001
R573 VSS.n304 VSS.n300 0.001
R574 VSS.n277 VSS.n273 0.001
R575 VSS.n266 VSS.n262 0.001
R576 VSS.n294 VSS.n290 0.001
R577 VSS.n296 VSS.n295 0.001
R578 VSS.n295 VSS.n294 0.001
R579 VSS.n146 VSS.n66 0.001
R580 VSS VSS.n14 0.001
R581 VSS VSS.n192 0.001
R582 VSS VSS.n185 0.001
R583 VSS VSS.n20 0.001
R584 VSS VSS.n178 0.001
R585 VSS.n322 VSS 0.001
R586 VSS.n282 VSS.n277 0.001
R587 VSS.n321 VSS.n315 0.001
R588 VSS.n155 VSS.n36 0.001
R589 VSS.n140 VSS.n99 0.001
R590 VSS.n66 VSS.n62 0.001
R591 VSS.n298 VSS.n296 0.001
R592 VSS.n272 VSS.n266 0.001
R593 VSS.n310 VSS.n304 0.001
R594 VSS.n90 VSS.n84 0.001
R595 VSS.n178 VSS.n177 0.001
R596 VSS.n158 VSS.n28 0.001
R597 VSS.n42 VSS.n38 0.001
R598 VSS.n217 VSS.n216 0.001
R599 VSS.n14 VSS.n13 0.001
R600 VSS.n223 VSS.n222 0.001
R601 VSS.n110 VSS.n106 0.001
R602 VSS.n192 VSS.n191 0.001
R603 VSS.n48 VSS.n44 0.001
R604 VSS.n272 VSS.n271 0.001
R605 VSS.n322 VSS.n4 0.001
R606 VSS.n310 VSS.n309 0.001
R607 VSS.n158 VSS.n23 0.001
R608 VSS.n90 VSS.n89 0.001
R609 VSS.n116 VSS.n112 0.001
R610 VSS.n185 VSS.n184 0.001
R611 VSS.n54 VSS.n50 0.001
R612 VSS.n20 VSS.n16 0.001
R613 a_16803_n2942.t5 a_16803_n2942.t4 800.071
R614 a_16803_n2942.n2 a_16803_n2942.n1 659.097
R615 a_16803_n2942.n0 a_16803_n2942.t7 285.109
R616 a_16803_n2942.n1 a_16803_n2942.t5 193.602
R617 a_16803_n2942.n4 a_16803_n2942.n3 192.754
R618 a_16803_n2942.n0 a_16803_n2942.t6 160.666
R619 a_16803_n2942.n1 a_16803_n2942.n0 91.507
R620 a_16803_n2942.n3 a_16803_n2942.t1 28.568
R621 a_16803_n2942.t0 a_16803_n2942.n4 28.565
R622 a_16803_n2942.n4 a_16803_n2942.t2 28.565
R623 a_16803_n2942.n2 a_16803_n2942.t3 19.061
R624 a_16803_n2942.n3 a_16803_n2942.n2 1.005
R625 a_6818_316.n0 a_6818_316.t2 14.282
R626 a_6818_316.t1 a_6818_316.n0 14.282
R627 a_6818_316.n0 a_6818_316.n14 90.436
R628 a_6818_316.n10 a_6818_316.n13 50.575
R629 a_6818_316.n14 a_6818_316.n10 74.302
R630 a_6818_316.n13 a_6818_316.n12 157.665
R631 a_6818_316.n12 a_6818_316.t6 8.7
R632 a_6818_316.n12 a_6818_316.t0 8.7
R633 a_6818_316.n13 a_6818_316.n11 122.999
R634 a_6818_316.n11 a_6818_316.t7 14.282
R635 a_6818_316.n11 a_6818_316.t5 14.282
R636 a_6818_316.n10 a_6818_316.n9 90.416
R637 a_6818_316.n9 a_6818_316.t4 14.282
R638 a_6818_316.n9 a_6818_316.t3 14.282
R639 a_6818_316.n1 a_6818_316.t12 220.285
R640 a_6818_316.n14 a_6818_316.n1 3509.5
R641 a_6818_316.n1 a_6818_316.n8 61.538
R642 a_6818_316.n8 a_6818_316.n3 465.933
R643 a_6818_316.n8 a_6818_316.n7 163.88
R644 a_6818_316.n7 a_6818_316.n6 6.615
R645 a_6818_316.n6 a_6818_316.t11 93.989
R646 a_6818_316.n7 a_6818_316.n5 97.816
R647 a_6818_316.n5 a_6818_316.t15 80.333
R648 a_6818_316.n5 a_6818_316.t9 394.151
R649 a_6818_316.t9 a_6818_316.n4 269.523
R650 a_6818_316.n4 a_6818_316.t17 160.666
R651 a_6818_316.n4 a_6818_316.t14 269.523
R652 a_6818_316.n6 a_6818_316.t16 198.043
R653 a_6818_316.n3 a_6818_316.t19 294.653
R654 a_6818_316.n3 a_6818_316.t18 111.663
R655 a_6818_316.t12 a_6818_316.t8 415.315
R656 a_6818_316.t8 a_6818_316.n2 214.335
R657 a_6818_316.n2 a_6818_316.t13 80.333
R658 a_6818_316.n2 a_6818_316.t10 214.335
R659 a_32246_4888.n0 a_32246_4888.t8 214.335
R660 a_32246_4888.t10 a_32246_4888.n0 214.335
R661 a_32246_4888.n1 a_32246_4888.t10 143.851
R662 a_32246_4888.n1 a_32246_4888.t7 135.658
R663 a_32246_4888.n0 a_32246_4888.t9 80.333
R664 a_32246_4888.n2 a_32246_4888.t4 28.565
R665 a_32246_4888.n2 a_32246_4888.t3 28.565
R666 a_32246_4888.n4 a_32246_4888.t2 28.565
R667 a_32246_4888.n4 a_32246_4888.t6 28.565
R668 a_32246_4888.t0 a_32246_4888.n7 28.565
R669 a_32246_4888.n7 a_32246_4888.t5 28.565
R670 a_32246_4888.n6 a_32246_4888.t1 9.714
R671 a_32246_4888.n7 a_32246_4888.n6 1.003
R672 a_32246_4888.n5 a_32246_4888.n3 0.833
R673 a_32246_4888.n3 a_32246_4888.n2 0.653
R674 a_32246_4888.n5 a_32246_4888.n4 0.653
R675 a_32246_4888.n6 a_32246_4888.n5 0.341
R676 a_32246_4888.n3 a_32246_4888.n1 0.032
R677 VDD.t71 VDD.t304 2079.61
R678 VDD.t6 VDD.t795 2079.61
R679 VDD.t1119 VDD.t1275 2079.61
R680 VDD.t341 VDD.t20 2079.61
R681 VDD.t449 VDD.t1115 2079.61
R682 VDD.t102 VDD.t1435 2079.61
R683 VDD.t276 VDD.t472 2079.61
R684 VDD.t1232 VDD.t1230 2079.61
R685 VDD.n138 VDD.n137 1412.62
R686 VDD.n749 VDD.n748 1412.62
R687 VDD.n332 VDD.n331 1412.59
R688 VDD.n533 VDD.n521 1408.41
R689 VDD.n815 VDD.n814 1404.25
R690 VDD.n271 VDD.n270 1239.11
R691 VDD.n661 VDD.n660 1235.85
R692 VDD.n203 VDD.n202 1235.85
R693 VDD.n641 VDD.n635 1033.13
R694 VDD.n499 VDD.n498 1033.13
R695 VDD.n717 VDD.n716 1033.13
R696 VDD.n760 VDD.n754 1033.13
R697 VDD.n172 VDD.n168 1033.13
R698 VDD.n837 VDD.n831 1033.12
R699 VDD.n626 VDD.n622 1029.22
R700 VDD.n229 VDD.n225 1029.22
R701 VDD.n112 VDD.n111 1029.21
R702 VDD.n958 VDD.n957 1029.21
R703 VDD.n297 VDD.n293 1025.3
R704 VDD.n486 VDD.n482 1025.3
R705 VDD.t1567 VDD.t314 999.845
R706 VDD.t760 VDD.t816 999.845
R707 VDD.t1105 VDD.t1123 999.845
R708 VDD.t870 VDD.t1551 999.845
R709 VDD.t1035 VDD.t814 999.845
R710 VDD.t533 VDD.t1626 999.845
R711 VDD.t381 VDD.t197 999.845
R712 VDD.t95 VDD.t1236 999.845
R713 VDD.n182 VDD.n176 880.922
R714 VDD.n704 VDD.n698 874.857
R715 VDD.n100 VDD.n94 874.857
R716 VDD.n786 VDD.n782 874.804
R717 VDD.n1022 VDD.n1016 871.811
R718 VDD.n312 VDD.n306 871.81
R719 VDD.n928 VDD.n927 871.81
R720 VDD.n248 VDD.n243 871.809
R721 VDD.n988 VDD.n987 871.808
R722 VDD.n594 VDD.n593 871.808
R723 VDD.n671 VDD.n670 871.808
R724 VDD.n795 VDD.n794 871.808
R725 VDD.n979 VDD.n978 809.201
R726 VDD.n599 VDD.n598 805.926
R727 VDD.n686 VDD.n685 805.926
R728 VDD.n845 VDD.n844 805.925
R729 VDD.n918 VDD.n917 802.647
R730 VDD.n948 VDD.n947 687.118
R731 VDD.n1010 VDD.n1008 687.068
R732 VDD.n766 VDD.n764 684.693
R733 VDD.n435 VDD.n434 600.209
R734 VDD.n457 VDD.n364 600.209
R735 VDD.n377 VDD.n376 600.207
R736 VDD.n409 VDD.n408 600.207
R737 VDD.n69 VDD.n68 491.958
R738 VDD.n692 VDD.t347 479.007
R739 VDD.n771 VDD.t457 479.007
R740 VDD.n999 VDD.t523 479.006
R741 VDD.n604 VDD.t1543 479.006
R742 VDD.n939 VDD.t246 479.006
R743 VDD.n972 VDD.t324 479.006
R744 VDD.n850 VDD.t878 424.731
R745 VDD.t1334 VDD.t1338 422.41
R746 VDD.t826 VDD.t398 422.41
R747 VDD.t1125 VDD.t499 422.41
R748 VDD.t1557 VDD.t1161 422.41
R749 VDD.t1311 VDD.t1291 422.41
R750 VDD.t379 VDD.t1188 422.41
R751 VDD.t113 VDD.t944 422.41
R752 VDD.t1019 VDD.t801 422.41
R753 VDD.n910 VDD.t1216 422.363
R754 VDD.t720 VDD.t716 394.32
R755 VDD.t964 VDD.t290 394.32
R756 VDD.t1087 VDD.t115 394.32
R757 VDD.t357 VDD.t1198 394.32
R758 VDD.t718 VDD.t551 352.102
R759 VDD.t968 VDD.t1390 352.102
R760 VDD.t1089 VDD.t443 352.102
R761 VDD.t1200 VDD.t672 352.102
R762 VDD.t1157 VDD.t1522 345.987
R763 VDD.t1522 VDD.t1567 345.987
R764 VDD.t314 VDD.t480 345.987
R765 VDD.t480 VDD.t71 345.987
R766 VDD.t1324 VDD.t1344 345.987
R767 VDD.t1338 VDD.t1324 345.987
R768 VDD.t421 VDD.t1063 345.987
R769 VDD.t1061 VDD.t421 345.987
R770 VDD.t86 VDD.t1061 345.987
R771 VDD.t1043 VDD.t86 345.987
R772 VDD.t571 VDD.t1328 345.987
R773 VDD.t1328 VDD.t1326 345.987
R774 VDD.t1326 VDD.t1336 345.987
R775 VDD.t318 VDD.t316 345.987
R776 VDD.t320 VDD.t318 345.987
R777 VDD.t1340 VDD.t320 345.987
R778 VDD.t1332 VDD.t1340 345.987
R779 VDD.t1330 VDD.t300 345.987
R780 VDD.t300 VDD.t850 345.987
R781 VDD.t850 VDD.t478 345.987
R782 VDD.t1289 VDD.t1285 345.987
R783 VDD.t1287 VDD.t1289 345.987
R784 VDD.t387 VDD.t1287 345.987
R785 VDD.t336 VDD.t387 345.987
R786 VDD.t334 VDD.t1242 345.987
R787 VDD.t1242 VDD.t1253 345.987
R788 VDD.t1253 VDD.t1238 345.987
R789 VDD.t732 VDD.t734 345.987
R790 VDD.t736 VDD.t732 345.987
R791 VDD.t36 VDD.t736 345.987
R792 VDD.t34 VDD.t36 345.987
R793 VDD.t32 VDD.t476 345.987
R794 VDD.t476 VDD.t926 345.987
R795 VDD.t926 VDD.t199 345.987
R796 VDD.t543 VDD.t545 345.987
R797 VDD.t1167 VDD.t543 345.987
R798 VDD.t1129 VDD.t1167 345.987
R799 VDD.t282 VDD.t1129 345.987
R800 VDD.t1486 VDD.t1607 345.987
R801 VDD.t1607 VDD.t1605 345.987
R802 VDD.t1605 VDD.t1433 345.987
R803 VDD.t752 VDD.t455 345.987
R804 VDD.t242 VDD.t752 345.987
R805 VDD.t742 VDD.t242 345.987
R806 VDD.t740 VDD.t742 345.987
R807 VDD.t758 VDD.t111 345.987
R808 VDD.t111 VDD.t109 345.987
R809 VDD.t109 VDD.t1127 345.987
R810 VDD.t1364 VDD.t1360 345.987
R811 VDD.t1362 VDD.t1364 345.987
R812 VDD.t146 VDD.t1362 345.987
R813 VDD.t142 VDD.t146 345.987
R814 VDD.t776 VDD.t706 345.987
R815 VDD.t706 VDD.t549 345.987
R816 VDD.t549 VDD.t547 345.987
R817 VDD.t1448 VDD.t1446 345.987
R818 VDD.t1500 VDD.t1448 345.987
R819 VDD.t789 VDD.t1500 345.987
R820 VDD.t1029 VDD.t789 345.987
R821 VDD.t153 VDD.t818 345.987
R822 VDD.t818 VDD.t810 345.987
R823 VDD.t810 VDD.t808 345.987
R824 VDD.t535 VDD.t44 345.987
R825 VDD.t44 VDD.t760 345.987
R826 VDD.t816 VDD.t806 345.987
R827 VDD.t806 VDD.t6 345.987
R828 VDD.t265 VDD.t1478 345.987
R829 VDD.t398 VDD.t265 345.987
R830 VDD.t427 VDD.t425 345.987
R831 VDD.t349 VDD.t427 345.987
R832 VDD.t0 VDD.t349 345.987
R833 VDD.t151 VDD.t0 345.987
R834 VDD.t787 VDD.t263 345.987
R835 VDD.t263 VDD.t1484 345.987
R836 VDD.t1484 VDD.t1482 345.987
R837 VDD.t148 VDD.t161 345.987
R838 VDD.t163 VDD.t148 345.987
R839 VDD.t267 VDD.t163 345.987
R840 VDD.t830 VDD.t267 345.987
R841 VDD.t828 VDD.t797 345.987
R842 VDD.t797 VDD.t8 345.987
R843 VDD.t8 VDD.t791 345.987
R844 VDD.t417 VDD.t48 345.987
R845 VDD.t123 VDD.t417 345.987
R846 VDD.t1005 VDD.t123 345.987
R847 VDD.t976 VDD.t1005 345.987
R848 VDD.t539 VDD.t1271 345.987
R849 VDD.t1271 VDD.t1283 345.987
R850 VDD.t1283 VDD.t1277 345.987
R851 VDD.t1190 VDD.t1194 345.987
R852 VDD.t1194 VDD.t1105 345.987
R853 VDD.t1123 VDD.t1279 345.987
R854 VDD.t1279 VDD.t1119 345.987
R855 VDD.t119 VDD.t501 345.987
R856 VDD.t499 VDD.t119 345.987
R857 VDD.t30 VDD.t666 345.987
R858 VDD.t1149 VDD.t30 345.987
R859 VDD.t585 VDD.t1149 345.987
R860 VDD.t660 VDD.t585 345.987
R861 VDD.t587 VDD.t696 345.987
R862 VDD.t696 VDD.t430 345.987
R863 VDD.t430 VDD.t557 345.987
R864 VDD.t1267 VDD.t1250 345.987
R865 VDD.t1248 VDD.t1267 345.987
R866 VDD.t238 VDD.t1248 345.987
R867 VDD.t1094 VDD.t238 345.987
R868 VDD.t559 VDD.t1269 345.987
R869 VDD.t1269 VDD.t1117 345.987
R870 VDD.t1117 VDD.t1281 345.987
R871 VDD.t1081 VDD.t1079 345.987
R872 VDD.t1103 VDD.t1081 345.987
R873 VDD.t602 VDD.t1103 345.987
R874 VDD.t842 VDD.t602 345.987
R875 VDD.t1559 VDD.t16 345.987
R876 VDD.t16 VDD.t1135 345.987
R877 VDD.t1135 VDD.t345 345.987
R878 VDD.t874 VDD.t953 345.987
R879 VDD.t953 VDD.t870 345.987
R880 VDD.t1551 VDD.t343 345.987
R881 VDD.t343 VDD.t341 345.987
R882 VDD.t187 VDD.t189 345.987
R883 VDD.t1161 VDD.t187 345.987
R884 VDD.t219 VDD.t217 345.987
R885 VDD.t832 VDD.t219 345.987
R886 VDD.t924 VDD.t832 345.987
R887 VDD.t844 VDD.t924 345.987
R888 VDD.t600 VDD.t1530 345.987
R889 VDD.t1530 VDD.t185 345.987
R890 VDD.t185 VDD.t1589 345.987
R891 VDD.t261 VDD.t193 345.987
R892 VDD.t195 VDD.t261 345.987
R893 VDD.t1163 VDD.t195 345.987
R894 VDD.t1587 VDD.t1163 345.987
R895 VDD.t1555 VDD.t1549 345.987
R896 VDD.t1549 VDD.t419 345.987
R897 VDD.t419 VDD.t1041 345.987
R898 VDD.t1352 VDD.t1358 345.987
R899 VDD.t1350 VDD.t1352 345.987
R900 VDD.t84 VDD.t1350 345.987
R901 VDD.t565 VDD.t84 345.987
R902 VDD.t567 VDD.t312 345.987
R903 VDD.t312 VDD.t69 345.987
R904 VDD.t69 VDD.t848 345.987
R905 VDD.t42 VDD.t1037 345.987
R906 VDD.t1037 VDD.t1035 345.987
R907 VDD.t814 VDD.t812 345.987
R908 VDD.t812 VDD.t449 345.987
R909 VDD.t1293 VDD.t1295 345.987
R910 VDD.t1291 VDD.t1293 345.987
R911 VDD.t1613 VDD.t1615 345.987
R912 VDD.t1585 VDD.t1613 345.987
R913 VDD.t738 VDD.t1585 345.987
R914 VDD.t355 VDD.t738 345.987
R915 VDD.t353 VDD.t1303 345.987
R916 VDD.t1303 VDD.t1301 345.987
R917 VDD.t1301 VDD.t1297 345.987
R918 VDD.t59 VDD.t211 345.987
R919 VDD.t57 VDD.t59 345.987
R920 VDD.t1307 VDD.t57 345.987
R921 VDD.t1305 VDD.t1307 345.987
R922 VDD.t1313 VDD.t490 345.987
R923 VDD.t490 VDD.t121 345.987
R924 VDD.t121 VDD.t492 345.987
R925 VDD.t484 VDD.t482 345.987
R926 VDD.t482 VDD.t533 345.987
R927 VDD.t1626 VDD.t1624 345.987
R928 VDD.t1624 VDD.t102 345.987
R929 VDD.t980 VDD.t982 345.987
R930 VDD.t1188 VDD.t980 345.987
R931 VDD.t1145 VDD.t1147 345.987
R932 VDD.t254 VDD.t1145 345.987
R933 VDD.t403 VDD.t254 345.987
R934 VDD.t205 VDD.t403 345.987
R935 VDD.t284 VDD.t676 345.987
R936 VDD.t676 VDD.t972 345.987
R937 VDD.t972 VDD.t970 345.987
R938 VDD.t127 VDD.t132 345.987
R939 VDD.t125 VDD.t127 345.987
R940 VDD.t377 VDD.t125 345.987
R941 VDD.t525 VDD.t377 345.987
R942 VDD.t674 VDD.t593 345.987
R943 VDD.t593 VDD.t591 345.987
R944 VDD.t591 VDD.t710 345.987
R945 VDD.t620 VDD.t383 345.987
R946 VDD.t383 VDD.t381 345.987
R947 VDD.t197 VDD.t82 345.987
R948 VDD.t82 VDD.t276 345.987
R949 VDD.t894 VDD.t892 345.987
R950 VDD.t944 VDD.t894 345.987
R951 VDD.t1055 VDD.t1386 345.987
R952 VDD.t1053 VDD.t1055 345.987
R953 VDD.t63 VDD.t1053 345.987
R954 VDD.t463 VDD.t63 345.987
R955 VDD.t918 VDD.t1169 345.987
R956 VDD.t1169 VDD.t1003 345.987
R957 VDD.t1003 VDD.t1001 345.987
R958 VDD.t140 VDD.t159 345.987
R959 VDD.t138 VDD.t140 345.987
R960 VDD.t860 VDD.t138 345.987
R961 VDD.t858 VDD.t860 345.987
R962 VDD.t946 VDD.t80 345.987
R963 VDD.t80 VDD.t474 345.987
R964 VDD.t474 VDD.t928 345.987
R965 VDD.t99 VDD.t97 345.987
R966 VDD.t97 VDD.t95 345.987
R967 VDD.t1236 VDD.t1234 345.987
R968 VDD.t1234 VDD.t1232 345.987
R969 VDD.t803 VDD.t914 345.987
R970 VDD.t801 VDD.t803 345.987
R971 VDD.t1057 VDD.t1059 345.987
R972 VDD.t423 VDD.t1057 345.987
R973 VDD.t38 VDD.t423 345.987
R974 VDD.t330 VDD.t38 345.987
R975 VDD.t326 VDD.t961 345.987
R976 VDD.t961 VDD.t1013 345.987
R977 VDD.t1013 VDD.t799 345.987
R978 VDD.t466 VDD.t468 345.987
R979 VDD.t1553 VDD.t466 345.987
R980 VDD.t912 VDD.t1553 345.987
R981 VDD.t910 VDD.t912 345.987
R982 VDD.t1017 VDD.t1257 345.987
R983 VDD.t1257 VDD.t1261 345.987
R984 VDD.t1261 VDD.t1240 345.987
R985 VDD.n68 VDD.t776 343.055
R986 VDD.t555 VDD.t1157 312.28
R987 VDD.t1093 VDD.t535 312.28
R988 VDD.t1610 VDD.t1190 312.28
R989 VDD.t429 VDD.t874 312.28
R990 VDD.t1156 VDD.t42 312.28
R991 VDD.t465 VDD.t484 312.28
R992 VDD.t1223 VDD.t620 312.28
R993 VDD.t984 VDD.t99 312.28
R994 VDD.n498 VDD.t571 240.432
R995 VDD.n482 VDD.t1330 240.432
R996 VDD.n927 VDD.t334 240.432
R997 VDD.n957 VDD.t32 240.432
R998 VDD.n987 VDD.t1486 240.432
R999 VDD.n1016 VDD.t758 240.432
R1000 VDD.n593 VDD.t153 240.432
R1001 VDD.n635 VDD.t787 240.432
R1002 VDD.n622 VDD.t828 240.432
R1003 VDD.n670 VDD.t539 240.432
R1004 VDD.n716 VDD.t587 240.432
R1005 VDD.n698 VDD.t559 240.432
R1006 VDD.n754 VDD.t1559 240.432
R1007 VDD.n794 VDD.t600 240.432
R1008 VDD.n782 VDD.t1555 240.432
R1009 VDD.n831 VDD.t567 240.432
R1010 VDD.n111 VDD.t353 240.432
R1011 VDD.n94 VDD.t1313 240.432
R1012 VDD.n176 VDD.t284 240.432
R1013 VDD.n168 VDD.t674 240.432
R1014 VDD.n243 VDD.t918 240.432
R1015 VDD.n225 VDD.t946 240.432
R1016 VDD.n306 VDD.t326 240.432
R1017 VDD.n293 VDD.t1017 240.432
R1018 VDD.t10 VDD.t563 218.264
R1019 VDD.t683 VDD.t1113 218.264
R1020 VDD.t715 VDD.t656 218.264
R1021 VDD.t1514 VDD.t920 218.264
R1022 VDD.t705 VDD.t1083 218.264
R1023 VDD.t748 VDD.t405 218.264
R1024 VDD.t489 VDD.t67 218.264
R1025 VDD.t1066 VDD.t40 218.264
R1026 VDD.t563 VDD.t203 213.931
R1027 VDD.t203 VDD.t88 213.931
R1028 VDD.t1212 VDD.t1210 213.931
R1029 VDD.t1210 VDD.t360 213.931
R1030 VDD.t360 VDD.t359 213.931
R1031 VDD.t359 VDD.t885 213.931
R1032 VDD.t822 VDD.t1206 213.931
R1033 VDD.t1206 VDD.t1074 213.931
R1034 VDD.t1074 VDD.t1073 213.931
R1035 VDD.t1073 VDD.t884 213.931
R1036 VDD.t991 VDD.t993 213.931
R1037 VDD.t993 VDD.t497 213.931
R1038 VDD.t497 VDD.t496 213.931
R1039 VDD.t496 VDD.t1048 213.931
R1040 VDD.t215 VDD.t664 213.931
R1041 VDD.t664 VDD.t1068 213.931
R1042 VDD.t1068 VDD.t1067 213.931
R1043 VDD.t1067 VDD.t1070 213.931
R1044 VDD.t1496 VDD.t507 213.931
R1045 VDD.t507 VDD.t725 213.931
R1046 VDD.t725 VDD.t724 213.931
R1047 VDD.t724 VDD.t308 213.931
R1048 VDD.t1139 VDD.t1137 213.931
R1049 VDD.t1137 VDD.t309 213.931
R1050 VDD.t309 VDD.t310 213.931
R1051 VDD.t310 VDD.t311 213.931
R1052 VDD.t1226 VDD.t1228 213.931
R1053 VDD.t1228 VDD.t435 213.931
R1054 VDD.t435 VDD.t438 213.931
R1055 VDD.t438 VDD.t437 213.931
R1056 VDD.t1244 VDD.t1265 213.931
R1057 VDD.t1265 VDD.t108 213.931
R1058 VDD.t108 VDD.t1108 213.931
R1059 VDD.t1108 VDD.t1107 213.931
R1060 VDD.t934 VDD.t295 213.931
R1061 VDD.t295 VDD.t165 213.931
R1062 VDD.t165 VDD.t150 213.931
R1063 VDD.t150 VDD.t166 213.931
R1064 VDD.t999 VDD.t712 213.931
R1065 VDD.t712 VDD.t1505 213.931
R1066 VDD.t1505 VDD.t498 213.931
R1067 VDD.t498 VDD.t1504 213.931
R1068 VDD.t1113 VDD.t1031 213.931
R1069 VDD.t1031 VDD.t1109 213.931
R1070 VDD.t681 VDD.t1603 213.931
R1071 VDD.t1603 VDD.t995 213.931
R1072 VDD.t995 VDD.t704 213.931
R1073 VDD.t704 VDD.t996 213.931
R1074 VDD.t1454 VDD.t1450 213.931
R1075 VDD.t1450 VDD.t606 213.931
R1076 VDD.t606 VDD.t79 213.931
R1077 VDD.t79 VDD.t605 213.931
R1078 VDD.t656 VDD.t658 213.931
R1079 VDD.t658 VDD.t541 213.931
R1080 VDD.t1318 VDD.t1322 213.931
R1081 VDD.t1322 VDD.t1612 213.931
R1082 VDD.t1612 VDD.t1611 213.931
R1083 VDD.t1611 VDD.t1441 213.931
R1084 VDD.t1599 VDD.t1214 213.931
R1085 VDD.t1214 VDD.t1246 213.931
R1086 VDD.t1246 VDD.t1247 213.931
R1087 VDD.t1247 VDD.t436 213.931
R1088 VDD.t920 VDD.t840 213.931
R1089 VDD.t840 VDD.t770 213.931
R1090 VDD.t1354 VDD.t1356 213.931
R1091 VDD.t1356 VDD.t1377 213.931
R1092 VDD.t1377 VDD.t1378 213.931
R1093 VDD.t1378 VDD.t1379 213.931
R1094 VDD.t505 VDD.t1096 213.931
R1095 VDD.t1096 VDD.t307 213.931
R1096 VDD.t307 VDD.t299 213.931
R1097 VDD.t299 VDD.t306 213.931
R1098 VDD.t1083 VDD.t1563 213.931
R1099 VDD.t1563 VDD.t1561 213.931
R1100 VDD.t405 VDD.t1569 213.931
R1101 VDD.t1569 VDD.t401 213.931
R1102 VDD.t67 VDD.t65 213.931
R1103 VDD.t65 VDD.t461 213.931
R1104 VDD.t40 VDD.t391 213.931
R1105 VDD.t391 VDD.t389 213.931
R1106 VDD.t1317 VDD.t1439 205.749
R1107 VDD.t129 VDD.t768 205.749
R1108 VDD.t271 VDD.t1474 205.749
R1109 VDD.t687 VDD.t628 205.749
R1110 VDD.t1439 VDD.t1437 197.707
R1111 VDD.t1437 VDD.t1581 197.707
R1112 VDD.t768 VDD.t766 197.707
R1113 VDD.t766 VDD.t1027 197.707
R1114 VDD.t716 VDD.t553 197.707
R1115 VDD.t1474 VDD.t1510 197.707
R1116 VDD.t1510 VDD.t1508 197.707
R1117 VDD.t290 VDD.t288 197.707
R1118 VDD.t628 VDD.t634 197.707
R1119 VDD.t634 VDD.t626 197.707
R1120 VDD.t115 VDD.t1085 197.707
R1121 VDD.t1198 VDD.t1196 197.707
R1122 VDD.t22 VDD.t684 196.666
R1123 VDD.t24 VDD.t22 196.666
R1124 VDD.t654 VDD.t24 196.666
R1125 VDD.t730 VDD.t654 196.666
R1126 VDD.t652 VDD.t730 196.666
R1127 VDD.t272 VDD.t1534 196.666
R1128 VDD.t1534 VDD.t213 196.666
R1129 VDD.t836 VDD.t834 196.666
R1130 VDD.t292 VDD.t836 196.666
R1131 VDD.t1183 VDD.t292 196.666
R1132 VDD.t1380 VDD.t1183 196.666
R1133 VDD.t820 VDD.t1380 196.666
R1134 VDD.t746 VDD.t375 196.666
R1135 VDD.t375 VDD.t1456 196.666
R1136 VDD.t236 VDD.t1618 196.666
R1137 VDD.t234 VDD.t236 196.666
R1138 VDD.t1591 VDD.t234 196.666
R1139 VDD.t274 VDD.t1591 196.666
R1140 VDD.t1464 VDD.t274 196.666
R1141 VDD.t1622 VDD.t459 196.666
R1142 VDD.t459 VDD.t974 196.666
R1143 VDD.t517 VDD.t519 196.666
R1144 VDD.t515 VDD.t517 196.666
R1145 VDD.t373 VDD.t515 196.666
R1146 VDD.t744 VDD.t373 196.666
R1147 VDD.t1460 VDD.t744 196.666
R1148 VDD.t728 VDD.t726 196.666
R1149 VDD.t726 VDD.t708 196.666
R1150 VDD.t1515 VDD.t1517 196.666
R1151 VDD.t985 VDD.t1515 196.666
R1152 VDD.t365 VDD.t985 196.666
R1153 VDD.t363 VDD.t365 196.666
R1154 VDD.t361 VDD.t363 196.666
R1155 VDD.t1153 VDD.t1151 196.666
R1156 VDD.t1151 VDD.t1011 196.666
R1157 VDD.t1368 VDD.t1366 196.666
R1158 VDD.t1620 VDD.t1368 196.666
R1159 VDD.t942 VDD.t1620 196.666
R1160 VDD.t782 VDD.t942 196.666
R1161 VDD.t868 VDD.t782 196.666
R1162 VDD.t1462 VDD.t231 196.666
R1163 VDD.t231 VDD.t1593 196.666
R1164 VDD.t1131 VDD.t1547 196.666
R1165 VDD.t1545 VDD.t1131 196.666
R1166 VDD.t385 VDD.t1545 196.666
R1167 VDD.t1071 VDD.t385 196.666
R1168 VDD.t229 VDD.t1071 196.666
R1169 VDD.t179 VDD.t722 196.666
R1170 VDD.t722 VDD.t1077 196.666
R1171 VDD.t1176 VDD.t1178 196.666
R1172 VDD.t908 VDD.t1176 196.666
R1173 VDD.t784 VDD.t908 196.666
R1174 VDD.t866 VDD.t784 196.666
R1175 VDD.t900 VDD.t866 196.666
R1176 VDD.t144 VDD.t774 196.666
R1177 VDD.t774 VDD.t225 196.666
R1178 VDD.t157 VDD.t155 196.666
R1179 VDD.t1033 VDD.t157 196.666
R1180 VDD.t1458 VDD.t1033 196.666
R1181 VDD.t371 VDD.t1458 196.666
R1182 VDD.t134 VDD.t371 196.666
R1183 VDD.t864 VDD.t862 196.666
R1184 VDD.t862 VDD.t780 196.666
R1185 VDD.t906 VDD.t904 196.666
R1186 VDD.t50 VDD.t906 196.666
R1187 VDD.t756 VDD.t50 196.666
R1188 VDD.t646 VDD.t756 196.666
R1189 VDD.t644 VDD.t646 196.666
R1190 VDD.t1415 VDD.t1392 196.666
R1191 VDD.t1392 VDD.t1403 196.666
R1192 VDD.t167 VDD.t171 196.666
R1193 VDD.t169 VDD.t167 196.666
R1194 VDD.t1075 VDD.t169 196.666
R1195 VDD.t1577 VDD.t1075 196.666
R1196 VDD.t1575 VDD.t1577 196.666
R1197 VDD.t854 VDD.t778 196.666
R1198 VDD.t778 VDD.t227 196.666
R1199 VDD.t1429 VDD.t1431 196.666
R1200 VDD.t1421 VDD.t1429 196.666
R1201 VDD.t1401 VDD.t1421 196.666
R1202 VDD.t1399 VDD.t1401 196.666
R1203 VDD.t1397 VDD.t1399 196.666
R1204 VDD.t940 VDD.t938 196.666
R1205 VDD.t938 VDD.t902 196.666
R1206 VDD.t75 VDD.t77 196.666
R1207 VDD.t73 VDD.t75 196.666
R1208 VDD.t688 VDD.t73 196.666
R1209 VDD.t1025 VDD.t688 196.666
R1210 VDD.t1023 VDD.t1025 196.666
R1211 VDD.t579 VDD.t577 196.666
R1212 VDD.t577 VDD.t720 196.666
R1213 VDD.t1372 VDD.t1370 196.666
R1214 VDD.t1374 VDD.t1372 196.666
R1215 VDD.t1512 VDD.t1374 196.666
R1216 VDD.t173 VDD.t1512 196.666
R1217 VDD.t177 VDD.t173 196.666
R1218 VDD.t1388 VDD.t966 196.666
R1219 VDD.t966 VDD.t964 196.666
R1220 VDD.t1423 VDD.t1425 196.666
R1221 VDD.t1427 VDD.t1423 196.666
R1222 VDD.t1413 VDD.t1427 196.666
R1223 VDD.t1405 VDD.t1413 196.666
R1224 VDD.t1417 VDD.t1405 196.666
R1225 VDD.t1009 VDD.t1470 196.666
R1226 VDD.t1470 VDD.t181 196.666
R1227 VDD.t616 VDD.t618 196.666
R1228 VDD.t614 VDD.t616 196.666
R1229 VDD.t636 VDD.t614 196.666
R1230 VDD.t632 VDD.t636 196.666
R1231 VDD.t640 VDD.t632 196.666
R1232 VDD.t1091 VDD.t441 196.666
R1233 VDD.t441 VDD.t1087 196.666
R1234 VDD.t648 VDD.t650 196.666
R1235 VDD.t191 VDD.t648 196.666
R1236 VDD.t415 VDD.t191 196.666
R1237 VDD.t882 VDD.t415 196.666
R1238 VDD.t880 VDD.t882 196.666
R1239 VDD.t1202 VDD.t1133 196.666
R1240 VDD.t1133 VDD.t357 196.666
R1241 VDD.t1100 VDD.t1174 196.666
R1242 VDD.t1098 VDD.t1100 196.666
R1243 VDD.t1384 VDD.t1098 196.666
R1244 VDD.t612 VDD.t1384 196.666
R1245 VDD.t1185 VDD.t612 196.666
R1246 VDD.t223 VDD.t221 196.666
R1247 VDD.t221 VDD.t856 196.666
R1248 VDD.t890 VDD.t395 196.666
R1249 VDD.t583 VDD.t890 196.666
R1250 VDD.t1411 VDD.t583 196.666
R1251 VDD.t1409 VDD.t1411 196.666
R1252 VDD.t1407 VDD.t1409 196.666
R1253 VDD.t1628 VDD.t1382 196.666
R1254 VDD.t1382 VDD.t1630 196.666
R1255 VDD.t1502 VDD.t1466 192.281
R1256 VDD.t1216 VDD.t1221 192.281
R1257 VDD.t1216 VDD.t1219 192.281
R1258 VDD.t838 VDD.t1021 192.281
R1259 VDD.t246 VDD.t248 192.281
R1260 VDD.t246 VDD.t244 192.281
R1261 VDD.t28 VDD.t1046 192.281
R1262 VDD.t324 VDD.t694 192.281
R1263 VDD.t324 VDD.t322 192.281
R1264 VDD.t486 VDD.t1595 192.281
R1265 VDD.t523 VDD.t447 192.281
R1266 VDD.t523 VDD.t521 192.281
R1267 VDD.t1442 VDD.t1172 192.281
R1268 VDD.t1543 VDD.t1476 192.281
R1269 VDD.t1543 VDD.t1541 192.281
R1270 VDD.t509 VDD.t932 192.281
R1271 VDD.t347 VDD.t1051 192.281
R1272 VDD.t347 VDD.t1049 192.281
R1273 VDD.t286 VDD.t411 192.281
R1274 VDD.t457 VDD.t513 192.281
R1275 VDD.t457 VDD.t511 192.281
R1276 VDD.t252 VDD.t250 192.281
R1277 VDD.t878 VDD.t409 192.281
R1278 VDD.t878 VDD.t407 192.281
R1279 VDD.n916 VDD.t1468 169.468
R1280 VDD.n946 VDD.t55 169.468
R1281 VDD.n977 VDD.t26 169.468
R1282 VDD.n1007 VDD.t1506 169.468
R1283 VDD.n597 VDD.t1444 169.468
R1284 VDD.n684 VDD.t930 169.468
R1285 VDD.n763 VDD.t413 169.468
R1286 VDD.n843 VDD.t445 169.468
R1287 VDD.n521 VDD.n520 142.5
R1288 VDD.n660 VDD.n659 142.5
R1289 VDD.n748 VDD.n747 142.5
R1290 VDD.n814 VDD.n813 142.5
R1291 VDD.n137 VDD.n136 142.5
R1292 VDD.n202 VDD.n201 142.5
R1293 VDD.n270 VDD.n269 142.5
R1294 VDD.n331 VDD.n330 142.5
R1295 VDD.t1216 VDD.t822 135.973
R1296 VDD.t246 VDD.t215 135.973
R1297 VDD.t324 VDD.t1139 135.973
R1298 VDD.t523 VDD.t1244 135.973
R1299 VDD.t1543 VDD.t999 135.973
R1300 VDD.t347 VDD.t1454 135.973
R1301 VDD.t457 VDD.t1599 135.973
R1302 VDD.t878 VDD.t505 135.973
R1303 VDD.n916 VDD.t1212 110.591
R1304 VDD.n946 VDD.t991 110.591
R1305 VDD.n977 VDD.t1496 110.591
R1306 VDD.n1007 VDD.t1226 110.591
R1307 VDD.n597 VDD.t934 110.591
R1308 VDD.n684 VDD.t681 110.591
R1309 VDD.n763 VDD.t1318 110.591
R1310 VDD.n843 VDD.t1354 110.591
R1311 VDD.n498 VDD.t1043 105.555
R1312 VDD.n482 VDD.t1332 105.555
R1313 VDD.n927 VDD.t336 105.555
R1314 VDD.n957 VDD.t34 105.555
R1315 VDD.n987 VDD.t282 105.555
R1316 VDD.n1016 VDD.t740 105.555
R1317 VDD.n593 VDD.t1029 105.555
R1318 VDD.n635 VDD.t151 105.555
R1319 VDD.n622 VDD.t830 105.555
R1320 VDD.n670 VDD.t976 105.555
R1321 VDD.n716 VDD.t660 105.555
R1322 VDD.n698 VDD.t1094 105.555
R1323 VDD.n754 VDD.t842 105.555
R1324 VDD.n794 VDD.t844 105.555
R1325 VDD.n782 VDD.t1587 105.555
R1326 VDD.n831 VDD.t565 105.555
R1327 VDD.n111 VDD.t355 105.555
R1328 VDD.n94 VDD.t1305 105.555
R1329 VDD.n176 VDD.t205 105.555
R1330 VDD.n168 VDD.t525 105.555
R1331 VDD.n243 VDD.t463 105.555
R1332 VDD.n225 VDD.t858 105.555
R1333 VDD.n306 VDD.t330 105.555
R1334 VDD.n293 VDD.t910 105.555
R1335 VDD.t1208 VDD.n916 103.339
R1336 VDD.t989 VDD.n946 103.339
R1337 VDD.t1498 VDD.n977 103.339
R1338 VDD.t1224 VDD.n1007 103.339
R1339 VDD.t297 VDD.n597 103.339
R1340 VDD.t1601 VDD.n684 103.339
R1341 VDD.t1320 VDD.n763 103.339
R1342 VDD.t1348 VDD.n843 103.339
R1343 VDD.t1216 VDD.t824 77.958
R1344 VDD.t246 VDD.t662 77.958
R1345 VDD.t324 VDD.t936 77.958
R1346 VDD.t523 VDD.t1263 77.958
R1347 VDD.t1543 VDD.t997 77.958
R1348 VDD.t347 VDD.t1452 77.958
R1349 VDD.t457 VDD.t1597 77.958
R1350 VDD.t878 VDD.t503 77.958
R1351 VDD.t611 VDD.t1342 53.244
R1352 VDD.t1520 VDD.t555 53.244
R1353 VDD.t94 VDD.t1480 53.244
R1354 VDD.t537 VDD.t1093 53.244
R1355 VDD.t233 VDD.t432 53.244
R1356 VDD.t1141 VDD.t1610 53.244
R1357 VDD.t452 VDD.t258 53.244
R1358 VDD.t951 VDD.t429 53.244
R1359 VDD.t751 VDD.t1299 53.244
R1360 VDD.t896 VDD.t1156 53.244
R1361 VDD.t886 VDD.t678 53.244
R1362 VDD.t527 VDD.t465 53.244
R1363 VDD.t958 VDD.t104 53.244
R1364 VDD.t1524 VDD.t1223 53.244
R1365 VDD.t394 VDD.t959 53.244
R1366 VDD.t1490 VDD.t984 53.244
R1367 VDD.t1346 VDD.n516 47.617
R1368 VDD.t1342 VDD.n517 47.617
R1369 VDD.n519 VDD.t183 47.617
R1370 VDD.n518 VDD.t1520 47.617
R1371 VDD.t269 VDD.n655 47.617
R1372 VDD.t1480 VDD.n656 47.617
R1373 VDD.n658 VDD.t762 47.617
R1374 VDD.n657 VDD.t537 47.617
R1375 VDD.t698 VDD.n743 47.617
R1376 VDD.t432 VDD.n744 47.617
R1377 VDD.n746 VDD.t1192 47.617
R1378 VDD.n745 VDD.t1141 47.617
R1379 VDD.t1165 VDD.n809 47.617
R1380 VDD.t258 VDD.n810 47.617
R1381 VDD.n812 VDD.t872 47.617
R1382 VDD.n811 VDD.t951 47.617
R1383 VDD.t1309 VDD.n132 47.617
R1384 VDD.t1299 VDD.n133 47.617
R1385 VDD.n135 VDD.t898 47.617
R1386 VDD.n134 VDD.t896 47.617
R1387 VDD.t978 VDD.n197 47.617
R1388 VDD.t678 VDD.n198 47.617
R1389 VDD.n200 VDD.t529 47.617
R1390 VDD.n199 VDD.t527 47.617
R1391 VDD.t106 VDD.n265 47.617
R1392 VDD.t104 VDD.n266 47.617
R1393 VDD.n268 VDD.t1526 47.617
R1394 VDD.n267 VDD.t1524 47.617
R1395 VDD.t1015 VDD.n326 47.617
R1396 VDD.t959 VDD.n327 47.617
R1397 VDD.n329 VDD.t1492 47.617
R1398 VDD.n328 VDD.t1490 47.617
R1399 VDD.t1045 VDD.t852 47.617
R1400 VDD.t260 VDD.t302 47.617
R1401 VDD.t889 VDD.t569 47.617
R1402 VDD.t680 VDD.t90 47.617
R1403 VDD.t11 VDD.t201 47.617
R1404 VDD.t1533 VDD.t793 47.617
R1405 VDD.t1528 VDD.t1181 47.617
R1406 VDD.t1529 VDD.t1111 47.617
R1407 VDD.t597 VDD.t4 47.617
R1408 VDD.t598 VDD.t2 47.617
R1409 VDD.t1394 VDD.t1273 47.617
R1410 VDD.t1395 VDD.t1121 47.617
R1411 VDD.t1396 VDD.t608 47.617
R1412 VDD.t876 VDD.t1007 47.617
R1413 VDD.t714 VDD.t668 47.617
R1414 VDD.t1102 VDD.t1039 47.617
R1415 VDD.t642 VDD.t18 47.617
R1416 VDD.t643 VDD.t772 47.617
R1417 VDD.t494 VDD.t922 47.617
R1418 VDD.t495 VDD.t846 47.617
R1419 VDD.t1580 VDD.t1538 47.617
R1420 VDD.t1579 VDD.t1536 47.617
R1421 VDD.t607 VDD.t369 47.617
R1422 VDD.t888 VDD.t367 47.617
R1423 VDD.t887 VDD.t351 47.617
R1424 VDD.t556 VDD.t702 47.617
R1425 VDD.t1180 VDD.t700 47.617
R1426 VDD.t805 VDD.t209 47.617
R1427 VDD.t750 VDD.t207 47.617
R1428 VDD.t749 VDD.t1488 47.617
R1429 VDD.t963 VDD.t280 47.617
R1430 VDD.t47 VDD.t278 47.617
R1431 VDD.t46 VDD.t916 47.617
R1432 VDD.t1252 VDD.t14 47.617
R1433 VDD.t1315 VDD.t12 47.617
R1434 VDD.t786 VDD.t1255 47.617
R1435 VDD.t590 VDD.t1259 47.617
R1436 VDD.t589 VDD.t332 47.617
R1437 VDD.t1065 VDD.t328 47.617
R1438 VDD.t604 VDD.t339 47.617
R1439 VDD.n917 VDD.t1208 47.137
R1440 VDD.n947 VDD.t989 47.137
R1441 VDD.n978 VDD.t1498 47.137
R1442 VDD.n1008 VDD.t1224 47.137
R1443 VDD.n598 VDD.t297 47.137
R1444 VDD.n685 VDD.t1601 47.137
R1445 VDD.n764 VDD.t1320 47.137
R1446 VDD.n844 VDD.t1348 47.137
R1447 VDD.t561 VDD.t950 45.992
R1448 VDD.t581 VDD.t949 45.992
R1449 VDD.t131 VDD.t575 45.992
R1450 VDD.t130 VDD.t573 45.992
R1451 VDD.t1571 VDD.t61 45.992
R1452 VDD.t1573 VDD.t877 45.992
R1453 VDD.t1617 VDD.t175 45.992
R1454 VDD.t338 VDD.t1472 45.992
R1455 VDD.t439 VDD.t1187 45.992
R1456 VDD.t117 VDD.t754 45.992
R1457 VDD.t1160 VDD.t624 45.992
R1458 VDD.t1159 VDD.t638 45.992
R1459 VDD.t670 VDD.t1218 45.992
R1460 VDD.t1204 VDD.t1540 45.992
R1461 VDD.t1316 VDD.t692 45.992
R1462 VDD.t1376 VDD.t690 45.992
R1463 VDD.n517 VDD.t1346 44.495
R1464 VDD.t1565 VDD.n519 44.495
R1465 VDD.t183 VDD.n518 44.495
R1466 VDD.n516 VDD.t1334 44.495
R1467 VDD.n656 VDD.t269 44.495
R1468 VDD.t764 VDD.n658 44.495
R1469 VDD.t762 VDD.n657 44.495
R1470 VDD.n655 VDD.t826 44.495
R1471 VDD.n744 VDD.t698 44.495
R1472 VDD.t1143 VDD.n746 44.495
R1473 VDD.t1192 VDD.n745 44.495
R1474 VDD.n743 VDD.t1125 44.495
R1475 VDD.n810 VDD.t1165 44.495
R1476 VDD.t955 VDD.n812 44.495
R1477 VDD.t872 VDD.n811 44.495
R1478 VDD.n809 VDD.t1557 44.495
R1479 VDD.n133 VDD.t1309 44.495
R1480 VDD.t595 VDD.n135 44.495
R1481 VDD.t898 VDD.n134 44.495
R1482 VDD.n132 VDD.t1311 44.495
R1483 VDD.n198 VDD.t978 44.495
R1484 VDD.t531 VDD.n200 44.495
R1485 VDD.t529 VDD.n199 44.495
R1486 VDD.n197 VDD.t379 44.495
R1487 VDD.n266 VDD.t106 44.495
R1488 VDD.t622 VDD.n268 44.495
R1489 VDD.t1526 VDD.n267 44.495
R1490 VDD.n265 VDD.t113 44.495
R1491 VDD.n327 VDD.t1015 44.495
R1492 VDD.t1494 VDD.n329 44.495
R1493 VDD.t1492 VDD.n328 44.495
R1494 VDD.n326 VDD.t1019 44.495
R1495 VDD.t304 VDD.t1045 44.494
R1496 VDD.t852 VDD.t260 44.494
R1497 VDD.t302 VDD.t889 44.494
R1498 VDD.t569 VDD.t680 44.494
R1499 VDD.t90 VDD.t11 44.494
R1500 VDD.t201 VDD.t10 44.494
R1501 VDD.t795 VDD.t1533 44.494
R1502 VDD.t793 VDD.t1528 44.494
R1503 VDD.t1181 VDD.t1529 44.494
R1504 VDD.t1111 VDD.t597 44.494
R1505 VDD.t4 VDD.t598 44.494
R1506 VDD.t2 VDD.t683 44.494
R1507 VDD.t1275 VDD.t1394 44.494
R1508 VDD.t1273 VDD.t1395 44.494
R1509 VDD.t1121 VDD.t1396 44.494
R1510 VDD.t608 VDD.t876 44.494
R1511 VDD.t1007 VDD.t714 44.494
R1512 VDD.t668 VDD.t715 44.494
R1513 VDD.t20 VDD.t1102 44.494
R1514 VDD.t1039 VDD.t642 44.494
R1515 VDD.t18 VDD.t643 44.494
R1516 VDD.t772 VDD.t494 44.494
R1517 VDD.t922 VDD.t495 44.494
R1518 VDD.t846 VDD.t1514 44.494
R1519 VDD.t1115 VDD.t1580 44.494
R1520 VDD.t1538 VDD.t1579 44.494
R1521 VDD.t1536 VDD.t607 44.494
R1522 VDD.t369 VDD.t888 44.494
R1523 VDD.t367 VDD.t887 44.494
R1524 VDD.t351 VDD.t705 44.494
R1525 VDD.t1435 VDD.t556 44.494
R1526 VDD.t702 VDD.t1180 44.494
R1527 VDD.t700 VDD.t805 44.494
R1528 VDD.t209 VDD.t750 44.494
R1529 VDD.t207 VDD.t749 44.494
R1530 VDD.t1488 VDD.t748 44.494
R1531 VDD.t472 VDD.t963 44.494
R1532 VDD.t280 VDD.t47 44.494
R1533 VDD.t278 VDD.t46 44.494
R1534 VDD.t916 VDD.t1252 44.494
R1535 VDD.t14 VDD.t1315 44.494
R1536 VDD.t12 VDD.t489 44.494
R1537 VDD.t1230 VDD.t786 44.494
R1538 VDD.t1255 VDD.t590 44.494
R1539 VDD.t1259 VDD.t589 44.494
R1540 VDD.t332 VDD.t1065 44.494
R1541 VDD.t328 VDD.t604 44.494
R1542 VDD.t339 VDD.t1066 44.494
R1543 VDD.t950 VDD.t718 42.976
R1544 VDD.t949 VDD.t561 42.976
R1545 VDD.t948 VDD.t581 42.976
R1546 VDD.t136 VDD.t131 42.976
R1547 VDD.t575 VDD.t130 42.976
R1548 VDD.t573 VDD.t129 42.976
R1549 VDD.t61 VDD.t968 42.976
R1550 VDD.t877 VDD.t1571 42.976
R1551 VDD.t62 VDD.t1573 42.976
R1552 VDD.t256 VDD.t1617 42.976
R1553 VDD.t175 VDD.t338 42.976
R1554 VDD.t1472 VDD.t271 42.976
R1555 VDD.t1187 VDD.t1089 42.976
R1556 VDD.t754 VDD.t439 42.976
R1557 VDD.t755 VDD.t117 42.976
R1558 VDD.t630 VDD.t1160 42.976
R1559 VDD.t624 VDD.t1159 42.976
R1560 VDD.t638 VDD.t687 42.976
R1561 VDD.t1218 VDD.t1200 42.976
R1562 VDD.t1540 VDD.t670 42.976
R1563 VDD.t294 VDD.t1204 42.976
R1564 VDD.t1583 VDD.t1316 42.976
R1565 VDD.t692 VDD.t1376 42.976
R1566 VDD.t690 VDD.t1317 42.976
R1567 VDD.n434 VDD.t136 37.698
R1568 VDD.n376 VDD.t256 37.698
R1569 VDD.n408 VDD.t630 37.698
R1570 VDD.n364 VDD.t1583 37.698
R1571 VDD.n16 VDD.t214 30.163
R1572 VDD.n7 VDD.t1457 30.163
R1573 VDD.n491 VDD.t1337 30.163
R1574 VDD.n479 VDD.t479 30.163
R1575 VDD.n924 VDD.t1239 30.163
R1576 VDD.n953 VDD.t200 30.163
R1577 VDD.n984 VDD.t1434 30.163
R1578 VDD.n1019 VDD.t1128 30.163
R1579 VDD.n62 VDD.t548 30.163
R1580 VDD.n884 VDD.t975 30.163
R1581 VDD.n893 VDD.t709 30.163
R1582 VDD.n59 VDD.t1012 30.163
R1583 VDD.n50 VDD.t1594 30.163
R1584 VDD.n41 VDD.t1078 30.163
R1585 VDD.n590 VDD.t809 30.163
R1586 VDD.n32 VDD.t226 30.163
R1587 VDD.n638 VDD.t1483 30.163
R1588 VDD.n629 VDD.t792 30.163
R1589 VDD.n667 VDD.t1278 30.163
R1590 VDD.n713 VDD.t558 30.163
R1591 VDD.n701 VDD.t1282 30.163
R1592 VDD.n757 VDD.t346 30.163
R1593 VDD.n791 VDD.t1590 30.163
R1594 VDD.n779 VDD.t1042 30.163
R1595 VDD.n834 VDD.t849 30.163
R1596 VDD.n24 VDD.t781 30.163
R1597 VDD.n115 VDD.t1298 30.163
R1598 VDD.n97 VDD.t493 30.163
R1599 VDD.n179 VDD.t971 30.163
R1600 VDD.n165 VDD.t711 30.163
R1601 VDD.n240 VDD.t1002 30.163
R1602 VDD.n232 VDD.t929 30.163
R1603 VDD.n309 VDD.t800 30.163
R1604 VDD.n300 VDD.t1241 30.163
R1605 VDD.n475 VDD.t1404 30.163
R1606 VDD.n466 VDD.t228 30.163
R1607 VDD.n352 VDD.t903 30.163
R1608 VDD.n448 VDD.t358 30.163
R1609 VDD.n443 VDD.t721 30.163
R1610 VDD.n385 VDD.t965 30.163
R1611 VDD.n417 VDD.t182 30.163
R1612 VDD.n395 VDD.t1088 30.163
R1613 VDD.n872 VDD.t857 30.163
R1614 VDD.n881 VDD.t1631 30.163
R1615 VDD.n520 VDD.t611 28.957
R1616 VDD.n659 VDD.t94 28.957
R1617 VDD.n747 VDD.t233 28.957
R1618 VDD.n813 VDD.t452 28.957
R1619 VDD.n136 VDD.t751 28.957
R1620 VDD.n201 VDD.t886 28.957
R1621 VDD.n269 VDD.t958 28.957
R1622 VDD.n330 VDD.t394 28.957
R1623 VDD.n523 VDD.t1158 28.664
R1624 VDD.n528 VDD.t1339 28.664
R1625 VDD.n505 VDD.t564 28.664
R1626 VDD.n510 VDD.t72 28.664
R1627 VDD.n609 VDD.t536 28.664
R1628 VDD.n614 VDD.t399 28.664
R1629 VDD.n644 VDD.t1114 28.664
R1630 VDD.n649 VDD.t7 28.664
R1631 VDD.n733 VDD.t1191 28.664
R1632 VDD.n738 VDD.t500 28.664
R1633 VDD.n720 VDD.t657 28.664
R1634 VDD.n725 VDD.t1120 28.664
R1635 VDD.n817 VDD.t875 28.664
R1636 VDD.n822 VDD.t1162 28.664
R1637 VDD.n798 VDD.t921 28.664
R1638 VDD.n803 VDD.t342 28.664
R1639 VDD.n84 VDD.t43 28.664
R1640 VDD.n89 VDD.t1292 28.664
R1641 VDD.n121 VDD.t1084 28.664
R1642 VDD.n126 VDD.t450 28.664
R1643 VDD.n150 VDD.t485 28.664
R1644 VDD.n155 VDD.t1189 28.664
R1645 VDD.n186 VDD.t406 28.664
R1646 VDD.n191 VDD.t103 28.664
R1647 VDD.n215 VDD.t621 28.664
R1648 VDD.n220 VDD.t945 28.664
R1649 VDD.n254 VDD.t68 28.664
R1650 VDD.n259 VDD.t277 28.664
R1651 VDD.n334 VDD.t100 28.664
R1652 VDD.n339 VDD.t802 28.664
R1653 VDD.n315 VDD.t41 28.664
R1654 VDD.n320 VDD.t1233 28.664
R1655 VDD.n359 VDD.t1440 28.664
R1656 VDD.n354 VDD.t673 28.664
R1657 VDD.n429 VDD.t769 28.664
R1658 VDD.n424 VDD.t552 28.664
R1659 VDD.n371 VDD.t1475 28.664
R1660 VDD.n366 VDD.t1391 28.664
R1661 VDD.n403 VDD.t629 28.664
R1662 VDD.n398 VDD.t444 28.664
R1663 VDD.n278 VDD.t1467 28.57
R1664 VDD.n285 VDD.t1222 28.57
R1665 VDD.n210 VDD.t1022 28.57
R1666 VDD.n934 VDD.t249 28.57
R1667 VDD.n145 VDD.t1047 28.57
R1668 VDD.n966 VDD.t695 28.57
R1669 VDD.n78 VDD.t1596 28.57
R1670 VDD.n994 VDD.t448 28.57
R1671 VDD.n580 VDD.t1173 28.57
R1672 VDD.n573 VDD.t1477 28.57
R1673 VDD.n677 VDD.t933 28.57
R1674 VDD.n563 VDD.t1052 28.57
R1675 VDD.n553 VDD.t412 28.57
R1676 VDD.n546 VDD.t514 28.57
R1677 VDD.n536 VDD.t251 28.57
R1678 VDD.n854 VDD.t410 28.57
R1679 VDD.n15 VDD.t273 28.565
R1680 VDD.n15 VDD.t1535 28.565
R1681 VDD.n10 VDD.t685 28.565
R1682 VDD.n10 VDD.t23 28.565
R1683 VDD.n11 VDD.t25 28.565
R1684 VDD.n11 VDD.t655 28.565
R1685 VDD.n13 VDD.t731 28.565
R1686 VDD.n13 VDD.t653 28.565
R1687 VDD.n6 VDD.t747 28.565
R1688 VDD.n6 VDD.t376 28.565
R1689 VDD.n1 VDD.t835 28.565
R1690 VDD.n1 VDD.t837 28.565
R1691 VDD.n2 VDD.t293 28.565
R1692 VDD.n2 VDD.t1184 28.565
R1693 VDD.n4 VDD.t1381 28.565
R1694 VDD.n4 VDD.t821 28.565
R1695 VDD.n524 VDD.t1523 28.565
R1696 VDD.n524 VDD.t1568 28.565
R1697 VDD.n529 VDD.t1345 28.565
R1698 VDD.n529 VDD.t1325 28.565
R1699 VDD.n506 VDD.t204 28.565
R1700 VDD.n506 VDD.t89 28.565
R1701 VDD.n511 VDD.t315 28.565
R1702 VDD.n511 VDD.t481 28.565
R1703 VDD.n490 VDD.t1329 28.565
R1704 VDD.n490 VDD.t1327 28.565
R1705 VDD.n494 VDD.t1064 28.565
R1706 VDD.n494 VDD.t422 28.565
R1707 VDD.n495 VDD.t1062 28.565
R1708 VDD.n495 VDD.t87 28.565
R1709 VDD.n489 VDD.t1044 28.565
R1710 VDD.n489 VDD.t572 28.565
R1711 VDD.n478 VDD.t301 28.565
R1712 VDD.n478 VDD.t851 28.565
R1713 VDD.n483 VDD.t317 28.565
R1714 VDD.n483 VDD.t319 28.565
R1715 VDD.n484 VDD.t321 28.565
R1716 VDD.n484 VDD.t1341 28.565
R1717 VDD.n477 VDD.t1333 28.565
R1718 VDD.n477 VDD.t1331 28.565
R1719 VDD.n923 VDD.t1243 28.565
R1720 VDD.n923 VDD.t1254 28.565
R1721 VDD.n273 VDD.t1286 28.565
R1722 VDD.n273 VDD.t1290 28.565
R1723 VDD.n274 VDD.t1288 28.565
R1724 VDD.n274 VDD.t388 28.565
R1725 VDD.n922 VDD.t337 28.565
R1726 VDD.n922 VDD.t335 28.565
R1727 VDD.n277 VDD.t1503 28.565
R1728 VDD.n277 VDD.t1469 28.565
R1729 VDD.n284 VDD.t1217 28.565
R1730 VDD.n284 VDD.t1220 28.565
R1731 VDD.n209 VDD.t839 28.565
R1732 VDD.n209 VDD.t56 28.565
R1733 VDD.n933 VDD.t247 28.565
R1734 VDD.n933 VDD.t245 28.565
R1735 VDD.n952 VDD.t477 28.565
R1736 VDD.n952 VDD.t927 28.565
R1737 VDD.n205 VDD.t735 28.565
R1738 VDD.n205 VDD.t733 28.565
R1739 VDD.n206 VDD.t737 28.565
R1740 VDD.n206 VDD.t37 28.565
R1741 VDD.n951 VDD.t35 28.565
R1742 VDD.n951 VDD.t33 28.565
R1743 VDD.n144 VDD.t29 28.565
R1744 VDD.n144 VDD.t27 28.565
R1745 VDD.n965 VDD.t325 28.565
R1746 VDD.n965 VDD.t323 28.565
R1747 VDD.n983 VDD.t1608 28.565
R1748 VDD.n983 VDD.t1606 28.565
R1749 VDD.n140 VDD.t546 28.565
R1750 VDD.n140 VDD.t544 28.565
R1751 VDD.n141 VDD.t1168 28.565
R1752 VDD.n141 VDD.t1130 28.565
R1753 VDD.n982 VDD.t283 28.565
R1754 VDD.n982 VDD.t1487 28.565
R1755 VDD.n77 VDD.t487 28.565
R1756 VDD.n77 VDD.t1507 28.565
R1757 VDD.n993 VDD.t524 28.565
R1758 VDD.n993 VDD.t522 28.565
R1759 VDD.n1018 VDD.t112 28.565
R1760 VDD.n1018 VDD.t110 28.565
R1761 VDD.n73 VDD.t456 28.565
R1762 VDD.n73 VDD.t753 28.565
R1763 VDD.n74 VDD.t243 28.565
R1764 VDD.n74 VDD.t743 28.565
R1765 VDD.n1017 VDD.t741 28.565
R1766 VDD.n1017 VDD.t759 28.565
R1767 VDD.n61 VDD.t707 28.565
R1768 VDD.n61 VDD.t550 28.565
R1769 VDD.n63 VDD.t1361 28.565
R1770 VDD.n63 VDD.t1365 28.565
R1771 VDD.n64 VDD.t1363 28.565
R1772 VDD.n64 VDD.t147 28.565
R1773 VDD.n66 VDD.t143 28.565
R1774 VDD.n66 VDD.t777 28.565
R1775 VDD.n883 VDD.t1623 28.565
R1776 VDD.n883 VDD.t460 28.565
R1777 VDD.n885 VDD.t1619 28.565
R1778 VDD.n885 VDD.t237 28.565
R1779 VDD.n886 VDD.t235 28.565
R1780 VDD.n886 VDD.t1592 28.565
R1781 VDD.n888 VDD.t275 28.565
R1782 VDD.n888 VDD.t1465 28.565
R1783 VDD.n892 VDD.t729 28.565
R1784 VDD.n892 VDD.t727 28.565
R1785 VDD.n894 VDD.t520 28.565
R1786 VDD.n894 VDD.t518 28.565
R1787 VDD.n895 VDD.t516 28.565
R1788 VDD.n895 VDD.t374 28.565
R1789 VDD.n897 VDD.t745 28.565
R1790 VDD.n897 VDD.t1461 28.565
R1791 VDD.n58 VDD.t1154 28.565
R1792 VDD.n58 VDD.t1152 28.565
R1793 VDD.n53 VDD.t1518 28.565
R1794 VDD.n53 VDD.t1516 28.565
R1795 VDD.n54 VDD.t986 28.565
R1796 VDD.n54 VDD.t366 28.565
R1797 VDD.n56 VDD.t364 28.565
R1798 VDD.n56 VDD.t362 28.565
R1799 VDD.n49 VDD.t1463 28.565
R1800 VDD.n49 VDD.t232 28.565
R1801 VDD.n44 VDD.t1367 28.565
R1802 VDD.n44 VDD.t1369 28.565
R1803 VDD.n45 VDD.t1621 28.565
R1804 VDD.n45 VDD.t943 28.565
R1805 VDD.n47 VDD.t783 28.565
R1806 VDD.n47 VDD.t869 28.565
R1807 VDD.n40 VDD.t180 28.565
R1808 VDD.n40 VDD.t723 28.565
R1809 VDD.n35 VDD.t1548 28.565
R1810 VDD.n35 VDD.t1132 28.565
R1811 VDD.n36 VDD.t1546 28.565
R1812 VDD.n36 VDD.t386 28.565
R1813 VDD.n38 VDD.t1072 28.565
R1814 VDD.n38 VDD.t230 28.565
R1815 VDD.n589 VDD.t819 28.565
R1816 VDD.n589 VDD.t811 28.565
R1817 VDD.n584 VDD.t1447 28.565
R1818 VDD.n584 VDD.t1449 28.565
R1819 VDD.n585 VDD.t1501 28.565
R1820 VDD.n585 VDD.t790 28.565
R1821 VDD.n588 VDD.t1030 28.565
R1822 VDD.n588 VDD.t154 28.565
R1823 VDD.n31 VDD.t145 28.565
R1824 VDD.n31 VDD.t775 28.565
R1825 VDD.n26 VDD.t1179 28.565
R1826 VDD.n26 VDD.t1177 28.565
R1827 VDD.n27 VDD.t909 28.565
R1828 VDD.n27 VDD.t785 28.565
R1829 VDD.n29 VDD.t867 28.565
R1830 VDD.n29 VDD.t901 28.565
R1831 VDD.n579 VDD.t1443 28.565
R1832 VDD.n579 VDD.t1445 28.565
R1833 VDD.n572 VDD.t1544 28.565
R1834 VDD.n572 VDD.t1542 28.565
R1835 VDD.n610 VDD.t45 28.565
R1836 VDD.n610 VDD.t761 28.565
R1837 VDD.n615 VDD.t1479 28.565
R1838 VDD.n615 VDD.t266 28.565
R1839 VDD.n645 VDD.t1032 28.565
R1840 VDD.n645 VDD.t1110 28.565
R1841 VDD.n650 VDD.t817 28.565
R1842 VDD.n650 VDD.t807 28.565
R1843 VDD.n637 VDD.t264 28.565
R1844 VDD.n637 VDD.t1485 28.565
R1845 VDD.n619 VDD.t426 28.565
R1846 VDD.n619 VDD.t428 28.565
R1847 VDD.n620 VDD.t350 28.565
R1848 VDD.n620 VDD.t1 28.565
R1849 VDD.n636 VDD.t152 28.565
R1850 VDD.n636 VDD.t788 28.565
R1851 VDD.n628 VDD.t798 28.565
R1852 VDD.n628 VDD.t9 28.565
R1853 VDD.n623 VDD.t162 28.565
R1854 VDD.n623 VDD.t149 28.565
R1855 VDD.n624 VDD.t164 28.565
R1856 VDD.n624 VDD.t268 28.565
R1857 VDD.n627 VDD.t831 28.565
R1858 VDD.n627 VDD.t829 28.565
R1859 VDD.n666 VDD.t1272 28.565
R1860 VDD.n666 VDD.t1284 28.565
R1861 VDD.n568 VDD.t49 28.565
R1862 VDD.n568 VDD.t418 28.565
R1863 VDD.n569 VDD.t124 28.565
R1864 VDD.n569 VDD.t1006 28.565
R1865 VDD.n665 VDD.t977 28.565
R1866 VDD.n665 VDD.t540 28.565
R1867 VDD.n676 VDD.t510 28.565
R1868 VDD.n676 VDD.t931 28.565
R1869 VDD.n562 VDD.t348 28.565
R1870 VDD.n562 VDD.t1050 28.565
R1871 VDD.n734 VDD.t1195 28.565
R1872 VDD.n734 VDD.t1106 28.565
R1873 VDD.n739 VDD.t502 28.565
R1874 VDD.n739 VDD.t120 28.565
R1875 VDD.n721 VDD.t659 28.565
R1876 VDD.n721 VDD.t542 28.565
R1877 VDD.n726 VDD.t1124 28.565
R1878 VDD.n726 VDD.t1280 28.565
R1879 VDD.n712 VDD.t697 28.565
R1880 VDD.n712 VDD.t431 28.565
R1881 VDD.n695 VDD.t667 28.565
R1882 VDD.n695 VDD.t31 28.565
R1883 VDD.n696 VDD.t1150 28.565
R1884 VDD.n696 VDD.t586 28.565
R1885 VDD.n711 VDD.t661 28.565
R1886 VDD.n711 VDD.t588 28.565
R1887 VDD.n700 VDD.t1270 28.565
R1888 VDD.n700 VDD.t1118 28.565
R1889 VDD.n705 VDD.t1251 28.565
R1890 VDD.n705 VDD.t1268 28.565
R1891 VDD.n706 VDD.t1249 28.565
R1892 VDD.n706 VDD.t239 28.565
R1893 VDD.n699 VDD.t1095 28.565
R1894 VDD.n699 VDD.t560 28.565
R1895 VDD.n756 VDD.t17 28.565
R1896 VDD.n756 VDD.t1136 28.565
R1897 VDD.n558 VDD.t1080 28.565
R1898 VDD.n558 VDD.t1082 28.565
R1899 VDD.n559 VDD.t1104 28.565
R1900 VDD.n559 VDD.t603 28.565
R1901 VDD.n755 VDD.t843 28.565
R1902 VDD.n755 VDD.t1560 28.565
R1903 VDD.n552 VDD.t287 28.565
R1904 VDD.n552 VDD.t414 28.565
R1905 VDD.n545 VDD.t458 28.565
R1906 VDD.n545 VDD.t512 28.565
R1907 VDD.n818 VDD.t954 28.565
R1908 VDD.n818 VDD.t871 28.565
R1909 VDD.n823 VDD.t190 28.565
R1910 VDD.n823 VDD.t188 28.565
R1911 VDD.n799 VDD.t841 28.565
R1912 VDD.n799 VDD.t771 28.565
R1913 VDD.n804 VDD.t1552 28.565
R1914 VDD.n804 VDD.t344 28.565
R1915 VDD.n790 VDD.t1531 28.565
R1916 VDD.n790 VDD.t186 28.565
R1917 VDD.n774 VDD.t218 28.565
R1918 VDD.n774 VDD.t220 28.565
R1919 VDD.n775 VDD.t833 28.565
R1920 VDD.n775 VDD.t925 28.565
R1921 VDD.n789 VDD.t845 28.565
R1922 VDD.n789 VDD.t601 28.565
R1923 VDD.n778 VDD.t1550 28.565
R1924 VDD.n778 VDD.t420 28.565
R1925 VDD.n783 VDD.t194 28.565
R1926 VDD.n783 VDD.t262 28.565
R1927 VDD.n784 VDD.t196 28.565
R1928 VDD.n784 VDD.t1164 28.565
R1929 VDD.n777 VDD.t1588 28.565
R1930 VDD.n777 VDD.t1556 28.565
R1931 VDD.n833 VDD.t313 28.565
R1932 VDD.n833 VDD.t70 28.565
R1933 VDD.n541 VDD.t1359 28.565
R1934 VDD.n541 VDD.t1353 28.565
R1935 VDD.n542 VDD.t1351 28.565
R1936 VDD.n542 VDD.t85 28.565
R1937 VDD.n832 VDD.t566 28.565
R1938 VDD.n832 VDD.t568 28.565
R1939 VDD.n535 VDD.t253 28.565
R1940 VDD.n535 VDD.t446 28.565
R1941 VDD.n853 VDD.t879 28.565
R1942 VDD.n853 VDD.t408 28.565
R1943 VDD.n23 VDD.t865 28.565
R1944 VDD.n23 VDD.t863 28.565
R1945 VDD.n18 VDD.t156 28.565
R1946 VDD.n18 VDD.t158 28.565
R1947 VDD.n19 VDD.t1034 28.565
R1948 VDD.n19 VDD.t1459 28.565
R1949 VDD.n21 VDD.t372 28.565
R1950 VDD.n21 VDD.t135 28.565
R1951 VDD.n85 VDD.t1038 28.565
R1952 VDD.n85 VDD.t1036 28.565
R1953 VDD.n90 VDD.t1296 28.565
R1954 VDD.n90 VDD.t1294 28.565
R1955 VDD.n122 VDD.t1564 28.565
R1956 VDD.n122 VDD.t1562 28.565
R1957 VDD.n127 VDD.t815 28.565
R1958 VDD.n127 VDD.t813 28.565
R1959 VDD.n114 VDD.t1304 28.565
R1960 VDD.n114 VDD.t1302 28.565
R1961 VDD.n107 VDD.t1616 28.565
R1962 VDD.n107 VDD.t1614 28.565
R1963 VDD.n108 VDD.t1586 28.565
R1964 VDD.n108 VDD.t739 28.565
R1965 VDD.n113 VDD.t356 28.565
R1966 VDD.n113 VDD.t354 28.565
R1967 VDD.n96 VDD.t491 28.565
R1968 VDD.n96 VDD.t122 28.565
R1969 VDD.n101 VDD.t212 28.565
R1970 VDD.n101 VDD.t60 28.565
R1971 VDD.n102 VDD.t58 28.565
R1972 VDD.n102 VDD.t1308 28.565
R1973 VDD.n95 VDD.t1306 28.565
R1974 VDD.n95 VDD.t1314 28.565
R1975 VDD.n151 VDD.t483 28.565
R1976 VDD.n151 VDD.t534 28.565
R1977 VDD.n156 VDD.t983 28.565
R1978 VDD.n156 VDD.t981 28.565
R1979 VDD.n187 VDD.t1570 28.565
R1980 VDD.n187 VDD.t402 28.565
R1981 VDD.n192 VDD.t1627 28.565
R1982 VDD.n192 VDD.t1625 28.565
R1983 VDD.n178 VDD.t677 28.565
R1984 VDD.n178 VDD.t973 28.565
R1985 VDD.n160 VDD.t1148 28.565
R1986 VDD.n160 VDD.t1146 28.565
R1987 VDD.n161 VDD.t255 28.565
R1988 VDD.n161 VDD.t404 28.565
R1989 VDD.n177 VDD.t206 28.565
R1990 VDD.n177 VDD.t285 28.565
R1991 VDD.n164 VDD.t594 28.565
R1992 VDD.n164 VDD.t592 28.565
R1993 VDD.n169 VDD.t133 28.565
R1994 VDD.n169 VDD.t128 28.565
R1995 VDD.n170 VDD.t126 28.565
R1996 VDD.n170 VDD.t378 28.565
R1997 VDD.n163 VDD.t526 28.565
R1998 VDD.n163 VDD.t675 28.565
R1999 VDD.n216 VDD.t384 28.565
R2000 VDD.n216 VDD.t382 28.565
R2001 VDD.n221 VDD.t893 28.565
R2002 VDD.n221 VDD.t895 28.565
R2003 VDD.n255 VDD.t66 28.565
R2004 VDD.n255 VDD.t462 28.565
R2005 VDD.n260 VDD.t198 28.565
R2006 VDD.n260 VDD.t83 28.565
R2007 VDD.n239 VDD.t1170 28.565
R2008 VDD.n239 VDD.t1004 28.565
R2009 VDD.n244 VDD.t1387 28.565
R2010 VDD.n244 VDD.t1056 28.565
R2011 VDD.n245 VDD.t1054 28.565
R2012 VDD.n245 VDD.t64 28.565
R2013 VDD.n238 VDD.t464 28.565
R2014 VDD.n238 VDD.t919 28.565
R2015 VDD.n231 VDD.t81 28.565
R2016 VDD.n231 VDD.t475 28.565
R2017 VDD.n226 VDD.t160 28.565
R2018 VDD.n226 VDD.t141 28.565
R2019 VDD.n227 VDD.t139 28.565
R2020 VDD.n227 VDD.t861 28.565
R2021 VDD.n230 VDD.t859 28.565
R2022 VDD.n230 VDD.t947 28.565
R2023 VDD.n335 VDD.t98 28.565
R2024 VDD.n335 VDD.t96 28.565
R2025 VDD.n340 VDD.t915 28.565
R2026 VDD.n340 VDD.t804 28.565
R2027 VDD.n316 VDD.t392 28.565
R2028 VDD.n316 VDD.t390 28.565
R2029 VDD.n321 VDD.t1237 28.565
R2030 VDD.n321 VDD.t1235 28.565
R2031 VDD.n308 VDD.t962 28.565
R2032 VDD.n308 VDD.t1014 28.565
R2033 VDD.n290 VDD.t1060 28.565
R2034 VDD.n290 VDD.t1058 28.565
R2035 VDD.n291 VDD.t424 28.565
R2036 VDD.n291 VDD.t39 28.565
R2037 VDD.n307 VDD.t331 28.565
R2038 VDD.n307 VDD.t327 28.565
R2039 VDD.n299 VDD.t1258 28.565
R2040 VDD.n299 VDD.t1262 28.565
R2041 VDD.n294 VDD.t469 28.565
R2042 VDD.n294 VDD.t467 28.565
R2043 VDD.n295 VDD.t1554 28.565
R2044 VDD.n295 VDD.t913 28.565
R2045 VDD.n298 VDD.t911 28.565
R2046 VDD.n298 VDD.t1018 28.565
R2047 VDD.n474 VDD.t1416 28.565
R2048 VDD.n474 VDD.t1393 28.565
R2049 VDD.n469 VDD.t905 28.565
R2050 VDD.n469 VDD.t907 28.565
R2051 VDD.n470 VDD.t51 28.565
R2052 VDD.n470 VDD.t757 28.565
R2053 VDD.n472 VDD.t647 28.565
R2054 VDD.n472 VDD.t645 28.565
R2055 VDD.n465 VDD.t855 28.565
R2056 VDD.n465 VDD.t779 28.565
R2057 VDD.n460 VDD.t172 28.565
R2058 VDD.n460 VDD.t168 28.565
R2059 VDD.n461 VDD.t170 28.565
R2060 VDD.n461 VDD.t1076 28.565
R2061 VDD.n463 VDD.t1578 28.565
R2062 VDD.n463 VDD.t1576 28.565
R2063 VDD.n351 VDD.t941 28.565
R2064 VDD.n351 VDD.t939 28.565
R2065 VDD.n346 VDD.t1432 28.565
R2066 VDD.n346 VDD.t1430 28.565
R2067 VDD.n347 VDD.t1422 28.565
R2068 VDD.n347 VDD.t1402 28.565
R2069 VDD.n349 VDD.t1400 28.565
R2070 VDD.n349 VDD.t1398 28.565
R2071 VDD.n360 VDD.t1438 28.565
R2072 VDD.n360 VDD.t1582 28.565
R2073 VDD.n355 VDD.t1199 28.565
R2074 VDD.n355 VDD.t1197 28.565
R2075 VDD.n447 VDD.t1203 28.565
R2076 VDD.n447 VDD.t1134 28.565
R2077 VDD.n449 VDD.t651 28.565
R2078 VDD.n449 VDD.t649 28.565
R2079 VDD.n450 VDD.t192 28.565
R2080 VDD.n450 VDD.t416 28.565
R2081 VDD.n452 VDD.t883 28.565
R2082 VDD.n452 VDD.t881 28.565
R2083 VDD.n430 VDD.t767 28.565
R2084 VDD.n430 VDD.t1028 28.565
R2085 VDD.n425 VDD.t717 28.565
R2086 VDD.n425 VDD.t554 28.565
R2087 VDD.n442 VDD.t580 28.565
R2088 VDD.n442 VDD.t578 28.565
R2089 VDD.n437 VDD.t78 28.565
R2090 VDD.n437 VDD.t76 28.565
R2091 VDD.n438 VDD.t74 28.565
R2092 VDD.n438 VDD.t689 28.565
R2093 VDD.n440 VDD.t1026 28.565
R2094 VDD.n440 VDD.t1024 28.565
R2095 VDD.n372 VDD.t1511 28.565
R2096 VDD.n372 VDD.t1509 28.565
R2097 VDD.n367 VDD.t291 28.565
R2098 VDD.n367 VDD.t289 28.565
R2099 VDD.n384 VDD.t1389 28.565
R2100 VDD.n384 VDD.t967 28.565
R2101 VDD.n379 VDD.t1371 28.565
R2102 VDD.n379 VDD.t1373 28.565
R2103 VDD.n380 VDD.t1375 28.565
R2104 VDD.n380 VDD.t1513 28.565
R2105 VDD.n382 VDD.t174 28.565
R2106 VDD.n382 VDD.t178 28.565
R2107 VDD.n404 VDD.t635 28.565
R2108 VDD.n404 VDD.t627 28.565
R2109 VDD.n399 VDD.t116 28.565
R2110 VDD.n399 VDD.t1086 28.565
R2111 VDD.n416 VDD.t1010 28.565
R2112 VDD.n416 VDD.t1471 28.565
R2113 VDD.n411 VDD.t1426 28.565
R2114 VDD.n411 VDD.t1424 28.565
R2115 VDD.n412 VDD.t1428 28.565
R2116 VDD.n412 VDD.t1414 28.565
R2117 VDD.n414 VDD.t1406 28.565
R2118 VDD.n414 VDD.t1418 28.565
R2119 VDD.n394 VDD.t1092 28.565
R2120 VDD.n394 VDD.t442 28.565
R2121 VDD.n389 VDD.t619 28.565
R2122 VDD.n389 VDD.t617 28.565
R2123 VDD.n390 VDD.t615 28.565
R2124 VDD.n390 VDD.t637 28.565
R2125 VDD.n392 VDD.t633 28.565
R2126 VDD.n392 VDD.t641 28.565
R2127 VDD.n871 VDD.t224 28.565
R2128 VDD.n871 VDD.t222 28.565
R2129 VDD.n866 VDD.t1175 28.565
R2130 VDD.n866 VDD.t1101 28.565
R2131 VDD.n867 VDD.t1099 28.565
R2132 VDD.n867 VDD.t1385 28.565
R2133 VDD.n869 VDD.t613 28.565
R2134 VDD.n869 VDD.t1186 28.565
R2135 VDD.n880 VDD.t1629 28.565
R2136 VDD.n880 VDD.t1383 28.565
R2137 VDD.n875 VDD.t396 28.565
R2138 VDD.n875 VDD.t891 28.565
R2139 VDD.n876 VDD.t584 28.565
R2140 VDD.n876 VDD.t1412 28.565
R2141 VDD.n878 VDD.t1410 28.565
R2142 VDD.n878 VDD.t1408 28.565
R2143 VDD.n520 VDD.t1565 23.418
R2144 VDD.n659 VDD.t764 23.418
R2145 VDD.n747 VDD.t1143 23.418
R2146 VDD.n813 VDD.t955 23.418
R2147 VDD.n136 VDD.t595 23.418
R2148 VDD.n201 VDD.t531 23.418
R2149 VDD.n269 VDD.t622 23.418
R2150 VDD.n330 VDD.t1494 23.418
R2151 VDD.n9 VDD.t272 23.317
R2152 VDD.n0 VDD.t746 23.317
R2153 VDD.n890 VDD.t1622 23.317
R2154 VDD.n899 VDD.t728 23.317
R2155 VDD.n52 VDD.t1153 23.317
R2156 VDD.n43 VDD.t1462 23.317
R2157 VDD.n34 VDD.t179 23.317
R2158 VDD.n25 VDD.t144 23.317
R2159 VDD.n17 VDD.t864 23.317
R2160 VDD.n468 VDD.t1415 23.317
R2161 VDD.n459 VDD.t854 23.317
R2162 VDD.n345 VDD.t940 23.317
R2163 VDD.n378 VDD.t1388 23.317
R2164 VDD.n410 VDD.t1009 23.317
R2165 VDD.n388 VDD.t1091 23.317
R2166 VDD.n865 VDD.t223 23.317
R2167 VDD.n874 VDD.t1628 23.317
R2168 VDD.n436 VDD.t579 23.316
R2169 VDD.n454 VDD.t1202 23.316
R2170 VDD.n916 VDD.t1502 22.813
R2171 VDD.n946 VDD.t838 22.813
R2172 VDD.n977 VDD.t28 22.813
R2173 VDD.n1007 VDD.t486 22.813
R2174 VDD.n597 VDD.t1442 22.813
R2175 VDD.n684 VDD.t509 22.813
R2176 VDD.n763 VDD.t286 22.813
R2177 VDD.n843 VDD.t252 22.813
R2178 VDD.n17 VDD.t134 20.186
R2179 VDD.n436 VDD.t1023 20.186
R2180 VDD.n454 VDD.t880 20.186
R2181 VDD.n9 VDD.t652 20.183
R2182 VDD.n0 VDD.t820 20.183
R2183 VDD.n890 VDD.t1464 20.183
R2184 VDD.n899 VDD.t1460 20.183
R2185 VDD.n52 VDD.t361 20.183
R2186 VDD.n43 VDD.t868 20.183
R2187 VDD.n34 VDD.t229 20.183
R2188 VDD.n25 VDD.t900 20.183
R2189 VDD.n468 VDD.t644 20.183
R2190 VDD.n459 VDD.t1575 20.183
R2191 VDD.n345 VDD.t1397 20.183
R2192 VDD.n378 VDD.t177 20.183
R2193 VDD.n410 VDD.t1417 20.183
R2194 VDD.n388 VDD.t640 20.183
R2195 VDD.n865 VDD.t1185 20.183
R2196 VDD.n874 VDD.t1407 20.183
R2197 VDD.n523 VDD.t1521 14.284
R2198 VDD.n528 VDD.t1335 14.284
R2199 VDD.n505 VDD.t202 14.284
R2200 VDD.n510 VDD.t305 14.284
R2201 VDD.n279 VDD.t1209 14.284
R2202 VDD.n286 VDD.t825 14.284
R2203 VDD.n211 VDD.t990 14.284
R2204 VDD.n935 VDD.t663 14.284
R2205 VDD.n146 VDD.t1499 14.284
R2206 VDD.n967 VDD.t937 14.284
R2207 VDD.n79 VDD.t1225 14.284
R2208 VDD.n995 VDD.t1264 14.284
R2209 VDD.n581 VDD.t298 14.284
R2210 VDD.n574 VDD.t998 14.284
R2211 VDD.n609 VDD.t538 14.284
R2212 VDD.n614 VDD.t827 14.284
R2213 VDD.n644 VDD.t3 14.284
R2214 VDD.n649 VDD.t796 14.284
R2215 VDD.n678 VDD.t1602 14.284
R2216 VDD.n564 VDD.t1453 14.284
R2217 VDD.n733 VDD.t1142 14.284
R2218 VDD.n738 VDD.t1126 14.284
R2219 VDD.n720 VDD.t669 14.284
R2220 VDD.n725 VDD.t1276 14.284
R2221 VDD.n554 VDD.t1321 14.284
R2222 VDD.n547 VDD.t1598 14.284
R2223 VDD.n817 VDD.t952 14.284
R2224 VDD.n822 VDD.t1558 14.284
R2225 VDD.n798 VDD.t847 14.284
R2226 VDD.n803 VDD.t21 14.284
R2227 VDD.n537 VDD.t1349 14.284
R2228 VDD.n855 VDD.t504 14.284
R2229 VDD.n84 VDD.t897 14.284
R2230 VDD.n89 VDD.t1312 14.284
R2231 VDD.n121 VDD.t352 14.284
R2232 VDD.n126 VDD.t1116 14.284
R2233 VDD.n150 VDD.t528 14.284
R2234 VDD.n155 VDD.t380 14.284
R2235 VDD.n186 VDD.t1489 14.284
R2236 VDD.n191 VDD.t1436 14.284
R2237 VDD.n215 VDD.t1525 14.284
R2238 VDD.n220 VDD.t114 14.284
R2239 VDD.n254 VDD.t13 14.284
R2240 VDD.n259 VDD.t473 14.284
R2241 VDD.n334 VDD.t1491 14.284
R2242 VDD.n339 VDD.t1020 14.284
R2243 VDD.n315 VDD.t340 14.284
R2244 VDD.n320 VDD.t1231 14.284
R2245 VDD.n359 VDD.t691 14.284
R2246 VDD.n354 VDD.t1201 14.284
R2247 VDD.n429 VDD.t574 14.284
R2248 VDD.n424 VDD.t719 14.284
R2249 VDD.n371 VDD.t1473 14.284
R2250 VDD.n366 VDD.t969 14.284
R2251 VDD.n403 VDD.t639 14.284
R2252 VDD.n398 VDD.t1090 14.284
R2253 VDD.n522 VDD.t1566 14.282
R2254 VDD.n522 VDD.t184 14.282
R2255 VDD.n527 VDD.t1347 14.282
R2256 VDD.n527 VDD.t1343 14.282
R2257 VDD.n504 VDD.t570 14.282
R2258 VDD.n504 VDD.t91 14.282
R2259 VDD.n509 VDD.t853 14.282
R2260 VDD.n509 VDD.t303 14.282
R2261 VDD.n276 VDD.t1213 14.282
R2262 VDD.n276 VDD.t1211 14.282
R2263 VDD.n283 VDD.t823 14.282
R2264 VDD.n283 VDD.t1207 14.282
R2265 VDD.n208 VDD.t992 14.282
R2266 VDD.n208 VDD.t994 14.282
R2267 VDD.n932 VDD.t216 14.282
R2268 VDD.n932 VDD.t665 14.282
R2269 VDD.n143 VDD.t1497 14.282
R2270 VDD.n143 VDD.t508 14.282
R2271 VDD.n964 VDD.t1140 14.282
R2272 VDD.n964 VDD.t1138 14.282
R2273 VDD.n76 VDD.t1227 14.282
R2274 VDD.n76 VDD.t1229 14.282
R2275 VDD.n992 VDD.t1245 14.282
R2276 VDD.n992 VDD.t1266 14.282
R2277 VDD.n578 VDD.t935 14.282
R2278 VDD.n578 VDD.t296 14.282
R2279 VDD.n571 VDD.t1000 14.282
R2280 VDD.n571 VDD.t713 14.282
R2281 VDD.n608 VDD.t765 14.282
R2282 VDD.n608 VDD.t763 14.282
R2283 VDD.n613 VDD.t270 14.282
R2284 VDD.n613 VDD.t1481 14.282
R2285 VDD.n643 VDD.t1112 14.282
R2286 VDD.n643 VDD.t5 14.282
R2287 VDD.n648 VDD.t794 14.282
R2288 VDD.n648 VDD.t1182 14.282
R2289 VDD.n675 VDD.t682 14.282
R2290 VDD.n675 VDD.t1604 14.282
R2291 VDD.n561 VDD.t1455 14.282
R2292 VDD.n561 VDD.t1451 14.282
R2293 VDD.n732 VDD.t1144 14.282
R2294 VDD.n732 VDD.t1193 14.282
R2295 VDD.n737 VDD.t699 14.282
R2296 VDD.n737 VDD.t433 14.282
R2297 VDD.n719 VDD.t609 14.282
R2298 VDD.n719 VDD.t1008 14.282
R2299 VDD.n724 VDD.t1274 14.282
R2300 VDD.n724 VDD.t1122 14.282
R2301 VDD.n551 VDD.t1319 14.282
R2302 VDD.n551 VDD.t1323 14.282
R2303 VDD.n544 VDD.t1600 14.282
R2304 VDD.n544 VDD.t1215 14.282
R2305 VDD.n816 VDD.t956 14.282
R2306 VDD.n816 VDD.t873 14.282
R2307 VDD.n821 VDD.t1166 14.282
R2308 VDD.n821 VDD.t259 14.282
R2309 VDD.n797 VDD.t773 14.282
R2310 VDD.n797 VDD.t923 14.282
R2311 VDD.n802 VDD.t1040 14.282
R2312 VDD.n802 VDD.t19 14.282
R2313 VDD.n534 VDD.t1355 14.282
R2314 VDD.n534 VDD.t1357 14.282
R2315 VDD.n852 VDD.t506 14.282
R2316 VDD.n852 VDD.t1097 14.282
R2317 VDD.n83 VDD.t596 14.282
R2318 VDD.n83 VDD.t899 14.282
R2319 VDD.n88 VDD.t1310 14.282
R2320 VDD.n88 VDD.t1300 14.282
R2321 VDD.n120 VDD.t370 14.282
R2322 VDD.n120 VDD.t368 14.282
R2323 VDD.n125 VDD.t1539 14.282
R2324 VDD.n125 VDD.t1537 14.282
R2325 VDD.n149 VDD.t532 14.282
R2326 VDD.n149 VDD.t530 14.282
R2327 VDD.n154 VDD.t979 14.282
R2328 VDD.n154 VDD.t679 14.282
R2329 VDD.n185 VDD.t210 14.282
R2330 VDD.n185 VDD.t208 14.282
R2331 VDD.n190 VDD.t703 14.282
R2332 VDD.n190 VDD.t701 14.282
R2333 VDD.n214 VDD.t623 14.282
R2334 VDD.n214 VDD.t1527 14.282
R2335 VDD.n219 VDD.t107 14.282
R2336 VDD.n219 VDD.t105 14.282
R2337 VDD.n253 VDD.t917 14.282
R2338 VDD.n253 VDD.t15 14.282
R2339 VDD.n258 VDD.t281 14.282
R2340 VDD.n258 VDD.t279 14.282
R2341 VDD.n333 VDD.t1495 14.282
R2342 VDD.n333 VDD.t1493 14.282
R2343 VDD.n338 VDD.t1016 14.282
R2344 VDD.n338 VDD.t960 14.282
R2345 VDD.n314 VDD.t333 14.282
R2346 VDD.n314 VDD.t329 14.282
R2347 VDD.n319 VDD.t1256 14.282
R2348 VDD.n319 VDD.t1260 14.282
R2349 VDD.n358 VDD.t1584 14.282
R2350 VDD.n358 VDD.t693 14.282
R2351 VDD.n353 VDD.t671 14.282
R2352 VDD.n353 VDD.t1205 14.282
R2353 VDD.n428 VDD.t137 14.282
R2354 VDD.n428 VDD.t576 14.282
R2355 VDD.n423 VDD.t562 14.282
R2356 VDD.n423 VDD.t582 14.282
R2357 VDD.n370 VDD.t257 14.282
R2358 VDD.n370 VDD.t176 14.282
R2359 VDD.n365 VDD.t1572 14.282
R2360 VDD.n365 VDD.t1574 14.282
R2361 VDD.n402 VDD.t631 14.282
R2362 VDD.n402 VDD.t625 14.282
R2363 VDD.n397 VDD.t440 14.282
R2364 VDD.n397 VDD.t118 14.282
R2365 VDD.n434 VDD.t948 8.293
R2366 VDD.n376 VDD.t62 8.293
R2367 VDD.n408 VDD.t755 8.293
R2368 VDD.n364 VDD.t294 8.293
R2369 VDD.n516 VDD.t1532 4.524
R2370 VDD.n517 VDD.t610 4.524
R2371 VDD.n519 VDD.t599 4.524
R2372 VDD.n518 VDD.t434 4.524
R2373 VDD.n655 VDD.t92 4.524
R2374 VDD.n656 VDD.t93 4.524
R2375 VDD.n658 VDD.t240 4.524
R2376 VDD.n657 VDD.t241 4.524
R2377 VDD.n743 VDD.t488 4.524
R2378 VDD.n744 VDD.t1171 4.524
R2379 VDD.n746 VDD.t397 4.524
R2380 VDD.n745 VDD.t1609 4.524
R2381 VDD.n809 VDD.t453 4.524
R2382 VDD.n810 VDD.t454 4.524
R2383 VDD.n812 VDD.t52 4.524
R2384 VDD.n811 VDD.t53 4.524
R2385 VDD.n132 VDD.t1069 4.524
R2386 VDD.n133 VDD.t400 4.524
R2387 VDD.n135 VDD.t1155 4.524
R2388 VDD.n134 VDD.t1519 4.524
R2389 VDD.n197 VDD.t471 4.524
R2390 VDD.n198 VDD.t470 4.524
R2391 VDD.n200 VDD.t1420 4.524
R2392 VDD.n199 VDD.t1419 4.524
R2393 VDD.n265 VDD.t957 4.524
R2394 VDD.n266 VDD.t451 4.524
R2395 VDD.n268 VDD.t54 4.524
R2396 VDD.n267 VDD.t101 4.524
R2397 VDD.n326 VDD.t686 4.524
R2398 VDD.n327 VDD.t393 4.524
R2399 VDD.n329 VDD.t988 4.524
R2400 VDD.n328 VDD.t987 4.524
R2401 VDD.n363 VDD.n362 4.331
R2402 VDD.n433 VDD.n432 4.331
R2403 VDD.n375 VDD.n374 4.331
R2404 VDD.n407 VDD.n406 4.331
R2405 VDD.n532 VDD.n526 4.276
R2406 VDD.n514 VDD.n508 4.276
R2407 VDD.n618 VDD.n612 4.276
R2408 VDD.n653 VDD.n647 4.276
R2409 VDD.n742 VDD.n736 4.276
R2410 VDD.n729 VDD.n723 4.276
R2411 VDD.n826 VDD.n820 4.276
R2412 VDD.n807 VDD.n801 4.276
R2413 VDD.n93 VDD.n87 4.276
R2414 VDD.n130 VDD.n124 4.276
R2415 VDD.n159 VDD.n153 4.276
R2416 VDD.n195 VDD.n189 4.276
R2417 VDD.n224 VDD.n218 4.276
R2418 VDD.n263 VDD.n257 4.276
R2419 VDD.n343 VDD.n337 4.276
R2420 VDD.n324 VDD.n318 4.276
R2421 VDD.n68 VDD.t142 2.932
R2422 VDD.n525 VDD.n524 2.451
R2423 VDD.n507 VDD.n506 2.451
R2424 VDD.n611 VDD.n610 2.451
R2425 VDD.n646 VDD.n645 2.451
R2426 VDD.n735 VDD.n734 2.451
R2427 VDD.n722 VDD.n721 2.451
R2428 VDD.n819 VDD.n818 2.451
R2429 VDD.n800 VDD.n799 2.451
R2430 VDD.n86 VDD.n85 2.451
R2431 VDD.n123 VDD.n122 2.451
R2432 VDD.n152 VDD.n151 2.451
R2433 VDD.n188 VDD.n187 2.451
R2434 VDD.n217 VDD.n216 2.451
R2435 VDD.n256 VDD.n255 2.451
R2436 VDD.n336 VDD.n335 2.451
R2437 VDD.n317 VDD.n316 2.451
R2438 VDD.n361 VDD.n360 2.451
R2439 VDD.n431 VDD.n430 2.451
R2440 VDD.n373 VDD.n372 2.451
R2441 VDD.n405 VDD.n404 2.451
R2442 VDD.n530 VDD.n529 2.449
R2443 VDD.n512 VDD.n511 2.449
R2444 VDD.n616 VDD.n615 2.449
R2445 VDD.n651 VDD.n650 2.449
R2446 VDD.n740 VDD.n739 2.449
R2447 VDD.n727 VDD.n726 2.449
R2448 VDD.n824 VDD.n823 2.449
R2449 VDD.n805 VDD.n804 2.449
R2450 VDD.n91 VDD.n90 2.449
R2451 VDD.n128 VDD.n127 2.449
R2452 VDD.n157 VDD.n156 2.449
R2453 VDD.n193 VDD.n192 2.449
R2454 VDD.n222 VDD.n221 2.449
R2455 VDD.n261 VDD.n260 2.449
R2456 VDD.n341 VDD.n340 2.449
R2457 VDD.n322 VDD.n321 2.449
R2458 VDD.n356 VDD.n355 2.449
R2459 VDD.n426 VDD.n425 2.449
R2460 VDD.n368 VDD.n367 2.449
R2461 VDD.n400 VDD.n399 2.449
R2462 VDD.n279 VDD.n278 2.195
R2463 VDD.n286 VDD.n285 2.195
R2464 VDD.n211 VDD.n210 2.195
R2465 VDD.n935 VDD.n934 2.195
R2466 VDD.n146 VDD.n145 2.195
R2467 VDD.n967 VDD.n966 2.195
R2468 VDD.n79 VDD.n78 2.195
R2469 VDD.n995 VDD.n994 2.195
R2470 VDD.n581 VDD.n580 2.195
R2471 VDD.n574 VDD.n573 2.195
R2472 VDD.n678 VDD.n677 2.195
R2473 VDD.n564 VDD.n563 2.195
R2474 VDD.n554 VDD.n553 2.195
R2475 VDD.n547 VDD.n546 2.195
R2476 VDD.n537 VDD.n536 2.195
R2477 VDD.n855 VDD.n854 2.195
R2478 VDD.n287 VDD.n283 1.72
R2479 VDD.n936 VDD.n932 1.72
R2480 VDD.n968 VDD.n964 1.72
R2481 VDD.n996 VDD.n992 1.72
R2482 VDD.n575 VDD.n571 1.72
R2483 VDD.n565 VDD.n561 1.72
R2484 VDD.n548 VDD.n544 1.72
R2485 VDD.n856 VDD.n852 1.72
R2486 VDD.n280 VDD.n276 1.698
R2487 VDD.n212 VDD.n208 1.698
R2488 VDD.n147 VDD.n143 1.698
R2489 VDD.n80 VDD.n76 1.698
R2490 VDD.n582 VDD.n578 1.698
R2491 VDD.n679 VDD.n675 1.698
R2492 VDD.n555 VDD.n551 1.698
R2493 VDD.n538 VDD.n534 1.698
R2494 VDD.n278 VDD.n277 1.651
R2495 VDD.n285 VDD.n284 1.651
R2496 VDD.n210 VDD.n209 1.651
R2497 VDD.n934 VDD.n933 1.651
R2498 VDD.n145 VDD.n144 1.651
R2499 VDD.n966 VDD.n965 1.651
R2500 VDD.n78 VDD.n77 1.651
R2501 VDD.n994 VDD.n993 1.651
R2502 VDD.n580 VDD.n579 1.651
R2503 VDD.n573 VDD.n572 1.651
R2504 VDD.n677 VDD.n676 1.651
R2505 VDD.n563 VDD.n562 1.651
R2506 VDD.n553 VDD.n552 1.651
R2507 VDD.n546 VDD.n545 1.651
R2508 VDD.n536 VDD.n535 1.651
R2509 VDD.n854 VDD.n853 1.651
R2510 VDD.n12 VDD.n10 1.564
R2511 VDD.n3 VDD.n1 1.564
R2512 VDD.n496 VDD.n494 1.564
R2513 VDD.n485 VDD.n483 1.564
R2514 VDD.n275 VDD.n273 1.564
R2515 VDD.n207 VDD.n205 1.564
R2516 VDD.n142 VDD.n140 1.564
R2517 VDD.n75 VDD.n73 1.564
R2518 VDD.n65 VDD.n63 1.564
R2519 VDD.n887 VDD.n885 1.564
R2520 VDD.n896 VDD.n894 1.564
R2521 VDD.n55 VDD.n53 1.564
R2522 VDD.n46 VDD.n44 1.564
R2523 VDD.n37 VDD.n35 1.564
R2524 VDD.n586 VDD.n584 1.564
R2525 VDD.n28 VDD.n26 1.564
R2526 VDD.n621 VDD.n619 1.564
R2527 VDD.n625 VDD.n623 1.564
R2528 VDD.n570 VDD.n568 1.564
R2529 VDD.n697 VDD.n695 1.564
R2530 VDD.n707 VDD.n705 1.564
R2531 VDD.n560 VDD.n558 1.564
R2532 VDD.n776 VDD.n774 1.564
R2533 VDD.n785 VDD.n783 1.564
R2534 VDD.n543 VDD.n541 1.564
R2535 VDD.n20 VDD.n18 1.564
R2536 VDD.n109 VDD.n107 1.564
R2537 VDD.n103 VDD.n101 1.564
R2538 VDD.n162 VDD.n160 1.564
R2539 VDD.n171 VDD.n169 1.564
R2540 VDD.n246 VDD.n244 1.564
R2541 VDD.n228 VDD.n226 1.564
R2542 VDD.n292 VDD.n290 1.564
R2543 VDD.n296 VDD.n294 1.564
R2544 VDD.n471 VDD.n469 1.564
R2545 VDD.n462 VDD.n460 1.564
R2546 VDD.n348 VDD.n346 1.564
R2547 VDD.n451 VDD.n449 1.564
R2548 VDD.n439 VDD.n437 1.564
R2549 VDD.n381 VDD.n379 1.564
R2550 VDD.n413 VDD.n411 1.564
R2551 VDD.n391 VDD.n389 1.564
R2552 VDD.n868 VDD.n866 1.564
R2553 VDD.n877 VDD.n875 1.564
R2554 VDD.n903 VDD.n902 1.496
R2555 VDD.n902 VDD.n901 1.232
R2556 VDD.n72 VDD.n71 1.224
R2557 VDD.n418 VDD.n8 1.212
R2558 VDD.n1031 VDD.n1030 1.054
R2559 VDD.n1032 VDD.n1031 1.031
R2560 VDD.n526 VDD.n522 0.922
R2561 VDD.n531 VDD.n527 0.922
R2562 VDD.n508 VDD.n504 0.922
R2563 VDD.n513 VDD.n509 0.922
R2564 VDD.n612 VDD.n608 0.922
R2565 VDD.n617 VDD.n613 0.922
R2566 VDD.n647 VDD.n643 0.922
R2567 VDD.n652 VDD.n648 0.922
R2568 VDD.n736 VDD.n732 0.922
R2569 VDD.n741 VDD.n737 0.922
R2570 VDD.n723 VDD.n719 0.922
R2571 VDD.n728 VDD.n724 0.922
R2572 VDD.n820 VDD.n816 0.922
R2573 VDD.n825 VDD.n821 0.922
R2574 VDD.n801 VDD.n797 0.922
R2575 VDD.n806 VDD.n802 0.922
R2576 VDD.n87 VDD.n83 0.922
R2577 VDD.n92 VDD.n88 0.922
R2578 VDD.n124 VDD.n120 0.922
R2579 VDD.n129 VDD.n125 0.922
R2580 VDD.n153 VDD.n149 0.922
R2581 VDD.n158 VDD.n154 0.922
R2582 VDD.n189 VDD.n185 0.922
R2583 VDD.n194 VDD.n190 0.922
R2584 VDD.n218 VDD.n214 0.922
R2585 VDD.n223 VDD.n219 0.922
R2586 VDD.n257 VDD.n253 0.922
R2587 VDD.n262 VDD.n258 0.922
R2588 VDD.n337 VDD.n333 0.922
R2589 VDD.n342 VDD.n338 0.922
R2590 VDD.n318 VDD.n314 0.922
R2591 VDD.n323 VDD.n319 0.922
R2592 VDD.n362 VDD.n358 0.922
R2593 VDD.n357 VDD.n353 0.922
R2594 VDD.n432 VDD.n428 0.922
R2595 VDD.n427 VDD.n423 0.922
R2596 VDD.n374 VDD.n370 0.922
R2597 VDD.n369 VDD.n365 0.922
R2598 VDD.n406 VDD.n402 0.922
R2599 VDD.n401 VDD.n397 0.922
R2600 VDD.n525 VDD.n523 0.921
R2601 VDD.n530 VDD.n528 0.921
R2602 VDD.n507 VDD.n505 0.921
R2603 VDD.n512 VDD.n510 0.921
R2604 VDD.n611 VDD.n609 0.921
R2605 VDD.n616 VDD.n614 0.921
R2606 VDD.n646 VDD.n644 0.921
R2607 VDD.n651 VDD.n649 0.921
R2608 VDD.n735 VDD.n733 0.921
R2609 VDD.n740 VDD.n738 0.921
R2610 VDD.n722 VDD.n720 0.921
R2611 VDD.n727 VDD.n725 0.921
R2612 VDD.n819 VDD.n817 0.921
R2613 VDD.n824 VDD.n822 0.921
R2614 VDD.n800 VDD.n798 0.921
R2615 VDD.n805 VDD.n803 0.921
R2616 VDD.n86 VDD.n84 0.921
R2617 VDD.n91 VDD.n89 0.921
R2618 VDD.n123 VDD.n121 0.921
R2619 VDD.n128 VDD.n126 0.921
R2620 VDD.n152 VDD.n150 0.921
R2621 VDD.n157 VDD.n155 0.921
R2622 VDD.n188 VDD.n186 0.921
R2623 VDD.n193 VDD.n191 0.921
R2624 VDD.n217 VDD.n215 0.921
R2625 VDD.n222 VDD.n220 0.921
R2626 VDD.n256 VDD.n254 0.921
R2627 VDD.n261 VDD.n259 0.921
R2628 VDD.n336 VDD.n334 0.921
R2629 VDD.n341 VDD.n339 0.921
R2630 VDD.n317 VDD.n315 0.921
R2631 VDD.n322 VDD.n320 0.921
R2632 VDD.n361 VDD.n359 0.921
R2633 VDD.n356 VDD.n354 0.921
R2634 VDD.n431 VDD.n429 0.921
R2635 VDD.n426 VDD.n424 0.921
R2636 VDD.n373 VDD.n371 0.921
R2637 VDD.n368 VDD.n366 0.921
R2638 VDD.n405 VDD.n403 0.921
R2639 VDD.n400 VDD.n398 0.921
R2640 VDD.n14 VDD.n12 0.85
R2641 VDD.n5 VDD.n3 0.85
R2642 VDD.n67 VDD.n65 0.85
R2643 VDD.n889 VDD.n887 0.85
R2644 VDD.n898 VDD.n896 0.85
R2645 VDD.n57 VDD.n55 0.85
R2646 VDD.n48 VDD.n46 0.85
R2647 VDD.n39 VDD.n37 0.85
R2648 VDD.n30 VDD.n28 0.85
R2649 VDD.n22 VDD.n20 0.85
R2650 VDD.n473 VDD.n471 0.85
R2651 VDD.n464 VDD.n462 0.85
R2652 VDD.n350 VDD.n348 0.85
R2653 VDD.n453 VDD.n451 0.85
R2654 VDD.n441 VDD.n439 0.85
R2655 VDD.n383 VDD.n381 0.85
R2656 VDD.n415 VDD.n413 0.85
R2657 VDD.n393 VDD.n391 0.85
R2658 VDD.n870 VDD.n868 0.85
R2659 VDD.n879 VDD.n877 0.85
R2660 VDD.n280 VDD.n279 0.806
R2661 VDD.n212 VDD.n211 0.806
R2662 VDD.n147 VDD.n146 0.806
R2663 VDD.n80 VDD.n79 0.806
R2664 VDD.n582 VDD.n581 0.806
R2665 VDD.n679 VDD.n678 0.806
R2666 VDD.n555 VDD.n554 0.806
R2667 VDD.n538 VDD.n537 0.806
R2668 VDD.n287 VDD.n286 0.778
R2669 VDD.n936 VDD.n935 0.778
R2670 VDD.n968 VDD.n967 0.778
R2671 VDD.n996 VDD.n995 0.778
R2672 VDD.n575 VDD.n574 0.778
R2673 VDD.n565 VDD.n564 0.778
R2674 VDD.n548 VDD.n547 0.778
R2675 VDD.n856 VDD.n855 0.778
R2676 VDD.n16 VDD.n15 0.747
R2677 VDD.n12 VDD.n11 0.747
R2678 VDD.n14 VDD.n13 0.747
R2679 VDD.n7 VDD.n6 0.747
R2680 VDD.n3 VDD.n2 0.747
R2681 VDD.n5 VDD.n4 0.747
R2682 VDD.n491 VDD.n490 0.747
R2683 VDD.n496 VDD.n495 0.747
R2684 VDD.n479 VDD.n478 0.747
R2685 VDD.n485 VDD.n484 0.747
R2686 VDD.n924 VDD.n923 0.747
R2687 VDD.n275 VDD.n274 0.747
R2688 VDD.n953 VDD.n952 0.747
R2689 VDD.n207 VDD.n206 0.747
R2690 VDD.n984 VDD.n983 0.747
R2691 VDD.n142 VDD.n141 0.747
R2692 VDD.n1019 VDD.n1018 0.747
R2693 VDD.n75 VDD.n74 0.747
R2694 VDD.n62 VDD.n61 0.747
R2695 VDD.n65 VDD.n64 0.747
R2696 VDD.n67 VDD.n66 0.747
R2697 VDD.n884 VDD.n883 0.747
R2698 VDD.n887 VDD.n886 0.747
R2699 VDD.n889 VDD.n888 0.747
R2700 VDD.n893 VDD.n892 0.747
R2701 VDD.n896 VDD.n895 0.747
R2702 VDD.n898 VDD.n897 0.747
R2703 VDD.n59 VDD.n58 0.747
R2704 VDD.n55 VDD.n54 0.747
R2705 VDD.n57 VDD.n56 0.747
R2706 VDD.n50 VDD.n49 0.747
R2707 VDD.n46 VDD.n45 0.747
R2708 VDD.n48 VDD.n47 0.747
R2709 VDD.n41 VDD.n40 0.747
R2710 VDD.n37 VDD.n36 0.747
R2711 VDD.n39 VDD.n38 0.747
R2712 VDD.n590 VDD.n589 0.747
R2713 VDD.n586 VDD.n585 0.747
R2714 VDD.n32 VDD.n31 0.747
R2715 VDD.n28 VDD.n27 0.747
R2716 VDD.n30 VDD.n29 0.747
R2717 VDD.n638 VDD.n637 0.747
R2718 VDD.n621 VDD.n620 0.747
R2719 VDD.n629 VDD.n628 0.747
R2720 VDD.n625 VDD.n624 0.747
R2721 VDD.n667 VDD.n666 0.747
R2722 VDD.n570 VDD.n569 0.747
R2723 VDD.n713 VDD.n712 0.747
R2724 VDD.n697 VDD.n696 0.747
R2725 VDD.n701 VDD.n700 0.747
R2726 VDD.n707 VDD.n706 0.747
R2727 VDD.n757 VDD.n756 0.747
R2728 VDD.n560 VDD.n559 0.747
R2729 VDD.n791 VDD.n790 0.747
R2730 VDD.n776 VDD.n775 0.747
R2731 VDD.n779 VDD.n778 0.747
R2732 VDD.n785 VDD.n784 0.747
R2733 VDD.n834 VDD.n833 0.747
R2734 VDD.n543 VDD.n542 0.747
R2735 VDD.n24 VDD.n23 0.747
R2736 VDD.n20 VDD.n19 0.747
R2737 VDD.n22 VDD.n21 0.747
R2738 VDD.n115 VDD.n114 0.747
R2739 VDD.n109 VDD.n108 0.747
R2740 VDD.n97 VDD.n96 0.747
R2741 VDD.n103 VDD.n102 0.747
R2742 VDD.n179 VDD.n178 0.747
R2743 VDD.n162 VDD.n161 0.747
R2744 VDD.n165 VDD.n164 0.747
R2745 VDD.n171 VDD.n170 0.747
R2746 VDD.n240 VDD.n239 0.747
R2747 VDD.n246 VDD.n245 0.747
R2748 VDD.n232 VDD.n231 0.747
R2749 VDD.n228 VDD.n227 0.747
R2750 VDD.n309 VDD.n308 0.747
R2751 VDD.n292 VDD.n291 0.747
R2752 VDD.n300 VDD.n299 0.747
R2753 VDD.n296 VDD.n295 0.747
R2754 VDD.n475 VDD.n474 0.747
R2755 VDD.n471 VDD.n470 0.747
R2756 VDD.n473 VDD.n472 0.747
R2757 VDD.n466 VDD.n465 0.747
R2758 VDD.n462 VDD.n461 0.747
R2759 VDD.n464 VDD.n463 0.747
R2760 VDD.n352 VDD.n351 0.747
R2761 VDD.n348 VDD.n347 0.747
R2762 VDD.n350 VDD.n349 0.747
R2763 VDD.n448 VDD.n447 0.747
R2764 VDD.n451 VDD.n450 0.747
R2765 VDD.n453 VDD.n452 0.747
R2766 VDD.n443 VDD.n442 0.747
R2767 VDD.n439 VDD.n438 0.747
R2768 VDD.n441 VDD.n440 0.747
R2769 VDD.n385 VDD.n384 0.747
R2770 VDD.n381 VDD.n380 0.747
R2771 VDD.n383 VDD.n382 0.747
R2772 VDD.n417 VDD.n416 0.747
R2773 VDD.n413 VDD.n412 0.747
R2774 VDD.n415 VDD.n414 0.747
R2775 VDD.n395 VDD.n394 0.747
R2776 VDD.n391 VDD.n390 0.747
R2777 VDD.n393 VDD.n392 0.747
R2778 VDD.n872 VDD.n871 0.747
R2779 VDD.n868 VDD.n867 0.747
R2780 VDD.n870 VDD.n869 0.747
R2781 VDD.n881 VDD.n880 0.747
R2782 VDD.n877 VDD.n876 0.747
R2783 VDD.n879 VDD.n878 0.747
R2784 VDD.n493 VDD.n489 0.689
R2785 VDD.n481 VDD.n477 0.689
R2786 VDD.n926 VDD.n922 0.689
R2787 VDD.n955 VDD.n951 0.689
R2788 VDD.n986 VDD.n982 0.689
R2789 VDD.n1021 VDD.n1017 0.689
R2790 VDD.n592 VDD.n588 0.689
R2791 VDD.n640 VDD.n636 0.689
R2792 VDD.n631 VDD.n627 0.689
R2793 VDD.n669 VDD.n665 0.689
R2794 VDD.n715 VDD.n711 0.689
R2795 VDD.n703 VDD.n699 0.689
R2796 VDD.n759 VDD.n755 0.689
R2797 VDD.n793 VDD.n789 0.689
R2798 VDD.n781 VDD.n777 0.689
R2799 VDD.n836 VDD.n832 0.689
R2800 VDD.n117 VDD.n113 0.689
R2801 VDD.n99 VDD.n95 0.689
R2802 VDD.n181 VDD.n177 0.689
R2803 VDD.n167 VDD.n163 0.689
R2804 VDD.n242 VDD.n238 0.689
R2805 VDD.n234 VDD.n230 0.689
R2806 VDD.n311 VDD.n307 0.689
R2807 VDD.n302 VDD.n298 0.689
R2808 VDD.n526 VDD.n525 0.686
R2809 VDD.n531 VDD.n530 0.686
R2810 VDD.n508 VDD.n507 0.686
R2811 VDD.n513 VDD.n512 0.686
R2812 VDD.n612 VDD.n611 0.686
R2813 VDD.n617 VDD.n616 0.686
R2814 VDD.n647 VDD.n646 0.686
R2815 VDD.n652 VDD.n651 0.686
R2816 VDD.n736 VDD.n735 0.686
R2817 VDD.n741 VDD.n740 0.686
R2818 VDD.n723 VDD.n722 0.686
R2819 VDD.n728 VDD.n727 0.686
R2820 VDD.n820 VDD.n819 0.686
R2821 VDD.n825 VDD.n824 0.686
R2822 VDD.n801 VDD.n800 0.686
R2823 VDD.n806 VDD.n805 0.686
R2824 VDD.n87 VDD.n86 0.686
R2825 VDD.n92 VDD.n91 0.686
R2826 VDD.n124 VDD.n123 0.686
R2827 VDD.n129 VDD.n128 0.686
R2828 VDD.n153 VDD.n152 0.686
R2829 VDD.n158 VDD.n157 0.686
R2830 VDD.n189 VDD.n188 0.686
R2831 VDD.n194 VDD.n193 0.686
R2832 VDD.n218 VDD.n217 0.686
R2833 VDD.n223 VDD.n222 0.686
R2834 VDD.n257 VDD.n256 0.686
R2835 VDD.n262 VDD.n261 0.686
R2836 VDD.n337 VDD.n336 0.686
R2837 VDD.n342 VDD.n341 0.686
R2838 VDD.n318 VDD.n317 0.686
R2839 VDD.n323 VDD.n322 0.686
R2840 VDD.n362 VDD.n361 0.686
R2841 VDD.n357 VDD.n356 0.686
R2842 VDD.n432 VDD.n431 0.686
R2843 VDD.n427 VDD.n426 0.686
R2844 VDD.n374 VDD.n373 0.686
R2845 VDD.n369 VDD.n368 0.686
R2846 VDD.n406 VDD.n405 0.686
R2847 VDD.n401 VDD.n400 0.686
R2848 VDD.n492 VDD.n491 0.571
R2849 VDD.n480 VDD.n479 0.571
R2850 VDD.n985 VDD.n984 0.571
R2851 VDD.n591 VDD.n590 0.571
R2852 VDD.n630 VDD.n629 0.571
R2853 VDD.n668 VDD.n667 0.571
R2854 VDD.n714 VDD.n713 0.571
R2855 VDD.n792 VDD.n791 0.571
R2856 VDD.n780 VDD.n779 0.571
R2857 VDD.n116 VDD.n115 0.571
R2858 VDD.n166 VDD.n165 0.571
R2859 VDD.n241 VDD.n240 0.571
R2860 VDD.n233 VDD.n232 0.571
R2861 VDD.n301 VDD.n300 0.571
R2862 VDD.n925 VDD.n924 0.57
R2863 VDD.n639 VDD.n638 0.57
R2864 VDD.n758 VDD.n757 0.57
R2865 VDD.n310 VDD.n309 0.57
R2866 VDD.n954 VDD.n953 0.569
R2867 VDD.n1020 VDD.n1019 0.569
R2868 VDD.n702 VDD.n701 0.569
R2869 VDD.n835 VDD.n834 0.569
R2870 VDD.n98 VDD.n97 0.569
R2871 VDD.n180 VDD.n179 0.569
R2872 VDD VDD.n8 0.557
R2873 VDD.n446 VDD.n445 0.476
R2874 VDD.n840 VDD.n543 0.452
R2875 VDD.n921 VDD.n275 0.452
R2876 VDD.n642 VDD.n621 0.452
R2877 VDD.n184 VDD.n162 0.452
R2878 VDD.n950 VDD.n207 0.452
R2879 VDD.n1014 VDD.n75 0.452
R2880 VDD.n761 VDD.n560 0.452
R2881 VDD.n313 VDD.n292 0.452
R2882 VDD.n708 VDD.n707 0.452
R2883 VDD.n104 VDD.n103 0.452
R2884 VDD.n981 VDD.n142 0.451
R2885 VDD.n595 VDD.n586 0.451
R2886 VDD.n672 VDD.n570 0.451
R2887 VDD.n718 VDD.n697 0.451
R2888 VDD.n796 VDD.n776 0.451
R2889 VDD.n486 VDD.n485 0.451
R2890 VDD.n786 VDD.n785 0.451
R2891 VDD.n626 VDD.n625 0.45
R2892 VDD.n297 VDD.n296 0.45
R2893 VDD.n229 VDD.n228 0.45
R2894 VDD.n172 VDD.n171 0.449
R2895 VDD.n110 VDD.n109 0.449
R2896 VDD.n422 VDD.n421 0.424
R2897 VDD.n497 VDD.n496 0.419
R2898 VDD.n247 VDD.n246 0.419
R2899 VDD.n282 VDD.n281 0.4
R2900 VDD.n289 VDD.n288 0.4
R2901 VDD.n970 VDD.n969 0.4
R2902 VDD.n82 VDD.n81 0.4
R2903 VDD.n577 VDD.n576 0.4
R2904 VDD.n681 VDD.n680 0.4
R2905 VDD.n567 VDD.n566 0.4
R2906 VDD.n557 VDD.n556 0.4
R2907 VDD.n550 VDD.n549 0.4
R2908 VDD.n540 VDD.n539 0.4
R2909 VDD.n858 VDD.n857 0.4
R2910 VDD VDD.n1032 0.367
R2911 VDD.n863 VDD.n862 0.303
R2912 VDD.n905 VDD.n904 0.286
R2913 VDD.n904 VDD.n903 0.283
R2914 VDD.n446 VDD.n422 0.273
R2915 VDD.n488 VDD.n487 0.271
R2916 VDD.n788 VDD.n787 0.271
R2917 VDD.n237 VDD.n236 0.271
R2918 VDD.n634 VDD.n633 0.271
R2919 VDD.n106 VDD.n105 0.271
R2920 VDD.n175 VDD.n174 0.271
R2921 VDD.n305 VDD.n304 0.271
R2922 VDD.n710 VDD.n709 0.271
R2923 VDD.n445 VDD.n435 0.252
R2924 VDD.n752 VDD.n751 0.244
R2925 VDD.n420 VDD.n419 0.233
R2926 VDD.n282 VDD.n280 0.23
R2927 VDD.n213 VDD.n212 0.23
R2928 VDD.n148 VDD.n147 0.23
R2929 VDD.n82 VDD.n80 0.23
R2930 VDD.n583 VDD.n582 0.23
R2931 VDD.n681 VDD.n679 0.23
R2932 VDD.n557 VDD.n555 0.23
R2933 VDD.n540 VDD.n538 0.23
R2934 VDD.n1028 VDD.n1027 0.228
R2935 VDD.n289 VDD.n287 0.218
R2936 VDD.n937 VDD.n936 0.218
R2937 VDD.n970 VDD.n968 0.218
R2938 VDD.n997 VDD.n996 0.218
R2939 VDD.n577 VDD.n575 0.218
R2940 VDD.n567 VDD.n565 0.218
R2941 VDD.n550 VDD.n548 0.218
R2942 VDD.n858 VDD.n856 0.218
R2943 VDD.n1032 VDD.n16 0.208
R2944 VDD.n8 VDD.n7 0.208
R2945 VDD.n70 VDD.n62 0.208
R2946 VDD.n891 VDD.n884 0.208
R2947 VDD.n900 VDD.n893 0.208
R2948 VDD.n60 VDD.n59 0.208
R2949 VDD.n51 VDD.n50 0.208
R2950 VDD.n42 VDD.n41 0.208
R2951 VDD.n33 VDD.n32 0.208
R2952 VDD.n1031 VDD.n24 0.208
R2953 VDD.n476 VDD.n475 0.208
R2954 VDD.n467 VDD.n466 0.208
R2955 VDD.n458 VDD.n352 0.208
R2956 VDD.n455 VDD.n448 0.208
R2957 VDD.n444 VDD.n443 0.208
R2958 VDD.n386 VDD.n385 0.208
R2959 VDD.n419 VDD.n417 0.208
R2960 VDD.n396 VDD.n395 0.208
R2961 VDD.n873 VDD.n872 0.208
R2962 VDD.n882 VDD.n881 0.208
R2963 VDD.n363 VDD.n357 0.203
R2964 VDD.n433 VDD.n427 0.203
R2965 VDD.n375 VDD.n369 0.203
R2966 VDD.n407 VDD.n401 0.203
R2967 VDD.n1032 VDD.n14 0.195
R2968 VDD.n8 VDD.n5 0.195
R2969 VDD.n70 VDD.n67 0.195
R2970 VDD.n891 VDD.n889 0.195
R2971 VDD.n900 VDD.n898 0.195
R2972 VDD.n60 VDD.n57 0.195
R2973 VDD.n51 VDD.n48 0.195
R2974 VDD.n42 VDD.n39 0.195
R2975 VDD.n33 VDD.n30 0.195
R2976 VDD.n1031 VDD.n22 0.195
R2977 VDD.n476 VDD.n473 0.195
R2978 VDD.n467 VDD.n464 0.195
R2979 VDD.n458 VDD.n350 0.195
R2980 VDD.n455 VDD.n453 0.195
R2981 VDD.n444 VDD.n441 0.195
R2982 VDD.n386 VDD.n383 0.195
R2983 VDD.n419 VDD.n415 0.195
R2984 VDD.n396 VDD.n393 0.195
R2985 VDD.n873 VDD.n870 0.195
R2986 VDD.n882 VDD.n879 0.195
R2987 VDD.n387 VDD.n377 0.195
R2988 VDD.n458 VDD.n457 0.193
R2989 VDD.n664 VDD.n663 0.186
R2990 VDD.n961 VDD.n960 0.186
R2991 VDD.n864 VDD.n863 0.185
R2992 VDD.n753 VDD.n752 0.185
R2993 VDD.n930 VDD.n929 0.184
R2994 VDD.n829 VDD.n828 0.182
R2995 VDD.n673 VDD.n672 0.182
R2996 VDD.n841 VDD.n840 0.182
R2997 VDD.n990 VDD.n989 0.18
R2998 VDD.n532 VDD.n531 0.179
R2999 VDD.n514 VDD.n513 0.179
R3000 VDD.n618 VDD.n617 0.179
R3001 VDD.n653 VDD.n652 0.179
R3002 VDD.n742 VDD.n741 0.179
R3003 VDD.n729 VDD.n728 0.179
R3004 VDD.n826 VDD.n825 0.179
R3005 VDD.n807 VDD.n806 0.179
R3006 VDD.n1026 VDD.n72 0.179
R3007 VDD.n93 VDD.n92 0.179
R3008 VDD.n130 VDD.n129 0.179
R3009 VDD.n159 VDD.n158 0.179
R3010 VDD.n195 VDD.n194 0.179
R3011 VDD.n224 VDD.n223 0.179
R3012 VDD.n263 VDD.n262 0.179
R3013 VDD.n343 VDD.n342 0.179
R3014 VDD.n324 VDD.n323 0.179
R3015 VDD.n1014 VDD.n1013 0.177
R3016 VDD.n981 VDD.n980 0.176
R3017 VDD.n332 VDD.n325 0.175
R3018 VDD.n203 VDD.n196 0.175
R3019 VDD.n271 VDD.n264 0.175
R3020 VDD.n661 VDD.n654 0.175
R3021 VDD.n138 VDD.n131 0.175
R3022 VDD.n533 VDD.n515 0.175
R3023 VDD.n815 VDD.n808 0.174
R3024 VDD.n950 VDD.n949 0.174
R3025 VDD.n921 VDD.n920 0.173
R3026 VDD.n1027 VDD.n51 0.17
R3027 VDD.n828 VDD.n827 0.168
R3028 VDD.n731 VDD.n730 0.168
R3029 VDD.n1030 VDD.n33 0.167
R3030 VDD.n72 VDD.n60 0.167
R3031 VDD.n1028 VDD.n42 0.166
R3032 VDD.n762 VDD.n761 0.164
R3033 VDD.n654 VDD.n642 0.162
R3034 VDD.n730 VDD.n718 0.162
R3035 VDD.n808 VDD.n796 0.162
R3036 VDD.n196 VDD.n184 0.162
R3037 VDD.n325 VDD.n313 0.162
R3038 VDD.n515 VDD.n503 0.161
R3039 VDD.n131 VDD.n119 0.161
R3040 VDD.n264 VDD.n252 0.161
R3041 VDD.n596 VDD.n595 0.16
R3042 VDD.n663 VDD.n662 0.155
R3043 VDD.n515 VDD.n514 0.142
R3044 VDD.n654 VDD.n653 0.142
R3045 VDD.n730 VDD.n729 0.142
R3046 VDD.n808 VDD.n807 0.142
R3047 VDD.n131 VDD.n130 0.142
R3048 VDD.n196 VDD.n195 0.142
R3049 VDD.n264 VDD.n263 0.142
R3050 VDD.n325 VDD.n324 0.142
R3051 VDD.n1029 VDD.n1028 0.137
R3052 VDD.n421 VDD.n420 0.131
R3053 VDD.n860 VDD.n533 0.128
R3054 VDD.n990 VDD.n139 0.128
R3055 VDD.n961 VDD.n204 0.128
R3056 VDD.n930 VDD.n272 0.128
R3057 VDD.n906 VDD.n344 0.128
R3058 VDD.n662 VDD.n618 0.125
R3059 VDD.n750 VDD.n742 0.125
R3060 VDD.n139 VDD.n93 0.125
R3061 VDD.n204 VDD.n159 0.125
R3062 VDD.n272 VDD.n224 0.125
R3063 VDD.n344 VDD.n343 0.125
R3064 VDD.n533 VDD.n532 0.124
R3065 VDD.n827 VDD.n826 0.123
R3066 VDD.n903 VDD.n882 0.114
R3067 VDD.n457 VDD.n456 0.114
R3068 VDD.n904 VDD.n873 0.113
R3069 VDD.n1026 VDD.n1025 0.105
R3070 VDD.n862 VDD.n476 0.1
R3071 VDD.n863 VDD.n467 0.1
R3072 VDD.n973 VDD.n963 0.098
R3073 VDD.n687 VDD.n674 0.098
R3074 VDD.n692 VDD.n691 0.097
R3075 VDD.n766 VDD.n765 0.097
R3076 VDD.n771 VDD.n770 0.097
R3077 VDD.n850 VDD.n849 0.097
R3078 VDD.n910 VDD.n909 0.095
R3079 VDD.n604 VDD.n603 0.095
R3080 VDD.n1010 VDD.n1009 0.093
R3081 VDD.n848 VDD.n847 0.086
R3082 VDD.n690 VDD.n689 0.085
R3083 VDD.n1005 VDD.n1004 0.082
R3084 VDD.n976 VDD.n975 0.082
R3085 VDD.n945 VDD.n944 0.081
R3086 VDD.n914 VDD.n913 0.081
R3087 VDD.n769 VDD.n768 0.077
R3088 VDD.n601 VDD.n600 0.076
R3089 VDD.n456 VDD.n446 0.068
R3090 VDD.n422 VDD.n387 0.061
R3091 VDD.n862 VDD.n861 0.057
R3092 VDD.n387 VDD.n386 0.055
R3093 VDD.n419 VDD.n418 0.053
R3094 VDD.n445 VDD.n444 0.053
R3095 VDD.n864 VDD.n458 0.051
R3096 VDD.n906 VDD.n905 0.048
R3097 VDD.n861 VDD.n860 0.044
R3098 VDD.n501 VDD.n500 0.043
R3099 VDD.n250 VDD.n249 0.042
R3100 VDD.n838 VDD.n830 0.042
R3101 VDD.n1011 VDD.n1006 0.042
R3102 VDD.n605 VDD.n602 0.042
R3103 VDD.n1023 VDD.n1015 0.041
R3104 VDD.n911 VDD.n908 0.041
R3105 VDD.n942 VDD.n941 0.041
R3106 VDD.n958 VDD.n956 0.04
R3107 VDD.n1002 VDD.n1001 0.04
R3108 VDD.n421 VDD.n396 0.039
R3109 VDD.n456 VDD.n455 0.037
R3110 VDD.n905 VDD.n864 0.032
R3111 VDD.n499 VDD.n497 0.03
R3112 VDD.n248 VDD.n247 0.03
R3113 VDD.n457 VDD.n363 0.03
R3114 VDD.n435 VDD.n433 0.03
R3115 VDD.n377 VDD.n375 0.03
R3116 VDD.n409 VDD.n407 0.03
R3117 VDD.n907 VDD.n906 0.026
R3118 VDD.n962 VDD.n961 0.026
R3119 VDD.n991 VDD.n990 0.026
R3120 VDD.n860 VDD.n859 0.025
R3121 VDD.n931 VDD.n930 0.025
R3122 VDD.n663 VDD.n607 0.022
R3123 VDD.n828 VDD.n773 0.022
R3124 VDD.n859 VDD.n858 0.021
R3125 VDD.n836 VDD.n835 0.021
R3126 VDD.n945 VDD.n213 0.02
R3127 VDD.n976 VDD.n148 0.02
R3128 VDD.n694 VDD.n567 0.02
R3129 VDD.n768 VDD.n557 0.02
R3130 VDD.n773 VDD.n550 0.02
R3131 VDD.n914 VDD.n282 0.02
R3132 VDD.n907 VDD.n289 0.02
R3133 VDD.n607 VDD.n577 0.02
R3134 VDD.n847 VDD.n540 0.02
R3135 VDD.n1005 VDD.n82 0.02
R3136 VDD.n926 VDD.n925 0.02
R3137 VDD.n955 VDD.n954 0.02
R3138 VDD.n1021 VDD.n1020 0.02
R3139 VDD.n640 VDD.n639 0.02
R3140 VDD.n703 VDD.n702 0.02
R3141 VDD.n759 VDD.n758 0.02
R3142 VDD.n99 VDD.n98 0.02
R3143 VDD.n181 VDD.n180 0.02
R3144 VDD.n311 VDD.n310 0.02
R3145 VDD.n481 VDD.n480 0.019
R3146 VDD.n986 VDD.n985 0.019
R3147 VDD.n592 VDD.n591 0.019
R3148 VDD.n631 VDD.n630 0.019
R3149 VDD.n669 VDD.n668 0.019
R3150 VDD.n715 VDD.n714 0.019
R3151 VDD.n793 VDD.n792 0.019
R3152 VDD.n781 VDD.n780 0.019
R3153 VDD.n302 VDD.n301 0.019
R3154 VDD.n600 VDD.n583 0.019
R3155 VDD.n493 VDD.n492 0.018
R3156 VDD.n117 VDD.n116 0.018
R3157 VDD.n167 VDD.n166 0.018
R3158 VDD.n242 VDD.n241 0.018
R3159 VDD.n234 VDD.n233 0.018
R3160 VDD.n752 VDD.n694 0.016
R3161 VDD.n502 VDD.n493 0.011
R3162 VDD.n486 VDD.n481 0.011
R3163 VDD.n938 VDD.n937 0.011
R3164 VDD.n971 VDD.n970 0.011
R3165 VDD.n988 VDD.n986 0.011
R3166 VDD.n998 VDD.n997 0.011
R3167 VDD.n594 VDD.n592 0.011
R3168 VDD.n632 VDD.n631 0.011
R3169 VDD.n671 VDD.n669 0.011
R3170 VDD.n682 VDD.n681 0.011
R3171 VDD.n717 VDD.n715 0.011
R3172 VDD.n760 VDD.n759 0.011
R3173 VDD.n795 VDD.n793 0.011
R3174 VDD.n786 VDD.n781 0.011
R3175 VDD.n1027 VDD.n1026 0.011
R3176 VDD.n118 VDD.n117 0.011
R3177 VDD.n173 VDD.n167 0.011
R3178 VDD.n251 VDD.n242 0.011
R3179 VDD.n235 VDD.n234 0.011
R3180 VDD.n312 VDD.n311 0.011
R3181 VDD.n303 VDD.n302 0.011
R3182 VDD.n928 VDD.n926 0.01
R3183 VDD.n641 VDD.n640 0.01
R3184 VDD.n704 VDD.n703 0.01
R3185 VDD.n100 VDD.n99 0.01
R3186 VDD.n182 VDD.n181 0.01
R3187 VDD.n1011 VDD.n1010 0.009
R3188 VDD.n958 VDD.n955 0.009
R3189 VDD.n1022 VDD.n1021 0.009
R3190 VDD.n1030 VDD.n1029 0.009
R3191 VDD.n837 VDD.n836 0.008
R3192 VDD.n972 VDD.n971 0.007
R3193 VDD.n1003 VDD.n1000 0.007
R3194 VDD.n751 VDD.n731 0.006
R3195 VDD.n911 VDD.n910 0.005
R3196 VDD.n683 VDD.n682 0.005
R3197 VDD.n940 VDD.n938 0.005
R3198 VDD.n605 VDD.n604 0.005
R3199 VDD.n838 VDD.n837 0.003
R3200 VDD.n173 VDD.n172 0.003
R3201 VDD.n943 VDD.n940 0.003
R3202 VDD.n1003 VDD.n1002 0.003
R3203 VDD.n501 VDD.n499 0.002
R3204 VDD.n118 VDD.n112 0.002
R3205 VDD.n235 VDD.n229 0.002
R3206 VDD.n632 VDD.n626 0.002
R3207 VDD.n303 VDD.n297 0.002
R3208 VDD.n919 VDD.n918 0.002
R3209 VDD.n420 VDD.n409 0.001
R3210 VDD.n973 VDD.n972 0.001
R3211 VDD.n1023 VDD.n1022 0.001
R3212 VDD.n250 VDD.n248 0.001
R3213 VDD.n751 VDD.n750 0.001
R3214 VDD.n1000 VDD.n998 0.001
R3215 VDD.n687 VDD.n686 0.001
R3216 VDD.n606 VDD.n605 0.001
R3217 VDD.n943 VDD.n942 0.001
R3218 VDD.n693 VDD.n692 0.001
R3219 VDD.n708 VDD.n704 0.001
R3220 VDD.n767 VDD.n766 0.001
R3221 VDD.n772 VDD.n771 0.001
R3222 VDD.n851 VDD.n850 0.001
R3223 VDD.n104 VDD.n100 0.001
R3224 VDD.n183 VDD.n182 0.001
R3225 VDD.n750 VDD.n749 0.001
R3226 VDD.n901 VDD.n900 0.001
R3227 VDD.n902 VDD.n891 0.001
R3228 VDD.n71 VDD.n70 0.001
R3229 VDD.n139 VDD.n138 0.001
R3230 VDD.n662 VDD.n661 0.001
R3231 VDD.n204 VDD.n203 0.001
R3232 VDD.n272 VDD.n271 0.001
R3233 VDD.n918 VDD.n915 0.001
R3234 VDD.n845 VDD.n842 0.001
R3235 VDD.n846 VDD.n845 0.001
R3236 VDD.n502 VDD.n501 0.001
R3237 VDD.n940 VDD.n939 0.001
R3238 VDD.n1031 VDD.n17 0.001
R3239 VDD.n1032 VDD.n9 0.001
R3240 VDD.n8 VDD.n0 0.001
R3241 VDD.n891 VDD.n890 0.001
R3242 VDD.n900 VDD.n899 0.001
R3243 VDD.n60 VDD.n52 0.001
R3244 VDD.n51 VDD.n43 0.001
R3245 VDD.n42 VDD.n34 0.001
R3246 VDD.n33 VDD.n25 0.001
R3247 VDD.n476 VDD.n468 0.001
R3248 VDD.n467 VDD.n459 0.001
R3249 VDD.n458 VDD.n345 0.001
R3250 VDD.n386 VDD.n378 0.001
R3251 VDD.n419 VDD.n410 0.001
R3252 VDD.n396 VDD.n388 0.001
R3253 VDD.n873 VDD.n865 0.001
R3254 VDD.n882 VDD.n874 0.001
R3255 VDD.n444 VDD.n436 0.001
R3256 VDD.n455 VDD.n454 0.001
R3257 VDD.n70 VDD.n69 0.001
R3258 VDD.n112 VDD.n110 0.001
R3259 VDD.n1000 VDD.n999 0.001
R3260 VDD.n846 VDD.n841 0.001
R3261 VDD.n839 VDD.n829 0.001
R3262 VDD.n689 VDD.n688 0.001
R3263 VDD.n1003 VDD.n991 0.001
R3264 VDD.n1013 VDD.n1012 0.001
R3265 VDD.n1025 VDD.n1024 0.001
R3266 VDD.n943 VDD.n931 0.001
R3267 VDD.n960 VDD.n959 0.001
R3268 VDD.n913 VDD.n912 0.001
R3269 VDD.n920 VDD.n919 0.001
R3270 VDD.n606 VDD.n601 0.001
R3271 VDD.n686 VDD.n683 0.001
R3272 VDD.n503 VDD.n502 0.001
R3273 VDD.n119 VDD.n118 0.001
R3274 VDD.n252 VDD.n251 0.001
R3275 VDD.n1012 VDD.n1011 0.001
R3276 VDD.n709 VDD.n708 0.001
R3277 VDD.n105 VDD.n104 0.001
R3278 VDD.n851 VDD.n848 0.001
R3279 VDD.n693 VDD.n690 0.001
R3280 VDD.n929 VDD.n928 0.001
R3281 VDD.n487 VDD.n486 0.001
R3282 VDD.n633 VDD.n632 0.001
R3283 VDD.n787 VDD.n786 0.001
R3284 VDD.n688 VDD.n673 0.001
R3285 VDD.n671 VDD.n664 0.001
R3286 VDD.n975 VDD.n974 0.001
R3287 VDD.n989 VDD.n988 0.001
R3288 VDD.n304 VDD.n303 0.001
R3289 VDD.n174 VDD.n173 0.001
R3290 VDD.n236 VDD.n235 0.001
R3291 VDD.n772 VDD.n769 0.001
R3292 VDD.n767 VDD.n762 0.001
R3293 VDD.n760 VDD.n753 0.001
R3294 VDD.n594 VDD.n587 0.001
R3295 VDD.n839 VDD.n838 0.001
R3296 VDD.n980 VDD.n979 0.001
R3297 VDD.n949 VDD.n948 0.001
R3298 VDD.n944 VDD.n943 0.001
R3299 VDD.n1004 VDD.n1003 0.001
R3300 VDD.n183 VDD.n175 0.001
R3301 VDD.n641 VDD.n634 0.001
R3302 VDD.n312 VDD.n305 0.001
R3303 VDD.n717 VDD.n710 0.001
R3304 VDD.n795 VDD.n788 0.001
R3305 VDD.n502 VDD.n488 0.001
R3306 VDD.n118 VDD.n106 0.001
R3307 VDD.n251 VDD.n237 0.001
R3308 VDD.n599 VDD.n596 0.001
R3309 VDD.n859 VDD.n851 0.001
R3310 VDD.n344 VDD.n332 0.001
R3311 VDD.n912 VDD.n911 0.001
R3312 VDD.n827 VDD.n815 0.001
R3313 VDD.n251 VDD.n250 0.001
R3314 VDD.n974 VDD.n962 0.001
R3315 VDD.n1024 VDD.n1023 0.001
R3316 VDD.n672 VDD.n671 0.001
R3317 VDD.n988 VDD.n981 0.001
R3318 VDD.n928 VDD.n921 0.001
R3319 VDD.n761 VDD.n760 0.001
R3320 VDD.n1024 VDD.n1014 0.001
R3321 VDD.n959 VDD.n950 0.001
R3322 VDD.n595 VDD.n594 0.001
R3323 VDD.n313 VDD.n312 0.001
R3324 VDD.n840 VDD.n839 0.001
R3325 VDD.n718 VDD.n717 0.001
R3326 VDD.n796 VDD.n795 0.001
R3327 VDD.n642 VDD.n641 0.001
R3328 VDD.n184 VDD.n183 0.001
R3329 VDD.n979 VDD.n976 0.001
R3330 VDD.n948 VDD.n945 0.001
R3331 VDD.n847 VDD.n846 0.001
R3332 VDD.n912 VDD.n907 0.001
R3333 VDD.n919 VDD.n914 0.001
R3334 VDD.n1012 VDD.n1005 0.001
R3335 VDD.n773 VDD.n772 0.001
R3336 VDD.n768 VDD.n767 0.001
R3337 VDD.n607 VDD.n606 0.001
R3338 VDD.n694 VDD.n693 0.001
R3339 VDD.n600 VDD.n599 0.001
R3340 VDD.n959 VDD.n958 0.001
R3341 VDD.n974 VDD.n973 0.001
R3342 VDD.n688 VDD.n687 0.001
R3343 a_12822_1097.n2 a_12822_1097.t6 318.922
R3344 a_12822_1097.n1 a_12822_1097.t7 273.935
R3345 a_12822_1097.n1 a_12822_1097.t4 273.935
R3346 a_12822_1097.n2 a_12822_1097.t5 269.116
R3347 a_12822_1097.n4 a_12822_1097.n0 193.227
R3348 a_12822_1097.t6 a_12822_1097.n1 179.142
R3349 a_12822_1097.n3 a_12822_1097.n2 106.999
R3350 a_12822_1097.t0 a_12822_1097.n4 28.568
R3351 a_12822_1097.n0 a_12822_1097.t2 28.565
R3352 a_12822_1097.n0 a_12822_1097.t3 28.565
R3353 a_12822_1097.n3 a_12822_1097.t1 18.149
R3354 a_12822_1097.n4 a_12822_1097.n3 3.726
R3355 a_13249_404.t0 a_13249_404.n0 14.282
R3356 a_13249_404.n0 a_13249_404.t10 14.282
R3357 a_13249_404.n0 a_13249_404.n9 0.999
R3358 a_13249_404.n6 a_13249_404.n8 0.575
R3359 a_13249_404.n9 a_13249_404.n6 0.2
R3360 a_13249_404.n9 a_13249_404.t5 16.058
R3361 a_13249_404.n8 a_13249_404.n7 0.999
R3362 a_13249_404.n7 a_13249_404.t3 14.282
R3363 a_13249_404.n7 a_13249_404.t1 14.282
R3364 a_13249_404.n8 a_13249_404.t2 16.058
R3365 a_13249_404.n6 a_13249_404.n4 0.227
R3366 a_13249_404.n4 a_13249_404.n5 1.511
R3367 a_13249_404.n5 a_13249_404.t8 14.282
R3368 a_13249_404.n5 a_13249_404.t11 14.282
R3369 a_13249_404.n4 a_13249_404.n1 0.669
R3370 a_13249_404.n1 a_13249_404.n2 0.001
R3371 a_13249_404.n1 a_13249_404.n3 267.767
R3372 a_13249_404.n3 a_13249_404.t6 14.282
R3373 a_13249_404.n3 a_13249_404.t7 14.282
R3374 a_13249_404.n2 a_13249_404.t9 14.282
R3375 a_13249_404.n2 a_13249_404.t4 14.282
R3376 a_13367_404.n0 a_13367_404.t4 14.282
R3377 a_13367_404.t0 a_13367_404.n0 14.282
R3378 a_13367_404.n0 a_13367_404.n16 90.416
R3379 a_13367_404.n16 a_13367_404.n15 50.575
R3380 a_13367_404.n16 a_13367_404.n12 74.302
R3381 a_13367_404.n15 a_13367_404.n14 157.665
R3382 a_13367_404.n14 a_13367_404.t1 8.7
R3383 a_13367_404.n14 a_13367_404.t6 8.7
R3384 a_13367_404.n15 a_13367_404.n13 122.999
R3385 a_13367_404.n13 a_13367_404.t2 14.282
R3386 a_13367_404.n13 a_13367_404.t3 14.282
R3387 a_13367_404.n12 a_13367_404.n11 90.436
R3388 a_13367_404.n11 a_13367_404.t7 14.282
R3389 a_13367_404.n11 a_13367_404.t5 14.282
R3390 a_13367_404.n12 a_13367_404.n1 216.635
R3391 a_13367_404.n1 a_13367_404.n3 16.411
R3392 a_13367_404.n3 a_13367_404.t10 198.921
R3393 a_13367_404.t10 a_13367_404.t8 415.315
R3394 a_13367_404.t8 a_13367_404.n10 214.335
R3395 a_13367_404.n10 a_13367_404.t18 80.333
R3396 a_13367_404.n10 a_13367_404.t14 214.335
R3397 a_13367_404.n3 a_13367_404.n9 861.987
R3398 a_13367_404.n9 a_13367_404.n4 560.726
R3399 a_13367_404.n9 a_13367_404.n8 65.07
R3400 a_13367_404.n8 a_13367_404.n7 6.615
R3401 a_13367_404.n7 a_13367_404.t16 93.989
R3402 a_13367_404.n8 a_13367_404.n6 97.816
R3403 a_13367_404.n6 a_13367_404.t12 80.333
R3404 a_13367_404.n6 a_13367_404.t19 394.151
R3405 a_13367_404.t19 a_13367_404.n5 269.523
R3406 a_13367_404.n5 a_13367_404.t13 160.666
R3407 a_13367_404.n5 a_13367_404.t21 269.523
R3408 a_13367_404.n7 a_13367_404.t20 198.043
R3409 a_13367_404.n4 a_13367_404.t11 294.653
R3410 a_13367_404.n4 a_13367_404.t15 111.663
R3411 a_13367_404.n1 a_13367_404.t22 217.716
R3412 a_13367_404.t22 a_13367_404.t23 415.315
R3413 a_13367_404.t23 a_13367_404.n2 214.335
R3414 a_13367_404.n2 a_13367_404.t17 80.333
R3415 a_13367_404.n2 a_13367_404.t9 214.335
R3416 a_16227_42.n0 a_16227_42.t8 214.335
R3417 a_16227_42.t10 a_16227_42.n0 214.335
R3418 a_16227_42.n1 a_16227_42.t10 143.851
R3419 a_16227_42.n1 a_16227_42.t9 135.658
R3420 a_16227_42.n0 a_16227_42.t7 80.333
R3421 a_16227_42.n2 a_16227_42.t2 28.565
R3422 a_16227_42.n2 a_16227_42.t6 28.565
R3423 a_16227_42.n4 a_16227_42.t5 28.565
R3424 a_16227_42.n4 a_16227_42.t3 28.565
R3425 a_16227_42.t0 a_16227_42.n7 28.565
R3426 a_16227_42.n7 a_16227_42.t1 28.565
R3427 a_16227_42.n6 a_16227_42.t4 9.714
R3428 a_16227_42.n7 a_16227_42.n6 1.003
R3429 a_16227_42.n5 a_16227_42.n3 0.833
R3430 a_16227_42.n3 a_16227_42.n2 0.653
R3431 a_16227_42.n5 a_16227_42.n4 0.653
R3432 a_16227_42.n6 a_16227_42.n5 0.341
R3433 a_16227_42.n3 a_16227_42.n1 0.032
R3434 a_16817_n395.t6 a_16817_n395.t7 574.43
R3435 a_16817_n395.n0 a_16817_n395.t5 285.109
R3436 a_16817_n395.n2 a_16817_n395.n1 197.217
R3437 a_16817_n395.n4 a_16817_n395.n3 192.754
R3438 a_16817_n395.n0 a_16817_n395.t4 160.666
R3439 a_16817_n395.n1 a_16817_n395.t6 160.666
R3440 a_16817_n395.n1 a_16817_n395.n0 114.829
R3441 a_16817_n395.n3 a_16817_n395.t2 28.568
R3442 a_16817_n395.t3 a_16817_n395.n4 28.565
R3443 a_16817_n395.n4 a_16817_n395.t1 28.565
R3444 a_16817_n395.n2 a_16817_n395.t0 18.838
R3445 a_16817_n395.n3 a_16817_n395.n2 1.129
R3446 a_2969_1600.n16 a_2969_1600.n15 3522.62
R3447 a_2969_1600.n7 a_2969_1600.n6 501.28
R3448 a_2969_1600.t17 a_2969_1600.t13 437.233
R3449 a_2969_1600.t19 a_2969_1600.t11 415.315
R3450 a_2969_1600.t4 a_2969_1600.n4 313.873
R3451 a_2969_1600.n6 a_2969_1600.t18 294.986
R3452 a_2969_1600.n3 a_2969_1600.t6 272.288
R3453 a_2969_1600.n7 a_2969_1600.t14 236.01
R3454 a_2969_1600.n10 a_2969_1600.t17 216.627
R3455 a_2969_1600.n8 a_2969_1600.t19 216.111
R3456 a_2969_1600.n9 a_2969_1600.t7 214.686
R3457 a_2969_1600.t13 a_2969_1600.n9 214.686
R3458 a_2969_1600.n2 a_2969_1600.t15 214.335
R3459 a_2969_1600.t11 a_2969_1600.n2 214.335
R3460 a_2969_1600.n17 a_2969_1600.n0 192.754
R3461 a_2969_1600.n5 a_2969_1600.t4 190.152
R3462 a_2969_1600.n5 a_2969_1600.t5 190.152
R3463 a_2969_1600.n3 a_2969_1600.t16 160.666
R3464 a_2969_1600.n4 a_2969_1600.t9 160.666
R3465 a_2969_1600.n8 a_2969_1600.n7 148.428
R3466 a_2969_1600.n6 a_2969_1600.t10 110.859
R3467 a_2969_1600.n4 a_2969_1600.n3 96.129
R3468 a_2969_1600.n9 a_2969_1600.t8 80.333
R3469 a_2969_1600.n2 a_2969_1600.t12 80.333
R3470 a_2969_1600.t14 a_2969_1600.n5 80.333
R3471 a_2969_1600.t1 a_2969_1600.n17 28.568
R3472 a_2969_1600.n0 a_2969_1600.t2 28.565
R3473 a_2969_1600.n0 a_2969_1600.t3 28.565
R3474 a_2969_1600.n16 a_2969_1600.t0 18.522
R3475 a_2969_1600.n15 a_2969_1600.n14 5.25
R3476 a_2969_1600.n14 a_2969_1600.n13 3.293
R3477 a_2969_1600.n10 a_2969_1600.n8 2.923
R3478 a_2969_1600.n17 a_2969_1600.n16 1.168
R3479 a_2969_1600.n11 a_2969_1600.n10 0.708
R3480 a_2969_1600.n14 a_2969_1600.n12 0.681
R3481 a_2969_1600.n12 a_2969_1600.n1 0.003
R3482 a_2969_1600.n12 a_2969_1600.n11 0.001
R3483 a_7112_290.n1 a_7112_290.t6 318.922
R3484 a_7112_290.n0 a_7112_290.t7 274.739
R3485 a_7112_290.n0 a_7112_290.t5 274.739
R3486 a_7112_290.n1 a_7112_290.t4 269.116
R3487 a_7112_290.t6 a_7112_290.n0 179.946
R3488 a_7112_290.n2 a_7112_290.n1 105.178
R3489 a_7112_290.n3 a_7112_290.t2 29.444
R3490 a_7112_290.n4 a_7112_290.t1 28.565
R3491 a_7112_290.t3 a_7112_290.n4 28.565
R3492 a_7112_290.n2 a_7112_290.t0 18.145
R3493 a_7112_290.n3 a_7112_290.n2 2.878
R3494 a_7112_290.n4 a_7112_290.n3 0.764
R3495 a_13367_n328.t0 a_13367_n328.t1 380.209
R3496 a_19826_n3212.n8 a_19826_n3212.n7 861.987
R3497 a_19826_n3212.n7 a_19826_n3212.n6 560.726
R3498 a_19826_n3212.t6 a_19826_n3212.t7 415.315
R3499 a_19826_n3212.t16 a_19826_n3212.t9 415.315
R3500 a_19826_n3212.n3 a_19826_n3212.t4 394.151
R3501 a_19826_n3212.n6 a_19826_n3212.t18 294.653
R3502 a_19826_n3212.n2 a_19826_n3212.t8 269.523
R3503 a_19826_n3212.t4 a_19826_n3212.n2 269.523
R3504 a_19826_n3212.n10 a_19826_n3212.t6 217.716
R3505 a_19826_n3212.n9 a_19826_n3212.t10 214.335
R3506 a_19826_n3212.t7 a_19826_n3212.n9 214.335
R3507 a_19826_n3212.n1 a_19826_n3212.t11 214.335
R3508 a_19826_n3212.t9 a_19826_n3212.n1 214.335
R3509 a_19826_n3212.n8 a_19826_n3212.t16 198.921
R3510 a_19826_n3212.n4 a_19826_n3212.t12 198.043
R3511 a_19826_n3212.n2 a_19826_n3212.t13 160.666
R3512 a_19826_n3212.n6 a_19826_n3212.t14 111.663
R3513 a_19826_n3212.n5 a_19826_n3212.n3 97.816
R3514 a_19826_n3212.n4 a_19826_n3212.t5 93.989
R3515 a_19826_n3212.n9 a_19826_n3212.t17 80.333
R3516 a_19826_n3212.n3 a_19826_n3212.t15 80.333
R3517 a_19826_n3212.n1 a_19826_n3212.t19 80.333
R3518 a_19826_n3212.n7 a_19826_n3212.n5 65.07
R3519 a_19826_n3212.t0 a_19826_n3212.n12 28.57
R3520 a_19826_n3212.n0 a_19826_n3212.t2 28.565
R3521 a_19826_n3212.n0 a_19826_n3212.t1 28.565
R3522 a_19826_n3212.n12 a_19826_n3212.t3 17.638
R3523 a_19826_n3212.n10 a_19826_n3212.n8 16.411
R3524 a_19826_n3212.n11 a_19826_n3212.n10 7.315
R3525 a_19826_n3212.n5 a_19826_n3212.n4 6.615
R3526 a_19826_n3212.n11 a_19826_n3212.n0 0.69
R3527 a_19826_n3212.n12 a_19826_n3212.n11 0.6
R3528 a_24630_404.t0 a_24630_404.n7 16.058
R3529 a_24630_404.n7 a_24630_404.n5 0.575
R3530 a_24630_404.n5 a_24630_404.n9 0.2
R3531 a_24630_404.n9 a_24630_404.t11 16.058
R3532 a_24630_404.n9 a_24630_404.n8 0.999
R3533 a_24630_404.n8 a_24630_404.t10 14.282
R3534 a_24630_404.n8 a_24630_404.t2 14.282
R3535 a_24630_404.n7 a_24630_404.n6 0.999
R3536 a_24630_404.n6 a_24630_404.t1 14.282
R3537 a_24630_404.n6 a_24630_404.t8 14.282
R3538 a_24630_404.n5 a_24630_404.n3 0.227
R3539 a_24630_404.n3 a_24630_404.n4 1.511
R3540 a_24630_404.n4 a_24630_404.t7 14.282
R3541 a_24630_404.n4 a_24630_404.t5 14.282
R3542 a_24630_404.n3 a_24630_404.n0 0.669
R3543 a_24630_404.n0 a_24630_404.n1 0.001
R3544 a_24630_404.n0 a_24630_404.n2 267.767
R3545 a_24630_404.n2 a_24630_404.t9 14.282
R3546 a_24630_404.n2 a_24630_404.t4 14.282
R3547 a_24630_404.n1 a_24630_404.t6 14.282
R3548 a_24630_404.n1 a_24630_404.t3 14.282
R3549 a_7414_n7824.n7 a_7414_n7824.n6 861.987
R3550 a_7414_n7824.n6 a_7414_n7824.n5 560.726
R3551 a_7414_n7824.t8 a_7414_n7824.t11 415.315
R3552 a_7414_n7824.t10 a_7414_n7824.t15 415.315
R3553 a_7414_n7824.n2 a_7414_n7824.t12 394.151
R3554 a_7414_n7824.n5 a_7414_n7824.t9 294.653
R3555 a_7414_n7824.n1 a_7414_n7824.t18 269.523
R3556 a_7414_n7824.t12 a_7414_n7824.n1 269.523
R3557 a_7414_n7824.n9 a_7414_n7824.t8 217.716
R3558 a_7414_n7824.n8 a_7414_n7824.t19 214.335
R3559 a_7414_n7824.t11 a_7414_n7824.n8 214.335
R3560 a_7414_n7824.n0 a_7414_n7824.t6 214.335
R3561 a_7414_n7824.t15 a_7414_n7824.n0 214.335
R3562 a_7414_n7824.n7 a_7414_n7824.t10 198.921
R3563 a_7414_n7824.n3 a_7414_n7824.t5 198.043
R3564 a_7414_n7824.n12 a_7414_n7824.n11 192.754
R3565 a_7414_n7824.n1 a_7414_n7824.t17 160.666
R3566 a_7414_n7824.n5 a_7414_n7824.t14 111.663
R3567 a_7414_n7824.n4 a_7414_n7824.n2 97.816
R3568 a_7414_n7824.n3 a_7414_n7824.t4 93.989
R3569 a_7414_n7824.n8 a_7414_n7824.t13 80.333
R3570 a_7414_n7824.n2 a_7414_n7824.t7 80.333
R3571 a_7414_n7824.n0 a_7414_n7824.t16 80.333
R3572 a_7414_n7824.n6 a_7414_n7824.n4 65.07
R3573 a_7414_n7824.t1 a_7414_n7824.n12 28.568
R3574 a_7414_n7824.n11 a_7414_n7824.t3 28.565
R3575 a_7414_n7824.n11 a_7414_n7824.t2 28.565
R3576 a_7414_n7824.n10 a_7414_n7824.t0 18.827
R3577 a_7414_n7824.n9 a_7414_n7824.n7 16.411
R3578 a_7414_n7824.n4 a_7414_n7824.n3 6.615
R3579 a_7414_n7824.n10 a_7414_n7824.n9 4.997
R3580 a_7414_n7824.n12 a_7414_n7824.n10 1.105
R3581 a_10918_n4773.n1 a_10918_n4773.t6 318.922
R3582 a_10918_n4773.n0 a_10918_n4773.t5 273.935
R3583 a_10918_n4773.n0 a_10918_n4773.t7 273.935
R3584 a_10918_n4773.n1 a_10918_n4773.t4 269.116
R3585 a_10918_n4773.n4 a_10918_n4773.n3 193.227
R3586 a_10918_n4773.t6 a_10918_n4773.n0 179.142
R3587 a_10918_n4773.n2 a_10918_n4773.n1 106.999
R3588 a_10918_n4773.n3 a_10918_n4773.t2 28.568
R3589 a_10918_n4773.n4 a_10918_n4773.t1 28.565
R3590 a_10918_n4773.t3 a_10918_n4773.n4 28.565
R3591 a_10918_n4773.n2 a_10918_n4773.t0 18.149
R3592 a_10918_n4773.n3 a_10918_n4773.n2 3.726
R3593 a_18543_3168.n0 a_18543_3168.t5 14.282
R3594 a_18543_3168.n0 a_18543_3168.t1 14.282
R3595 a_18543_3168.n1 a_18543_3168.t4 14.282
R3596 a_18543_3168.n1 a_18543_3168.t3 14.282
R3597 a_18543_3168.n3 a_18543_3168.t2 14.282
R3598 a_18543_3168.t0 a_18543_3168.n3 14.282
R3599 a_18543_3168.n3 a_18543_3168.n2 2.546
R3600 a_18543_3168.n2 a_18543_3168.n1 2.367
R3601 a_18543_3168.n2 a_18543_3168.n0 0.001
R3602 a_18425_3168.t6 a_18425_3168.n2 404.877
R3603 a_18425_3168.n1 a_18425_3168.t5 210.902
R3604 a_18425_3168.n3 a_18425_3168.t6 136.943
R3605 a_18425_3168.n2 a_18425_3168.n1 107.801
R3606 a_18425_3168.n1 a_18425_3168.t8 80.333
R3607 a_18425_3168.n2 a_18425_3168.t7 80.333
R3608 a_18425_3168.n0 a_18425_3168.t4 17.4
R3609 a_18425_3168.n0 a_18425_3168.t0 17.4
R3610 a_18425_3168.n4 a_18425_3168.t1 15.032
R3611 a_18425_3168.n5 a_18425_3168.t2 14.282
R3612 a_18425_3168.t3 a_18425_3168.n5 14.282
R3613 a_18425_3168.n5 a_18425_3168.n4 1.65
R3614 a_18425_3168.n3 a_18425_3168.n0 0.672
R3615 a_18425_3168.n4 a_18425_3168.n3 0.665
R3616 a_3029_1626.n4 a_3029_1626.t8 214.335
R3617 a_3029_1626.t7 a_3029_1626.n4 214.335
R3618 a_3029_1626.n5 a_3029_1626.t7 143.851
R3619 a_3029_1626.n5 a_3029_1626.t9 135.658
R3620 a_3029_1626.n4 a_3029_1626.t10 80.333
R3621 a_3029_1626.n0 a_3029_1626.t5 28.565
R3622 a_3029_1626.n0 a_3029_1626.t6 28.565
R3623 a_3029_1626.n2 a_3029_1626.t2 28.565
R3624 a_3029_1626.n2 a_3029_1626.t4 28.565
R3625 a_3029_1626.t0 a_3029_1626.n7 28.565
R3626 a_3029_1626.n7 a_3029_1626.t1 28.565
R3627 a_3029_1626.n1 a_3029_1626.t3 9.714
R3628 a_3029_1626.n1 a_3029_1626.n0 1.003
R3629 a_3029_1626.n6 a_3029_1626.n3 0.833
R3630 a_3029_1626.n3 a_3029_1626.n2 0.653
R3631 a_3029_1626.n7 a_3029_1626.n6 0.653
R3632 a_3029_1626.n3 a_3029_1626.n1 0.341
R3633 a_3029_1626.n6 a_3029_1626.n5 0.032
R3634 a_3619_1189.t4 a_3619_1189.t5 574.43
R3635 a_3619_1189.n0 a_3619_1189.t6 285.109
R3636 a_3619_1189.n2 a_3619_1189.n1 211.136
R3637 a_3619_1189.n4 a_3619_1189.n3 192.754
R3638 a_3619_1189.n0 a_3619_1189.t7 160.666
R3639 a_3619_1189.n1 a_3619_1189.t4 160.666
R3640 a_3619_1189.n1 a_3619_1189.n0 114.829
R3641 a_3619_1189.n3 a_3619_1189.t2 28.568
R3642 a_3619_1189.n4 a_3619_1189.t1 28.565
R3643 a_3619_1189.t3 a_3619_1189.n4 28.565
R3644 a_3619_1189.n2 a_3619_1189.t0 19.084
R3645 a_3619_1189.n3 a_3619_1189.n2 1.051
R3646 a_30337_n7043.n1 a_30337_n7043.t6 318.922
R3647 a_30337_n7043.n0 a_30337_n7043.t5 273.935
R3648 a_30337_n7043.n0 a_30337_n7043.t7 273.935
R3649 a_30337_n7043.n1 a_30337_n7043.t4 269.116
R3650 a_30337_n7043.n4 a_30337_n7043.n3 193.227
R3651 a_30337_n7043.t6 a_30337_n7043.n0 179.142
R3652 a_30337_n7043.n2 a_30337_n7043.n1 106.999
R3653 a_30337_n7043.n3 a_30337_n7043.t3 28.568
R3654 a_30337_n7043.n4 a_30337_n7043.t1 28.565
R3655 a_30337_n7043.t0 a_30337_n7043.n4 28.565
R3656 a_30337_n7043.n2 a_30337_n7043.t2 18.149
R3657 a_30337_n7043.n3 a_30337_n7043.n2 3.726
R3658 a_30882_n8468.t0 a_30882_n8468.t1 380.209
R3659 Y[3].n4 Y[3].n2 157.665
R3660 Y[3] Y[3].n6 145.563
R3661 Y[3].n4 Y[3].n3 122.999
R3662 Y[3].n6 Y[3].n0 90.436
R3663 Y[3].n5 Y[3].n1 90.416
R3664 Y[3].n6 Y[3].n5 74.302
R3665 Y[3].n5 Y[3].n4 50.575
R3666 Y[3].n0 Y[3].t3 14.282
R3667 Y[3].n0 Y[3].t2 14.282
R3668 Y[3].n1 Y[3].t1 14.282
R3669 Y[3].n1 Y[3].t7 14.282
R3670 Y[3].n3 Y[3].t4 14.282
R3671 Y[3].n3 Y[3].t5 14.282
R3672 Y[3].n2 Y[3].t0 8.7
R3673 Y[3].n2 Y[3].t6 8.7
R3674 a_11771_3236.t6 a_11771_3236.n2 404.877
R3675 a_11771_3236.n1 a_11771_3236.t8 210.902
R3676 a_11771_3236.n3 a_11771_3236.t6 136.943
R3677 a_11771_3236.n2 a_11771_3236.n1 107.801
R3678 a_11771_3236.n1 a_11771_3236.t5 80.333
R3679 a_11771_3236.n2 a_11771_3236.t7 80.333
R3680 a_11771_3236.n0 a_11771_3236.t0 17.4
R3681 a_11771_3236.n0 a_11771_3236.t4 17.4
R3682 a_11771_3236.n4 a_11771_3236.t3 15.032
R3683 a_11771_3236.n5 a_11771_3236.t2 14.282
R3684 a_11771_3236.t1 a_11771_3236.n5 14.282
R3685 a_11771_3236.n5 a_11771_3236.n4 1.65
R3686 a_11771_3236.n3 a_11771_3236.n0 0.672
R3687 a_11771_3236.n4 a_11771_3236.n3 0.665
R3688 a_12035_2653.t4 a_12035_2653.t6 800.071
R3689 a_12035_2653.n3 a_12035_2653.n2 672.951
R3690 a_12035_2653.n1 a_12035_2653.t5 285.109
R3691 a_12035_2653.n2 a_12035_2653.t4 193.602
R3692 a_12035_2653.n1 a_12035_2653.t7 160.666
R3693 a_12035_2653.n2 a_12035_2653.n1 91.507
R3694 a_12035_2653.n0 a_12035_2653.t2 28.57
R3695 a_12035_2653.n4 a_12035_2653.t1 28.565
R3696 a_12035_2653.t3 a_12035_2653.n4 28.565
R3697 a_12035_2653.n0 a_12035_2653.t0 17.638
R3698 a_12035_2653.n4 a_12035_2653.n3 0.69
R3699 a_12035_2653.n3 a_12035_2653.n0 0.6
R3700 a_25042_n2632.t6 a_25042_n2632.n2 404.877
R3701 a_25042_n2632.n1 a_25042_n2632.t5 210.902
R3702 a_25042_n2632.n3 a_25042_n2632.t6 136.943
R3703 a_25042_n2632.n2 a_25042_n2632.n1 107.801
R3704 a_25042_n2632.n1 a_25042_n2632.t8 80.333
R3705 a_25042_n2632.n2 a_25042_n2632.t7 80.333
R3706 a_25042_n2632.n0 a_25042_n2632.t4 17.4
R3707 a_25042_n2632.n0 a_25042_n2632.t2 17.4
R3708 a_25042_n2632.n4 a_25042_n2632.t3 15.032
R3709 a_25042_n2632.n5 a_25042_n2632.t1 14.282
R3710 a_25042_n2632.t0 a_25042_n2632.n5 14.282
R3711 a_25042_n2632.n5 a_25042_n2632.n4 1.65
R3712 a_25042_n2632.n3 a_25042_n2632.n0 0.672
R3713 a_25042_n2632.n4 a_25042_n2632.n3 0.665
R3714 a_25306_n3215.t7 a_25306_n3215.t6 800.071
R3715 a_25306_n3215.n3 a_25306_n3215.n2 672.951
R3716 a_25306_n3215.n1 a_25306_n3215.t5 285.109
R3717 a_25306_n3215.n2 a_25306_n3215.t7 193.602
R3718 a_25306_n3215.n1 a_25306_n3215.t4 160.666
R3719 a_25306_n3215.n2 a_25306_n3215.n1 91.507
R3720 a_25306_n3215.n0 a_25306_n3215.t2 28.57
R3721 a_25306_n3215.t3 a_25306_n3215.n4 28.565
R3722 a_25306_n3215.n4 a_25306_n3215.t1 28.565
R3723 a_25306_n3215.n0 a_25306_n3215.t0 17.638
R3724 a_25306_n3215.n4 a_25306_n3215.n3 0.69
R3725 a_25306_n3215.n3 a_25306_n3215.n0 0.6
R3726 a_11463_n5466.n0 a_11463_n5466.n12 122.999
R3727 a_11463_n5466.n0 a_11463_n5466.t1 14.282
R3728 a_11463_n5466.t0 a_11463_n5466.n0 14.282
R3729 a_11463_n5466.n12 a_11463_n5466.n10 50.575
R3730 a_11463_n5466.n10 a_11463_n5466.n8 74.302
R3731 a_11463_n5466.n12 a_11463_n5466.n11 157.665
R3732 a_11463_n5466.n11 a_11463_n5466.t2 8.7
R3733 a_11463_n5466.n11 a_11463_n5466.t5 8.7
R3734 a_11463_n5466.n10 a_11463_n5466.n9 90.416
R3735 a_11463_n5466.n9 a_11463_n5466.t3 14.282
R3736 a_11463_n5466.n9 a_11463_n5466.t6 14.282
R3737 a_11463_n5466.n8 a_11463_n5466.n7 90.436
R3738 a_11463_n5466.n7 a_11463_n5466.t7 14.282
R3739 a_11463_n5466.n7 a_11463_n5466.t4 14.282
R3740 a_11463_n5466.n8 a_11463_n5466.n1 342.688
R3741 a_11463_n5466.n1 a_11463_n5466.n6 126.566
R3742 a_11463_n5466.n6 a_11463_n5466.t9 294.653
R3743 a_11463_n5466.n6 a_11463_n5466.t10 111.663
R3744 a_11463_n5466.n1 a_11463_n5466.n5 552.333
R3745 a_11463_n5466.n5 a_11463_n5466.n4 6.615
R3746 a_11463_n5466.n4 a_11463_n5466.t15 93.989
R3747 a_11463_n5466.n5 a_11463_n5466.n3 97.816
R3748 a_11463_n5466.n3 a_11463_n5466.t8 80.333
R3749 a_11463_n5466.n3 a_11463_n5466.t11 394.151
R3750 a_11463_n5466.t11 a_11463_n5466.n2 269.523
R3751 a_11463_n5466.n2 a_11463_n5466.t12 160.666
R3752 a_11463_n5466.n2 a_11463_n5466.t13 269.523
R3753 a_11463_n5466.n4 a_11463_n5466.t14 198.043
R3754 a_12816_n4773.n1 a_12816_n4773.t5 318.922
R3755 a_12816_n4773.n0 a_12816_n4773.t7 273.935
R3756 a_12816_n4773.n0 a_12816_n4773.t6 273.935
R3757 a_12816_n4773.n1 a_12816_n4773.t4 269.116
R3758 a_12816_n4773.n4 a_12816_n4773.n3 193.227
R3759 a_12816_n4773.t5 a_12816_n4773.n0 179.142
R3760 a_12816_n4773.n2 a_12816_n4773.n1 106.999
R3761 a_12816_n4773.n3 a_12816_n4773.t2 28.568
R3762 a_12816_n4773.t3 a_12816_n4773.n4 28.565
R3763 a_12816_n4773.n4 a_12816_n4773.t1 28.565
R3764 a_12816_n4773.n2 a_12816_n4773.t0 18.149
R3765 a_12816_n4773.n3 a_12816_n4773.n2 3.726
R3766 A[0].t10 A[0].t1 437.233
R3767 A[0].t9 A[0].t2 415.315
R3768 A[0].t8 A[0].t12 415.315
R3769 A[0].t11 A[0].t4 415.315
R3770 A[0].n5 A[0].t8 221.468
R3771 A[0].n2 A[0].t10 219.798
R3772 A[0].n2 A[0].t9 217.276
R3773 A[0].n5 A[0].t11 217.129
R3774 A[0].n1 A[0].t7 214.686
R3775 A[0].t1 A[0].n1 214.686
R3776 A[0].n0 A[0].t0 214.335
R3777 A[0].t2 A[0].n0 214.335
R3778 A[0].n3 A[0].t14 214.335
R3779 A[0].t12 A[0].n3 214.335
R3780 A[0].n4 A[0].t6 214.335
R3781 A[0].t4 A[0].n4 214.335
R3782 A[0].n1 A[0].t15 80.333
R3783 A[0].n0 A[0].t3 80.333
R3784 A[0].n3 A[0].t13 80.333
R3785 A[0].n4 A[0].t5 80.333
R3786 A[0].n6 A[0].n5 54.612
R3787 A[0].n6 A[0].n2 49.781
R3788 A[0] A[0].n6 4.509
R3789 a_28645_5296.n0 a_28645_5296.t8 214.335
R3790 a_28645_5296.t10 a_28645_5296.n0 214.335
R3791 a_28645_5296.n1 a_28645_5296.t10 143.851
R3792 a_28645_5296.n1 a_28645_5296.t9 135.658
R3793 a_28645_5296.n0 a_28645_5296.t7 80.333
R3794 a_28645_5296.n2 a_28645_5296.t3 28.565
R3795 a_28645_5296.n2 a_28645_5296.t1 28.565
R3796 a_28645_5296.n4 a_28645_5296.t2 28.565
R3797 a_28645_5296.n4 a_28645_5296.t5 28.565
R3798 a_28645_5296.n7 a_28645_5296.t6 28.565
R3799 a_28645_5296.t0 a_28645_5296.n7 28.565
R3800 a_28645_5296.n6 a_28645_5296.t4 9.714
R3801 a_28645_5296.n7 a_28645_5296.n6 1.003
R3802 a_28645_5296.n5 a_28645_5296.n3 0.833
R3803 a_28645_5296.n3 a_28645_5296.n2 0.653
R3804 a_28645_5296.n5 a_28645_5296.n4 0.653
R3805 a_28645_5296.n6 a_28645_5296.n5 0.341
R3806 a_28645_5296.n3 a_28645_5296.n1 0.032
R3807 a_26302_n2628.n0 a_26302_n2628.t0 14.282
R3808 a_26302_n2628.n0 a_26302_n2628.t5 14.282
R3809 a_26302_n2628.n1 a_26302_n2628.t1 14.282
R3810 a_26302_n2628.n1 a_26302_n2628.t2 14.282
R3811 a_26302_n2628.n3 a_26302_n2628.t4 14.282
R3812 a_26302_n2628.t3 a_26302_n2628.n3 14.282
R3813 a_26302_n2628.n3 a_26302_n2628.n2 2.546
R3814 a_26302_n2628.n2 a_26302_n2628.n1 2.367
R3815 a_26302_n2628.n2 a_26302_n2628.n0 0.001
R3816 a_23425_n2941.t7 a_23425_n2941.t6 800.071
R3817 a_23425_n2941.n3 a_23425_n2941.n2 659.097
R3818 a_23425_n2941.n1 a_23425_n2941.t5 285.109
R3819 a_23425_n2941.n2 a_23425_n2941.t7 193.602
R3820 a_23425_n2941.n4 a_23425_n2941.n0 192.754
R3821 a_23425_n2941.n1 a_23425_n2941.t4 160.666
R3822 a_23425_n2941.n2 a_23425_n2941.n1 91.507
R3823 a_23425_n2941.t0 a_23425_n2941.n4 28.568
R3824 a_23425_n2941.n0 a_23425_n2941.t3 28.565
R3825 a_23425_n2941.n0 a_23425_n2941.t2 28.565
R3826 a_23425_n2941.n3 a_23425_n2941.t1 19.061
R3827 a_23425_n2941.n4 a_23425_n2941.n3 1.005
R3828 a_25160_n2632.n0 a_25160_n2632.t2 14.282
R3829 a_25160_n2632.n0 a_25160_n2632.t1 14.282
R3830 a_25160_n2632.n1 a_25160_n2632.t3 14.282
R3831 a_25160_n2632.n1 a_25160_n2632.t4 14.282
R3832 a_25160_n2632.t0 a_25160_n2632.n3 14.282
R3833 a_25160_n2632.n3 a_25160_n2632.t5 14.282
R3834 a_25160_n2632.n3 a_25160_n2632.n2 2.546
R3835 a_25160_n2632.n2 a_25160_n2632.n1 2.367
R3836 a_25160_n2632.n2 a_25160_n2632.n0 0.001
R3837 a_18689_2585.t7 a_18689_2585.t6 800.071
R3838 a_18689_2585.n3 a_18689_2585.n2 672.951
R3839 a_18689_2585.n1 a_18689_2585.t4 285.109
R3840 a_18689_2585.n2 a_18689_2585.t7 193.602
R3841 a_18689_2585.n1 a_18689_2585.t5 160.666
R3842 a_18689_2585.n2 a_18689_2585.n1 91.507
R3843 a_18689_2585.n0 a_18689_2585.t2 28.57
R3844 a_18689_2585.t3 a_18689_2585.n4 28.565
R3845 a_18689_2585.n4 a_18689_2585.t1 28.565
R3846 a_18689_2585.n0 a_18689_2585.t0 17.638
R3847 a_18689_2585.n4 a_18689_2585.n3 0.69
R3848 a_18689_2585.n3 a_18689_2585.n0 0.6
R3849 a_19685_3172.n0 a_19685_3172.t1 14.282
R3850 a_19685_3172.n0 a_19685_3172.t4 14.282
R3851 a_19685_3172.n1 a_19685_3172.t3 14.282
R3852 a_19685_3172.n1 a_19685_3172.t2 14.282
R3853 a_19685_3172.n3 a_19685_3172.t5 14.282
R3854 a_19685_3172.t0 a_19685_3172.n3 14.282
R3855 a_19685_3172.n3 a_19685_3172.n2 2.546
R3856 a_19685_3172.n2 a_19685_3172.n1 2.367
R3857 a_19685_3172.n2 a_19685_3172.n0 0.001
R3858 a_16232_1646.n0 a_16232_1646.t9 214.335
R3859 a_16232_1646.t7 a_16232_1646.n0 214.335
R3860 a_16232_1646.n1 a_16232_1646.t7 143.851
R3861 a_16232_1646.n1 a_16232_1646.t8 135.658
R3862 a_16232_1646.n0 a_16232_1646.t10 80.333
R3863 a_16232_1646.n2 a_16232_1646.t4 28.565
R3864 a_16232_1646.n2 a_16232_1646.t3 28.565
R3865 a_16232_1646.n4 a_16232_1646.t5 28.565
R3866 a_16232_1646.n4 a_16232_1646.t1 28.565
R3867 a_16232_1646.t0 a_16232_1646.n7 28.565
R3868 a_16232_1646.n7 a_16232_1646.t6 28.565
R3869 a_16232_1646.n6 a_16232_1646.t2 9.714
R3870 a_16232_1646.n7 a_16232_1646.n6 1.003
R3871 a_16232_1646.n5 a_16232_1646.n3 0.833
R3872 a_16232_1646.n3 a_16232_1646.n2 0.653
R3873 a_16232_1646.n5 a_16232_1646.n4 0.653
R3874 a_16232_1646.n6 a_16232_1646.n5 0.341
R3875 a_16232_1646.n3 a_16232_1646.n1 0.032
R3876 A[1].n6 A[1].n4 1494.07
R3877 A[1].t13 A[1].t3 437.233
R3878 A[1].t14 A[1].t0 437.233
R3879 A[1].t8 A[1].t11 437.233
R3880 A[1].t15 A[1].t7 415.315
R3881 A[1].n3 A[1].t14 224.833
R3882 A[1].n4 A[1].t15 219.944
R3883 A[1].n6 A[1].t8 217.054
R3884 A[1].n3 A[1].t13 216.198
R3885 A[1].n2 A[1].t1 214.686
R3886 A[1].t3 A[1].n2 214.686
R3887 A[1].n1 A[1].t5 214.686
R3888 A[1].t0 A[1].n1 214.686
R3889 A[1].n5 A[1].t4 214.686
R3890 A[1].t11 A[1].n5 214.686
R3891 A[1].n0 A[1].t12 214.335
R3892 A[1].t7 A[1].n0 214.335
R3893 A[1].n0 A[1].t10 80.333
R3894 A[1].n2 A[1].t2 80.333
R3895 A[1].n1 A[1].t9 80.333
R3896 A[1].n5 A[1].t6 80.333
R3897 A[1].n4 A[1].n3 34.046
R3898 A[1] A[1].n6 0.788
R3899 a_28640_n308.n4 a_28640_n308.t10 214.335
R3900 a_28640_n308.t9 a_28640_n308.n4 214.335
R3901 a_28640_n308.n5 a_28640_n308.t9 143.851
R3902 a_28640_n308.n5 a_28640_n308.t7 135.658
R3903 a_28640_n308.n4 a_28640_n308.t8 80.333
R3904 a_28640_n308.n0 a_28640_n308.t1 28.565
R3905 a_28640_n308.n0 a_28640_n308.t2 28.565
R3906 a_28640_n308.n2 a_28640_n308.t5 28.565
R3907 a_28640_n308.n2 a_28640_n308.t3 28.565
R3908 a_28640_n308.t4 a_28640_n308.n7 28.565
R3909 a_28640_n308.n7 a_28640_n308.t6 28.565
R3910 a_28640_n308.n1 a_28640_n308.t0 9.714
R3911 a_28640_n308.n1 a_28640_n308.n0 1.003
R3912 a_28640_n308.n6 a_28640_n308.n3 0.833
R3913 a_28640_n308.n3 a_28640_n308.n2 0.653
R3914 a_28640_n308.n7 a_28640_n308.n6 0.653
R3915 a_28640_n308.n3 a_28640_n308.n1 0.341
R3916 a_28640_n308.n6 a_28640_n308.n5 0.032
R3917 B[1].n5 B[1].t3 1361.95
R3918 B[1].n4 B[1].t13 1211.76
R3919 B[1].n5 B[1].t10 561.041
R3920 B[1].t3 B[1].t8 437.233
R3921 B[1].t10 B[1].t11 437.233
R3922 B[1].t13 B[1].t14 415.315
R3923 B[1].t2 B[1].t0 415.315
R3924 B[1].n4 B[1].t2 219.359
R3925 B[1].n0 B[1].t1 214.686
R3926 B[1].t8 B[1].n0 214.686
R3927 B[1].n1 B[1].t4 214.686
R3928 B[1].t11 B[1].n1 214.686
R3929 B[1].n2 B[1].t9 214.335
R3930 B[1].t14 B[1].n2 214.335
R3931 B[1].n3 B[1].t6 214.335
R3932 B[1].t0 B[1].n3 214.335
R3933 B[1].n0 B[1].t7 80.333
R3934 B[1].n1 B[1].t15 80.333
R3935 B[1].n2 B[1].t5 80.333
R3936 B[1].n3 B[1].t12 80.333
R3937 B[1].n5 B[1].n4 1.018
R3938 B[1] B[1].n5 0.23
R3939 a_125_3543.n0 a_125_3543.t10 214.335
R3940 a_125_3543.t7 a_125_3543.n0 214.335
R3941 a_125_3543.n1 a_125_3543.t7 143.851
R3942 a_125_3543.n1 a_125_3543.t8 135.658
R3943 a_125_3543.n0 a_125_3543.t9 80.333
R3944 a_125_3543.n2 a_125_3543.t5 28.565
R3945 a_125_3543.n2 a_125_3543.t4 28.565
R3946 a_125_3543.n4 a_125_3543.t6 28.565
R3947 a_125_3543.n4 a_125_3543.t1 28.565
R3948 a_125_3543.n7 a_125_3543.t2 28.565
R3949 a_125_3543.t3 a_125_3543.n7 28.565
R3950 a_125_3543.n6 a_125_3543.t0 9.714
R3951 a_125_3543.n7 a_125_3543.n6 1.003
R3952 a_125_3543.n5 a_125_3543.n3 0.833
R3953 a_125_3543.n3 a_125_3543.n2 0.653
R3954 a_125_3543.n5 a_125_3543.n4 0.653
R3955 a_125_3543.n6 a_125_3543.n5 0.341
R3956 a_125_3543.n3 a_125_3543.n1 0.032
R3957 a_18123_336.t0 a_18123_336.n0 14.282
R3958 a_18123_336.n0 a_18123_336.t3 14.282
R3959 a_18123_336.n0 a_18123_336.n12 90.416
R3960 a_18123_336.n12 a_18123_336.n11 50.575
R3961 a_18123_336.n12 a_18123_336.n8 74.302
R3962 a_18123_336.n11 a_18123_336.n10 157.665
R3963 a_18123_336.n10 a_18123_336.t5 8.7
R3964 a_18123_336.n10 a_18123_336.t7 8.7
R3965 a_18123_336.n11 a_18123_336.n9 122.999
R3966 a_18123_336.n9 a_18123_336.t6 14.282
R3967 a_18123_336.n9 a_18123_336.t1 14.282
R3968 a_18123_336.n8 a_18123_336.n7 90.436
R3969 a_18123_336.n7 a_18123_336.t2 14.282
R3970 a_18123_336.n7 a_18123_336.t4 14.282
R3971 a_18123_336.n8 a_18123_336.n1 342.688
R3972 a_18123_336.n1 a_18123_336.n6 126.566
R3973 a_18123_336.n6 a_18123_336.t12 294.653
R3974 a_18123_336.n6 a_18123_336.t15 111.663
R3975 a_18123_336.n1 a_18123_336.n5 552.333
R3976 a_18123_336.n5 a_18123_336.n4 6.615
R3977 a_18123_336.n4 a_18123_336.t9 93.989
R3978 a_18123_336.n5 a_18123_336.n3 97.816
R3979 a_18123_336.n3 a_18123_336.t14 80.333
R3980 a_18123_336.n3 a_18123_336.t8 394.151
R3981 a_18123_336.t8 a_18123_336.n2 269.523
R3982 a_18123_336.n2 a_18123_336.t13 160.666
R3983 a_18123_336.n2 a_18123_336.t10 269.523
R3984 a_18123_336.n4 a_18123_336.t11 198.043
R3985 a_19903_336.n0 a_19903_336.t1 14.282
R3986 a_19903_336.t0 a_19903_336.n0 14.282
R3987 a_19903_336.n0 a_19903_336.n9 0.999
R3988 a_19903_336.n9 a_19903_336.n6 0.575
R3989 a_19903_336.n6 a_19903_336.n8 0.2
R3990 a_19903_336.n8 a_19903_336.t5 16.058
R3991 a_19903_336.n8 a_19903_336.n7 0.999
R3992 a_19903_336.n7 a_19903_336.t4 14.282
R3993 a_19903_336.n7 a_19903_336.t6 14.282
R3994 a_19903_336.n9 a_19903_336.t3 16.058
R3995 a_19903_336.n6 a_19903_336.n4 0.227
R3996 a_19903_336.n4 a_19903_336.n5 1.511
R3997 a_19903_336.n5 a_19903_336.t9 14.282
R3998 a_19903_336.n5 a_19903_336.t7 14.282
R3999 a_19903_336.n4 a_19903_336.n1 0.669
R4000 a_19903_336.n1 a_19903_336.n2 0.001
R4001 a_19903_336.n1 a_19903_336.n3 267.767
R4002 a_19903_336.n3 a_19903_336.t10 14.282
R4003 a_19903_336.n3 a_19903_336.t11 14.282
R4004 a_19903_336.n2 a_19903_336.t8 14.282
R4005 a_19903_336.n2 a_19903_336.t2 14.282
R4006 a_16822_1209.t6 a_16822_1209.t7 574.43
R4007 a_16822_1209.n0 a_16822_1209.t4 285.109
R4008 a_16822_1209.n2 a_16822_1209.n1 211.136
R4009 a_16822_1209.n4 a_16822_1209.n3 192.754
R4010 a_16822_1209.n0 a_16822_1209.t5 160.666
R4011 a_16822_1209.n1 a_16822_1209.t6 160.666
R4012 a_16822_1209.n1 a_16822_1209.n0 114.829
R4013 a_16822_1209.n3 a_16822_1209.t2 28.568
R4014 a_16822_1209.n4 a_16822_1209.t1 28.565
R4015 a_16822_1209.t3 a_16822_1209.n4 28.565
R4016 a_16822_1209.n2 a_16822_1209.t0 19.084
R4017 a_16822_1209.n3 a_16822_1209.n2 1.051
R4018 a_7379_5006.n5 a_7379_5006.n4 535.449
R4019 a_7379_5006.t14 a_7379_5006.t15 437.233
R4020 a_7379_5006.t6 a_7379_5006.t12 437.233
R4021 a_7379_5006.t17 a_7379_5006.n2 313.873
R4022 a_7379_5006.n4 a_7379_5006.t13 294.986
R4023 a_7379_5006.n1 a_7379_5006.t18 272.288
R4024 a_7379_5006.n5 a_7379_5006.t11 245.184
R4025 a_7379_5006.n7 a_7379_5006.t6 218.628
R4026 a_7379_5006.n9 a_7379_5006.t14 217.024
R4027 a_7379_5006.n8 a_7379_5006.t10 214.686
R4028 a_7379_5006.t15 a_7379_5006.n8 214.686
R4029 a_7379_5006.n6 a_7379_5006.t4 214.686
R4030 a_7379_5006.t12 a_7379_5006.n6 214.686
R4031 a_7379_5006.n11 a_7379_5006.n0 192.754
R4032 a_7379_5006.n3 a_7379_5006.t17 190.152
R4033 a_7379_5006.n3 a_7379_5006.t19 190.152
R4034 a_7379_5006.n1 a_7379_5006.t8 160.666
R4035 a_7379_5006.n2 a_7379_5006.t9 160.666
R4036 a_7379_5006.n4 a_7379_5006.t7 110.859
R4037 a_7379_5006.n2 a_7379_5006.n1 96.129
R4038 a_7379_5006.n8 a_7379_5006.t5 80.333
R4039 a_7379_5006.t11 a_7379_5006.n3 80.333
R4040 a_7379_5006.n6 a_7379_5006.t16 80.333
R4041 a_7379_5006.t0 a_7379_5006.n11 28.568
R4042 a_7379_5006.n0 a_7379_5006.t1 28.565
R4043 a_7379_5006.n0 a_7379_5006.t2 28.565
R4044 a_7379_5006.n10 a_7379_5006.t3 18.819
R4045 a_7379_5006.n7 a_7379_5006.n5 14.9
R4046 a_7379_5006.n10 a_7379_5006.n9 2.96
R4047 a_7379_5006.n9 a_7379_5006.n7 2.599
R4048 a_7379_5006.n11 a_7379_5006.n10 1.098
R4049 a_9573_110.n4 a_9573_110.t8 214.335
R4050 a_9573_110.t7 a_9573_110.n4 214.335
R4051 a_9573_110.n5 a_9573_110.t7 143.851
R4052 a_9573_110.n5 a_9573_110.t9 135.658
R4053 a_9573_110.n4 a_9573_110.t10 80.333
R4054 a_9573_110.n0 a_9573_110.t2 28.565
R4055 a_9573_110.n0 a_9573_110.t4 28.565
R4056 a_9573_110.n2 a_9573_110.t1 28.565
R4057 a_9573_110.n2 a_9573_110.t3 28.565
R4058 a_9573_110.t0 a_9573_110.n7 28.565
R4059 a_9573_110.n7 a_9573_110.t6 28.565
R4060 a_9573_110.n1 a_9573_110.t5 9.714
R4061 a_9573_110.n1 a_9573_110.n0 1.003
R4062 a_9573_110.n6 a_9573_110.n3 0.833
R4063 a_9573_110.n3 a_9573_110.n2 0.653
R4064 a_9573_110.n7 a_9573_110.n6 0.653
R4065 a_9573_110.n3 a_9573_110.n1 0.341
R4066 a_9573_110.n6 a_9573_110.n5 0.032
R4067 a_20016_n5465.t0 a_20016_n5465.n0 14.282
R4068 a_20016_n5465.n0 a_20016_n5465.t4 14.282
R4069 a_20016_n5465.n0 a_20016_n5465.n15 90.416
R4070 a_20016_n5465.n15 a_20016_n5465.n14 50.575
R4071 a_20016_n5465.n15 a_20016_n5465.n11 74.302
R4072 a_20016_n5465.n14 a_20016_n5465.n13 157.665
R4073 a_20016_n5465.n13 a_20016_n5465.t5 8.7
R4074 a_20016_n5465.n13 a_20016_n5465.t7 8.7
R4075 a_20016_n5465.n14 a_20016_n5465.n12 122.999
R4076 a_20016_n5465.n12 a_20016_n5465.t6 14.282
R4077 a_20016_n5465.n12 a_20016_n5465.t1 14.282
R4078 a_20016_n5465.n11 a_20016_n5465.n10 90.436
R4079 a_20016_n5465.n10 a_20016_n5465.t2 14.282
R4080 a_20016_n5465.n10 a_20016_n5465.t3 14.282
R4081 a_20016_n5465.n11 a_20016_n5465.n9 220.49
R4082 a_20016_n5465.n9 a_20016_n5465.n2 2.599
R4083 a_20016_n5465.n2 a_20016_n5465.t11 218.628
R4084 a_20016_n5465.t11 a_20016_n5465.t12 437.233
R4085 a_20016_n5465.t12 a_20016_n5465.n8 214.686
R4086 a_20016_n5465.n8 a_20016_n5465.t15 80.333
R4087 a_20016_n5465.n8 a_20016_n5465.t9 214.686
R4088 a_20016_n5465.n2 a_20016_n5465.n3 14.9
R4089 a_20016_n5465.n3 a_20016_n5465.n7 535.449
R4090 a_20016_n5465.n7 a_20016_n5465.t22 294.986
R4091 a_20016_n5465.n7 a_20016_n5465.t14 110.859
R4092 a_20016_n5465.n3 a_20016_n5465.t17 245.184
R4093 a_20016_n5465.t17 a_20016_n5465.n6 80.333
R4094 a_20016_n5465.n6 a_20016_n5465.t18 190.152
R4095 a_20016_n5465.n6 a_20016_n5465.t16 190.152
R4096 a_20016_n5465.t16 a_20016_n5465.n5 313.873
R4097 a_20016_n5465.n5 a_20016_n5465.t23 160.666
R4098 a_20016_n5465.n5 a_20016_n5465.n4 96.129
R4099 a_20016_n5465.n4 a_20016_n5465.t21 160.666
R4100 a_20016_n5465.n4 a_20016_n5465.t13 272.288
R4101 a_20016_n5465.n9 a_20016_n5465.t8 217.024
R4102 a_20016_n5465.t8 a_20016_n5465.t10 437.233
R4103 a_20016_n5465.t10 a_20016_n5465.n1 214.686
R4104 a_20016_n5465.n1 a_20016_n5465.t20 80.333
R4105 a_20016_n5465.n1 a_20016_n5465.t19 214.686
R4106 a_22835_n2504.n2 a_22835_n2504.t7 214.335
R4107 a_22835_n2504.t9 a_22835_n2504.n2 214.335
R4108 a_22835_n2504.n3 a_22835_n2504.t9 143.851
R4109 a_22835_n2504.n3 a_22835_n2504.t8 135.658
R4110 a_22835_n2504.n2 a_22835_n2504.t10 80.333
R4111 a_22835_n2504.n4 a_22835_n2504.t2 28.565
R4112 a_22835_n2504.n4 a_22835_n2504.t1 28.565
R4113 a_22835_n2504.n0 a_22835_n2504.t4 28.565
R4114 a_22835_n2504.n0 a_22835_n2504.t5 28.565
R4115 a_22835_n2504.t0 a_22835_n2504.n7 28.565
R4116 a_22835_n2504.n7 a_22835_n2504.t6 28.565
R4117 a_22835_n2504.n1 a_22835_n2504.t3 9.714
R4118 a_22835_n2504.n1 a_22835_n2504.n0 1.003
R4119 a_22835_n2504.n6 a_22835_n2504.n5 0.833
R4120 a_22835_n2504.n5 a_22835_n2504.n4 0.653
R4121 a_22835_n2504.n7 a_22835_n2504.n6 0.653
R4122 a_22835_n2504.n6 a_22835_n2504.n1 0.341
R4123 a_22835_n2504.n5 a_22835_n2504.n3 0.032
R4124 a_23072_n3141.t0 a_23072_n3141.t1 17.4
R4125 a_2961_n4180.n6 a_2961_n4180.n5 501.28
R4126 a_2961_n4180.t10 a_2961_n4180.t14 437.233
R4127 a_2961_n4180.t19 a_2961_n4180.t6 415.315
R4128 a_2961_n4180.t16 a_2961_n4180.n3 313.873
R4129 a_2961_n4180.n5 a_2961_n4180.t7 294.986
R4130 a_2961_n4180.n2 a_2961_n4180.t12 272.288
R4131 a_2961_n4180.n6 a_2961_n4180.t17 236.01
R4132 a_2961_n4180.n9 a_2961_n4180.t10 216.627
R4133 a_2961_n4180.n7 a_2961_n4180.t19 216.111
R4134 a_2961_n4180.n8 a_2961_n4180.t11 214.686
R4135 a_2961_n4180.t14 a_2961_n4180.n8 214.686
R4136 a_2961_n4180.n1 a_2961_n4180.t9 214.335
R4137 a_2961_n4180.t6 a_2961_n4180.n1 214.335
R4138 a_2961_n4180.n4 a_2961_n4180.t16 190.152
R4139 a_2961_n4180.n4 a_2961_n4180.t18 190.152
R4140 a_2961_n4180.n2 a_2961_n4180.t4 160.666
R4141 a_2961_n4180.n3 a_2961_n4180.t5 160.666
R4142 a_2961_n4180.n7 a_2961_n4180.n6 148.428
R4143 a_2961_n4180.n5 a_2961_n4180.t15 110.859
R4144 a_2961_n4180.n3 a_2961_n4180.n2 96.129
R4145 a_2961_n4180.n8 a_2961_n4180.t13 80.333
R4146 a_2961_n4180.n1 a_2961_n4180.t8 80.333
R4147 a_2961_n4180.t17 a_2961_n4180.n4 80.333
R4148 a_2961_n4180.n0 a_2961_n4180.t2 28.57
R4149 a_2961_n4180.t0 a_2961_n4180.n11 28.565
R4150 a_2961_n4180.n11 a_2961_n4180.t3 28.565
R4151 a_2961_n4180.n0 a_2961_n4180.t1 17.638
R4152 a_2961_n4180.n10 a_2961_n4180.n9 7.04
R4153 a_2961_n4180.n9 a_2961_n4180.n7 2.923
R4154 a_2961_n4180.n11 a_2961_n4180.n10 0.69
R4155 a_2961_n4180.n10 a_2961_n4180.n0 0.6
R4156 a_6692_n5464.n0 a_6692_n5464.t5 14.282
R4157 a_6692_n5464.t0 a_6692_n5464.n0 14.282
R4158 a_6692_n5464.n0 a_6692_n5464.n9 0.999
R4159 a_6692_n5464.n6 a_6692_n5464.n8 0.575
R4160 a_6692_n5464.n9 a_6692_n5464.n6 0.2
R4161 a_6692_n5464.n9 a_6692_n5464.t8 16.058
R4162 a_6692_n5464.n8 a_6692_n5464.n7 0.999
R4163 a_6692_n5464.n7 a_6692_n5464.t11 14.282
R4164 a_6692_n5464.n7 a_6692_n5464.t9 14.282
R4165 a_6692_n5464.n8 a_6692_n5464.t10 16.058
R4166 a_6692_n5464.n6 a_6692_n5464.n4 0.227
R4167 a_6692_n5464.n4 a_6692_n5464.n5 1.511
R4168 a_6692_n5464.n5 a_6692_n5464.t6 14.282
R4169 a_6692_n5464.n5 a_6692_n5464.t7 14.282
R4170 a_6692_n5464.n4 a_6692_n5464.n1 0.669
R4171 a_6692_n5464.n1 a_6692_n5464.n2 0.001
R4172 a_6692_n5464.n1 a_6692_n5464.n3 267.767
R4173 a_6692_n5464.n3 a_6692_n5464.t4 14.282
R4174 a_6692_n5464.n3 a_6692_n5464.t3 14.282
R4175 a_6692_n5464.n2 a_6692_n5464.t1 14.282
R4176 a_6692_n5464.n2 a_6692_n5464.t2 14.282
R4177 a_19562_n2629.t8 a_19562_n2629.n2 404.877
R4178 a_19562_n2629.n1 a_19562_n2629.t7 210.902
R4179 a_19562_n2629.n3 a_19562_n2629.t8 136.943
R4180 a_19562_n2629.n2 a_19562_n2629.n1 107.801
R4181 a_19562_n2629.n1 a_19562_n2629.t6 80.333
R4182 a_19562_n2629.n2 a_19562_n2629.t5 80.333
R4183 a_19562_n2629.n0 a_19562_n2629.t0 17.4
R4184 a_19562_n2629.n0 a_19562_n2629.t4 17.4
R4185 a_19562_n2629.n4 a_19562_n2629.t3 15.032
R4186 a_19562_n2629.n5 a_19562_n2629.t2 14.282
R4187 a_19562_n2629.t1 a_19562_n2629.n5 14.282
R4188 a_19562_n2629.n5 a_19562_n2629.n4 1.65
R4189 a_19562_n2629.n3 a_19562_n2629.n0 0.672
R4190 a_19562_n2629.n4 a_19562_n2629.n3 0.665
R4191 a_32248_n2698.n0 a_32248_n2698.t10 214.335
R4192 a_32248_n2698.t8 a_32248_n2698.n0 214.335
R4193 a_32248_n2698.n1 a_32248_n2698.t8 143.851
R4194 a_32248_n2698.n1 a_32248_n2698.t7 135.658
R4195 a_32248_n2698.n0 a_32248_n2698.t9 80.333
R4196 a_32248_n2698.n2 a_32248_n2698.t2 28.565
R4197 a_32248_n2698.n2 a_32248_n2698.t4 28.565
R4198 a_32248_n2698.n4 a_32248_n2698.t3 28.565
R4199 a_32248_n2698.n4 a_32248_n2698.t6 28.565
R4200 a_32248_n2698.n7 a_32248_n2698.t5 28.565
R4201 a_32248_n2698.t1 a_32248_n2698.n7 28.565
R4202 a_32248_n2698.n6 a_32248_n2698.t0 9.714
R4203 a_32248_n2698.n7 a_32248_n2698.n6 1.003
R4204 a_32248_n2698.n5 a_32248_n2698.n3 0.833
R4205 a_32248_n2698.n3 a_32248_n2698.n2 0.653
R4206 a_32248_n2698.n5 a_32248_n2698.n4 0.653
R4207 a_32248_n2698.n6 a_32248_n2698.n5 0.341
R4208 a_32248_n2698.n3 a_32248_n2698.n1 0.032
R4209 a_22789_n4180.n4 a_22789_n4180.n3 501.28
R4210 a_22789_n4180.t8 a_22789_n4180.t10 437.233
R4211 a_22789_n4180.t11 a_22789_n4180.t14 415.315
R4212 a_22789_n4180.t6 a_22789_n4180.n1 313.873
R4213 a_22789_n4180.n3 a_22789_n4180.t18 294.986
R4214 a_22789_n4180.n0 a_22789_n4180.t9 272.288
R4215 a_22789_n4180.n4 a_22789_n4180.t7 236.01
R4216 a_22789_n4180.n8 a_22789_n4180.t8 216.627
R4217 a_22789_n4180.n6 a_22789_n4180.t11 216.069
R4218 a_22789_n4180.n7 a_22789_n4180.t5 214.686
R4219 a_22789_n4180.t10 a_22789_n4180.n7 214.686
R4220 a_22789_n4180.n5 a_22789_n4180.t17 214.335
R4221 a_22789_n4180.t14 a_22789_n4180.n5 214.335
R4222 a_22789_n4180.n11 a_22789_n4180.n10 192.754
R4223 a_22789_n4180.n2 a_22789_n4180.t6 190.152
R4224 a_22789_n4180.n2 a_22789_n4180.t19 190.152
R4225 a_22789_n4180.n0 a_22789_n4180.t13 160.666
R4226 a_22789_n4180.n1 a_22789_n4180.t15 160.666
R4227 a_22789_n4180.n6 a_22789_n4180.n4 148.384
R4228 a_22789_n4180.n3 a_22789_n4180.t4 110.859
R4229 a_22789_n4180.n1 a_22789_n4180.n0 96.129
R4230 a_22789_n4180.n7 a_22789_n4180.t12 80.333
R4231 a_22789_n4180.n5 a_22789_n4180.t16 80.333
R4232 a_22789_n4180.t7 a_22789_n4180.n2 80.333
R4233 a_22789_n4180.n9 a_22789_n4180.n8 47.31
R4234 a_22789_n4180.n10 a_22789_n4180.t1 28.568
R4235 a_22789_n4180.n11 a_22789_n4180.t2 28.565
R4236 a_22789_n4180.t3 a_22789_n4180.n11 28.565
R4237 a_22789_n4180.n9 a_22789_n4180.t0 18.466
R4238 a_22789_n4180.n8 a_22789_n4180.n6 2.697
R4239 a_22789_n4180.n10 a_22789_n4180.n9 1.161
R4240 a_13361_n5466.t0 a_13361_n5466.n0 14.282
R4241 a_13361_n5466.n0 a_13361_n5466.t1 14.282
R4242 a_13361_n5466.n0 a_13361_n5466.n13 90.436
R4243 a_13361_n5466.n9 a_13361_n5466.n12 50.575
R4244 a_13361_n5466.n13 a_13361_n5466.n9 74.302
R4245 a_13361_n5466.n12 a_13361_n5466.n11 157.665
R4246 a_13361_n5466.n11 a_13361_n5466.t2 8.7
R4247 a_13361_n5466.n11 a_13361_n5466.t6 8.7
R4248 a_13361_n5466.n12 a_13361_n5466.n10 122.999
R4249 a_13361_n5466.n10 a_13361_n5466.t4 14.282
R4250 a_13361_n5466.n10 a_13361_n5466.t3 14.282
R4251 a_13361_n5466.n9 a_13361_n5466.n8 90.416
R4252 a_13361_n5466.n8 a_13361_n5466.t5 14.282
R4253 a_13361_n5466.n8 a_13361_n5466.t7 14.282
R4254 a_13361_n5466.n13 a_13361_n5466.n1 1712.43
R4255 a_13361_n5466.n1 a_13361_n5466.t15 217.826
R4256 a_13361_n5466.n1 a_13361_n5466.n6 133.839
R4257 a_13361_n5466.t15 a_13361_n5466.t17 437.233
R4258 a_13361_n5466.t17 a_13361_n5466.n7 214.686
R4259 a_13361_n5466.n7 a_13361_n5466.t16 80.333
R4260 a_13361_n5466.n7 a_13361_n5466.t14 214.686
R4261 a_13361_n5466.n6 a_13361_n5466.n2 563.136
R4262 a_13361_n5466.n6 a_13361_n5466.t10 178.973
R4263 a_13361_n5466.t10 a_13361_n5466.n5 80.333
R4264 a_13361_n5466.n5 a_13361_n5466.t11 190.152
R4265 a_13361_n5466.n5 a_13361_n5466.t9 190.152
R4266 a_13361_n5466.t9 a_13361_n5466.n4 313.873
R4267 a_13361_n5466.n4 a_13361_n5466.t13 160.666
R4268 a_13361_n5466.n4 a_13361_n5466.n3 96.129
R4269 a_13361_n5466.n3 a_13361_n5466.t19 160.666
R4270 a_13361_n5466.n3 a_13361_n5466.t18 272.288
R4271 a_13361_n5466.n2 a_13361_n5466.t12 294.986
R4272 a_13361_n5466.n2 a_13361_n5466.t8 110.859
R4273 a_31176_n7762.n1 a_31176_n7762.t6 318.922
R4274 a_31176_n7762.n0 a_31176_n7762.t5 274.739
R4275 a_31176_n7762.n0 a_31176_n7762.t7 274.739
R4276 a_31176_n7762.n1 a_31176_n7762.t4 269.116
R4277 a_31176_n7762.t6 a_31176_n7762.n0 179.946
R4278 a_31176_n7762.n2 a_31176_n7762.n1 107.263
R4279 a_31176_n7762.n3 a_31176_n7762.t1 29.444
R4280 a_31176_n7762.n4 a_31176_n7762.t2 28.565
R4281 a_31176_n7762.t3 a_31176_n7762.n4 28.565
R4282 a_31176_n7762.n2 a_31176_n7762.t0 18.145
R4283 a_31176_n7762.n3 a_31176_n7762.n2 2.878
R4284 a_31176_n7762.n4 a_31176_n7762.n3 0.764
R4285 a_24740_n5464.n0 a_24740_n5464.t6 14.282
R4286 a_24740_n5464.t0 a_24740_n5464.n0 14.282
R4287 a_24740_n5464.n0 a_24740_n5464.n12 90.416
R4288 a_24740_n5464.n12 a_24740_n5464.n11 50.575
R4289 a_24740_n5464.n12 a_24740_n5464.n8 74.302
R4290 a_24740_n5464.n11 a_24740_n5464.n10 157.665
R4291 a_24740_n5464.n10 a_24740_n5464.t2 8.7
R4292 a_24740_n5464.n10 a_24740_n5464.t4 8.7
R4293 a_24740_n5464.n11 a_24740_n5464.n9 122.999
R4294 a_24740_n5464.n9 a_24740_n5464.t7 14.282
R4295 a_24740_n5464.n9 a_24740_n5464.t3 14.282
R4296 a_24740_n5464.n8 a_24740_n5464.n7 90.436
R4297 a_24740_n5464.n7 a_24740_n5464.t1 14.282
R4298 a_24740_n5464.n7 a_24740_n5464.t5 14.282
R4299 a_24740_n5464.n8 a_24740_n5464.n1 342.688
R4300 a_24740_n5464.n1 a_24740_n5464.n6 126.566
R4301 a_24740_n5464.n6 a_24740_n5464.t14 294.653
R4302 a_24740_n5464.n6 a_24740_n5464.t15 111.663
R4303 a_24740_n5464.n1 a_24740_n5464.n5 552.333
R4304 a_24740_n5464.n5 a_24740_n5464.n4 6.615
R4305 a_24740_n5464.n4 a_24740_n5464.t12 93.989
R4306 a_24740_n5464.n5 a_24740_n5464.n3 97.816
R4307 a_24740_n5464.n3 a_24740_n5464.t13 80.333
R4308 a_24740_n5464.n3 a_24740_n5464.t8 394.151
R4309 a_24740_n5464.t8 a_24740_n5464.n2 269.523
R4310 a_24740_n5464.n2 a_24740_n5464.t9 160.666
R4311 a_24740_n5464.n2 a_24740_n5464.t10 269.523
R4312 a_24740_n5464.n4 a_24740_n5464.t11 198.043
R4313 a_26520_n5464.n0 a_26520_n5464.t1 14.282
R4314 a_26520_n5464.t0 a_26520_n5464.n0 14.282
R4315 a_26520_n5464.n0 a_26520_n5464.n9 0.999
R4316 a_26520_n5464.n6 a_26520_n5464.n8 0.575
R4317 a_26520_n5464.n9 a_26520_n5464.n6 0.2
R4318 a_26520_n5464.n9 a_26520_n5464.t8 16.058
R4319 a_26520_n5464.n8 a_26520_n5464.n7 0.999
R4320 a_26520_n5464.n7 a_26520_n5464.t10 14.282
R4321 a_26520_n5464.n7 a_26520_n5464.t11 14.282
R4322 a_26520_n5464.n8 a_26520_n5464.t9 16.058
R4323 a_26520_n5464.n6 a_26520_n5464.n4 0.227
R4324 a_26520_n5464.n4 a_26520_n5464.n5 1.511
R4325 a_26520_n5464.n5 a_26520_n5464.t4 14.282
R4326 a_26520_n5464.n5 a_26520_n5464.t3 14.282
R4327 a_26520_n5464.n4 a_26520_n5464.n1 0.669
R4328 a_26520_n5464.n1 a_26520_n5464.n2 0.001
R4329 a_26520_n5464.n1 a_26520_n5464.n3 267.767
R4330 a_26520_n5464.n3 a_26520_n5464.t6 14.282
R4331 a_26520_n5464.n3 a_26520_n5464.t5 14.282
R4332 a_26520_n5464.n2 a_26520_n5464.t2 14.282
R4333 a_26520_n5464.n2 a_26520_n5464.t7 14.282
R4334 a_715_3106.n4 a_715_3106.n3 535.449
R4335 a_715_3106.t16 a_715_3106.t18 437.233
R4336 a_715_3106.t11 a_715_3106.t14 437.233
R4337 a_715_3106.t10 a_715_3106.n1 313.873
R4338 a_715_3106.n3 a_715_3106.t9 294.986
R4339 a_715_3106.n0 a_715_3106.t19 272.288
R4340 a_715_3106.n4 a_715_3106.t4 245.184
R4341 a_715_3106.n6 a_715_3106.t11 218.628
R4342 a_715_3106.n8 a_715_3106.t16 217.024
R4343 a_715_3106.n7 a_715_3106.t5 214.686
R4344 a_715_3106.t18 a_715_3106.n7 214.686
R4345 a_715_3106.n5 a_715_3106.t7 214.686
R4346 a_715_3106.t14 a_715_3106.n5 214.686
R4347 a_715_3106.n11 a_715_3106.n10 192.754
R4348 a_715_3106.n2 a_715_3106.t10 190.152
R4349 a_715_3106.n2 a_715_3106.t17 190.152
R4350 a_715_3106.n0 a_715_3106.t8 160.666
R4351 a_715_3106.n1 a_715_3106.t13 160.666
R4352 a_715_3106.n3 a_715_3106.t15 110.859
R4353 a_715_3106.n1 a_715_3106.n0 96.129
R4354 a_715_3106.n7 a_715_3106.t6 80.333
R4355 a_715_3106.t4 a_715_3106.n2 80.333
R4356 a_715_3106.n5 a_715_3106.t12 80.333
R4357 a_715_3106.n10 a_715_3106.t1 28.568
R4358 a_715_3106.n11 a_715_3106.t2 28.565
R4359 a_715_3106.t3 a_715_3106.n11 28.565
R4360 a_715_3106.n9 a_715_3106.t0 18.726
R4361 a_715_3106.n6 a_715_3106.n4 14.9
R4362 a_715_3106.n8 a_715_3106.n6 2.599
R4363 a_715_3106.n9 a_715_3106.n8 2.514
R4364 a_715_3106.n10 a_715_3106.n9 1.123
R4365 a_29301_n2665.n5 a_29301_n2665.n4 465.933
R4366 a_29301_n2665.t15 a_29301_n2665.t7 415.315
R4367 a_29301_n2665.n1 a_29301_n2665.t8 394.151
R4368 a_29301_n2665.n4 a_29301_n2665.t9 294.653
R4369 a_29301_n2665.n0 a_29301_n2665.t4 269.523
R4370 a_29301_n2665.t8 a_29301_n2665.n0 269.523
R4371 a_29301_n2665.n7 a_29301_n2665.t15 220.285
R4372 a_29301_n2665.n6 a_29301_n2665.t13 214.335
R4373 a_29301_n2665.t7 a_29301_n2665.n6 214.335
R4374 a_29301_n2665.n2 a_29301_n2665.t11 198.043
R4375 a_29301_n2665.n10 a_29301_n2665.n9 192.754
R4376 a_29301_n2665.n5 a_29301_n2665.n3 163.88
R4377 a_29301_n2665.n0 a_29301_n2665.t6 160.666
R4378 a_29301_n2665.n4 a_29301_n2665.t14 111.663
R4379 a_29301_n2665.n3 a_29301_n2665.n1 97.816
R4380 a_29301_n2665.n2 a_29301_n2665.t12 93.989
R4381 a_29301_n2665.n6 a_29301_n2665.t5 80.333
R4382 a_29301_n2665.n1 a_29301_n2665.t10 80.333
R4383 a_29301_n2665.n7 a_29301_n2665.n5 61.538
R4384 a_29301_n2665.n9 a_29301_n2665.t2 28.568
R4385 a_29301_n2665.n10 a_29301_n2665.t1 28.565
R4386 a_29301_n2665.t0 a_29301_n2665.n10 28.565
R4387 a_29301_n2665.n8 a_29301_n2665.t3 18.824
R4388 a_29301_n2665.n3 a_29301_n2665.n2 6.615
R4389 a_29301_n2665.n8 a_29301_n2665.n7 5.5
R4390 a_29301_n2665.n9 a_29301_n2665.n8 1.105
R4391 a_30764_107.n5 a_30764_107.n7 0.575
R4392 a_30764_107.n9 a_30764_107.n5 0.2
R4393 a_30764_107.t3 a_30764_107.n9 16.058
R4394 a_30764_107.n9 a_30764_107.n8 0.999
R4395 a_30764_107.n8 a_30764_107.t4 14.282
R4396 a_30764_107.n8 a_30764_107.t7 14.282
R4397 a_30764_107.n7 a_30764_107.n6 0.999
R4398 a_30764_107.n6 a_30764_107.t6 14.282
R4399 a_30764_107.n6 a_30764_107.t11 14.282
R4400 a_30764_107.n7 a_30764_107.t5 16.058
R4401 a_30764_107.n5 a_30764_107.n3 0.227
R4402 a_30764_107.n3 a_30764_107.n4 1.511
R4403 a_30764_107.n4 a_30764_107.t0 14.282
R4404 a_30764_107.n4 a_30764_107.t1 14.282
R4405 a_30764_107.n3 a_30764_107.n0 0.669
R4406 a_30764_107.n0 a_30764_107.n1 0.001
R4407 a_30764_107.n0 a_30764_107.n2 267.767
R4408 a_30764_107.n2 a_30764_107.t9 14.282
R4409 a_30764_107.n2 a_30764_107.t8 14.282
R4410 a_30764_107.n1 a_30764_107.t2 14.282
R4411 a_30764_107.n1 a_30764_107.t10 14.282
R4412 a_29305_n8580.n6 a_29305_n8580.n5 465.933
R4413 a_29305_n8580.t9 a_29305_n8580.t12 415.315
R4414 a_29305_n8580.n2 a_29305_n8580.t10 394.151
R4415 a_29305_n8580.n5 a_29305_n8580.t5 294.653
R4416 a_29305_n8580.n1 a_29305_n8580.t15 269.523
R4417 a_29305_n8580.t10 a_29305_n8580.n1 269.523
R4418 a_29305_n8580.n8 a_29305_n8580.t9 220.285
R4419 a_29305_n8580.n7 a_29305_n8580.t4 214.335
R4420 a_29305_n8580.t12 a_29305_n8580.n7 214.335
R4421 a_29305_n8580.n3 a_29305_n8580.t14 198.043
R4422 a_29305_n8580.n10 a_29305_n8580.n0 192.754
R4423 a_29305_n8580.n6 a_29305_n8580.n4 163.88
R4424 a_29305_n8580.n1 a_29305_n8580.t11 160.666
R4425 a_29305_n8580.n5 a_29305_n8580.t8 111.663
R4426 a_29305_n8580.n4 a_29305_n8580.n2 97.816
R4427 a_29305_n8580.n3 a_29305_n8580.t6 93.989
R4428 a_29305_n8580.n7 a_29305_n8580.t13 80.333
R4429 a_29305_n8580.n2 a_29305_n8580.t7 80.333
R4430 a_29305_n8580.n8 a_29305_n8580.n6 61.538
R4431 a_29305_n8580.t0 a_29305_n8580.n10 28.568
R4432 a_29305_n8580.n0 a_29305_n8580.t3 28.565
R4433 a_29305_n8580.n0 a_29305_n8580.t2 28.565
R4434 a_29305_n8580.n9 a_29305_n8580.t1 18.824
R4435 a_29305_n8580.n4 a_29305_n8580.n3 6.615
R4436 a_29305_n8580.n9 a_29305_n8580.n8 2.736
R4437 a_29305_n8580.n10 a_29305_n8580.n9 1.105
R4438 a_32248_n7046.n4 a_32248_n7046.t9 214.335
R4439 a_32248_n7046.t7 a_32248_n7046.n4 214.335
R4440 a_32248_n7046.n5 a_32248_n7046.t7 143.851
R4441 a_32248_n7046.n5 a_32248_n7046.t10 135.658
R4442 a_32248_n7046.n4 a_32248_n7046.t8 80.333
R4443 a_32248_n7046.n0 a_32248_n7046.t5 28.565
R4444 a_32248_n7046.n0 a_32248_n7046.t6 28.565
R4445 a_32248_n7046.n2 a_32248_n7046.t1 28.565
R4446 a_32248_n7046.n2 a_32248_n7046.t4 28.565
R4447 a_32248_n7046.t2 a_32248_n7046.n7 28.565
R4448 a_32248_n7046.n7 a_32248_n7046.t0 28.565
R4449 a_32248_n7046.n1 a_32248_n7046.t3 9.714
R4450 a_32248_n7046.n1 a_32248_n7046.n0 1.003
R4451 a_32248_n7046.n6 a_32248_n7046.n3 0.833
R4452 a_32248_n7046.n3 a_32248_n7046.n2 0.653
R4453 a_32248_n7046.n7 a_32248_n7046.n6 0.653
R4454 a_32248_n7046.n3 a_32248_n7046.n1 0.341
R4455 a_32248_n7046.n6 a_32248_n7046.n5 0.032
R4456 a_22844_n5758.n0 a_22844_n5758.t8 214.335
R4457 a_22844_n5758.t10 a_22844_n5758.n0 214.335
R4458 a_22844_n5758.n1 a_22844_n5758.t10 143.851
R4459 a_22844_n5758.n1 a_22844_n5758.t9 135.658
R4460 a_22844_n5758.n0 a_22844_n5758.t7 80.333
R4461 a_22844_n5758.n2 a_22844_n5758.t4 28.565
R4462 a_22844_n5758.n2 a_22844_n5758.t5 28.565
R4463 a_22844_n5758.n4 a_22844_n5758.t6 28.565
R4464 a_22844_n5758.n4 a_22844_n5758.t2 28.565
R4465 a_22844_n5758.n7 a_22844_n5758.t1 28.565
R4466 a_22844_n5758.t3 a_22844_n5758.n7 28.565
R4467 a_22844_n5758.n6 a_22844_n5758.t0 9.714
R4468 a_22844_n5758.n7 a_22844_n5758.n6 1.003
R4469 a_22844_n5758.n5 a_22844_n5758.n3 0.833
R4470 a_22844_n5758.n3 a_22844_n5758.n2 0.653
R4471 a_22844_n5758.n5 a_22844_n5758.n4 0.653
R4472 a_22844_n5758.n6 a_22844_n5758.n5 0.341
R4473 a_22844_n5758.n3 a_22844_n5758.n1 0.032
R4474 a_23434_n6195.t5 a_23434_n6195.t4 574.43
R4475 a_23434_n6195.n0 a_23434_n6195.t7 285.109
R4476 a_23434_n6195.n2 a_23434_n6195.n1 197.217
R4477 a_23434_n6195.n4 a_23434_n6195.n3 192.754
R4478 a_23434_n6195.n0 a_23434_n6195.t6 160.666
R4479 a_23434_n6195.n1 a_23434_n6195.t5 160.666
R4480 a_23434_n6195.n1 a_23434_n6195.n0 114.829
R4481 a_23434_n6195.n3 a_23434_n6195.t2 28.568
R4482 a_23434_n6195.t3 a_23434_n6195.n4 28.565
R4483 a_23434_n6195.n4 a_23434_n6195.t1 28.565
R4484 a_23434_n6195.n2 a_23434_n6195.t0 18.838
R4485 a_23434_n6195.n3 a_23434_n6195.n2 1.129
R4486 a_16172_1620.n17 a_16172_1620.n16 538.835
R4487 a_16172_1620.n9 a_16172_1620.n8 501.28
R4488 a_16172_1620.t9 a_16172_1620.t8 437.233
R4489 a_16172_1620.t11 a_16172_1620.t17 415.315
R4490 a_16172_1620.t14 a_16172_1620.n6 313.873
R4491 a_16172_1620.n8 a_16172_1620.t19 294.986
R4492 a_16172_1620.n5 a_16172_1620.t4 272.288
R4493 a_16172_1620.n9 a_16172_1620.t6 236.01
R4494 a_16172_1620.n12 a_16172_1620.t9 216.627
R4495 a_16172_1620.n10 a_16172_1620.t11 216.111
R4496 a_16172_1620.n11 a_16172_1620.t13 214.686
R4497 a_16172_1620.t8 a_16172_1620.n11 214.686
R4498 a_16172_1620.n4 a_16172_1620.t15 214.335
R4499 a_16172_1620.t17 a_16172_1620.n4 214.335
R4500 a_16172_1620.n19 a_16172_1620.n18 192.754
R4501 a_16172_1620.n7 a_16172_1620.t14 190.152
R4502 a_16172_1620.n7 a_16172_1620.t7 190.152
R4503 a_16172_1620.n5 a_16172_1620.t16 160.666
R4504 a_16172_1620.n6 a_16172_1620.t18 160.666
R4505 a_16172_1620.n10 a_16172_1620.n9 148.428
R4506 a_16172_1620.n8 a_16172_1620.t10 110.859
R4507 a_16172_1620.n6 a_16172_1620.n5 96.129
R4508 a_16172_1620.n11 a_16172_1620.t5 80.333
R4509 a_16172_1620.n4 a_16172_1620.t12 80.333
R4510 a_16172_1620.t6 a_16172_1620.n7 80.333
R4511 a_16172_1620.n18 a_16172_1620.t1 28.568
R4512 a_16172_1620.n19 a_16172_1620.t2 28.565
R4513 a_16172_1620.t3 a_16172_1620.n19 28.565
R4514 a_16172_1620.n17 a_16172_1620.t0 18.514
R4515 a_16172_1620.n16 a_16172_1620.n15 4.161
R4516 a_16172_1620.n12 a_16172_1620.n10 2.923
R4517 a_16172_1620.n18 a_16172_1620.n17 1.177
R4518 a_16172_1620.n13 a_16172_1620.n12 0.707
R4519 a_16172_1620.n15 a_16172_1620.n14 0.078
R4520 a_16172_1620.n1 a_16172_1620.n0 0.045
R4521 a_16172_1620.n3 a_16172_1620.n2 0.006
R4522 a_16172_1620.n15 a_16172_1620.n1 0.003
R4523 a_16172_1620.n13 a_16172_1620.n3 0.002
R4524 a_16172_1620.n15 a_16172_1620.n13 0.001
R4525 a_13177_2657.n5 a_13177_2657.n4 535.449
R4526 a_13177_2657.t11 a_13177_2657.t18 437.233
R4527 a_13177_2657.t19 a_13177_2657.t4 437.233
R4528 a_13177_2657.t7 a_13177_2657.n2 313.873
R4529 a_13177_2657.n4 a_13177_2657.t14 294.986
R4530 a_13177_2657.n1 a_13177_2657.t8 272.288
R4531 a_13177_2657.n5 a_13177_2657.t6 245.184
R4532 a_13177_2657.n7 a_13177_2657.t19 218.628
R4533 a_13177_2657.n9 a_13177_2657.t11 217.024
R4534 a_13177_2657.n8 a_13177_2657.t12 214.686
R4535 a_13177_2657.t18 a_13177_2657.n8 214.686
R4536 a_13177_2657.n6 a_13177_2657.t15 214.686
R4537 a_13177_2657.t4 a_13177_2657.n6 214.686
R4538 a_13177_2657.n3 a_13177_2657.t7 190.152
R4539 a_13177_2657.n3 a_13177_2657.t10 190.152
R4540 a_13177_2657.n1 a_13177_2657.t9 160.666
R4541 a_13177_2657.n2 a_13177_2657.t16 160.666
R4542 a_13177_2657.n4 a_13177_2657.t5 110.859
R4543 a_13177_2657.n2 a_13177_2657.n1 96.129
R4544 a_13177_2657.n8 a_13177_2657.t13 80.333
R4545 a_13177_2657.t6 a_13177_2657.n3 80.333
R4546 a_13177_2657.n6 a_13177_2657.t17 80.333
R4547 a_13177_2657.n0 a_13177_2657.t2 28.57
R4548 a_13177_2657.n11 a_13177_2657.t3 28.565
R4549 a_13177_2657.t0 a_13177_2657.n11 28.565
R4550 a_13177_2657.n0 a_13177_2657.t1 17.638
R4551 a_13177_2657.n7 a_13177_2657.n5 14.9
R4552 a_13177_2657.n10 a_13177_2657.n9 8.819
R4553 a_13177_2657.n9 a_13177_2657.n7 2.599
R4554 a_13177_2657.n11 a_13177_2657.n10 0.69
R4555 a_13177_2657.n10 a_13177_2657.n0 0.6
R4556 a_16222_n5759.n4 a_16222_n5759.t10 214.335
R4557 a_16222_n5759.t8 a_16222_n5759.n4 214.335
R4558 a_16222_n5759.n5 a_16222_n5759.t8 143.851
R4559 a_16222_n5759.n5 a_16222_n5759.t7 135.658
R4560 a_16222_n5759.n4 a_16222_n5759.t9 80.333
R4561 a_16222_n5759.n0 a_16222_n5759.t1 28.565
R4562 a_16222_n5759.n0 a_16222_n5759.t2 28.565
R4563 a_16222_n5759.n2 a_16222_n5759.t6 28.565
R4564 a_16222_n5759.n2 a_16222_n5759.t3 28.565
R4565 a_16222_n5759.n7 a_16222_n5759.t5 28.565
R4566 a_16222_n5759.t4 a_16222_n5759.n7 28.565
R4567 a_16222_n5759.n1 a_16222_n5759.t0 9.714
R4568 a_16222_n5759.n1 a_16222_n5759.n0 1.003
R4569 a_16222_n5759.n6 a_16222_n5759.n3 0.833
R4570 a_16222_n5759.n3 a_16222_n5759.n2 0.653
R4571 a_16222_n5759.n7 a_16222_n5759.n6 0.653
R4572 a_16222_n5759.n3 a_16222_n5759.n1 0.341
R4573 a_16222_n5759.n6 a_16222_n5759.n5 0.032
R4574 a_3015_3276.n2 a_3015_3276.t7 214.335
R4575 a_3015_3276.t10 a_3015_3276.n2 214.335
R4576 a_3015_3276.n3 a_3015_3276.t10 143.851
R4577 a_3015_3276.n3 a_3015_3276.t9 135.658
R4578 a_3015_3276.n2 a_3015_3276.t8 80.333
R4579 a_3015_3276.n4 a_3015_3276.t5 28.565
R4580 a_3015_3276.n4 a_3015_3276.t6 28.565
R4581 a_3015_3276.n0 a_3015_3276.t2 28.565
R4582 a_3015_3276.n0 a_3015_3276.t3 28.565
R4583 a_3015_3276.t0 a_3015_3276.n7 28.565
R4584 a_3015_3276.n7 a_3015_3276.t1 28.565
R4585 a_3015_3276.n1 a_3015_3276.t4 9.714
R4586 a_3015_3276.n1 a_3015_3276.n0 1.003
R4587 a_3015_3276.n6 a_3015_3276.n5 0.833
R4588 a_3015_3276.n5 a_3015_3276.n4 0.653
R4589 a_3015_3276.n7 a_3015_3276.n6 0.653
R4590 a_3015_3276.n6 a_3015_3276.n1 0.341
R4591 a_3015_3276.n5 a_3015_3276.n3 0.032
R4592 a_3605_2839.t5 a_3605_2839.t4 800.071
R4593 a_3605_2839.n3 a_3605_2839.n2 659.097
R4594 a_3605_2839.n1 a_3605_2839.t6 285.109
R4595 a_3605_2839.n2 a_3605_2839.t5 193.602
R4596 a_3605_2839.n4 a_3605_2839.n0 192.754
R4597 a_3605_2839.n1 a_3605_2839.t7 160.666
R4598 a_3605_2839.n2 a_3605_2839.n1 91.507
R4599 a_3605_2839.t3 a_3605_2839.n4 28.568
R4600 a_3605_2839.n0 a_3605_2839.t2 28.565
R4601 a_3605_2839.n0 a_3605_2839.t1 28.565
R4602 a_3605_2839.n3 a_3605_2839.t0 19.061
R4603 a_3605_2839.n4 a_3605_2839.n3 1.005
R4604 a_4920_316.t1 a_4920_316.n0 14.282
R4605 a_4920_316.n0 a_4920_316.t6 14.282
R4606 a_4920_316.n0 a_4920_316.n12 90.416
R4607 a_4920_316.n12 a_4920_316.n11 50.575
R4608 a_4920_316.n12 a_4920_316.n8 74.302
R4609 a_4920_316.n11 a_4920_316.n10 157.665
R4610 a_4920_316.n10 a_4920_316.t3 8.7
R4611 a_4920_316.n10 a_4920_316.t0 8.7
R4612 a_4920_316.n11 a_4920_316.n9 122.999
R4613 a_4920_316.n9 a_4920_316.t4 14.282
R4614 a_4920_316.n9 a_4920_316.t2 14.282
R4615 a_4920_316.n8 a_4920_316.n7 90.436
R4616 a_4920_316.n7 a_4920_316.t5 14.282
R4617 a_4920_316.n7 a_4920_316.t7 14.282
R4618 a_4920_316.n8 a_4920_316.n1 342.688
R4619 a_4920_316.n1 a_4920_316.n6 126.566
R4620 a_4920_316.n6 a_4920_316.t10 294.653
R4621 a_4920_316.n6 a_4920_316.t11 111.663
R4622 a_4920_316.n1 a_4920_316.n5 552.333
R4623 a_4920_316.n5 a_4920_316.n4 6.615
R4624 a_4920_316.n4 a_4920_316.t9 93.989
R4625 a_4920_316.n5 a_4920_316.n3 97.816
R4626 a_4920_316.n3 a_4920_316.t15 80.333
R4627 a_4920_316.n3 a_4920_316.t8 394.151
R4628 a_4920_316.t8 a_4920_316.n2 269.523
R4629 a_4920_316.n2 a_4920_316.t13 160.666
R4630 a_4920_316.n2 a_4920_316.t14 269.523
R4631 a_4920_316.n4 a_4920_316.t12 198.043
R4632 a_6700_316.n0 a_6700_316.t4 14.282
R4633 a_6700_316.t3 a_6700_316.n0 14.282
R4634 a_6700_316.n0 a_6700_316.n9 0.999
R4635 a_6700_316.n9 a_6700_316.n6 0.575
R4636 a_6700_316.n6 a_6700_316.n8 0.2
R4637 a_6700_316.n8 a_6700_316.t7 16.058
R4638 a_6700_316.n8 a_6700_316.n7 0.999
R4639 a_6700_316.n7 a_6700_316.t5 14.282
R4640 a_6700_316.n7 a_6700_316.t6 14.282
R4641 a_6700_316.n9 a_6700_316.t8 16.058
R4642 a_6700_316.n6 a_6700_316.n4 0.227
R4643 a_6700_316.n4 a_6700_316.n5 1.511
R4644 a_6700_316.n5 a_6700_316.t2 14.282
R4645 a_6700_316.n5 a_6700_316.t1 14.282
R4646 a_6700_316.n4 a_6700_316.n1 0.669
R4647 a_6700_316.n1 a_6700_316.n2 0.001
R4648 a_6700_316.n1 a_6700_316.n3 267.767
R4649 a_6700_316.n3 a_6700_316.t9 14.282
R4650 a_6700_316.n3 a_6700_316.t10 14.282
R4651 a_6700_316.n2 a_6700_316.t0 14.282
R4652 a_6700_316.n2 a_6700_316.t11 14.282
R4653 a_3024_22.n0 a_3024_22.t9 214.335
R4654 a_3024_22.t10 a_3024_22.n0 214.335
R4655 a_3024_22.n1 a_3024_22.t10 143.851
R4656 a_3024_22.n1 a_3024_22.t8 135.658
R4657 a_3024_22.n0 a_3024_22.t7 80.333
R4658 a_3024_22.n2 a_3024_22.t4 28.565
R4659 a_3024_22.n2 a_3024_22.t5 28.565
R4660 a_3024_22.n4 a_3024_22.t6 28.565
R4661 a_3024_22.n4 a_3024_22.t0 28.565
R4662 a_3024_22.n7 a_3024_22.t1 28.565
R4663 a_3024_22.t2 a_3024_22.n7 28.565
R4664 a_3024_22.n6 a_3024_22.t3 9.714
R4665 a_3024_22.n7 a_3024_22.n6 1.003
R4666 a_3024_22.n5 a_3024_22.n3 0.833
R4667 a_3024_22.n3 a_3024_22.n2 0.653
R4668 a_3024_22.n5 a_3024_22.n4 0.653
R4669 a_3024_22.n6 a_3024_22.n5 0.341
R4670 a_3024_22.n3 a_3024_22.n1 0.032
R4671 a_3614_n415.t7 a_3614_n415.t4 574.43
R4672 a_3614_n415.n0 a_3614_n415.t6 285.109
R4673 a_3614_n415.n2 a_3614_n415.n1 197.217
R4674 a_3614_n415.n4 a_3614_n415.n3 192.754
R4675 a_3614_n415.n0 a_3614_n415.t5 160.666
R4676 a_3614_n415.n1 a_3614_n415.t7 160.666
R4677 a_3614_n415.n1 a_3614_n415.n0 114.829
R4678 a_3614_n415.n3 a_3614_n415.t2 28.568
R4679 a_3614_n415.t3 a_3614_n415.n4 28.565
R4680 a_3614_n415.n4 a_3614_n415.t1 28.565
R4681 a_3614_n415.n2 a_3614_n415.t0 18.838
R4682 a_3614_n415.n3 a_3614_n415.n2 1.129
R4683 a_707_521.n7 a_707_521.n6 861.987
R4684 a_707_521.n6 a_707_521.n5 560.726
R4685 a_707_521.t8 a_707_521.t19 415.315
R4686 a_707_521.t15 a_707_521.t9 415.315
R4687 a_707_521.n2 a_707_521.t12 394.151
R4688 a_707_521.n5 a_707_521.t17 294.653
R4689 a_707_521.n1 a_707_521.t6 269.523
R4690 a_707_521.t12 a_707_521.n1 269.523
R4691 a_707_521.n9 a_707_521.t8 217.716
R4692 a_707_521.n8 a_707_521.t10 214.335
R4693 a_707_521.t19 a_707_521.n8 214.335
R4694 a_707_521.n0 a_707_521.t11 214.335
R4695 a_707_521.t9 a_707_521.n0 214.335
R4696 a_707_521.n7 a_707_521.t15 198.921
R4697 a_707_521.n3 a_707_521.t5 198.043
R4698 a_707_521.n12 a_707_521.n11 192.754
R4699 a_707_521.n1 a_707_521.t13 160.666
R4700 a_707_521.n5 a_707_521.t4 111.663
R4701 a_707_521.n4 a_707_521.n2 97.816
R4702 a_707_521.n3 a_707_521.t16 93.989
R4703 a_707_521.n8 a_707_521.t14 80.333
R4704 a_707_521.n2 a_707_521.t7 80.333
R4705 a_707_521.n0 a_707_521.t18 80.333
R4706 a_707_521.n6 a_707_521.n4 65.07
R4707 a_707_521.n11 a_707_521.t3 28.568
R4708 a_707_521.t0 a_707_521.n12 28.565
R4709 a_707_521.n12 a_707_521.t2 28.565
R4710 a_707_521.n10 a_707_521.t1 18.825
R4711 a_707_521.n9 a_707_521.n7 16.411
R4712 a_707_521.n4 a_707_521.n3 6.615
R4713 a_707_521.n10 a_707_521.n9 2.757
R4714 a_707_521.n11 a_707_521.n10 1.105
R4715 a_4375_1009.n2 a_4375_1009.t5 318.922
R4716 a_4375_1009.n1 a_4375_1009.t7 273.935
R4717 a_4375_1009.n1 a_4375_1009.t4 273.935
R4718 a_4375_1009.n2 a_4375_1009.t6 269.116
R4719 a_4375_1009.n4 a_4375_1009.n0 193.227
R4720 a_4375_1009.t5 a_4375_1009.n1 179.142
R4721 a_4375_1009.n3 a_4375_1009.n2 106.999
R4722 a_4375_1009.t3 a_4375_1009.n4 28.568
R4723 a_4375_1009.n0 a_4375_1009.t2 28.565
R4724 a_4375_1009.n0 a_4375_1009.t1 28.565
R4725 a_4375_1009.n3 a_4375_1009.t0 18.149
R4726 a_4375_1009.n4 a_4375_1009.n3 3.726
R4727 a_10163_n327.t6 a_10163_n327.t7 574.43
R4728 a_10163_n327.n0 a_10163_n327.t5 285.109
R4729 a_10163_n327.n2 a_10163_n327.n1 197.217
R4730 a_10163_n327.n4 a_10163_n327.n3 192.754
R4731 a_10163_n327.n0 a_10163_n327.t4 160.666
R4732 a_10163_n327.n1 a_10163_n327.t6 160.666
R4733 a_10163_n327.n1 a_10163_n327.n0 114.829
R4734 a_10163_n327.n3 a_10163_n327.t2 28.568
R4735 a_10163_n327.n4 a_10163_n327.t1 28.565
R4736 a_10163_n327.t3 a_10163_n327.n4 28.565
R4737 a_10163_n327.n2 a_10163_n327.t0 18.838
R4738 a_10163_n327.n3 a_10163_n327.n2 1.129
R4739 B[2].t8 B[2].t3 437.233
R4740 B[2].t10 B[2].t6 437.233
R4741 B[2].t11 B[2].t12 415.315
R4742 B[2].t2 B[2].t14 415.315
R4743 B[2].n2 B[2].t2 240.379
R4744 B[2].n5 B[2].t10 227.856
R4745 B[2].n2 B[2].t11 218.339
R4746 B[2].n5 B[2].t8 218.225
R4747 B[2].n3 B[2].t0 214.686
R4748 B[2].t3 B[2].n3 214.686
R4749 B[2].n4 B[2].t4 214.686
R4750 B[2].t6 B[2].n4 214.686
R4751 B[2].n1 B[2].t13 214.335
R4752 B[2].t12 B[2].n1 214.335
R4753 B[2].n0 B[2].t9 214.335
R4754 B[2].t14 B[2].n0 214.335
R4755 B[2].n1 B[2].t7 80.333
R4756 B[2].n0 B[2].t15 80.333
R4757 B[2].n3 B[2].t1 80.333
R4758 B[2].n4 B[2].t5 80.333
R4759 B[2].n6 B[2].n2 28.897
R4760 B[2].n6 B[2].n5 7.414
R4761 B[2] B[2].n6 3.805
R4762 a_6824_n8261.n2 a_6824_n8261.t8 214.335
R4763 a_6824_n8261.t9 a_6824_n8261.n2 214.335
R4764 a_6824_n8261.n3 a_6824_n8261.t9 143.85
R4765 a_6824_n8261.n3 a_6824_n8261.t7 135.66
R4766 a_6824_n8261.n2 a_6824_n8261.t10 80.333
R4767 a_6824_n8261.n4 a_6824_n8261.t0 28.565
R4768 a_6824_n8261.n4 a_6824_n8261.t1 28.565
R4769 a_6824_n8261.n0 a_6824_n8261.t4 28.565
R4770 a_6824_n8261.n0 a_6824_n8261.t5 28.565
R4771 a_6824_n8261.t2 a_6824_n8261.n7 28.565
R4772 a_6824_n8261.n7 a_6824_n8261.t3 28.565
R4773 a_6824_n8261.n1 a_6824_n8261.t6 9.714
R4774 a_6824_n8261.n1 a_6824_n8261.n0 1.003
R4775 a_6824_n8261.n6 a_6824_n8261.n5 0.836
R4776 a_6824_n8261.n7 a_6824_n8261.n6 0.653
R4777 a_6824_n8261.n5 a_6824_n8261.n4 0.65
R4778 a_6824_n8261.n6 a_6824_n8261.n1 0.341
R4779 a_6824_n8261.n5 a_6824_n8261.n3 0.032
R4780 a_32248_797.n0 a_32248_797.t7 214.335
R4781 a_32248_797.t9 a_32248_797.n0 214.335
R4782 a_32248_797.n1 a_32248_797.t9 143.851
R4783 a_32248_797.n1 a_32248_797.t10 135.658
R4784 a_32248_797.n0 a_32248_797.t8 80.333
R4785 a_32248_797.n2 a_32248_797.t0 28.565
R4786 a_32248_797.n2 a_32248_797.t2 28.565
R4787 a_32248_797.n4 a_32248_797.t1 28.565
R4788 a_32248_797.n4 a_32248_797.t6 28.565
R4789 a_32248_797.n7 a_32248_797.t5 28.565
R4790 a_32248_797.t4 a_32248_797.n7 28.565
R4791 a_32248_797.n6 a_32248_797.t3 9.714
R4792 a_32248_797.n7 a_32248_797.n6 1.003
R4793 a_32248_797.n5 a_32248_797.n3 0.833
R4794 a_32248_797.n3 a_32248_797.n2 0.653
R4795 a_32248_797.n5 a_32248_797.n4 0.653
R4796 a_32248_797.n6 a_32248_797.n5 0.341
R4797 a_32248_797.n3 a_32248_797.n1 0.032
R4798 a_31176_81.n1 a_31176_81.t4 318.922
R4799 a_31176_81.n0 a_31176_81.t6 274.739
R4800 a_31176_81.n0 a_31176_81.t5 274.739
R4801 a_31176_81.n1 a_31176_81.t7 269.116
R4802 a_31176_81.t4 a_31176_81.n0 179.946
R4803 a_31176_81.n2 a_31176_81.n1 107.263
R4804 a_31176_81.n3 a_31176_81.t1 29.444
R4805 a_31176_81.t0 a_31176_81.n4 28.565
R4806 a_31176_81.n4 a_31176_81.t3 28.565
R4807 a_31176_81.n2 a_31176_81.t2 18.145
R4808 a_31176_81.n3 a_31176_81.n2 2.878
R4809 a_31176_81.n4 a_31176_81.n3 0.764
R4810 Y[1].n4 Y[1].n2 157.665
R4811 Y[1] Y[1].n6 145.596
R4812 Y[1].n4 Y[1].n3 122.999
R4813 Y[1].n6 Y[1].n0 90.436
R4814 Y[1].n5 Y[1].n1 90.416
R4815 Y[1].n6 Y[1].n5 74.302
R4816 Y[1].n5 Y[1].n4 50.575
R4817 Y[1].n0 Y[1].t4 14.282
R4818 Y[1].n0 Y[1].t5 14.282
R4819 Y[1].n1 Y[1].t3 14.282
R4820 Y[1].n1 Y[1].t7 14.282
R4821 Y[1].n3 Y[1].t2 14.282
R4822 Y[1].n3 Y[1].t1 14.282
R4823 Y[1].n2 Y[1].t0 8.7
R4824 Y[1].n2 Y[1].t6 8.7
R4825 a_20617_n7831.n7 a_20617_n7831.n6 861.987
R4826 a_20617_n7831.n6 a_20617_n7831.n5 560.726
R4827 a_20617_n7831.t5 a_20617_n7831.t13 415.315
R4828 a_20617_n7831.t7 a_20617_n7831.t9 415.315
R4829 a_20617_n7831.n2 a_20617_n7831.t8 394.151
R4830 a_20617_n7831.n5 a_20617_n7831.t4 294.653
R4831 a_20617_n7831.n1 a_20617_n7831.t12 269.523
R4832 a_20617_n7831.t8 a_20617_n7831.n1 269.523
R4833 a_20617_n7831.n9 a_20617_n7831.t5 217.716
R4834 a_20617_n7831.n8 a_20617_n7831.t15 214.335
R4835 a_20617_n7831.t13 a_20617_n7831.n8 214.335
R4836 a_20617_n7831.n0 a_20617_n7831.t18 214.335
R4837 a_20617_n7831.t9 a_20617_n7831.n0 214.335
R4838 a_20617_n7831.n7 a_20617_n7831.t7 198.921
R4839 a_20617_n7831.n3 a_20617_n7831.t16 198.043
R4840 a_20617_n7831.n12 a_20617_n7831.n11 192.754
R4841 a_20617_n7831.n1 a_20617_n7831.t10 160.666
R4842 a_20617_n7831.n5 a_20617_n7831.t6 111.663
R4843 a_20617_n7831.n4 a_20617_n7831.n2 97.816
R4844 a_20617_n7831.n3 a_20617_n7831.t17 93.989
R4845 a_20617_n7831.n8 a_20617_n7831.t14 80.333
R4846 a_20617_n7831.n2 a_20617_n7831.t19 80.333
R4847 a_20617_n7831.n0 a_20617_n7831.t11 80.333
R4848 a_20617_n7831.n6 a_20617_n7831.n4 65.07
R4849 a_20617_n7831.n11 a_20617_n7831.t3 28.568
R4850 a_20617_n7831.n12 a_20617_n7831.t1 28.565
R4851 a_20617_n7831.t0 a_20617_n7831.n12 28.565
R4852 a_20617_n7831.n10 a_20617_n7831.t2 18.827
R4853 a_20617_n7831.n9 a_20617_n7831.n7 16.411
R4854 a_20617_n7831.n4 a_20617_n7831.n3 6.615
R4855 a_20617_n7831.n10 a_20617_n7831.n9 4.58
R4856 a_20617_n7831.n11 a_20617_n7831.n10 1.105
R4857 a_24976_n6196.t0 a_24976_n6196.t1 17.4
R4858 a_16218_3296.n2 a_16218_3296.t7 214.335
R4859 a_16218_3296.t10 a_16218_3296.n2 214.335
R4860 a_16218_3296.n3 a_16218_3296.t10 143.851
R4861 a_16218_3296.n3 a_16218_3296.t9 135.658
R4862 a_16218_3296.n2 a_16218_3296.t8 80.333
R4863 a_16218_3296.n4 a_16218_3296.t6 28.565
R4864 a_16218_3296.n4 a_16218_3296.t5 28.565
R4865 a_16218_3296.n0 a_16218_3296.t3 28.565
R4866 a_16218_3296.n0 a_16218_3296.t1 28.565
R4867 a_16218_3296.n7 a_16218_3296.t4 28.565
R4868 a_16218_3296.t0 a_16218_3296.n7 28.565
R4869 a_16218_3296.n1 a_16218_3296.t2 9.714
R4870 a_16218_3296.n1 a_16218_3296.n0 1.003
R4871 a_16218_3296.n6 a_16218_3296.n5 0.833
R4872 a_16218_3296.n5 a_16218_3296.n4 0.653
R4873 a_16218_3296.n7 a_16218_3296.n6 0.653
R4874 a_16218_3296.n6 a_16218_3296.n1 0.341
R4875 a_16218_3296.n5 a_16218_3296.n3 0.032
R4876 a_11469_404.n0 a_11469_404.n12 122.999
R4877 a_11469_404.n0 a_11469_404.t3 14.282
R4878 a_11469_404.t2 a_11469_404.n0 14.282
R4879 a_11469_404.n12 a_11469_404.n10 50.575
R4880 a_11469_404.n10 a_11469_404.n8 74.302
R4881 a_11469_404.n12 a_11469_404.n11 157.665
R4882 a_11469_404.n11 a_11469_404.t0 8.7
R4883 a_11469_404.n11 a_11469_404.t1 8.7
R4884 a_11469_404.n10 a_11469_404.n9 90.416
R4885 a_11469_404.n9 a_11469_404.t4 14.282
R4886 a_11469_404.n9 a_11469_404.t7 14.282
R4887 a_11469_404.n8 a_11469_404.n7 90.436
R4888 a_11469_404.n7 a_11469_404.t6 14.282
R4889 a_11469_404.n7 a_11469_404.t5 14.282
R4890 a_11469_404.n8 a_11469_404.n1 342.688
R4891 a_11469_404.n1 a_11469_404.n6 126.566
R4892 a_11469_404.n6 a_11469_404.t13 294.653
R4893 a_11469_404.n6 a_11469_404.t9 111.663
R4894 a_11469_404.n1 a_11469_404.n5 552.333
R4895 a_11469_404.n5 a_11469_404.n4 6.615
R4896 a_11469_404.n4 a_11469_404.t12 93.989
R4897 a_11469_404.n5 a_11469_404.n3 97.816
R4898 a_11469_404.n3 a_11469_404.t10 80.333
R4899 a_11469_404.n3 a_11469_404.t14 394.151
R4900 a_11469_404.t14 a_11469_404.n2 269.523
R4901 a_11469_404.n2 a_11469_404.t11 160.666
R4902 a_11469_404.n2 a_11469_404.t15 269.523
R4903 a_11469_404.n4 a_11469_404.t8 198.043
R4904 a_26932_n5490.n1 a_26932_n5490.t6 318.922
R4905 a_26932_n5490.n0 a_26932_n5490.t7 274.739
R4906 a_26932_n5490.n0 a_26932_n5490.t4 274.739
R4907 a_26932_n5490.n1 a_26932_n5490.t5 269.116
R4908 a_26932_n5490.t6 a_26932_n5490.n0 179.946
R4909 a_26932_n5490.n2 a_26932_n5490.n1 105.178
R4910 a_26932_n5490.n3 a_26932_n5490.t1 29.444
R4911 a_26932_n5490.n4 a_26932_n5490.t2 28.565
R4912 a_26932_n5490.t3 a_26932_n5490.n4 28.565
R4913 a_26932_n5490.n2 a_26932_n5490.t0 18.145
R4914 a_26932_n5490.n3 a_26932_n5490.n2 2.878
R4915 a_26932_n5490.n4 a_26932_n5490.n3 0.764
R4916 Y[5] Y[5].n6 214.948
R4917 Y[5].n4 Y[5].n2 157.665
R4918 Y[5].n4 Y[5].n3 122.999
R4919 Y[5].n6 Y[5].n0 90.436
R4920 Y[5].n5 Y[5].n1 90.416
R4921 Y[5].n6 Y[5].n5 74.302
R4922 Y[5].n5 Y[5].n4 50.575
R4923 Y[5].n0 Y[5].t2 14.282
R4924 Y[5].n0 Y[5].t1 14.282
R4925 Y[5].n1 Y[5].t0 14.282
R4926 Y[5].n1 Y[5].t7 14.282
R4927 Y[5].n3 Y[5].t6 14.282
R4928 Y[5].n3 Y[5].t5 14.282
R4929 Y[5].n2 Y[5].t3 8.7
R4930 Y[5].n2 Y[5].t4 8.7
R4931 a_9512_n4182.n6 a_9512_n4182.n5 501.28
R4932 a_9512_n4182.t10 a_9512_n4182.t14 437.233
R4933 a_9512_n4182.t12 a_9512_n4182.t13 415.315
R4934 a_9512_n4182.t11 a_9512_n4182.n3 313.873
R4935 a_9512_n4182.n5 a_9512_n4182.t5 294.986
R4936 a_9512_n4182.n2 a_9512_n4182.t15 272.288
R4937 a_9512_n4182.n6 a_9512_n4182.t17 236.01
R4938 a_9512_n4182.n9 a_9512_n4182.t10 216.627
R4939 a_9512_n4182.n7 a_9512_n4182.t12 216.111
R4940 a_9512_n4182.n8 a_9512_n4182.t7 214.686
R4941 a_9512_n4182.t14 a_9512_n4182.n8 214.686
R4942 a_9512_n4182.n1 a_9512_n4182.t4 214.335
R4943 a_9512_n4182.t13 a_9512_n4182.n1 214.335
R4944 a_9512_n4182.n11 a_9512_n4182.n0 192.754
R4945 a_9512_n4182.n4 a_9512_n4182.t11 190.152
R4946 a_9512_n4182.n4 a_9512_n4182.t18 190.152
R4947 a_9512_n4182.n2 a_9512_n4182.t16 160.666
R4948 a_9512_n4182.n3 a_9512_n4182.t6 160.666
R4949 a_9512_n4182.n7 a_9512_n4182.n6 148.428
R4950 a_9512_n4182.n5 a_9512_n4182.t9 110.859
R4951 a_9512_n4182.n10 a_9512_n4182.n9 102.569
R4952 a_9512_n4182.n3 a_9512_n4182.n2 96.129
R4953 a_9512_n4182.n8 a_9512_n4182.t8 80.333
R4954 a_9512_n4182.n1 a_9512_n4182.t19 80.333
R4955 a_9512_n4182.t17 a_9512_n4182.n4 80.333
R4956 a_9512_n4182.t3 a_9512_n4182.n11 28.568
R4957 a_9512_n4182.n0 a_9512_n4182.t2 28.565
R4958 a_9512_n4182.n0 a_9512_n4182.t1 28.565
R4959 a_9512_n4182.n10 a_9512_n4182.t0 18.523
R4960 a_9512_n4182.n9 a_9512_n4182.n7 2.923
R4961 a_9512_n4182.n11 a_9512_n4182.n10 1.167
R4962 a_16469_1009.t0 a_16469_1009.t1 17.4
R4963 a_22857_1714.n0 a_22857_1714.t8 214.335
R4964 a_22857_1714.t7 a_22857_1714.n0 214.335
R4965 a_22857_1714.n1 a_22857_1714.t7 143.851
R4966 a_22857_1714.n1 a_22857_1714.t9 135.658
R4967 a_22857_1714.n0 a_22857_1714.t10 80.333
R4968 a_22857_1714.n2 a_22857_1714.t1 28.565
R4969 a_22857_1714.n2 a_22857_1714.t0 28.565
R4970 a_22857_1714.n4 a_22857_1714.t2 28.565
R4971 a_22857_1714.n4 a_22857_1714.t4 28.565
R4972 a_22857_1714.t3 a_22857_1714.n7 28.565
R4973 a_22857_1714.n7 a_22857_1714.t5 28.565
R4974 a_22857_1714.n6 a_22857_1714.t6 9.714
R4975 a_22857_1714.n7 a_22857_1714.n6 1.003
R4976 a_22857_1714.n5 a_22857_1714.n3 0.833
R4977 a_22857_1714.n3 a_22857_1714.n2 0.653
R4978 a_22857_1714.n5 a_22857_1714.n4 0.653
R4979 a_22857_1714.n6 a_22857_1714.n5 0.341
R4980 a_22857_1714.n3 a_22857_1714.n1 0.032
R4981 a_23447_1277.t4 a_23447_1277.t5 574.43
R4982 a_23447_1277.n0 a_23447_1277.t6 285.109
R4983 a_23447_1277.n2 a_23447_1277.n1 211.136
R4984 a_23447_1277.n4 a_23447_1277.n3 192.754
R4985 a_23447_1277.n0 a_23447_1277.t7 160.666
R4986 a_23447_1277.n1 a_23447_1277.t4 160.666
R4987 a_23447_1277.n1 a_23447_1277.n0 114.829
R4988 a_23447_1277.n3 a_23447_1277.t2 28.568
R4989 a_23447_1277.n4 a_23447_1277.t1 28.565
R4990 a_23447_1277.t3 a_23447_1277.n4 28.565
R4991 a_23447_1277.n2 a_23447_1277.t0 19.084
R4992 a_23447_1277.n3 a_23447_1277.n2 1.051
R4993 a_24203_1097.n1 a_24203_1097.t7 318.922
R4994 a_24203_1097.n0 a_24203_1097.t5 273.935
R4995 a_24203_1097.n0 a_24203_1097.t4 273.935
R4996 a_24203_1097.n1 a_24203_1097.t6 269.116
R4997 a_24203_1097.n4 a_24203_1097.n3 193.227
R4998 a_24203_1097.t7 a_24203_1097.n0 179.142
R4999 a_24203_1097.n2 a_24203_1097.n1 106.999
R5000 a_24203_1097.n3 a_24203_1097.t2 28.568
R5001 a_24203_1097.n4 a_24203_1097.t1 28.565
R5002 a_24203_1097.t3 a_24203_1097.n4 28.565
R5003 a_24203_1097.n2 a_24203_1097.t0 18.149
R5004 a_24203_1097.n3 a_24203_1097.n2 3.726
R5005 a_10162_n4593.t7 a_10162_n4593.t4 574.43
R5006 a_10162_n4593.n0 a_10162_n4593.t5 285.109
R5007 a_10162_n4593.n2 a_10162_n4593.n1 211.136
R5008 a_10162_n4593.n4 a_10162_n4593.n3 192.754
R5009 a_10162_n4593.n0 a_10162_n4593.t6 160.666
R5010 a_10162_n4593.n1 a_10162_n4593.t7 160.666
R5011 a_10162_n4593.n1 a_10162_n4593.n0 114.829
R5012 a_10162_n4593.n3 a_10162_n4593.t3 28.568
R5013 a_10162_n4593.n4 a_10162_n4593.t2 28.565
R5014 a_10162_n4593.t0 a_10162_n4593.n4 28.565
R5015 a_10162_n4593.n2 a_10162_n4593.t1 19.084
R5016 a_10162_n4593.n3 a_10162_n4593.n2 1.051
R5017 a_12907_n2630.t6 a_12907_n2630.n3 404.877
R5018 a_12907_n2630.n2 a_12907_n2630.t8 210.902
R5019 a_12907_n2630.n4 a_12907_n2630.t6 136.943
R5020 a_12907_n2630.n3 a_12907_n2630.n2 107.801
R5021 a_12907_n2630.n2 a_12907_n2630.t7 80.333
R5022 a_12907_n2630.n3 a_12907_n2630.t5 80.333
R5023 a_12907_n2630.n1 a_12907_n2630.t4 17.4
R5024 a_12907_n2630.n1 a_12907_n2630.t0 17.4
R5025 a_12907_n2630.t1 a_12907_n2630.n5 15.032
R5026 a_12907_n2630.n0 a_12907_n2630.t3 14.282
R5027 a_12907_n2630.n0 a_12907_n2630.t2 14.282
R5028 a_12907_n2630.n5 a_12907_n2630.n0 1.65
R5029 a_12907_n2630.n4 a_12907_n2630.n1 0.672
R5030 a_12907_n2630.n5 a_12907_n2630.n4 0.665
R5031 a_13968_n7819.n7 a_13968_n7819.n6 861.987
R5032 a_13968_n7819.n6 a_13968_n7819.n5 560.726
R5033 a_13968_n7819.t6 a_13968_n7819.t9 415.315
R5034 a_13968_n7819.t19 a_13968_n7819.t8 415.315
R5035 a_13968_n7819.n2 a_13968_n7819.t4 394.151
R5036 a_13968_n7819.n5 a_13968_n7819.t13 294.653
R5037 a_13968_n7819.n1 a_13968_n7819.t7 269.523
R5038 a_13968_n7819.t4 a_13968_n7819.n1 269.523
R5039 a_13968_n7819.n9 a_13968_n7819.t6 217.716
R5040 a_13968_n7819.n8 a_13968_n7819.t11 214.335
R5041 a_13968_n7819.t9 a_13968_n7819.n8 214.335
R5042 a_13968_n7819.n0 a_13968_n7819.t15 214.335
R5043 a_13968_n7819.t8 a_13968_n7819.n0 214.335
R5044 a_13968_n7819.n7 a_13968_n7819.t19 198.921
R5045 a_13968_n7819.n3 a_13968_n7819.t12 198.043
R5046 a_13968_n7819.n12 a_13968_n7819.n11 192.754
R5047 a_13968_n7819.n1 a_13968_n7819.t5 160.666
R5048 a_13968_n7819.n5 a_13968_n7819.t18 111.663
R5049 a_13968_n7819.n4 a_13968_n7819.n2 97.816
R5050 a_13968_n7819.n3 a_13968_n7819.t16 93.989
R5051 a_13968_n7819.n8 a_13968_n7819.t10 80.333
R5052 a_13968_n7819.n2 a_13968_n7819.t17 80.333
R5053 a_13968_n7819.n0 a_13968_n7819.t14 80.333
R5054 a_13968_n7819.n6 a_13968_n7819.n4 65.07
R5055 a_13968_n7819.n11 a_13968_n7819.t2 28.568
R5056 a_13968_n7819.n12 a_13968_n7819.t1 28.565
R5057 a_13968_n7819.t0 a_13968_n7819.n12 28.565
R5058 a_13968_n7819.n10 a_13968_n7819.t3 18.826
R5059 a_13968_n7819.n9 a_13968_n7819.n7 16.411
R5060 a_13968_n7819.n4 a_13968_n7819.n3 6.615
R5061 a_13968_n7819.n10 a_13968_n7819.n9 5.027
R5062 a_13968_n7819.n11 a_13968_n7819.n10 1.101
R5063 a_18000_n5465.t0 a_18000_n5465.n0 14.282
R5064 a_18000_n5465.n0 a_18000_n5465.t1 14.282
R5065 a_18000_n5465.n0 a_18000_n5465.n9 0.999
R5066 a_18000_n5465.n6 a_18000_n5465.n8 0.575
R5067 a_18000_n5465.n9 a_18000_n5465.n6 0.2
R5068 a_18000_n5465.n9 a_18000_n5465.t9 16.058
R5069 a_18000_n5465.n8 a_18000_n5465.n7 0.999
R5070 a_18000_n5465.n7 a_18000_n5465.t11 14.282
R5071 a_18000_n5465.n7 a_18000_n5465.t10 14.282
R5072 a_18000_n5465.n8 a_18000_n5465.t8 16.058
R5073 a_18000_n5465.n6 a_18000_n5465.n4 0.227
R5074 a_18000_n5465.n4 a_18000_n5465.n5 1.511
R5075 a_18000_n5465.n5 a_18000_n5465.t4 14.282
R5076 a_18000_n5465.n5 a_18000_n5465.t3 14.282
R5077 a_18000_n5465.n4 a_18000_n5465.n1 0.669
R5078 a_18000_n5465.n1 a_18000_n5465.n2 0.001
R5079 a_18000_n5465.n1 a_18000_n5465.n3 267.767
R5080 a_18000_n5465.n3 a_18000_n5465.t6 14.282
R5081 a_18000_n5465.n3 a_18000_n5465.t5 14.282
R5082 a_18000_n5465.n2 a_18000_n5465.t2 14.282
R5083 a_18000_n5465.n2 a_18000_n5465.t7 14.282
R5084 a_704_n5517.n7 a_704_n5517.n6 861.987
R5085 a_704_n5517.n6 a_704_n5517.n5 560.726
R5086 a_704_n5517.t17 a_704_n5517.t19 415.315
R5087 a_704_n5517.t18 a_704_n5517.t7 415.315
R5088 a_704_n5517.n2 a_704_n5517.t6 394.151
R5089 a_704_n5517.n5 a_704_n5517.t14 294.653
R5090 a_704_n5517.n1 a_704_n5517.t5 269.523
R5091 a_704_n5517.t6 a_704_n5517.n1 269.523
R5092 a_704_n5517.n9 a_704_n5517.t17 217.716
R5093 a_704_n5517.n8 a_704_n5517.t11 214.335
R5094 a_704_n5517.t19 a_704_n5517.n8 214.335
R5095 a_704_n5517.n0 a_704_n5517.t9 214.335
R5096 a_704_n5517.t7 a_704_n5517.n0 214.335
R5097 a_704_n5517.n7 a_704_n5517.t18 198.921
R5098 a_704_n5517.n3 a_704_n5517.t12 198.043
R5099 a_704_n5517.n12 a_704_n5517.n11 192.754
R5100 a_704_n5517.n1 a_704_n5517.t4 160.666
R5101 a_704_n5517.n5 a_704_n5517.t16 111.663
R5102 a_704_n5517.n4 a_704_n5517.n2 97.816
R5103 a_704_n5517.n3 a_704_n5517.t13 93.989
R5104 a_704_n5517.n8 a_704_n5517.t10 80.333
R5105 a_704_n5517.n2 a_704_n5517.t15 80.333
R5106 a_704_n5517.n0 a_704_n5517.t8 80.333
R5107 a_704_n5517.n6 a_704_n5517.n4 65.07
R5108 a_704_n5517.n11 a_704_n5517.t3 28.568
R5109 a_704_n5517.n12 a_704_n5517.t2 28.565
R5110 a_704_n5517.t1 a_704_n5517.n12 28.565
R5111 a_704_n5517.n10 a_704_n5517.t0 18.825
R5112 a_704_n5517.n9 a_704_n5517.n7 16.411
R5113 a_704_n5517.n4 a_704_n5517.n3 6.615
R5114 a_704_n5517.n10 a_704_n5517.n9 2.988
R5115 a_704_n5517.n11 a_704_n5517.n10 1.105
R5116 a_4794_n5464.t0 a_4794_n5464.n0 14.282
R5117 a_4794_n5464.n0 a_4794_n5464.t10 14.282
R5118 a_4794_n5464.n0 a_4794_n5464.n9 0.999
R5119 a_4794_n5464.n6 a_4794_n5464.n8 0.575
R5120 a_4794_n5464.n9 a_4794_n5464.n6 0.2
R5121 a_4794_n5464.n9 a_4794_n5464.t11 16.058
R5122 a_4794_n5464.n8 a_4794_n5464.n7 0.999
R5123 a_4794_n5464.n7 a_4794_n5464.t2 14.282
R5124 a_4794_n5464.n7 a_4794_n5464.t3 14.282
R5125 a_4794_n5464.n8 a_4794_n5464.t1 16.058
R5126 a_4794_n5464.n6 a_4794_n5464.n4 0.227
R5127 a_4794_n5464.n4 a_4794_n5464.n5 1.511
R5128 a_4794_n5464.n5 a_4794_n5464.t7 14.282
R5129 a_4794_n5464.n5 a_4794_n5464.t9 14.282
R5130 a_4794_n5464.n4 a_4794_n5464.n1 0.669
R5131 a_4794_n5464.n1 a_4794_n5464.n2 0.001
R5132 a_4794_n5464.n1 a_4794_n5464.n3 267.767
R5133 a_4794_n5464.n3 a_4794_n5464.t6 14.282
R5134 a_4794_n5464.n3 a_4794_n5464.t4 14.282
R5135 a_4794_n5464.n2 a_4794_n5464.t8 14.282
R5136 a_4794_n5464.n2 a_4794_n5464.t5 14.282
R5137 a_22849_n4154.n0 a_22849_n4154.t8 214.335
R5138 a_22849_n4154.t10 a_22849_n4154.n0 214.335
R5139 a_22849_n4154.n1 a_22849_n4154.t10 143.851
R5140 a_22849_n4154.n1 a_22849_n4154.t9 135.658
R5141 a_22849_n4154.n0 a_22849_n4154.t7 80.333
R5142 a_22849_n4154.n2 a_22849_n4154.t4 28.565
R5143 a_22849_n4154.n2 a_22849_n4154.t5 28.565
R5144 a_22849_n4154.n4 a_22849_n4154.t6 28.565
R5145 a_22849_n4154.n4 a_22849_n4154.t1 28.565
R5146 a_22849_n4154.n7 a_22849_n4154.t0 28.565
R5147 a_22849_n4154.t2 a_22849_n4154.n7 28.565
R5148 a_22849_n4154.n6 a_22849_n4154.t3 9.714
R5149 a_22849_n4154.n7 a_22849_n4154.n6 1.003
R5150 a_22849_n4154.n5 a_22849_n4154.n3 0.833
R5151 a_22849_n4154.n3 a_22849_n4154.n2 0.653
R5152 a_22849_n4154.n5 a_22849_n4154.n4 0.653
R5153 a_22849_n4154.n6 a_22849_n4154.n5 0.341
R5154 a_22849_n4154.n3 a_22849_n4154.n1 0.032
R5155 a_23439_n4591.t4 a_23439_n4591.t6 574.43
R5156 a_23439_n4591.n0 a_23439_n4591.t7 285.109
R5157 a_23439_n4591.n2 a_23439_n4591.n1 211.136
R5158 a_23439_n4591.n4 a_23439_n4591.n3 192.754
R5159 a_23439_n4591.n0 a_23439_n4591.t5 160.666
R5160 a_23439_n4591.n1 a_23439_n4591.t4 160.666
R5161 a_23439_n4591.n1 a_23439_n4591.n0 114.829
R5162 a_23439_n4591.n3 a_23439_n4591.t2 28.568
R5163 a_23439_n4591.t3 a_23439_n4591.n4 28.565
R5164 a_23439_n4591.n4 a_23439_n4591.t1 28.565
R5165 a_23439_n4591.n2 a_23439_n4591.t0 19.084
R5166 a_23439_n4591.n3 a_23439_n4591.n2 1.051
R5167 a_13338_5442.n0 a_13338_5442.t7 214.335
R5168 a_13338_5442.t9 a_13338_5442.n0 214.335
R5169 a_13338_5442.n1 a_13338_5442.t9 143.851
R5170 a_13338_5442.n1 a_13338_5442.t10 135.658
R5171 a_13338_5442.n0 a_13338_5442.t8 80.333
R5172 a_13338_5442.n2 a_13338_5442.t3 28.565
R5173 a_13338_5442.n2 a_13338_5442.t5 28.565
R5174 a_13338_5442.n4 a_13338_5442.t4 28.565
R5175 a_13338_5442.n4 a_13338_5442.t2 28.565
R5176 a_13338_5442.n7 a_13338_5442.t6 28.565
R5177 a_13338_5442.t0 a_13338_5442.n7 28.565
R5178 a_13338_5442.n6 a_13338_5442.t1 9.714
R5179 a_13338_5442.n7 a_13338_5442.n6 1.003
R5180 a_13338_5442.n5 a_13338_5442.n3 0.833
R5181 a_13338_5442.n3 a_13338_5442.n2 0.653
R5182 a_13338_5442.n5 a_13338_5442.n4 0.653
R5183 a_13338_5442.n6 a_13338_5442.n5 0.341
R5184 a_13338_5442.n3 a_13338_5442.n1 0.032
R5185 a_13928_5005.n5 a_13928_5005.n4 535.449
R5186 a_13928_5005.t11 a_13928_5005.t13 437.233
R5187 a_13928_5005.t17 a_13928_5005.t16 437.233
R5188 a_13928_5005.t4 a_13928_5005.n2 313.873
R5189 a_13928_5005.n4 a_13928_5005.t10 294.986
R5190 a_13928_5005.n1 a_13928_5005.t14 272.288
R5191 a_13928_5005.n5 a_13928_5005.t5 245.184
R5192 a_13928_5005.n7 a_13928_5005.t17 218.628
R5193 a_13928_5005.n9 a_13928_5005.t11 217.024
R5194 a_13928_5005.n8 a_13928_5005.t6 214.686
R5195 a_13928_5005.t13 a_13928_5005.n8 214.686
R5196 a_13928_5005.n6 a_13928_5005.t9 214.686
R5197 a_13928_5005.t16 a_13928_5005.n6 214.686
R5198 a_13928_5005.n11 a_13928_5005.n0 192.754
R5199 a_13928_5005.n3 a_13928_5005.t4 190.152
R5200 a_13928_5005.n3 a_13928_5005.t18 190.152
R5201 a_13928_5005.n1 a_13928_5005.t7 160.666
R5202 a_13928_5005.n2 a_13928_5005.t15 160.666
R5203 a_13928_5005.n4 a_13928_5005.t8 110.859
R5204 a_13928_5005.n2 a_13928_5005.n1 96.129
R5205 a_13928_5005.n8 a_13928_5005.t19 80.333
R5206 a_13928_5005.t5 a_13928_5005.n3 80.333
R5207 a_13928_5005.n6 a_13928_5005.t12 80.333
R5208 a_13928_5005.t3 a_13928_5005.n11 28.568
R5209 a_13928_5005.n0 a_13928_5005.t2 28.565
R5210 a_13928_5005.n0 a_13928_5005.t1 28.565
R5211 a_13928_5005.n10 a_13928_5005.t0 20.07
R5212 a_13928_5005.n7 a_13928_5005.n5 14.9
R5213 a_13928_5005.n10 a_13928_5005.n9 3.139
R5214 a_13928_5005.n9 a_13928_5005.n7 2.599
R5215 a_13928_5005.n11 a_13928_5005.n10 1.101
R5216 a_10168_1277.t5 a_10168_1277.t6 574.43
R5217 a_10168_1277.n0 a_10168_1277.t7 285.109
R5218 a_10168_1277.n2 a_10168_1277.n1 211.136
R5219 a_10168_1277.n4 a_10168_1277.n3 192.754
R5220 a_10168_1277.n0 a_10168_1277.t4 160.666
R5221 a_10168_1277.n1 a_10168_1277.t5 160.666
R5222 a_10168_1277.n1 a_10168_1277.n0 114.829
R5223 a_10168_1277.n3 a_10168_1277.t2 28.568
R5224 a_10168_1277.t0 a_10168_1277.n4 28.565
R5225 a_10168_1277.n4 a_10168_1277.t3 28.565
R5226 a_10168_1277.n2 a_10168_1277.t1 19.084
R5227 a_10168_1277.n3 a_10168_1277.n2 1.051
R5228 a_13031_3240.n0 a_13031_3240.t5 14.282
R5229 a_13031_3240.n0 a_13031_3240.t2 14.282
R5230 a_13031_3240.n1 a_13031_3240.t4 14.282
R5231 a_13031_3240.n1 a_13031_3240.t3 14.282
R5232 a_13031_3240.n3 a_13031_3240.t1 14.282
R5233 a_13031_3240.t0 a_13031_3240.n3 14.282
R5234 a_13031_3240.n3 a_13031_3240.n2 2.546
R5235 a_13031_3240.n2 a_13031_3240.n1 2.367
R5236 a_13031_3240.n2 a_13031_3240.n0 0.001
R5237 a_12913_3240.t6 a_12913_3240.n2 404.877
R5238 a_12913_3240.n1 a_12913_3240.t8 210.902
R5239 a_12913_3240.n3 a_12913_3240.t6 136.943
R5240 a_12913_3240.n2 a_12913_3240.n1 107.801
R5241 a_12913_3240.n1 a_12913_3240.t5 80.333
R5242 a_12913_3240.n2 a_12913_3240.t7 80.333
R5243 a_12913_3240.n0 a_12913_3240.t4 17.4
R5244 a_12913_3240.n0 a_12913_3240.t0 17.4
R5245 a_12913_3240.n4 a_12913_3240.t2 15.032
R5246 a_12913_3240.n5 a_12913_3240.t1 14.282
R5247 a_12913_3240.t3 a_12913_3240.n5 14.282
R5248 a_12913_3240.n5 a_12913_3240.n4 1.65
R5249 a_12913_3240.n3 a_12913_3240.n0 0.672
R5250 a_12913_3240.n4 a_12913_3240.n3 0.665
R5251 a_20582_5026.n4 a_20582_5026.n3 535.449
R5252 a_20582_5026.t15 a_20582_5026.t13 437.233
R5253 a_20582_5026.t19 a_20582_5026.t4 437.233
R5254 a_20582_5026.t18 a_20582_5026.n1 313.873
R5255 a_20582_5026.n3 a_20582_5026.t17 294.986
R5256 a_20582_5026.n0 a_20582_5026.t5 272.288
R5257 a_20582_5026.n4 a_20582_5026.t8 245.184
R5258 a_20582_5026.n6 a_20582_5026.t19 218.628
R5259 a_20582_5026.n8 a_20582_5026.t15 217.024
R5260 a_20582_5026.n7 a_20582_5026.t10 214.686
R5261 a_20582_5026.t13 a_20582_5026.n7 214.686
R5262 a_20582_5026.n5 a_20582_5026.t7 214.686
R5263 a_20582_5026.t4 a_20582_5026.n5 214.686
R5264 a_20582_5026.n11 a_20582_5026.n10 192.754
R5265 a_20582_5026.n2 a_20582_5026.t18 190.152
R5266 a_20582_5026.n2 a_20582_5026.t14 190.152
R5267 a_20582_5026.n0 a_20582_5026.t12 160.666
R5268 a_20582_5026.n1 a_20582_5026.t6 160.666
R5269 a_20582_5026.n3 a_20582_5026.t9 110.859
R5270 a_20582_5026.n1 a_20582_5026.n0 96.129
R5271 a_20582_5026.n7 a_20582_5026.t16 80.333
R5272 a_20582_5026.t8 a_20582_5026.n2 80.333
R5273 a_20582_5026.n5 a_20582_5026.t11 80.333
R5274 a_20582_5026.n10 a_20582_5026.t2 28.568
R5275 a_20582_5026.n11 a_20582_5026.t3 28.565
R5276 a_20582_5026.t0 a_20582_5026.n11 28.565
R5277 a_20582_5026.n9 a_20582_5026.t1 18.823
R5278 a_20582_5026.n6 a_20582_5026.n4 14.9
R5279 a_20582_5026.n9 a_20582_5026.n8 3.074
R5280 a_20582_5026.n8 a_20582_5026.n6 2.599
R5281 a_20582_5026.n10 a_20582_5026.n9 1.105
R5282 a_22852_110.n2 a_22852_110.t7 214.335
R5283 a_22852_110.t9 a_22852_110.n2 214.335
R5284 a_22852_110.n3 a_22852_110.t9 143.851
R5285 a_22852_110.n3 a_22852_110.t10 135.658
R5286 a_22852_110.n2 a_22852_110.t8 80.333
R5287 a_22852_110.n4 a_22852_110.t6 28.565
R5288 a_22852_110.n4 a_22852_110.t5 28.565
R5289 a_22852_110.n0 a_22852_110.t0 28.565
R5290 a_22852_110.n0 a_22852_110.t1 28.565
R5291 a_22852_110.t4 a_22852_110.n7 28.565
R5292 a_22852_110.n7 a_22852_110.t2 28.565
R5293 a_22852_110.n1 a_22852_110.t3 9.714
R5294 a_22852_110.n1 a_22852_110.n0 1.003
R5295 a_22852_110.n6 a_22852_110.n5 0.833
R5296 a_22852_110.n5 a_22852_110.n4 0.653
R5297 a_22852_110.n7 a_22852_110.n6 0.653
R5298 a_22852_110.n6 a_22852_110.n1 0.341
R5299 a_22852_110.n5 a_22852_110.n3 0.032
R5300 a_26940_378.n1 a_26940_378.t4 318.922
R5301 a_26940_378.n0 a_26940_378.t5 274.739
R5302 a_26940_378.n0 a_26940_378.t6 274.739
R5303 a_26940_378.n1 a_26940_378.t7 269.116
R5304 a_26940_378.t4 a_26940_378.n0 179.946
R5305 a_26940_378.n2 a_26940_378.n1 105.178
R5306 a_26940_378.n3 a_26940_378.t3 29.444
R5307 a_26940_378.t0 a_26940_378.n4 28.565
R5308 a_26940_378.n4 a_26940_378.t2 28.565
R5309 a_26940_378.n2 a_26940_378.t1 18.145
R5310 a_26940_378.n3 a_26940_378.n2 2.878
R5311 a_26940_378.n4 a_26940_378.n3 0.764
R5312 a_26528_404.n0 a_26528_404.n9 1.511
R5313 a_26528_404.n0 a_26528_404.t10 14.282
R5314 a_26528_404.t0 a_26528_404.n0 14.282
R5315 a_26528_404.n9 a_26528_404.n5 0.227
R5316 a_26528_404.n9 a_26528_404.n6 0.669
R5317 a_26528_404.n6 a_26528_404.n7 0.001
R5318 a_26528_404.n6 a_26528_404.n8 267.767
R5319 a_26528_404.n8 a_26528_404.t9 14.282
R5320 a_26528_404.n8 a_26528_404.t7 14.282
R5321 a_26528_404.n7 a_26528_404.t11 14.282
R5322 a_26528_404.n7 a_26528_404.t8 14.282
R5323 a_26528_404.n5 a_26528_404.n2 0.575
R5324 a_26528_404.n5 a_26528_404.n4 0.2
R5325 a_26528_404.n4 a_26528_404.t5 16.058
R5326 a_26528_404.n4 a_26528_404.n3 0.999
R5327 a_26528_404.n3 a_26528_404.t6 14.282
R5328 a_26528_404.n3 a_26528_404.t4 14.282
R5329 a_26528_404.n2 a_26528_404.n1 0.999
R5330 a_26528_404.n1 a_26528_404.t1 14.282
R5331 a_26528_404.n1 a_26528_404.t3 14.282
R5332 a_26528_404.n2 a_26528_404.t2 16.058
R5333 Y[6] Y[6].n6 224.816
R5334 Y[6].n4 Y[6].n2 157.665
R5335 Y[6].n4 Y[6].n3 122.999
R5336 Y[6].n6 Y[6].n0 90.436
R5337 Y[6].n5 Y[6].n1 90.416
R5338 Y[6].n6 Y[6].n5 74.302
R5339 Y[6].n5 Y[6].n4 50.575
R5340 Y[6].n0 Y[6].t4 14.282
R5341 Y[6].n0 Y[6].t6 14.282
R5342 Y[6].n1 Y[6].t5 14.282
R5343 Y[6].n1 Y[6].t2 14.282
R5344 Y[6].n3 Y[6].t0 14.282
R5345 Y[6].n3 Y[6].t1 14.282
R5346 Y[6].n2 Y[6].t7 8.7
R5347 Y[6].n2 Y[6].t3 8.7
R5348 a_13378_n8256.n0 a_13378_n8256.t9 214.335
R5349 a_13378_n8256.t7 a_13378_n8256.n0 214.335
R5350 a_13378_n8256.n1 a_13378_n8256.t7 143.85
R5351 a_13378_n8256.n1 a_13378_n8256.t10 135.66
R5352 a_13378_n8256.n0 a_13378_n8256.t8 80.333
R5353 a_13378_n8256.n2 a_13378_n8256.t4 28.565
R5354 a_13378_n8256.n2 a_13378_n8256.t5 28.565
R5355 a_13378_n8256.n4 a_13378_n8256.t6 28.565
R5356 a_13378_n8256.n4 a_13378_n8256.t3 28.565
R5357 a_13378_n8256.t0 a_13378_n8256.n7 28.565
R5358 a_13378_n8256.n7 a_13378_n8256.t1 28.565
R5359 a_13378_n8256.n3 a_13378_n8256.t2 9.714
R5360 a_13378_n8256.n3 a_13378_n8256.n2 1.003
R5361 a_13378_n8256.n6 a_13378_n8256.n5 0.836
R5362 a_13378_n8256.n5 a_13378_n8256.n4 0.653
R5363 a_13378_n8256.n7 a_13378_n8256.n6 0.65
R5364 a_13378_n8256.n5 a_13378_n8256.n3 0.341
R5365 a_13378_n8256.n6 a_13378_n8256.n1 0.032
R5366 a_28640_2725.n2 a_28640_2725.t8 214.335
R5367 a_28640_2725.t7 a_28640_2725.n2 214.335
R5368 a_28640_2725.n3 a_28640_2725.t7 143.851
R5369 a_28640_2725.n3 a_28640_2725.t10 135.658
R5370 a_28640_2725.n2 a_28640_2725.t9 80.333
R5371 a_28640_2725.n4 a_28640_2725.t6 28.565
R5372 a_28640_2725.n4 a_28640_2725.t4 28.565
R5373 a_28640_2725.n0 a_28640_2725.t0 28.565
R5374 a_28640_2725.n0 a_28640_2725.t1 28.565
R5375 a_28640_2725.n7 a_28640_2725.t5 28.565
R5376 a_28640_2725.t2 a_28640_2725.n7 28.565
R5377 a_28640_2725.n1 a_28640_2725.t3 9.714
R5378 a_28640_2725.n1 a_28640_2725.n0 1.003
R5379 a_28640_2725.n6 a_28640_2725.n5 0.833
R5380 a_28640_2725.n5 a_28640_2725.n4 0.653
R5381 a_28640_2725.n7 a_28640_2725.n6 0.653
R5382 a_28640_2725.n6 a_28640_2725.n1 0.341
R5383 a_28640_2725.n5 a_28640_2725.n3 0.032
R5384 a_29230_2288.n4 a_29230_2288.n3 563.136
R5385 a_29230_2288.t14 a_29230_2288.t8 437.233
R5386 a_29230_2288.t15 a_29230_2288.n1 313.873
R5387 a_29230_2288.n3 a_29230_2288.t11 294.986
R5388 a_29230_2288.n0 a_29230_2288.t5 272.288
R5389 a_29230_2288.n6 a_29230_2288.t14 217.824
R5390 a_29230_2288.n5 a_29230_2288.t6 214.686
R5391 a_29230_2288.t8 a_29230_2288.n5 214.686
R5392 a_29230_2288.n9 a_29230_2288.n8 192.754
R5393 a_29230_2288.n2 a_29230_2288.t15 190.152
R5394 a_29230_2288.n2 a_29230_2288.t4 190.152
R5395 a_29230_2288.n4 a_29230_2288.t9 178.973
R5396 a_29230_2288.n0 a_29230_2288.t12 160.666
R5397 a_29230_2288.n1 a_29230_2288.t7 160.666
R5398 a_29230_2288.n6 a_29230_2288.n4 133.838
R5399 a_29230_2288.n3 a_29230_2288.t10 110.859
R5400 a_29230_2288.n1 a_29230_2288.n0 96.129
R5401 a_29230_2288.t9 a_29230_2288.n2 80.333
R5402 a_29230_2288.n5 a_29230_2288.t13 80.333
R5403 a_29230_2288.n8 a_29230_2288.t2 28.568
R5404 a_29230_2288.n9 a_29230_2288.t1 28.565
R5405 a_29230_2288.t3 a_29230_2288.n9 28.565
R5406 a_29230_2288.n7 a_29230_2288.t0 18.822
R5407 a_29230_2288.n7 a_29230_2288.n6 5.647
R5408 a_29230_2288.n8 a_29230_2288.n7 1.105
R5409 a_19992_5463.n0 a_19992_5463.t9 214.335
R5410 a_19992_5463.t7 a_19992_5463.n0 214.335
R5411 a_19992_5463.n1 a_19992_5463.t7 143.851
R5412 a_19992_5463.n1 a_19992_5463.t8 135.658
R5413 a_19992_5463.n0 a_19992_5463.t10 80.333
R5414 a_19992_5463.n2 a_19992_5463.t4 28.565
R5415 a_19992_5463.n2 a_19992_5463.t5 28.565
R5416 a_19992_5463.n4 a_19992_5463.t3 28.565
R5417 a_19992_5463.n4 a_19992_5463.t2 28.565
R5418 a_19992_5463.t0 a_19992_5463.n7 28.565
R5419 a_19992_5463.n7 a_19992_5463.t6 28.565
R5420 a_19992_5463.n6 a_19992_5463.t1 9.714
R5421 a_19992_5463.n7 a_19992_5463.n6 1.003
R5422 a_19992_5463.n5 a_19992_5463.n3 0.833
R5423 a_19992_5463.n3 a_19992_5463.n2 0.653
R5424 a_19992_5463.n5 a_19992_5463.n4 0.653
R5425 a_19992_5463.n6 a_19992_5463.n5 0.341
R5426 a_19992_5463.n3 a_19992_5463.n1 0.032
R5427 a_12029_n3217.t5 a_12029_n3217.t4 800.071
R5428 a_12029_n3217.n3 a_12029_n3217.n2 672.951
R5429 a_12029_n3217.n1 a_12029_n3217.t7 285.109
R5430 a_12029_n3217.n2 a_12029_n3217.t5 193.602
R5431 a_12029_n3217.n1 a_12029_n3217.t6 160.666
R5432 a_12029_n3217.n2 a_12029_n3217.n1 91.507
R5433 a_12029_n3217.t0 a_12029_n3217.n4 28.57
R5434 a_12029_n3217.n0 a_12029_n3217.t3 28.565
R5435 a_12029_n3217.n0 a_12029_n3217.t1 28.565
R5436 a_12029_n3217.n4 a_12029_n3217.t2 17.638
R5437 a_12029_n3217.n3 a_12029_n3217.n0 0.69
R5438 a_12029_n3217.n4 a_12029_n3217.n3 0.6
R5439 a_28711_n2228.n0 a_28711_n2228.t9 214.335
R5440 a_28711_n2228.t7 a_28711_n2228.n0 214.335
R5441 a_28711_n2228.n1 a_28711_n2228.t7 143.851
R5442 a_28711_n2228.n1 a_28711_n2228.t10 135.658
R5443 a_28711_n2228.n0 a_28711_n2228.t8 80.333
R5444 a_28711_n2228.n2 a_28711_n2228.t4 28.565
R5445 a_28711_n2228.n2 a_28711_n2228.t5 28.565
R5446 a_28711_n2228.n4 a_28711_n2228.t6 28.565
R5447 a_28711_n2228.n4 a_28711_n2228.t1 28.565
R5448 a_28711_n2228.n7 a_28711_n2228.t2 28.565
R5449 a_28711_n2228.t3 a_28711_n2228.n7 28.565
R5450 a_28711_n2228.n6 a_28711_n2228.t0 9.714
R5451 a_28711_n2228.n7 a_28711_n2228.n6 1.003
R5452 a_28711_n2228.n5 a_28711_n2228.n3 0.833
R5453 a_28711_n2228.n3 a_28711_n2228.n2 0.653
R5454 a_28711_n2228.n5 a_28711_n2228.n4 0.653
R5455 a_28711_n2228.n6 a_28711_n2228.n5 0.341
R5456 a_28711_n2228.n3 a_28711_n2228.n1 0.032
R5457 a_11763_378.n1 a_11763_378.t5 318.922
R5458 a_11763_378.n0 a_11763_378.t6 274.739
R5459 a_11763_378.n0 a_11763_378.t4 274.739
R5460 a_11763_378.n1 a_11763_378.t7 269.116
R5461 a_11763_378.t5 a_11763_378.n0 179.946
R5462 a_11763_378.n2 a_11763_378.n1 107.263
R5463 a_11763_378.n3 a_11763_378.t1 29.444
R5464 a_11763_378.t3 a_11763_378.n4 28.565
R5465 a_11763_378.n4 a_11763_378.t2 28.565
R5466 a_11763_378.n2 a_11763_378.t0 18.145
R5467 a_11763_378.n3 a_11763_378.n2 2.878
R5468 a_11763_378.n4 a_11763_378.n3 0.764
R5469 a_11351_404.n0 a_11351_404.n1 0.001
R5470 a_11351_404.t3 a_11351_404.n0 14.282
R5471 a_11351_404.n0 a_11351_404.t5 14.282
R5472 a_11351_404.n1 a_11351_404.n9 267.767
R5473 a_11351_404.n9 a_11351_404.t7 14.282
R5474 a_11351_404.n9 a_11351_404.t6 14.282
R5475 a_11351_404.n1 a_11351_404.n7 0.669
R5476 a_11351_404.n7 a_11351_404.n8 1.511
R5477 a_11351_404.n8 a_11351_404.t4 14.282
R5478 a_11351_404.n8 a_11351_404.t11 14.282
R5479 a_11351_404.n7 a_11351_404.n6 0.227
R5480 a_11351_404.n6 a_11351_404.n3 0.575
R5481 a_11351_404.n6 a_11351_404.n5 0.2
R5482 a_11351_404.n5 a_11351_404.t2 16.058
R5483 a_11351_404.n5 a_11351_404.n4 0.999
R5484 a_11351_404.n4 a_11351_404.t0 14.282
R5485 a_11351_404.n4 a_11351_404.t1 14.282
R5486 a_11351_404.n3 a_11351_404.n2 0.999
R5487 a_11351_404.n2 a_11351_404.t8 14.282
R5488 a_11351_404.n2 a_11351_404.t10 14.282
R5489 a_11351_404.n3 a_11351_404.t9 16.058
R5490 a_29230_n745.n4 a_29230_n745.n3 563.136
R5491 a_29230_n745.t5 a_29230_n745.t9 437.233
R5492 a_29230_n745.t10 a_29230_n745.n1 313.873
R5493 a_29230_n745.n3 a_29230_n745.t6 294.986
R5494 a_29230_n745.n0 a_29230_n745.t15 272.288
R5495 a_29230_n745.n6 a_29230_n745.t5 217.824
R5496 a_29230_n745.n5 a_29230_n745.t11 214.686
R5497 a_29230_n745.t9 a_29230_n745.n5 214.686
R5498 a_29230_n745.n9 a_29230_n745.n8 192.754
R5499 a_29230_n745.n2 a_29230_n745.t10 190.152
R5500 a_29230_n745.n2 a_29230_n745.t4 190.152
R5501 a_29230_n745.n4 a_29230_n745.t7 178.973
R5502 a_29230_n745.n0 a_29230_n745.t14 160.666
R5503 a_29230_n745.n1 a_29230_n745.t13 160.666
R5504 a_29230_n745.n6 a_29230_n745.n4 133.838
R5505 a_29230_n745.n3 a_29230_n745.t8 110.859
R5506 a_29230_n745.n1 a_29230_n745.n0 96.129
R5507 a_29230_n745.t7 a_29230_n745.n2 80.333
R5508 a_29230_n745.n5 a_29230_n745.t12 80.333
R5509 a_29230_n745.n8 a_29230_n745.t1 28.568
R5510 a_29230_n745.t3 a_29230_n745.n9 28.565
R5511 a_29230_n745.n9 a_29230_n745.t2 28.565
R5512 a_29230_n745.n7 a_29230_n745.t0 18.824
R5513 a_29230_n745.n7 a_29230_n745.n6 5.567
R5514 a_29230_n745.n8 a_29230_n745.n7 1.105
R5515 a_30762_4198.t6 a_30762_4198.n7 16.058
R5516 a_30762_4198.n7 a_30762_4198.n5 0.575
R5517 a_30762_4198.n5 a_30762_4198.n9 0.2
R5518 a_30762_4198.n9 a_30762_4198.t11 16.058
R5519 a_30762_4198.n9 a_30762_4198.n8 0.999
R5520 a_30762_4198.n8 a_30762_4198.t8 14.282
R5521 a_30762_4198.n8 a_30762_4198.t7 14.282
R5522 a_30762_4198.n7 a_30762_4198.n6 0.999
R5523 a_30762_4198.n6 a_30762_4198.t9 14.282
R5524 a_30762_4198.n6 a_30762_4198.t10 14.282
R5525 a_30762_4198.n5 a_30762_4198.n3 0.227
R5526 a_30762_4198.n3 a_30762_4198.n4 1.511
R5527 a_30762_4198.n4 a_30762_4198.t2 14.282
R5528 a_30762_4198.n4 a_30762_4198.t0 14.282
R5529 a_30762_4198.n3 a_30762_4198.n0 0.669
R5530 a_30762_4198.n0 a_30762_4198.n1 0.001
R5531 a_30762_4198.n0 a_30762_4198.n2 267.767
R5532 a_30762_4198.n2 a_30762_4198.t3 14.282
R5533 a_30762_4198.n2 a_30762_4198.t4 14.282
R5534 a_30762_4198.n1 a_30762_4198.t1 14.282
R5535 a_30762_4198.n1 a_30762_4198.t5 14.282
R5536 a_18412_n5491.n1 a_18412_n5491.t7 318.922
R5537 a_18412_n5491.n0 a_18412_n5491.t6 274.739
R5538 a_18412_n5491.n0 a_18412_n5491.t4 274.739
R5539 a_18412_n5491.n1 a_18412_n5491.t5 269.116
R5540 a_18412_n5491.t7 a_18412_n5491.n0 179.946
R5541 a_18412_n5491.n2 a_18412_n5491.n1 107.263
R5542 a_18412_n5491.n3 a_18412_n5491.t1 29.444
R5543 a_18412_n5491.t3 a_18412_n5491.n4 28.565
R5544 a_18412_n5491.n4 a_18412_n5491.t2 28.565
R5545 a_18412_n5491.n2 a_18412_n5491.t0 18.145
R5546 a_18412_n5491.n3 a_18412_n5491.n2 2.878
R5547 a_18412_n5491.n4 a_18412_n5491.n3 0.764
R5548 a_9567_n5760.n0 a_9567_n5760.t9 214.335
R5549 a_9567_n5760.t7 a_9567_n5760.n0 214.335
R5550 a_9567_n5760.n1 a_9567_n5760.t7 143.851
R5551 a_9567_n5760.n1 a_9567_n5760.t10 135.658
R5552 a_9567_n5760.n0 a_9567_n5760.t8 80.333
R5553 a_9567_n5760.n2 a_9567_n5760.t6 28.565
R5554 a_9567_n5760.n2 a_9567_n5760.t4 28.565
R5555 a_9567_n5760.n4 a_9567_n5760.t5 28.565
R5556 a_9567_n5760.n4 a_9567_n5760.t1 28.565
R5557 a_9567_n5760.t0 a_9567_n5760.n7 28.565
R5558 a_9567_n5760.n7 a_9567_n5760.t3 28.565
R5559 a_9567_n5760.n6 a_9567_n5760.t2 9.714
R5560 a_9567_n5760.n7 a_9567_n5760.n6 1.003
R5561 a_9567_n5760.n5 a_9567_n5760.n3 0.833
R5562 a_9567_n5760.n3 a_9567_n5760.n2 0.653
R5563 a_9567_n5760.n5 a_9567_n5760.n4 0.653
R5564 a_9567_n5760.n6 a_9567_n5760.n5 0.341
R5565 a_9567_n5760.n3 a_9567_n5760.n1 0.032
R5566 a_31174_4172.n1 a_31174_4172.t6 318.922
R5567 a_31174_4172.n0 a_31174_4172.t7 274.739
R5568 a_31174_4172.n0 a_31174_4172.t4 274.739
R5569 a_31174_4172.n1 a_31174_4172.t5 269.116
R5570 a_31174_4172.t6 a_31174_4172.n0 179.946
R5571 a_31174_4172.n2 a_31174_4172.n1 107.263
R5572 a_31174_4172.t3 a_31174_4172.n4 29.444
R5573 a_31174_4172.n3 a_31174_4172.t2 28.565
R5574 a_31174_4172.n3 a_31174_4172.t1 28.565
R5575 a_31174_4172.n2 a_31174_4172.t0 18.145
R5576 a_31174_4172.n4 a_31174_4172.n2 2.878
R5577 a_31174_4172.n4 a_31174_4172.n3 0.764
R5578 Y[2].n4 Y[2].n2 157.665
R5579 Y[2] Y[2].n6 145.593
R5580 Y[2].n4 Y[2].n3 122.999
R5581 Y[2].n6 Y[2].n0 90.436
R5582 Y[2].n5 Y[2].n1 90.416
R5583 Y[2].n6 Y[2].n5 74.302
R5584 Y[2].n5 Y[2].n4 50.575
R5585 Y[2].n0 Y[2].t7 14.282
R5586 Y[2].n0 Y[2].t6 14.282
R5587 Y[2].n1 Y[2].t5 14.282
R5588 Y[2].n1 Y[2].t4 14.282
R5589 Y[2].n3 Y[2].t3 14.282
R5590 Y[2].n3 Y[2].t2 14.282
R5591 Y[2].n2 Y[2].t0 8.7
R5592 Y[2].n2 Y[2].t1 8.7
R5593 A[3].n2 A[3].t10 2858.78
R5594 A[3].n6 A[3].n2 2573.2
R5595 A[3].t10 A[3].t11 437.233
R5596 A[3].t12 A[3].t13 415.315
R5597 A[3].t14 A[3].t3 415.315
R5598 A[3].t15 A[3].t8 415.315
R5599 A[3].n5 A[3].t15 238.523
R5600 A[3].n5 A[3].t14 217.897
R5601 A[3].n2 A[3].t12 217.528
R5602 A[3].n1 A[3].t6 214.686
R5603 A[3].t11 A[3].n1 214.686
R5604 A[3].n0 A[3].t7 214.335
R5605 A[3].t13 A[3].n0 214.335
R5606 A[3].n3 A[3].t5 214.335
R5607 A[3].t3 A[3].n3 214.335
R5608 A[3].n4 A[3].t1 214.335
R5609 A[3].t8 A[3].n4 214.335
R5610 A[3].n0 A[3].t0 80.333
R5611 A[3].n1 A[3].t2 80.333
R5612 A[3].n3 A[3].t4 80.333
R5613 A[3].n4 A[3].t9 80.333
R5614 A[3] A[3].n6 0.607
R5615 A[3].n6 A[3].n5 0.274
R5616 a_6789_5443.n0 a_6789_5443.t9 214.335
R5617 a_6789_5443.t7 a_6789_5443.n0 214.335
R5618 a_6789_5443.n1 a_6789_5443.t7 143.851
R5619 a_6789_5443.n1 a_6789_5443.t8 135.658
R5620 a_6789_5443.n0 a_6789_5443.t10 80.333
R5621 a_6789_5443.n2 a_6789_5443.t5 28.565
R5622 a_6789_5443.n2 a_6789_5443.t6 28.565
R5623 a_6789_5443.n4 a_6789_5443.t4 28.565
R5624 a_6789_5443.n4 a_6789_5443.t2 28.565
R5625 a_6789_5443.n7 a_6789_5443.t1 28.565
R5626 a_6789_5443.t3 a_6789_5443.n7 28.565
R5627 a_6789_5443.n6 a_6789_5443.t0 9.714
R5628 a_6789_5443.n7 a_6789_5443.n6 1.003
R5629 a_6789_5443.n5 a_6789_5443.n3 0.833
R5630 a_6789_5443.n3 a_6789_5443.n2 0.653
R5631 a_6789_5443.n5 a_6789_5443.n4 0.653
R5632 a_6789_5443.n6 a_6789_5443.n5 0.341
R5633 a_6789_5443.n3 a_6789_5443.n1 0.032
R5634 a_16808_2859.t4 a_16808_2859.t5 800.071
R5635 a_16808_2859.n3 a_16808_2859.n2 659.097
R5636 a_16808_2859.n1 a_16808_2859.t7 285.109
R5637 a_16808_2859.n2 a_16808_2859.t4 193.602
R5638 a_16808_2859.n4 a_16808_2859.n0 192.754
R5639 a_16808_2859.n1 a_16808_2859.t6 160.666
R5640 a_16808_2859.n2 a_16808_2859.n1 91.507
R5641 a_16808_2859.t3 a_16808_2859.n4 28.568
R5642 a_16808_2859.n0 a_16808_2859.t2 28.565
R5643 a_16808_2859.n0 a_16808_2859.t1 28.565
R5644 a_16808_2859.n3 a_16808_2859.t0 19.061
R5645 a_16808_2859.n4 a_16808_2859.n3 1.005
R5646 a_22843_3364.n0 a_22843_3364.t7 214.335
R5647 a_22843_3364.t9 a_22843_3364.n0 214.335
R5648 a_22843_3364.n1 a_22843_3364.t9 143.851
R5649 a_22843_3364.n1 a_22843_3364.t8 135.658
R5650 a_22843_3364.n0 a_22843_3364.t10 80.333
R5651 a_22843_3364.n2 a_22843_3364.t5 28.565
R5652 a_22843_3364.n2 a_22843_3364.t4 28.565
R5653 a_22843_3364.n4 a_22843_3364.t6 28.565
R5654 a_22843_3364.n4 a_22843_3364.t1 28.565
R5655 a_22843_3364.n7 a_22843_3364.t0 28.565
R5656 a_22843_3364.t2 a_22843_3364.n7 28.565
R5657 a_22843_3364.n6 a_22843_3364.t3 9.714
R5658 a_22843_3364.n7 a_22843_3364.n6 1.003
R5659 a_22843_3364.n5 a_22843_3364.n3 0.833
R5660 a_22843_3364.n3 a_22843_3364.n2 0.653
R5661 a_22843_3364.n5 a_22843_3364.n4 0.653
R5662 a_22843_3364.n6 a_22843_3364.n5 0.341
R5663 a_22843_3364.n3 a_22843_3364.n1 0.032
R5664 a_23433_2927.t6 a_23433_2927.t5 800.071
R5665 a_23433_2927.n3 a_23433_2927.n2 659.097
R5666 a_23433_2927.n1 a_23433_2927.t7 285.109
R5667 a_23433_2927.n2 a_23433_2927.t6 193.602
R5668 a_23433_2927.n4 a_23433_2927.n0 192.754
R5669 a_23433_2927.n1 a_23433_2927.t4 160.666
R5670 a_23433_2927.n2 a_23433_2927.n1 91.507
R5671 a_23433_2927.t3 a_23433_2927.n4 28.568
R5672 a_23433_2927.n0 a_23433_2927.t1 28.565
R5673 a_23433_2927.n0 a_23433_2927.t2 28.565
R5674 a_23433_2927.n3 a_23433_2927.t0 19.061
R5675 a_23433_2927.n4 a_23433_2927.n3 1.005
R5676 a_22797_1688.n6 a_22797_1688.n5 501.28
R5677 a_22797_1688.t5 a_22797_1688.t16 437.233
R5678 a_22797_1688.t12 a_22797_1688.t17 415.315
R5679 a_22797_1688.t10 a_22797_1688.n3 313.873
R5680 a_22797_1688.n5 a_22797_1688.t6 294.986
R5681 a_22797_1688.n2 a_22797_1688.t7 272.288
R5682 a_22797_1688.n6 a_22797_1688.t18 236.01
R5683 a_22797_1688.n9 a_22797_1688.t5 216.627
R5684 a_22797_1688.n7 a_22797_1688.t12 216.111
R5685 a_22797_1688.n8 a_22797_1688.t9 214.686
R5686 a_22797_1688.t16 a_22797_1688.n8 214.686
R5687 a_22797_1688.n1 a_22797_1688.t11 214.335
R5688 a_22797_1688.t17 a_22797_1688.n1 214.335
R5689 a_22797_1688.n4 a_22797_1688.t10 190.152
R5690 a_22797_1688.n4 a_22797_1688.t8 190.152
R5691 a_22797_1688.n2 a_22797_1688.t4 160.666
R5692 a_22797_1688.n3 a_22797_1688.t14 160.666
R5693 a_22797_1688.n7 a_22797_1688.n6 148.428
R5694 a_22797_1688.n5 a_22797_1688.t19 110.859
R5695 a_22797_1688.n3 a_22797_1688.n2 96.129
R5696 a_22797_1688.n8 a_22797_1688.t15 80.333
R5697 a_22797_1688.n1 a_22797_1688.t13 80.333
R5698 a_22797_1688.t18 a_22797_1688.n4 80.333
R5699 a_22797_1688.n0 a_22797_1688.t2 28.57
R5700 a_22797_1688.n11 a_22797_1688.t3 28.565
R5701 a_22797_1688.t0 a_22797_1688.n11 28.565
R5702 a_22797_1688.n0 a_22797_1688.t1 17.638
R5703 a_22797_1688.n10 a_22797_1688.n9 11.942
R5704 a_22797_1688.n9 a_22797_1688.n7 2.923
R5705 a_22797_1688.n11 a_22797_1688.n10 0.69
R5706 a_22797_1688.n10 a_22797_1688.n0 0.6
R5707 a_6273_1009.n1 a_6273_1009.t5 318.922
R5708 a_6273_1009.n0 a_6273_1009.t7 273.935
R5709 a_6273_1009.n0 a_6273_1009.t4 273.935
R5710 a_6273_1009.n1 a_6273_1009.t6 269.116
R5711 a_6273_1009.n4 a_6273_1009.n3 193.227
R5712 a_6273_1009.t5 a_6273_1009.n0 179.142
R5713 a_6273_1009.n2 a_6273_1009.n1 106.999
R5714 a_6273_1009.n3 a_6273_1009.t2 28.568
R5715 a_6273_1009.n4 a_6273_1009.t1 28.565
R5716 a_6273_1009.t3 a_6273_1009.n4 28.565
R5717 a_6273_1009.n2 a_6273_1009.t0 18.149
R5718 a_6273_1009.n3 a_6273_1009.n2 3.726
R5719 a_18359_n396.t0 a_18359_n396.t1 17.4
R5720 a_16450_n3142.t0 a_16450_n3142.t1 17.4
R5721 a_20310_n5491.n1 a_20310_n5491.t5 318.922
R5722 a_20310_n5491.n0 a_20310_n5491.t7 274.739
R5723 a_20310_n5491.n0 a_20310_n5491.t6 274.739
R5724 a_20310_n5491.n1 a_20310_n5491.t4 269.116
R5725 a_20310_n5491.t5 a_20310_n5491.n0 179.946
R5726 a_20310_n5491.n2 a_20310_n5491.n1 105.178
R5727 a_20310_n5491.t1 a_20310_n5491.n4 29.444
R5728 a_20310_n5491.n3 a_20310_n5491.t2 28.565
R5729 a_20310_n5491.n3 a_20310_n5491.t3 28.565
R5730 a_20310_n5491.n2 a_20310_n5491.t0 18.145
R5731 a_20310_n5491.n4 a_20310_n5491.n2 2.878
R5732 a_20310_n5491.n4 a_20310_n5491.n3 0.764
R5733 a_20016_n6197.t0 a_20016_n6197.t1 380.209
R5734 a_20315_310.n1 a_20315_310.t5 318.922
R5735 a_20315_310.n0 a_20315_310.t6 274.739
R5736 a_20315_310.n0 a_20315_310.t4 274.739
R5737 a_20315_310.n1 a_20315_310.t7 269.116
R5738 a_20315_310.t5 a_20315_310.n0 179.946
R5739 a_20315_310.n2 a_20315_310.n1 105.178
R5740 a_20315_310.n3 a_20315_310.t2 29.444
R5741 a_20315_310.t3 a_20315_310.n4 28.565
R5742 a_20315_310.n4 a_20315_310.t1 28.565
R5743 a_20315_310.n2 a_20315_310.t0 18.145
R5744 a_20315_310.n3 a_20315_310.n2 2.878
R5745 a_20315_310.n4 a_20315_310.n3 0.764
R5746 a_20021_336.t0 a_20021_336.n0 14.282
R5747 a_20021_336.n0 a_20021_336.t2 14.282
R5748 a_20021_336.n0 a_20021_336.n13 90.416
R5749 a_20021_336.n13 a_20021_336.n12 50.575
R5750 a_20021_336.n13 a_20021_336.n9 74.302
R5751 a_20021_336.n12 a_20021_336.n11 157.665
R5752 a_20021_336.n11 a_20021_336.t6 8.7
R5753 a_20021_336.n11 a_20021_336.t7 8.7
R5754 a_20021_336.n12 a_20021_336.n10 122.999
R5755 a_20021_336.n10 a_20021_336.t5 14.282
R5756 a_20021_336.n10 a_20021_336.t1 14.282
R5757 a_20021_336.n9 a_20021_336.n8 90.436
R5758 a_20021_336.n8 a_20021_336.t3 14.282
R5759 a_20021_336.n8 a_20021_336.t4 14.282
R5760 a_20021_336.n1 a_20021_336.t18 217.826
R5761 a_20021_336.n9 a_20021_336.n1 277.579
R5762 a_20021_336.n1 a_20021_336.n6 133.839
R5763 a_20021_336.t18 a_20021_336.t9 437.233
R5764 a_20021_336.t9 a_20021_336.n7 214.686
R5765 a_20021_336.n7 a_20021_336.t8 80.333
R5766 a_20021_336.n7 a_20021_336.t19 214.686
R5767 a_20021_336.n6 a_20021_336.n2 563.136
R5768 a_20021_336.n6 a_20021_336.t15 178.973
R5769 a_20021_336.t15 a_20021_336.n5 80.333
R5770 a_20021_336.n5 a_20021_336.t16 190.152
R5771 a_20021_336.n5 a_20021_336.t14 190.152
R5772 a_20021_336.t14 a_20021_336.n4 313.873
R5773 a_20021_336.n4 a_20021_336.t17 160.666
R5774 a_20021_336.n4 a_20021_336.n3 96.129
R5775 a_20021_336.n3 a_20021_336.t12 160.666
R5776 a_20021_336.n3 a_20021_336.t11 272.288
R5777 a_20021_336.n2 a_20021_336.t13 294.986
R5778 a_20021_336.n2 a_20021_336.t10 110.859
R5779 a_7054_n416.t0 a_7054_n416.t1 17.4
R5780 a_10157_n6197.t5 a_10157_n6197.t4 574.43
R5781 a_10157_n6197.n0 a_10157_n6197.t7 285.109
R5782 a_10157_n6197.n2 a_10157_n6197.n1 197.217
R5783 a_10157_n6197.n4 a_10157_n6197.n3 192.754
R5784 a_10157_n6197.n0 a_10157_n6197.t6 160.666
R5785 a_10157_n6197.n1 a_10157_n6197.t5 160.666
R5786 a_10157_n6197.n1 a_10157_n6197.n0 114.829
R5787 a_10157_n6197.n3 a_10157_n6197.t1 28.568
R5788 a_10157_n6197.n4 a_10157_n6197.t2 28.565
R5789 a_10157_n6197.t3 a_10157_n6197.n4 28.565
R5790 a_10157_n6197.n2 a_10157_n6197.t0 18.838
R5791 a_10157_n6197.n3 a_10157_n6197.n2 1.129
R5792 a_11765_n2634.t7 a_11765_n2634.n3 404.877
R5793 a_11765_n2634.n2 a_11765_n2634.t8 210.902
R5794 a_11765_n2634.n4 a_11765_n2634.t7 136.943
R5795 a_11765_n2634.n3 a_11765_n2634.n2 107.801
R5796 a_11765_n2634.n2 a_11765_n2634.t6 80.333
R5797 a_11765_n2634.n3 a_11765_n2634.t5 80.333
R5798 a_11765_n2634.n1 a_11765_n2634.t4 17.4
R5799 a_11765_n2634.n1 a_11765_n2634.t1 17.4
R5800 a_11765_n2634.t0 a_11765_n2634.n5 15.032
R5801 a_11765_n2634.n0 a_11765_n2634.t2 14.282
R5802 a_11765_n2634.n0 a_11765_n2634.t3 14.282
R5803 a_11765_n2634.n5 a_11765_n2634.n0 1.65
R5804 a_11765_n2634.n4 a_11765_n2634.n1 0.672
R5805 a_11765_n2634.n5 a_11765_n2634.n4 0.665
R5806 Y[0].n1 Y[0].n0 192.754
R5807 Y[0].n1 Y[0].t2 28.568
R5808 Y[0].n0 Y[0].t3 28.565
R5809 Y[0].n0 Y[0].t1 28.565
R5810 Y[0].n2 Y[0].t0 19.164
R5811 Y[0] Y[0].n2 1.564
R5812 Y[0].n2 Y[0].n1 1.101
R5813 a_5214_290.n1 a_5214_290.t5 318.922
R5814 a_5214_290.n0 a_5214_290.t6 274.739
R5815 a_5214_290.n0 a_5214_290.t4 274.739
R5816 a_5214_290.n1 a_5214_290.t7 269.116
R5817 a_5214_290.t5 a_5214_290.n0 179.946
R5818 a_5214_290.n2 a_5214_290.n1 107.263
R5819 a_5214_290.n3 a_5214_290.t1 29.444
R5820 a_5214_290.t3 a_5214_290.n4 28.565
R5821 a_5214_290.n4 a_5214_290.t2 28.565
R5822 a_5214_290.n2 a_5214_290.t0 18.145
R5823 a_5214_290.n3 a_5214_290.n2 2.878
R5824 a_5214_290.n4 a_5214_290.n3 0.764
R5825 a_6620_n3211.n8 a_6620_n3211.n7 861.987
R5826 a_6620_n3211.n7 a_6620_n3211.n6 560.726
R5827 a_6620_n3211.t8 a_6620_n3211.t10 415.315
R5828 a_6620_n3211.t18 a_6620_n3211.t13 415.315
R5829 a_6620_n3211.n3 a_6620_n3211.t5 394.151
R5830 a_6620_n3211.n6 a_6620_n3211.t4 294.653
R5831 a_6620_n3211.n2 a_6620_n3211.t9 269.523
R5832 a_6620_n3211.t5 a_6620_n3211.n2 269.523
R5833 a_6620_n3211.n10 a_6620_n3211.t8 217.716
R5834 a_6620_n3211.n9 a_6620_n3211.t16 214.335
R5835 a_6620_n3211.t10 a_6620_n3211.n9 214.335
R5836 a_6620_n3211.n1 a_6620_n3211.t12 214.335
R5837 a_6620_n3211.t13 a_6620_n3211.n1 214.335
R5838 a_6620_n3211.n8 a_6620_n3211.t18 198.921
R5839 a_6620_n3211.n4 a_6620_n3211.t11 198.043
R5840 a_6620_n3211.n2 a_6620_n3211.t17 160.666
R5841 a_6620_n3211.n6 a_6620_n3211.t14 111.663
R5842 a_6620_n3211.n5 a_6620_n3211.n3 97.816
R5843 a_6620_n3211.n4 a_6620_n3211.t6 93.989
R5844 a_6620_n3211.n9 a_6620_n3211.t19 80.333
R5845 a_6620_n3211.n3 a_6620_n3211.t15 80.333
R5846 a_6620_n3211.n1 a_6620_n3211.t7 80.333
R5847 a_6620_n3211.n7 a_6620_n3211.n5 65.07
R5848 a_6620_n3211.n0 a_6620_n3211.t1 28.57
R5849 a_6620_n3211.t0 a_6620_n3211.n12 28.565
R5850 a_6620_n3211.n12 a_6620_n3211.t2 28.565
R5851 a_6620_n3211.n0 a_6620_n3211.t3 17.638
R5852 a_6620_n3211.n10 a_6620_n3211.n8 16.411
R5853 a_6620_n3211.n11 a_6620_n3211.n10 8.712
R5854 a_6620_n3211.n5 a_6620_n3211.n4 6.615
R5855 a_6620_n3211.n12 a_6620_n3211.n11 0.69
R5856 a_6620_n3211.n11 a_6620_n3211.n0 0.6
R5857 a_11705_n328.t0 a_11705_n328.t1 17.4
R5858 a_13361_n6198.t0 a_13361_n6198.t1 380.209
R5859 a_19567_3172.t6 a_19567_3172.n2 404.877
R5860 a_19567_3172.n1 a_19567_3172.t8 210.902
R5861 a_19567_3172.n3 a_19567_3172.t6 136.943
R5862 a_19567_3172.n2 a_19567_3172.n1 107.801
R5863 a_19567_3172.n1 a_19567_3172.t5 80.333
R5864 a_19567_3172.n2 a_19567_3172.t7 80.333
R5865 a_19567_3172.n0 a_19567_3172.t0 17.4
R5866 a_19567_3172.n0 a_19567_3172.t1 17.4
R5867 a_19567_3172.n4 a_19567_3172.t2 15.032
R5868 a_19567_3172.t4 a_19567_3172.n5 14.282
R5869 a_19567_3172.n5 a_19567_3172.t3 14.282
R5870 a_19567_3172.n5 a_19567_3172.n4 1.65
R5871 a_19567_3172.n3 a_19567_3172.n0 0.672
R5872 a_19567_3172.n4 a_19567_3172.n3 0.665
R5873 a_16167_n4181.n6 a_16167_n4181.n5 501.28
R5874 a_16167_n4181.t19 a_16167_n4181.t4 437.233
R5875 a_16167_n4181.t5 a_16167_n4181.t8 415.315
R5876 a_16167_n4181.t7 a_16167_n4181.n3 313.873
R5877 a_16167_n4181.n5 a_16167_n4181.t17 294.986
R5878 a_16167_n4181.n2 a_16167_n4181.t11 272.288
R5879 a_16167_n4181.n6 a_16167_n4181.t14 236.01
R5880 a_16167_n4181.n9 a_16167_n4181.t19 216.627
R5881 a_16167_n4181.n7 a_16167_n4181.t5 216.111
R5882 a_16167_n4181.n8 a_16167_n4181.t15 214.686
R5883 a_16167_n4181.t4 a_16167_n4181.n8 214.686
R5884 a_16167_n4181.n1 a_16167_n4181.t10 214.335
R5885 a_16167_n4181.t8 a_16167_n4181.n1 214.335
R5886 a_16167_n4181.n4 a_16167_n4181.t7 190.152
R5887 a_16167_n4181.n4 a_16167_n4181.t13 190.152
R5888 a_16167_n4181.n2 a_16167_n4181.t12 160.666
R5889 a_16167_n4181.n3 a_16167_n4181.t18 160.666
R5890 a_16167_n4181.n7 a_16167_n4181.n6 148.428
R5891 a_16167_n4181.n5 a_16167_n4181.t6 110.859
R5892 a_16167_n4181.n3 a_16167_n4181.n2 96.129
R5893 a_16167_n4181.n8 a_16167_n4181.t16 80.333
R5894 a_16167_n4181.n1 a_16167_n4181.t9 80.333
R5895 a_16167_n4181.t14 a_16167_n4181.n4 80.333
R5896 a_16167_n4181.n0 a_16167_n4181.t2 28.57
R5897 a_16167_n4181.n11 a_16167_n4181.t1 28.565
R5898 a_16167_n4181.t3 a_16167_n4181.n11 28.565
R5899 a_16167_n4181.n0 a_16167_n4181.t0 17.638
R5900 a_16167_n4181.n10 a_16167_n4181.n9 6.64
R5901 a_16167_n4181.n9 a_16167_n4181.n7 2.923
R5902 a_16167_n4181.n11 a_16167_n4181.n10 0.69
R5903 a_16167_n4181.n10 a_16167_n4181.n0 0.6
R5904 a_24195_n4771.n2 a_24195_n4771.t7 318.922
R5905 a_24195_n4771.n1 a_24195_n4771.t5 273.935
R5906 a_24195_n4771.n1 a_24195_n4771.t4 273.935
R5907 a_24195_n4771.n2 a_24195_n4771.t6 269.116
R5908 a_24195_n4771.n4 a_24195_n4771.n0 193.227
R5909 a_24195_n4771.t7 a_24195_n4771.n1 179.142
R5910 a_24195_n4771.n3 a_24195_n4771.n2 106.999
R5911 a_24195_n4771.t3 a_24195_n4771.n4 28.568
R5912 a_24195_n4771.n0 a_24195_n4771.t1 28.565
R5913 a_24195_n4771.n0 a_24195_n4771.t2 28.565
R5914 a_24195_n4771.n3 a_24195_n4771.t0 18.149
R5915 a_24195_n4771.n4 a_24195_n4771.n3 3.726
R5916 a_6265_n4771.n1 a_6265_n4771.t5 318.922
R5917 a_6265_n4771.n0 a_6265_n4771.t7 273.935
R5918 a_6265_n4771.n0 a_6265_n4771.t6 273.935
R5919 a_6265_n4771.n1 a_6265_n4771.t4 269.116
R5920 a_6265_n4771.n4 a_6265_n4771.n3 193.227
R5921 a_6265_n4771.t5 a_6265_n4771.n0 179.142
R5922 a_6265_n4771.n2 a_6265_n4771.n1 106.999
R5923 a_6265_n4771.n3 a_6265_n4771.t2 28.568
R5924 a_6265_n4771.t0 a_6265_n4771.n4 28.565
R5925 a_6265_n4771.n4 a_6265_n4771.t3 28.565
R5926 a_6265_n4771.n2 a_6265_n4771.t1 18.149
R5927 a_6265_n4771.n3 a_6265_n4771.n2 3.726
R5928 a_6810_n6196.t0 a_6810_n6196.t1 380.209
R5929 a_6810_n5464.t1 a_6810_n5464.n0 14.282
R5930 a_6810_n5464.n0 a_6810_n5464.t7 14.282
R5931 a_6810_n5464.n0 a_6810_n5464.n15 90.436
R5932 a_6810_n5464.n11 a_6810_n5464.n14 50.575
R5933 a_6810_n5464.n15 a_6810_n5464.n11 74.302
R5934 a_6810_n5464.n14 a_6810_n5464.n13 157.665
R5935 a_6810_n5464.n13 a_6810_n5464.t5 8.7
R5936 a_6810_n5464.n13 a_6810_n5464.t0 8.7
R5937 a_6810_n5464.n14 a_6810_n5464.n12 122.999
R5938 a_6810_n5464.n12 a_6810_n5464.t2 14.282
R5939 a_6810_n5464.n12 a_6810_n5464.t4 14.282
R5940 a_6810_n5464.n11 a_6810_n5464.n10 90.416
R5941 a_6810_n5464.n10 a_6810_n5464.t3 14.282
R5942 a_6810_n5464.n10 a_6810_n5464.t6 14.282
R5943 a_6810_n5464.n15 a_6810_n5464.n9 220.358
R5944 a_6810_n5464.n9 a_6810_n5464.n2 2.596
R5945 a_6810_n5464.n2 a_6810_n5464.t18 218.628
R5946 a_6810_n5464.t18 a_6810_n5464.t21 437.233
R5947 a_6810_n5464.t21 a_6810_n5464.n8 214.686
R5948 a_6810_n5464.n8 a_6810_n5464.t20 80.333
R5949 a_6810_n5464.n8 a_6810_n5464.t19 214.686
R5950 a_6810_n5464.n2 a_6810_n5464.n3 14.9
R5951 a_6810_n5464.n3 a_6810_n5464.n7 535.449
R5952 a_6810_n5464.n7 a_6810_n5464.t15 294.986
R5953 a_6810_n5464.n7 a_6810_n5464.t22 110.859
R5954 a_6810_n5464.n3 a_6810_n5464.t12 245.184
R5955 a_6810_n5464.t12 a_6810_n5464.n6 80.333
R5956 a_6810_n5464.n6 a_6810_n5464.t13 190.152
R5957 a_6810_n5464.n6 a_6810_n5464.t23 190.152
R5958 a_6810_n5464.t23 a_6810_n5464.n5 313.873
R5959 a_6810_n5464.n5 a_6810_n5464.t9 160.666
R5960 a_6810_n5464.n5 a_6810_n5464.n4 96.129
R5961 a_6810_n5464.n4 a_6810_n5464.t11 160.666
R5962 a_6810_n5464.n4 a_6810_n5464.t10 272.288
R5963 a_6810_n5464.n9 a_6810_n5464.t14 217.023
R5964 a_6810_n5464.t14 a_6810_n5464.t17 437.233
R5965 a_6810_n5464.t17 a_6810_n5464.n1 214.686
R5966 a_6810_n5464.n1 a_6810_n5464.t16 80.333
R5967 a_6810_n5464.n1 a_6810_n5464.t8 214.686
R5968 a_9518_1688.n6 a_9518_1688.n5 501.28
R5969 a_9518_1688.t4 a_9518_1688.t18 437.233
R5970 a_9518_1688.t15 a_9518_1688.t13 415.315
R5971 a_9518_1688.t10 a_9518_1688.n3 313.873
R5972 a_9518_1688.n5 a_9518_1688.t8 294.986
R5973 a_9518_1688.n2 a_9518_1688.t7 272.288
R5974 a_9518_1688.n6 a_9518_1688.t16 236.01
R5975 a_9518_1688.n9 a_9518_1688.t4 216.627
R5976 a_9518_1688.n7 a_9518_1688.t15 216.111
R5977 a_9518_1688.n8 a_9518_1688.t12 214.686
R5978 a_9518_1688.t18 a_9518_1688.n8 214.686
R5979 a_9518_1688.n1 a_9518_1688.t5 214.335
R5980 a_9518_1688.t13 a_9518_1688.n1 214.335
R5981 a_9518_1688.n4 a_9518_1688.t10 190.152
R5982 a_9518_1688.n4 a_9518_1688.t11 190.152
R5983 a_9518_1688.n2 a_9518_1688.t19 160.666
R5984 a_9518_1688.n3 a_9518_1688.t14 160.666
R5985 a_9518_1688.n7 a_9518_1688.n6 148.428
R5986 a_9518_1688.n5 a_9518_1688.t17 110.859
R5987 a_9518_1688.n3 a_9518_1688.n2 96.129
R5988 a_9518_1688.n8 a_9518_1688.t6 80.333
R5989 a_9518_1688.n1 a_9518_1688.t9 80.333
R5990 a_9518_1688.t16 a_9518_1688.n4 80.333
R5991 a_9518_1688.t3 a_9518_1688.n11 28.57
R5992 a_9518_1688.n0 a_9518_1688.t1 28.565
R5993 a_9518_1688.n0 a_9518_1688.t2 28.565
R5994 a_9518_1688.n11 a_9518_1688.t0 17.638
R5995 a_9518_1688.n10 a_9518_1688.n9 12.318
R5996 a_9518_1688.n9 a_9518_1688.n7 2.923
R5997 a_9518_1688.n10 a_9518_1688.n0 0.69
R5998 a_9518_1688.n11 a_9518_1688.n10 0.6
R5999 a_688_n2757.n5 a_688_n2757.n4 535.449
R6000 a_688_n2757.t11 a_688_n2757.t13 437.233
R6001 a_688_n2757.t14 a_688_n2757.t18 437.233
R6002 a_688_n2757.t7 a_688_n2757.n2 313.873
R6003 a_688_n2757.n4 a_688_n2757.t16 294.986
R6004 a_688_n2757.n1 a_688_n2757.t4 272.288
R6005 a_688_n2757.n5 a_688_n2757.t8 245.184
R6006 a_688_n2757.n7 a_688_n2757.t14 218.628
R6007 a_688_n2757.n9 a_688_n2757.t11 217.026
R6008 a_688_n2757.n8 a_688_n2757.t15 214.686
R6009 a_688_n2757.t13 a_688_n2757.n8 214.686
R6010 a_688_n2757.n6 a_688_n2757.t19 214.686
R6011 a_688_n2757.t18 a_688_n2757.n6 214.686
R6012 a_688_n2757.n11 a_688_n2757.n0 192.754
R6013 a_688_n2757.n3 a_688_n2757.t7 190.152
R6014 a_688_n2757.n3 a_688_n2757.t9 190.152
R6015 a_688_n2757.n1 a_688_n2757.t5 160.666
R6016 a_688_n2757.n2 a_688_n2757.t10 160.666
R6017 a_688_n2757.n4 a_688_n2757.t6 110.859
R6018 a_688_n2757.n2 a_688_n2757.n1 96.129
R6019 a_688_n2757.n8 a_688_n2757.t12 80.333
R6020 a_688_n2757.t8 a_688_n2757.n3 80.333
R6021 a_688_n2757.n6 a_688_n2757.t17 80.333
R6022 a_688_n2757.t0 a_688_n2757.n11 28.568
R6023 a_688_n2757.n0 a_688_n2757.t1 28.565
R6024 a_688_n2757.n0 a_688_n2757.t3 28.565
R6025 a_688_n2757.n10 a_688_n2757.t2 18.722
R6026 a_688_n2757.n7 a_688_n2757.n5 14.9
R6027 a_688_n2757.n9 a_688_n2757.n7 2.603
R6028 a_688_n2757.n10 a_688_n2757.n9 2.382
R6029 a_688_n2757.n11 a_688_n2757.n10 1.281
R6030 a_19476_1029.n1 a_19476_1029.t5 318.922
R6031 a_19476_1029.n0 a_19476_1029.t6 273.935
R6032 a_19476_1029.n0 a_19476_1029.t4 273.935
R6033 a_19476_1029.n1 a_19476_1029.t7 269.116
R6034 a_19476_1029.n4 a_19476_1029.n3 193.227
R6035 a_19476_1029.t5 a_19476_1029.n0 179.142
R6036 a_19476_1029.n2 a_19476_1029.n1 106.999
R6037 a_19476_1029.n3 a_19476_1029.t2 28.568
R6038 a_19476_1029.n4 a_19476_1029.t1 28.565
R6039 a_19476_1029.t3 a_19476_1029.n4 28.565
R6040 a_19476_1029.n2 a_19476_1029.t0 18.149
R6041 a_19476_1029.n3 a_19476_1029.n2 3.726
R6042 a_3611_n4591.t4 a_3611_n4591.t7 574.43
R6043 a_3611_n4591.n0 a_3611_n4591.t6 285.109
R6044 a_3611_n4591.n2 a_3611_n4591.n1 211.136
R6045 a_3611_n4591.n4 a_3611_n4591.n3 192.754
R6046 a_3611_n4591.n0 a_3611_n4591.t5 160.666
R6047 a_3611_n4591.n1 a_3611_n4591.t4 160.666
R6048 a_3611_n4591.n1 a_3611_n4591.n0 114.829
R6049 a_3611_n4591.n3 a_3611_n4591.t3 28.568
R6050 a_3611_n4591.n4 a_3611_n4591.t2 28.565
R6051 a_3611_n4591.t1 a_3611_n4591.n4 28.565
R6052 a_3611_n4591.n2 a_3611_n4591.t0 19.084
R6053 a_3611_n4591.n3 a_3611_n4591.n2 1.051
R6054 a_6356_n2628.t5 a_6356_n2628.n2 404.877
R6055 a_6356_n2628.n1 a_6356_n2628.t8 210.902
R6056 a_6356_n2628.n3 a_6356_n2628.t5 136.943
R6057 a_6356_n2628.n2 a_6356_n2628.n1 107.801
R6058 a_6356_n2628.n1 a_6356_n2628.t7 80.333
R6059 a_6356_n2628.n2 a_6356_n2628.t6 80.333
R6060 a_6356_n2628.n0 a_6356_n2628.t4 17.4
R6061 a_6356_n2628.n0 a_6356_n2628.t2 17.4
R6062 a_6356_n2628.n4 a_6356_n2628.t3 15.032
R6063 a_6356_n2628.n5 a_6356_n2628.t1 14.282
R6064 a_6356_n2628.t0 a_6356_n2628.n5 14.282
R6065 a_6356_n2628.n5 a_6356_n2628.n4 1.65
R6066 a_6356_n2628.n3 a_6356_n2628.n0 0.672
R6067 a_6356_n2628.n4 a_6356_n2628.n3 0.665
R6068 a_6474_n2628.n1 a_6474_n2628.t5 14.282
R6069 a_6474_n2628.n1 a_6474_n2628.t0 14.282
R6070 a_6474_n2628.n0 a_6474_n2628.t1 14.282
R6071 a_6474_n2628.n0 a_6474_n2628.t2 14.282
R6072 a_6474_n2628.n3 a_6474_n2628.t4 14.282
R6073 a_6474_n2628.t3 a_6474_n2628.n3 14.282
R6074 a_6474_n2628.n2 a_6474_n2628.n0 2.546
R6075 a_6474_n2628.n3 a_6474_n2628.n2 2.367
R6076 a_6474_n2628.n2 a_6474_n2628.n1 0.001
R6077 a_3606_n6195.t4 a_3606_n6195.t7 574.43
R6078 a_3606_n6195.n0 a_3606_n6195.t6 285.109
R6079 a_3606_n6195.n2 a_3606_n6195.n1 197.217
R6080 a_3606_n6195.n4 a_3606_n6195.n3 192.754
R6081 a_3606_n6195.n0 a_3606_n6195.t5 160.666
R6082 a_3606_n6195.n1 a_3606_n6195.t4 160.666
R6083 a_3606_n6195.n1 a_3606_n6195.n0 114.829
R6084 a_3606_n6195.n3 a_3606_n6195.t2 28.568
R6085 a_3606_n6195.n4 a_3606_n6195.t1 28.565
R6086 a_3606_n6195.t0 a_3606_n6195.n4 28.565
R6087 a_3606_n6195.n2 a_3606_n6195.t3 18.838
R6088 a_3606_n6195.n3 a_3606_n6195.n2 1.129
R6089 a_5214_n2632.t6 a_5214_n2632.n3 404.877
R6090 a_5214_n2632.n2 a_5214_n2632.t8 210.902
R6091 a_5214_n2632.n4 a_5214_n2632.t6 136.943
R6092 a_5214_n2632.n3 a_5214_n2632.n2 107.801
R6093 a_5214_n2632.n2 a_5214_n2632.t7 80.333
R6094 a_5214_n2632.n3 a_5214_n2632.t5 80.333
R6095 a_5214_n2632.n1 a_5214_n2632.t4 17.4
R6096 a_5214_n2632.n1 a_5214_n2632.t0 17.4
R6097 a_5214_n2632.t1 a_5214_n2632.n5 15.032
R6098 a_5214_n2632.n0 a_5214_n2632.t2 14.282
R6099 a_5214_n2632.n0 a_5214_n2632.t3 14.282
R6100 a_5214_n2632.n5 a_5214_n2632.n0 1.65
R6101 a_5214_n2632.n4 a_5214_n2632.n1 0.672
R6102 a_5214_n2632.n5 a_5214_n2632.n4 0.665
R6103 a_5332_n2632.n1 a_5332_n2632.t5 14.282
R6104 a_5332_n2632.n1 a_5332_n2632.t0 14.282
R6105 a_5332_n2632.n0 a_5332_n2632.t1 14.282
R6106 a_5332_n2632.n0 a_5332_n2632.t2 14.282
R6107 a_5332_n2632.t3 a_5332_n2632.n3 14.282
R6108 a_5332_n2632.n3 a_5332_n2632.t4 14.282
R6109 a_5332_n2632.n2 a_5332_n2632.n0 2.546
R6110 a_5332_n2632.n3 a_5332_n2632.n2 2.367
R6111 a_5332_n2632.n2 a_5332_n2632.n1 0.001
R6112 a_25034_n5490.n1 a_25034_n5490.t5 318.922
R6113 a_25034_n5490.n0 a_25034_n5490.t4 274.739
R6114 a_25034_n5490.n0 a_25034_n5490.t6 274.739
R6115 a_25034_n5490.n1 a_25034_n5490.t7 269.116
R6116 a_25034_n5490.t5 a_25034_n5490.n0 179.946
R6117 a_25034_n5490.n2 a_25034_n5490.n1 107.263
R6118 a_25034_n5490.n3 a_25034_n5490.t1 29.444
R6119 a_25034_n5490.n4 a_25034_n5490.t2 28.565
R6120 a_25034_n5490.t3 a_25034_n5490.n4 28.565
R6121 a_25034_n5490.n2 a_25034_n5490.t0 18.145
R6122 a_25034_n5490.n3 a_25034_n5490.n2 2.878
R6123 a_25034_n5490.n4 a_25034_n5490.n3 0.764
R6124 a_24622_n5464.n2 a_24622_n5464.n0 267.767
R6125 a_24622_n5464.n6 a_24622_n5464.t7 16.058
R6126 a_24622_n5464.n8 a_24622_n5464.t0 16.058
R6127 a_24622_n5464.n1 a_24622_n5464.t5 14.282
R6128 a_24622_n5464.n1 a_24622_n5464.t9 14.282
R6129 a_24622_n5464.n0 a_24622_n5464.t3 14.282
R6130 a_24622_n5464.n0 a_24622_n5464.t4 14.282
R6131 a_24622_n5464.n3 a_24622_n5464.t10 14.282
R6132 a_24622_n5464.n3 a_24622_n5464.t11 14.282
R6133 a_24622_n5464.n5 a_24622_n5464.t8 14.282
R6134 a_24622_n5464.n5 a_24622_n5464.t6 14.282
R6135 a_24622_n5464.n9 a_24622_n5464.t1 14.282
R6136 a_24622_n5464.t2 a_24622_n5464.n9 14.282
R6137 a_24622_n5464.n4 a_24622_n5464.n3 1.511
R6138 a_24622_n5464.n6 a_24622_n5464.n5 0.999
R6139 a_24622_n5464.n9 a_24622_n5464.n8 0.999
R6140 a_24622_n5464.n4 a_24622_n5464.n2 0.669
R6141 a_24622_n5464.n7 a_24622_n5464.n6 0.575
R6142 a_24622_n5464.n7 a_24622_n5464.n4 0.227
R6143 a_24622_n5464.n8 a_24622_n5464.n7 0.2
R6144 a_24622_n5464.n2 a_24622_n5464.n1 0.001
R6145 a_11889_3236.n1 a_11889_3236.t5 14.282
R6146 a_11889_3236.n1 a_11889_3236.t1 14.282
R6147 a_11889_3236.n0 a_11889_3236.t2 14.282
R6148 a_11889_3236.n0 a_11889_3236.t0 14.282
R6149 a_11889_3236.n3 a_11889_3236.t4 14.282
R6150 a_11889_3236.t3 a_11889_3236.n3 14.282
R6151 a_11889_3236.n2 a_11889_3236.n0 2.546
R6152 a_11889_3236.n3 a_11889_3236.n2 2.367
R6153 a_11889_3236.n2 a_11889_3236.n1 0.001
R6154 a_28708_n5298.n4 a_28708_n5298.t10 214.335
R6155 a_28708_n5298.t8 a_28708_n5298.n4 214.335
R6156 a_28708_n5298.n5 a_28708_n5298.t8 143.851
R6157 a_28708_n5298.n5 a_28708_n5298.t7 135.658
R6158 a_28708_n5298.n4 a_28708_n5298.t9 80.333
R6159 a_28708_n5298.n0 a_28708_n5298.t1 28.565
R6160 a_28708_n5298.n0 a_28708_n5298.t2 28.565
R6161 a_28708_n5298.n2 a_28708_n5298.t5 28.565
R6162 a_28708_n5298.n2 a_28708_n5298.t0 28.565
R6163 a_28708_n5298.n7 a_28708_n5298.t6 28.565
R6164 a_28708_n5298.t4 a_28708_n5298.n7 28.565
R6165 a_28708_n5298.n1 a_28708_n5298.t3 9.714
R6166 a_28708_n5298.n1 a_28708_n5298.n0 1.003
R6167 a_28708_n5298.n6 a_28708_n5298.n3 0.833
R6168 a_28708_n5298.n3 a_28708_n5298.n2 0.653
R6169 a_28708_n5298.n7 a_28708_n5298.n6 0.653
R6170 a_28708_n5298.n3 a_28708_n5298.n1 0.341
R6171 a_28708_n5298.n6 a_28708_n5298.n5 0.032
R6172 a_10148_n2943.t5 a_10148_n2943.t4 800.071
R6173 a_10148_n2943.n2 a_10148_n2943.n1 659.097
R6174 a_10148_n2943.n0 a_10148_n2943.t7 285.109
R6175 a_10148_n2943.n1 a_10148_n2943.t5 193.602
R6176 a_10148_n2943.n4 a_10148_n2943.n3 192.754
R6177 a_10148_n2943.n0 a_10148_n2943.t6 160.666
R6178 a_10148_n2943.n1 a_10148_n2943.n0 91.507
R6179 a_10148_n2943.n3 a_10148_n2943.t1 28.568
R6180 a_10148_n2943.t0 a_10148_n2943.n4 28.565
R6181 a_10148_n2943.n4 a_10148_n2943.t2 28.565
R6182 a_10148_n2943.n2 a_10148_n2943.t3 19.061
R6183 a_10148_n2943.n3 a_10148_n2943.n2 1.005
R6184 a_13597_n6198.t0 a_13597_n6198.t1 17.4
R6185 a_4912_n5464.n0 a_4912_n5464.t4 14.282
R6186 a_4912_n5464.t0 a_4912_n5464.n0 14.282
R6187 a_4912_n5464.n0 a_4912_n5464.n12 90.416
R6188 a_4912_n5464.n12 a_4912_n5464.n11 50.575
R6189 a_4912_n5464.n12 a_4912_n5464.n8 74.302
R6190 a_4912_n5464.n11 a_4912_n5464.n10 157.665
R6191 a_4912_n5464.n10 a_4912_n5464.t1 8.7
R6192 a_4912_n5464.n10 a_4912_n5464.t5 8.7
R6193 a_4912_n5464.n11 a_4912_n5464.n9 122.999
R6194 a_4912_n5464.n9 a_4912_n5464.t2 14.282
R6195 a_4912_n5464.n9 a_4912_n5464.t3 14.282
R6196 a_4912_n5464.n8 a_4912_n5464.n7 90.436
R6197 a_4912_n5464.n7 a_4912_n5464.t6 14.282
R6198 a_4912_n5464.n7 a_4912_n5464.t7 14.282
R6199 a_4912_n5464.n8 a_4912_n5464.n1 342.688
R6200 a_4912_n5464.n1 a_4912_n5464.n6 126.566
R6201 a_4912_n5464.n6 a_4912_n5464.t8 294.653
R6202 a_4912_n5464.n6 a_4912_n5464.t10 111.663
R6203 a_4912_n5464.n1 a_4912_n5464.n5 552.333
R6204 a_4912_n5464.n5 a_4912_n5464.n4 6.615
R6205 a_4912_n5464.n4 a_4912_n5464.t15 93.989
R6206 a_4912_n5464.n5 a_4912_n5464.n3 97.816
R6207 a_4912_n5464.n3 a_4912_n5464.t9 80.333
R6208 a_4912_n5464.n3 a_4912_n5464.t12 394.151
R6209 a_4912_n5464.t12 a_4912_n5464.n2 269.523
R6210 a_4912_n5464.n2 a_4912_n5464.t13 160.666
R6211 a_4912_n5464.n2 a_4912_n5464.t11 269.523
R6212 a_4912_n5464.n4 a_4912_n5464.t14 198.043
R6213 a_7046_n6196.t0 a_7046_n6196.t1 17.4
R6214 A[2].n6 A[2].t1 3756.03
R6215 A[2].t10 A[2].t14 437.233
R6216 A[2].t1 A[2].t2 437.233
R6217 A[2].t8 A[2].t12 415.315
R6218 A[2].t7 A[2].t15 415.315
R6219 A[2].n5 A[2].t7 256.298
R6220 A[2].n3 A[2].t10 219.994
R6221 A[2].n3 A[2].t8 217.552
R6222 A[2].n1 A[2].t5 214.686
R6223 A[2].t14 A[2].n1 214.686
R6224 A[2].n0 A[2].t0 214.686
R6225 A[2].t2 A[2].n0 214.686
R6226 A[2].n2 A[2].t6 214.335
R6227 A[2].t12 A[2].n2 214.335
R6228 A[2].n4 A[2].t4 214.335
R6229 A[2].t15 A[2].n4 214.335
R6230 A[2].n2 A[2].t9 80.333
R6231 A[2].n1 A[2].t13 80.333
R6232 A[2].n4 A[2].t3 80.333
R6233 A[2].n0 A[2].t11 80.333
R6234 A[2].n5 A[2].n3 0.426
R6235 A[2] A[2].n6 0.373
R6236 A[2].n6 A[2].n5 0.09
R6237 a_16817_n4592.t4 a_16817_n4592.t5 574.43
R6238 a_16817_n4592.n0 a_16817_n4592.t7 285.109
R6239 a_16817_n4592.n2 a_16817_n4592.n1 211.136
R6240 a_16817_n4592.n4 a_16817_n4592.n3 192.754
R6241 a_16817_n4592.n0 a_16817_n4592.t6 160.666
R6242 a_16817_n4592.n1 a_16817_n4592.t4 160.666
R6243 a_16817_n4592.n1 a_16817_n4592.n0 114.829
R6244 a_16817_n4592.n3 a_16817_n4592.t3 28.568
R6245 a_16817_n4592.n4 a_16817_n4592.t2 28.565
R6246 a_16817_n4592.t1 a_16817_n4592.n4 28.565
R6247 a_16817_n4592.n2 a_16817_n4592.t0 19.084
R6248 a_16817_n4592.n3 a_16817_n4592.n2 1.051
R6249 a_19680_n2629.n1 a_19680_n2629.t2 14.282
R6250 a_19680_n2629.n1 a_19680_n2629.t3 14.282
R6251 a_19680_n2629.n0 a_19680_n2629.t4 14.282
R6252 a_19680_n2629.n0 a_19680_n2629.t5 14.282
R6253 a_19680_n2629.n3 a_19680_n2629.t1 14.282
R6254 a_19680_n2629.t0 a_19680_n2629.n3 14.282
R6255 a_19680_n2629.n2 a_19680_n2629.n0 2.546
R6256 a_19680_n2629.n3 a_19680_n2629.n2 2.367
R6257 a_19680_n2629.n2 a_19680_n2629.n1 0.001
R6258 a_3016_n5758.n0 a_3016_n5758.t10 214.335
R6259 a_3016_n5758.t8 a_3016_n5758.n0 214.335
R6260 a_3016_n5758.n1 a_3016_n5758.t8 143.851
R6261 a_3016_n5758.n1 a_3016_n5758.t7 135.658
R6262 a_3016_n5758.n0 a_3016_n5758.t9 80.333
R6263 a_3016_n5758.n2 a_3016_n5758.t4 28.565
R6264 a_3016_n5758.n2 a_3016_n5758.t5 28.565
R6265 a_3016_n5758.n4 a_3016_n5758.t6 28.565
R6266 a_3016_n5758.n4 a_3016_n5758.t2 28.565
R6267 a_3016_n5758.t3 a_3016_n5758.n7 28.565
R6268 a_3016_n5758.n7 a_3016_n5758.t1 28.565
R6269 a_3016_n5758.n6 a_3016_n5758.t0 9.714
R6270 a_3016_n5758.n7 a_3016_n5758.n6 1.003
R6271 a_3016_n5758.n5 a_3016_n5758.n3 0.833
R6272 a_3016_n5758.n3 a_3016_n5758.n2 0.653
R6273 a_3016_n5758.n5 a_3016_n5758.n4 0.653
R6274 a_3016_n5758.n6 a_3016_n5758.n5 0.341
R6275 a_3016_n5758.n3 a_3016_n5758.n1 0.032
R6276 a_5222_3148.t8 a_5222_3148.n2 404.877
R6277 a_5222_3148.n1 a_5222_3148.t5 210.902
R6278 a_5222_3148.n3 a_5222_3148.t8 136.943
R6279 a_5222_3148.n2 a_5222_3148.n1 107.801
R6280 a_5222_3148.n1 a_5222_3148.t6 80.333
R6281 a_5222_3148.n2 a_5222_3148.t7 80.333
R6282 a_5222_3148.n0 a_5222_3148.t0 17.4
R6283 a_5222_3148.n0 a_5222_3148.t1 17.4
R6284 a_5222_3148.n4 a_5222_3148.t4 15.032
R6285 a_5222_3148.t2 a_5222_3148.n5 14.282
R6286 a_5222_3148.n5 a_5222_3148.t3 14.282
R6287 a_5222_3148.n5 a_5222_3148.n4 1.65
R6288 a_5222_3148.n3 a_5222_3148.n0 0.672
R6289 a_5222_3148.n4 a_5222_3148.n3 0.665
R6290 a_18118_n5465.n0 a_18118_n5465.n12 122.999
R6291 a_18118_n5465.t1 a_18118_n5465.n0 14.282
R6292 a_18118_n5465.n0 a_18118_n5465.t4 14.282
R6293 a_18118_n5465.n12 a_18118_n5465.n10 50.575
R6294 a_18118_n5465.n10 a_18118_n5465.n8 74.302
R6295 a_18118_n5465.n12 a_18118_n5465.n11 157.665
R6296 a_18118_n5465.n11 a_18118_n5465.t2 8.7
R6297 a_18118_n5465.n11 a_18118_n5465.t0 8.7
R6298 a_18118_n5465.n10 a_18118_n5465.n9 90.416
R6299 a_18118_n5465.n9 a_18118_n5465.t3 14.282
R6300 a_18118_n5465.n9 a_18118_n5465.t6 14.282
R6301 a_18118_n5465.n8 a_18118_n5465.n7 90.436
R6302 a_18118_n5465.n7 a_18118_n5465.t5 14.282
R6303 a_18118_n5465.n7 a_18118_n5465.t7 14.282
R6304 a_18118_n5465.n8 a_18118_n5465.n1 342.688
R6305 a_18118_n5465.n1 a_18118_n5465.n6 126.566
R6306 a_18118_n5465.n6 a_18118_n5465.t14 294.653
R6307 a_18118_n5465.n6 a_18118_n5465.t15 111.663
R6308 a_18118_n5465.n1 a_18118_n5465.n5 552.333
R6309 a_18118_n5465.n5 a_18118_n5465.n4 6.615
R6310 a_18118_n5465.n4 a_18118_n5465.t11 93.989
R6311 a_18118_n5465.n5 a_18118_n5465.n3 97.816
R6312 a_18118_n5465.n3 a_18118_n5465.t12 80.333
R6313 a_18118_n5465.n3 a_18118_n5465.t8 394.151
R6314 a_18118_n5465.t8 a_18118_n5465.n2 269.523
R6315 a_18118_n5465.n2 a_18118_n5465.t9 160.666
R6316 a_18118_n5465.n2 a_18118_n5465.t13 269.523
R6317 a_18118_n5465.n4 a_18118_n5465.t10 198.043
R6318 a_19898_n5465.n0 a_19898_n5465.t1 14.282
R6319 a_19898_n5465.t0 a_19898_n5465.n0 14.282
R6320 a_19898_n5465.n0 a_19898_n5465.n9 0.999
R6321 a_19898_n5465.n9 a_19898_n5465.n6 0.575
R6322 a_19898_n5465.n6 a_19898_n5465.n8 0.2
R6323 a_19898_n5465.n8 a_19898_n5465.t10 16.058
R6324 a_19898_n5465.n8 a_19898_n5465.n7 0.999
R6325 a_19898_n5465.n7 a_19898_n5465.t9 14.282
R6326 a_19898_n5465.n7 a_19898_n5465.t11 14.282
R6327 a_19898_n5465.n9 a_19898_n5465.t8 16.058
R6328 a_19898_n5465.n6 a_19898_n5465.n4 0.227
R6329 a_19898_n5465.n4 a_19898_n5465.n5 1.511
R6330 a_19898_n5465.n5 a_19898_n5465.t4 14.282
R6331 a_19898_n5465.n5 a_19898_n5465.t3 14.282
R6332 a_19898_n5465.n4 a_19898_n5465.n1 0.669
R6333 a_19898_n5465.n1 a_19898_n5465.n2 0.001
R6334 a_19898_n5465.n1 a_19898_n5465.n3 267.767
R6335 a_19898_n5465.n3 a_19898_n5465.t6 14.282
R6336 a_19898_n5465.n3 a_19898_n5465.t5 14.282
R6337 a_19898_n5465.n2 a_19898_n5465.t2 14.282
R6338 a_19898_n5465.n2 a_19898_n5465.t7 14.282
R6339 a_30335_4891.n1 a_30335_4891.t4 318.922
R6340 a_30335_4891.n0 a_30335_4891.t7 273.935
R6341 a_30335_4891.n0 a_30335_4891.t5 273.935
R6342 a_30335_4891.n1 a_30335_4891.t6 269.116
R6343 a_30335_4891.n4 a_30335_4891.n3 193.227
R6344 a_30335_4891.t4 a_30335_4891.n0 179.142
R6345 a_30335_4891.n2 a_30335_4891.n1 106.999
R6346 a_30335_4891.n3 a_30335_4891.t1 28.568
R6347 a_30335_4891.n4 a_30335_4891.t2 28.565
R6348 a_30335_4891.t3 a_30335_4891.n4 28.565
R6349 a_30335_4891.n2 a_30335_4891.t0 18.149
R6350 a_30335_4891.n3 a_30335_4891.n2 3.726
R6351 a_18684_n3216.t5 a_18684_n3216.t6 800.071
R6352 a_18684_n3216.n3 a_18684_n3216.n2 672.951
R6353 a_18684_n3216.n1 a_18684_n3216.t4 285.109
R6354 a_18684_n3216.n2 a_18684_n3216.t5 193.602
R6355 a_18684_n3216.n1 a_18684_n3216.t7 160.666
R6356 a_18684_n3216.n2 a_18684_n3216.n1 91.507
R6357 a_18684_n3216.t0 a_18684_n3216.n4 28.57
R6358 a_18684_n3216.n0 a_18684_n3216.t3 28.565
R6359 a_18684_n3216.n0 a_18684_n3216.t2 28.565
R6360 a_18684_n3216.n4 a_18684_n3216.t1 17.638
R6361 a_18684_n3216.n3 a_18684_n3216.n0 0.69
R6362 a_18684_n3216.n4 a_18684_n3216.n3 0.6
R6363 a_29298_n5735.n5 a_29298_n5735.n4 465.933
R6364 a_29298_n5735.t15 a_29298_n5735.t6 415.315
R6365 a_29298_n5735.n1 a_29298_n5735.t4 394.151
R6366 a_29298_n5735.n4 a_29298_n5735.t10 294.653
R6367 a_29298_n5735.n0 a_29298_n5735.t9 269.523
R6368 a_29298_n5735.t4 a_29298_n5735.n0 269.523
R6369 a_29298_n5735.n7 a_29298_n5735.t15 220.285
R6370 a_29298_n5735.n6 a_29298_n5735.t11 214.335
R6371 a_29298_n5735.t6 a_29298_n5735.n6 214.335
R6372 a_29298_n5735.n2 a_29298_n5735.t8 198.043
R6373 a_29298_n5735.n10 a_29298_n5735.n9 192.754
R6374 a_29298_n5735.n5 a_29298_n5735.n3 163.88
R6375 a_29298_n5735.n0 a_29298_n5735.t5 160.666
R6376 a_29298_n5735.n4 a_29298_n5735.t14 111.663
R6377 a_29298_n5735.n3 a_29298_n5735.n1 97.816
R6378 a_29298_n5735.n2 a_29298_n5735.t12 93.989
R6379 a_29298_n5735.n6 a_29298_n5735.t7 80.333
R6380 a_29298_n5735.n1 a_29298_n5735.t13 80.333
R6381 a_29298_n5735.n7 a_29298_n5735.n5 61.538
R6382 a_29298_n5735.n9 a_29298_n5735.t1 28.568
R6383 a_29298_n5735.n10 a_29298_n5735.t2 28.565
R6384 a_29298_n5735.t3 a_29298_n5735.n10 28.565
R6385 a_29298_n5735.n8 a_29298_n5735.t0 18.824
R6386 a_29298_n5735.n3 a_29298_n5735.n2 6.615
R6387 a_29298_n5735.n8 a_29298_n5735.n7 4.769
R6388 a_29298_n5735.n9 a_29298_n5735.n8 1.105
R6389 a_30764_n3388.t0 a_30764_n3388.n0 14.282
R6390 a_30764_n3388.n0 a_30764_n3388.t8 14.282
R6391 a_30764_n3388.n0 a_30764_n3388.n9 0.999
R6392 a_30764_n3388.n6 a_30764_n3388.n8 0.575
R6393 a_30764_n3388.n9 a_30764_n3388.n6 0.2
R6394 a_30764_n3388.n9 a_30764_n3388.t1 16.058
R6395 a_30764_n3388.n8 a_30764_n3388.n7 0.999
R6396 a_30764_n3388.n7 a_30764_n3388.t4 14.282
R6397 a_30764_n3388.n7 a_30764_n3388.t2 14.282
R6398 a_30764_n3388.n8 a_30764_n3388.t3 16.058
R6399 a_30764_n3388.n6 a_30764_n3388.n4 0.227
R6400 a_30764_n3388.n4 a_30764_n3388.n5 1.511
R6401 a_30764_n3388.n5 a_30764_n3388.t11 14.282
R6402 a_30764_n3388.n5 a_30764_n3388.t10 14.282
R6403 a_30764_n3388.n4 a_30764_n3388.n1 0.669
R6404 a_30764_n3388.n1 a_30764_n3388.n2 0.001
R6405 a_30764_n3388.n1 a_30764_n3388.n3 267.767
R6406 a_30764_n3388.n3 a_30764_n3388.t6 14.282
R6407 a_30764_n3388.n3 a_30764_n3388.t5 14.282
R6408 a_30764_n3388.n2 a_30764_n3388.t9 14.282
R6409 a_30764_n3388.n2 a_30764_n3388.t7 14.282
R6410 a_30764_n7736.n2 a_30764_n7736.n0 267.767
R6411 a_30764_n7736.n6 a_30764_n7736.t11 16.058
R6412 a_30764_n7736.n4 a_30764_n7736.t3 16.058
R6413 a_30764_n7736.n5 a_30764_n7736.t9 14.282
R6414 a_30764_n7736.n5 a_30764_n7736.t10 14.282
R6415 a_30764_n7736.n3 a_30764_n7736.t4 14.282
R6416 a_30764_n7736.n3 a_30764_n7736.t5 14.282
R6417 a_30764_n7736.n1 a_30764_n7736.t7 14.282
R6418 a_30764_n7736.n1 a_30764_n7736.t0 14.282
R6419 a_30764_n7736.n0 a_30764_n7736.t8 14.282
R6420 a_30764_n7736.n0 a_30764_n7736.t6 14.282
R6421 a_30764_n7736.n9 a_30764_n7736.t1 14.282
R6422 a_30764_n7736.t2 a_30764_n7736.n9 14.282
R6423 a_30764_n7736.n9 a_30764_n7736.n8 1.511
R6424 a_30764_n7736.n6 a_30764_n7736.n5 0.999
R6425 a_30764_n7736.n4 a_30764_n7736.n3 0.999
R6426 a_30764_n7736.n8 a_30764_n7736.n2 0.669
R6427 a_30764_n7736.n7 a_30764_n7736.n6 0.575
R6428 a_30764_n7736.n8 a_30764_n7736.n7 0.227
R6429 a_30764_n7736.n7 a_30764_n7736.n4 0.2
R6430 a_30764_n7736.n2 a_30764_n7736.n1 0.001
R6431 a_4802_316.n8 a_4802_316.n0 267.767
R6432 a_4802_316.n4 a_4802_316.t9 16.058
R6433 a_4802_316.n2 a_4802_316.t8 16.058
R6434 a_4802_316.n3 a_4802_316.t11 14.282
R6435 a_4802_316.n3 a_4802_316.t10 14.282
R6436 a_4802_316.n1 a_4802_316.t7 14.282
R6437 a_4802_316.n1 a_4802_316.t6 14.282
R6438 a_4802_316.n6 a_4802_316.t0 14.282
R6439 a_4802_316.n6 a_4802_316.t1 14.282
R6440 a_4802_316.n0 a_4802_316.t4 14.282
R6441 a_4802_316.n0 a_4802_316.t5 14.282
R6442 a_4802_316.n9 a_4802_316.t3 14.282
R6443 a_4802_316.t2 a_4802_316.n9 14.282
R6444 a_4802_316.n7 a_4802_316.n6 1.511
R6445 a_4802_316.n4 a_4802_316.n3 0.999
R6446 a_4802_316.n2 a_4802_316.n1 0.999
R6447 a_4802_316.n8 a_4802_316.n7 0.669
R6448 a_4802_316.n5 a_4802_316.n4 0.575
R6449 a_4802_316.n7 a_4802_316.n5 0.227
R6450 a_4802_316.n5 a_4802_316.n2 0.2
R6451 a_4802_316.n9 a_4802_316.n8 0.001
R6452 a_9558_n2506.n0 a_9558_n2506.t9 214.335
R6453 a_9558_n2506.t7 a_9558_n2506.n0 214.335
R6454 a_9558_n2506.n1 a_9558_n2506.t7 143.851
R6455 a_9558_n2506.n1 a_9558_n2506.t10 135.658
R6456 a_9558_n2506.n0 a_9558_n2506.t8 80.333
R6457 a_9558_n2506.n2 a_9558_n2506.t4 28.565
R6458 a_9558_n2506.n2 a_9558_n2506.t5 28.565
R6459 a_9558_n2506.n4 a_9558_n2506.t6 28.565
R6460 a_9558_n2506.n4 a_9558_n2506.t1 28.565
R6461 a_9558_n2506.n7 a_9558_n2506.t2 28.565
R6462 a_9558_n2506.t3 a_9558_n2506.n7 28.565
R6463 a_9558_n2506.n6 a_9558_n2506.t0 9.714
R6464 a_9558_n2506.n7 a_9558_n2506.n6 1.003
R6465 a_9558_n2506.n5 a_9558_n2506.n3 0.833
R6466 a_9558_n2506.n3 a_9558_n2506.n2 0.653
R6467 a_9558_n2506.n5 a_9558_n2506.n4 0.653
R6468 a_9558_n2506.n6 a_9558_n2506.n5 0.341
R6469 a_9558_n2506.n3 a_9558_n2506.n1 0.032
R6470 a_32485_160.t0 a_32485_160.t1 17.4
R6471 a_11345_n5466.n5 a_11345_n5466.n7 0.575
R6472 a_11345_n5466.n9 a_11345_n5466.n5 0.2
R6473 a_11345_n5466.t6 a_11345_n5466.n9 16.058
R6474 a_11345_n5466.n9 a_11345_n5466.n8 0.999
R6475 a_11345_n5466.n8 a_11345_n5466.t10 14.282
R6476 a_11345_n5466.n8 a_11345_n5466.t11 14.282
R6477 a_11345_n5466.n7 a_11345_n5466.n6 0.999
R6478 a_11345_n5466.n6 a_11345_n5466.t4 14.282
R6479 a_11345_n5466.n6 a_11345_n5466.t3 14.282
R6480 a_11345_n5466.n7 a_11345_n5466.t5 16.058
R6481 a_11345_n5466.n5 a_11345_n5466.n3 0.227
R6482 a_11345_n5466.n3 a_11345_n5466.n4 1.511
R6483 a_11345_n5466.n4 a_11345_n5466.t9 14.282
R6484 a_11345_n5466.n4 a_11345_n5466.t8 14.282
R6485 a_11345_n5466.n3 a_11345_n5466.n0 0.669
R6486 a_11345_n5466.n0 a_11345_n5466.n1 0.001
R6487 a_11345_n5466.n0 a_11345_n5466.n2 267.767
R6488 a_11345_n5466.n2 a_11345_n5466.t0 14.282
R6489 a_11345_n5466.n2 a_11345_n5466.t2 14.282
R6490 a_11345_n5466.n1 a_11345_n5466.t7 14.282
R6491 a_11345_n5466.n1 a_11345_n5466.t1 14.282
R6492 a_13025_n2630.n0 a_13025_n2630.t4 14.282
R6493 a_13025_n2630.n0 a_13025_n2630.t3 14.282
R6494 a_13025_n2630.n1 a_13025_n2630.t0 14.282
R6495 a_13025_n2630.n1 a_13025_n2630.t1 14.282
R6496 a_13025_n2630.t2 a_13025_n2630.n3 14.282
R6497 a_13025_n2630.n3 a_13025_n2630.t5 14.282
R6498 a_13025_n2630.n2 a_13025_n2630.n0 2.546
R6499 a_13025_n2630.n2 a_13025_n2630.n1 2.367
R6500 a_13025_n2630.n3 a_13025_n2630.n2 0.001
R6501 a_26192_3240.t8 a_26192_3240.n2 404.877
R6502 a_26192_3240.n1 a_26192_3240.t7 210.902
R6503 a_26192_3240.n3 a_26192_3240.t8 136.943
R6504 a_26192_3240.n2 a_26192_3240.n1 107.801
R6505 a_26192_3240.n1 a_26192_3240.t5 80.333
R6506 a_26192_3240.n2 a_26192_3240.t6 80.333
R6507 a_26192_3240.n0 a_26192_3240.t4 17.4
R6508 a_26192_3240.n0 a_26192_3240.t0 17.4
R6509 a_26192_3240.n4 a_26192_3240.t3 15.032
R6510 a_26192_3240.n5 a_26192_3240.t2 14.282
R6511 a_26192_3240.t1 a_26192_3240.n5 14.282
R6512 a_26192_3240.n5 a_26192_3240.n4 1.65
R6513 a_26192_3240.n3 a_26192_3240.n0 0.672
R6514 a_26192_3240.n4 a_26192_3240.n3 0.665
R6515 Y[7].n0 Y[7].t2 28.57
R6516 Y[7].n1 Y[7].t1 28.565
R6517 Y[7].n1 Y[7].t3 28.565
R6518 Y[7].n0 Y[7].t0 17.638
R6519 Y[7] Y[7].n2 5.368
R6520 Y[7].n2 Y[7].n1 0.69
R6521 Y[7].n2 Y[7].n0 0.6
R6522 a_24748_404.t4 a_24748_404.n0 14.282
R6523 a_24748_404.n0 a_24748_404.t7 14.282
R6524 a_24748_404.n0 a_24748_404.n12 90.436
R6525 a_24748_404.n8 a_24748_404.n11 50.575
R6526 a_24748_404.n12 a_24748_404.n8 74.302
R6527 a_24748_404.n11 a_24748_404.n10 157.665
R6528 a_24748_404.n10 a_24748_404.t3 8.7
R6529 a_24748_404.n10 a_24748_404.t5 8.7
R6530 a_24748_404.n11 a_24748_404.n9 122.999
R6531 a_24748_404.n9 a_24748_404.t1 14.282
R6532 a_24748_404.n9 a_24748_404.t0 14.282
R6533 a_24748_404.n8 a_24748_404.n7 90.416
R6534 a_24748_404.n7 a_24748_404.t2 14.282
R6535 a_24748_404.n7 a_24748_404.t6 14.282
R6536 a_24748_404.n12 a_24748_404.n1 342.688
R6537 a_24748_404.n1 a_24748_404.n6 126.566
R6538 a_24748_404.n6 a_24748_404.t11 294.653
R6539 a_24748_404.n6 a_24748_404.t9 111.663
R6540 a_24748_404.n1 a_24748_404.n5 552.333
R6541 a_24748_404.n5 a_24748_404.n4 6.615
R6542 a_24748_404.n4 a_24748_404.t13 93.989
R6543 a_24748_404.n5 a_24748_404.n3 97.816
R6544 a_24748_404.n3 a_24748_404.t10 80.333
R6545 a_24748_404.n3 a_24748_404.t12 394.151
R6546 a_24748_404.t12 a_24748_404.n2 269.523
R6547 a_24748_404.n2 a_24748_404.t8 160.666
R6548 a_24748_404.n2 a_24748_404.t14 269.523
R6549 a_24748_404.n4 a_24748_404.t15 198.043
R6550 a_13243_n5466.n0 a_13243_n5466.t8 14.282
R6551 a_13243_n5466.t0 a_13243_n5466.n0 14.282
R6552 a_13243_n5466.n0 a_13243_n5466.n9 0.999
R6553 a_13243_n5466.n6 a_13243_n5466.n8 0.575
R6554 a_13243_n5466.n9 a_13243_n5466.n6 0.2
R6555 a_13243_n5466.n9 a_13243_n5466.t1 16.058
R6556 a_13243_n5466.n8 a_13243_n5466.n7 0.999
R6557 a_13243_n5466.n7 a_13243_n5466.t4 14.282
R6558 a_13243_n5466.n7 a_13243_n5466.t3 14.282
R6559 a_13243_n5466.n8 a_13243_n5466.t2 16.058
R6560 a_13243_n5466.n6 a_13243_n5466.n4 0.227
R6561 a_13243_n5466.n4 a_13243_n5466.n5 1.511
R6562 a_13243_n5466.n5 a_13243_n5466.t7 14.282
R6563 a_13243_n5466.n5 a_13243_n5466.t6 14.282
R6564 a_13243_n5466.n4 a_13243_n5466.n1 0.669
R6565 a_13243_n5466.n1 a_13243_n5466.n2 0.001
R6566 a_13243_n5466.n1 a_13243_n5466.n3 267.767
R6567 a_13243_n5466.n3 a_13243_n5466.t9 14.282
R6568 a_13243_n5466.n3 a_13243_n5466.t11 14.282
R6569 a_13243_n5466.n2 a_13243_n5466.t5 14.282
R6570 a_13243_n5466.n2 a_13243_n5466.t10 14.282
R6571 a_16227_n4155.n2 a_16227_n4155.t10 214.335
R6572 a_16227_n4155.t8 a_16227_n4155.n2 214.335
R6573 a_16227_n4155.n3 a_16227_n4155.t8 143.851
R6574 a_16227_n4155.n3 a_16227_n4155.t7 135.658
R6575 a_16227_n4155.n2 a_16227_n4155.t9 80.333
R6576 a_16227_n4155.n4 a_16227_n4155.t0 28.565
R6577 a_16227_n4155.n4 a_16227_n4155.t1 28.565
R6578 a_16227_n4155.n0 a_16227_n4155.t4 28.565
R6579 a_16227_n4155.n0 a_16227_n4155.t5 28.565
R6580 a_16227_n4155.t2 a_16227_n4155.n7 28.565
R6581 a_16227_n4155.n7 a_16227_n4155.t6 28.565
R6582 a_16227_n4155.n1 a_16227_n4155.t3 9.714
R6583 a_16227_n4155.n1 a_16227_n4155.n0 1.003
R6584 a_16227_n4155.n6 a_16227_n4155.n5 0.833
R6585 a_16227_n4155.n5 a_16227_n4155.n4 0.653
R6586 a_16227_n4155.n7 a_16227_n4155.n6 0.653
R6587 a_16227_n4155.n6 a_16227_n4155.n1 0.341
R6588 a_16227_n4155.n5 a_16227_n4155.n3 0.032
R6589 a_23094_1077.t0 a_23094_1077.t1 17.4
R6590 a_3021_n4154.n0 a_3021_n4154.t9 214.335
R6591 a_3021_n4154.t7 a_3021_n4154.n0 214.335
R6592 a_3021_n4154.n1 a_3021_n4154.t7 143.851
R6593 a_3021_n4154.n1 a_3021_n4154.t10 135.658
R6594 a_3021_n4154.n0 a_3021_n4154.t8 80.333
R6595 a_3021_n4154.n2 a_3021_n4154.t4 28.565
R6596 a_3021_n4154.n2 a_3021_n4154.t5 28.565
R6597 a_3021_n4154.n4 a_3021_n4154.t6 28.565
R6598 a_3021_n4154.n4 a_3021_n4154.t0 28.565
R6599 a_3021_n4154.n7 a_3021_n4154.t1 28.565
R6600 a_3021_n4154.t2 a_3021_n4154.n7 28.565
R6601 a_3021_n4154.n6 a_3021_n4154.t3 9.714
R6602 a_3021_n4154.n7 a_3021_n4154.n6 1.003
R6603 a_3021_n4154.n5 a_3021_n4154.n3 0.833
R6604 a_3021_n4154.n3 a_3021_n4154.n2 0.653
R6605 a_3021_n4154.n5 a_3021_n4154.n4 0.653
R6606 a_3021_n4154.n6 a_3021_n4154.n5 0.341
R6607 a_3021_n4154.n3 a_3021_n4154.n1 0.032
R6608 a_23086_n4791.t0 a_23086_n4791.t1 17.4
R6609 a_13655_n5492.n1 a_13655_n5492.t6 318.922
R6610 a_13655_n5492.n0 a_13655_n5492.t5 274.739
R6611 a_13655_n5492.n0 a_13655_n5492.t7 274.739
R6612 a_13655_n5492.n1 a_13655_n5492.t4 269.116
R6613 a_13655_n5492.t6 a_13655_n5492.n0 179.946
R6614 a_13655_n5492.n2 a_13655_n5492.n1 105.178
R6615 a_13655_n5492.n3 a_13655_n5492.t1 29.444
R6616 a_13655_n5492.n4 a_13655_n5492.t2 28.565
R6617 a_13655_n5492.t3 a_13655_n5492.n4 28.565
R6618 a_13655_n5492.n2 a_13655_n5492.t0 18.145
R6619 a_13655_n5492.n3 a_13655_n5492.n2 2.878
R6620 a_13655_n5492.n4 a_13655_n5492.n3 0.764
R6621 a_31118_n8468.t0 a_31118_n8468.t1 17.4
R6622 a_25050_3236.t6 a_25050_3236.n2 404.877
R6623 a_25050_3236.n1 a_25050_3236.t7 210.902
R6624 a_25050_3236.n3 a_25050_3236.t6 136.943
R6625 a_25050_3236.n2 a_25050_3236.n1 107.801
R6626 a_25050_3236.n1 a_25050_3236.t8 80.333
R6627 a_25050_3236.n2 a_25050_3236.t5 80.333
R6628 a_25050_3236.n0 a_25050_3236.t0 17.4
R6629 a_25050_3236.n0 a_25050_3236.t4 17.4
R6630 a_25050_3236.n4 a_25050_3236.t3 15.032
R6631 a_25050_3236.t1 a_25050_3236.n5 14.282
R6632 a_25050_3236.n5 a_25050_3236.t2 14.282
R6633 a_25050_3236.n5 a_25050_3236.n4 1.65
R6634 a_25050_3236.n3 a_25050_3236.n0 0.672
R6635 a_25050_3236.n4 a_25050_3236.n3 0.665
R6636 a_25314_2653.t7 a_25314_2653.t6 800.071
R6637 a_25314_2653.n3 a_25314_2653.n2 672.951
R6638 a_25314_2653.n1 a_25314_2653.t4 285.109
R6639 a_25314_2653.n2 a_25314_2653.t7 193.602
R6640 a_25314_2653.n1 a_25314_2653.t5 160.666
R6641 a_25314_2653.n2 a_25314_2653.n1 91.507
R6642 a_25314_2653.t3 a_25314_2653.n4 28.57
R6643 a_25314_2653.n0 a_25314_2653.t2 28.565
R6644 a_25314_2653.n0 a_25314_2653.t1 28.565
R6645 a_25314_2653.n4 a_25314_2653.t0 17.638
R6646 a_25314_2653.n3 a_25314_2653.n0 0.69
R6647 a_25314_2653.n4 a_25314_2653.n3 0.6
R6648 a_26882_n328.t0 a_26882_n328.t1 17.4
R6649 a_31118_n625.t0 a_31118_n625.t1 17.4
R6650 a_9564_3364.n0 a_9564_3364.t8 214.335
R6651 a_9564_3364.t7 a_9564_3364.n0 214.335
R6652 a_9564_3364.n1 a_9564_3364.t7 143.851
R6653 a_9564_3364.n1 a_9564_3364.t9 135.658
R6654 a_9564_3364.n0 a_9564_3364.t10 80.333
R6655 a_9564_3364.n2 a_9564_3364.t5 28.565
R6656 a_9564_3364.n2 a_9564_3364.t4 28.565
R6657 a_9564_3364.n4 a_9564_3364.t6 28.565
R6658 a_9564_3364.n4 a_9564_3364.t1 28.565
R6659 a_9564_3364.t3 a_9564_3364.n7 28.565
R6660 a_9564_3364.n7 a_9564_3364.t2 28.565
R6661 a_9564_3364.n6 a_9564_3364.t0 9.714
R6662 a_9564_3364.n7 a_9564_3364.n6 1.003
R6663 a_9564_3364.n5 a_9564_3364.n3 0.833
R6664 a_9564_3364.n3 a_9564_3364.n2 0.653
R6665 a_9564_3364.n5 a_9564_3364.n4 0.653
R6666 a_9564_3364.n6 a_9564_3364.n5 0.341
R6667 a_9564_3364.n3 a_9564_3364.n1 0.032
R6668 a_10154_2927.t7 a_10154_2927.t5 800.071
R6669 a_10154_2927.n2 a_10154_2927.n1 659.097
R6670 a_10154_2927.n0 a_10154_2927.t6 285.109
R6671 a_10154_2927.n1 a_10154_2927.t7 193.602
R6672 a_10154_2927.n4 a_10154_2927.n3 192.754
R6673 a_10154_2927.n0 a_10154_2927.t4 160.666
R6674 a_10154_2927.n1 a_10154_2927.n0 91.507
R6675 a_10154_2927.n3 a_10154_2927.t2 28.568
R6676 a_10154_2927.n4 a_10154_2927.t1 28.565
R6677 a_10154_2927.t3 a_10154_2927.n4 28.565
R6678 a_10154_2927.n2 a_10154_2927.t0 19.061
R6679 a_10154_2927.n3 a_10154_2927.n2 1.005
R6680 a_20027_n8268.n0 a_20027_n8268.t10 214.335
R6681 a_20027_n8268.t8 a_20027_n8268.n0 214.335
R6682 a_20027_n8268.n1 a_20027_n8268.t8 143.85
R6683 a_20027_n8268.n1 a_20027_n8268.t7 135.66
R6684 a_20027_n8268.n0 a_20027_n8268.t9 80.333
R6685 a_20027_n8268.n2 a_20027_n8268.t1 28.565
R6686 a_20027_n8268.n2 a_20027_n8268.t2 28.565
R6687 a_20027_n8268.n4 a_20027_n8268.t0 28.565
R6688 a_20027_n8268.n4 a_20027_n8268.t6 28.565
R6689 a_20027_n8268.t3 a_20027_n8268.n7 28.565
R6690 a_20027_n8268.n7 a_20027_n8268.t4 28.565
R6691 a_20027_n8268.n6 a_20027_n8268.t5 9.714
R6692 a_20027_n8268.n7 a_20027_n8268.n6 1.003
R6693 a_20027_n8268.n5 a_20027_n8268.n3 0.836
R6694 a_20027_n8268.n5 a_20027_n8268.n4 0.653
R6695 a_20027_n8268.n3 a_20027_n8268.n2 0.65
R6696 a_20027_n8268.n6 a_20027_n8268.n5 0.341
R6697 a_20027_n8268.n3 a_20027_n8268.n1 0.032
R6698 a_9578_1714.n0 a_9578_1714.t9 214.335
R6699 a_9578_1714.t7 a_9578_1714.n0 214.335
R6700 a_9578_1714.n1 a_9578_1714.t7 143.851
R6701 a_9578_1714.n1 a_9578_1714.t8 135.658
R6702 a_9578_1714.n0 a_9578_1714.t10 80.333
R6703 a_9578_1714.n2 a_9578_1714.t5 28.565
R6704 a_9578_1714.n2 a_9578_1714.t6 28.565
R6705 a_9578_1714.n4 a_9578_1714.t4 28.565
R6706 a_9578_1714.n4 a_9578_1714.t1 28.565
R6707 a_9578_1714.t3 a_9578_1714.n7 28.565
R6708 a_9578_1714.n7 a_9578_1714.t2 28.565
R6709 a_9578_1714.n6 a_9578_1714.t0 9.714
R6710 a_9578_1714.n7 a_9578_1714.n6 1.003
R6711 a_9578_1714.n5 a_9578_1714.n3 0.833
R6712 a_9578_1714.n3 a_9578_1714.n2 0.653
R6713 a_9578_1714.n5 a_9578_1714.n4 0.653
R6714 a_9578_1714.n6 a_9578_1714.n5 0.341
R6715 a_9578_1714.n3 a_9578_1714.n1 0.032
R6716 a_9815_1077.t0 a_9815_1077.t1 17.4
R6717 a_18417_310.n1 a_18417_310.t6 318.922
R6718 a_18417_310.n0 a_18417_310.t7 274.739
R6719 a_18417_310.n0 a_18417_310.t5 274.739
R6720 a_18417_310.n1 a_18417_310.t4 269.116
R6721 a_18417_310.t6 a_18417_310.n0 179.946
R6722 a_18417_310.n2 a_18417_310.n1 107.263
R6723 a_18417_310.n3 a_18417_310.t1 29.444
R6724 a_18417_310.n4 a_18417_310.t2 28.565
R6725 a_18417_310.t3 a_18417_310.n4 28.565
R6726 a_18417_310.n2 a_18417_310.t0 18.145
R6727 a_18417_310.n3 a_18417_310.n2 2.878
R6728 a_18417_310.n4 a_18417_310.n3 0.764
R6729 a_18123_n396.t0 a_18123_n396.t1 380.209
R6730 a_5206_n5490.n1 a_5206_n5490.t6 318.922
R6731 a_5206_n5490.n0 a_5206_n5490.t5 274.739
R6732 a_5206_n5490.n0 a_5206_n5490.t7 274.739
R6733 a_5206_n5490.n1 a_5206_n5490.t4 269.116
R6734 a_5206_n5490.t6 a_5206_n5490.n0 179.946
R6735 a_5206_n5490.n2 a_5206_n5490.n1 107.263
R6736 a_5206_n5490.n3 a_5206_n5490.t1 29.444
R6737 a_5206_n5490.n4 a_5206_n5490.t2 28.565
R6738 a_5206_n5490.t3 a_5206_n5490.n4 28.565
R6739 a_5206_n5490.n2 a_5206_n5490.t0 18.145
R6740 a_5206_n5490.n3 a_5206_n5490.n2 2.878
R6741 a_5206_n5490.n4 a_5206_n5490.n3 0.764
R6742 a_23081_n6395.t0 a_23081_n6395.t1 17.4
R6743 a_6364_3152.t5 a_6364_3152.n2 404.877
R6744 a_6364_3152.n1 a_6364_3152.t8 210.902
R6745 a_6364_3152.n3 a_6364_3152.t5 136.943
R6746 a_6364_3152.n2 a_6364_3152.n1 107.801
R6747 a_6364_3152.n1 a_6364_3152.t7 80.333
R6748 a_6364_3152.n2 a_6364_3152.t6 80.333
R6749 a_6364_3152.n0 a_6364_3152.t0 17.4
R6750 a_6364_3152.n0 a_6364_3152.t2 17.4
R6751 a_6364_3152.n4 a_6364_3152.t4 15.032
R6752 a_6364_3152.n5 a_6364_3152.t3 14.282
R6753 a_6364_3152.t1 a_6364_3152.n5 14.282
R6754 a_6364_3152.n5 a_6364_3152.n4 1.65
R6755 a_6364_3152.n3 a_6364_3152.n0 0.672
R6756 a_6364_3152.n4 a_6364_3152.n3 0.665
R6757 a_6482_3152.n0 a_6482_3152.t1 14.282
R6758 a_6482_3152.n0 a_6482_3152.t3 14.282
R6759 a_6482_3152.n1 a_6482_3152.t4 14.282
R6760 a_6482_3152.n1 a_6482_3152.t5 14.282
R6761 a_6482_3152.t0 a_6482_3152.n3 14.282
R6762 a_6482_3152.n3 a_6482_3152.t2 14.282
R6763 a_6482_3152.n2 a_6482_3152.n0 2.546
R6764 a_6482_3152.n2 a_6482_3152.n1 2.367
R6765 a_6482_3152.n3 a_6482_3152.n2 0.001
R6766 a_3252_2639.t0 a_3252_2639.t1 17.4
R6767 a_26093_n4771.n2 a_26093_n4771.t6 318.922
R6768 a_26093_n4771.n1 a_26093_n4771.t5 273.935
R6769 a_26093_n4771.n1 a_26093_n4771.t7 273.935
R6770 a_26093_n4771.n2 a_26093_n4771.t4 269.116
R6771 a_26093_n4771.n4 a_26093_n4771.n0 193.227
R6772 a_26093_n4771.t6 a_26093_n4771.n1 179.142
R6773 a_26093_n4771.n3 a_26093_n4771.n2 106.999
R6774 a_26093_n4771.t3 a_26093_n4771.n4 28.568
R6775 a_26093_n4771.n0 a_26093_n4771.t1 28.565
R6776 a_26093_n4771.n0 a_26093_n4771.t2 28.565
R6777 a_26093_n4771.n3 a_26093_n4771.t0 18.149
R6778 a_26093_n4771.n4 a_26093_n4771.n3 3.726
R6779 a_13575_4805.t0 a_13575_4805.t1 17.4
R6780 a_9572_n4156.n4 a_9572_n4156.t9 214.335
R6781 a_9572_n4156.t7 a_9572_n4156.n4 214.335
R6782 a_9572_n4156.n5 a_9572_n4156.t7 143.851
R6783 a_9572_n4156.n5 a_9572_n4156.t10 135.658
R6784 a_9572_n4156.n4 a_9572_n4156.t8 80.333
R6785 a_9572_n4156.n0 a_9572_n4156.t5 28.565
R6786 a_9572_n4156.n0 a_9572_n4156.t6 28.565
R6787 a_9572_n4156.n2 a_9572_n4156.t1 28.565
R6788 a_9572_n4156.n2 a_9572_n4156.t4 28.565
R6789 a_9572_n4156.t2 a_9572_n4156.n7 28.565
R6790 a_9572_n4156.n7 a_9572_n4156.t0 28.565
R6791 a_9572_n4156.n1 a_9572_n4156.t3 9.714
R6792 a_9572_n4156.n1 a_9572_n4156.n0 1.003
R6793 a_9572_n4156.n6 a_9572_n4156.n3 0.833
R6794 a_9572_n4156.n3 a_9572_n4156.n2 0.653
R6795 a_9572_n4156.n7 a_9572_n4156.n6 0.653
R6796 a_9572_n4156.n3 a_9572_n4156.n1 0.341
R6797 a_9572_n4156.n6 a_9572_n4156.n5 0.032
R6798 a_16812_n6196.t5 a_16812_n6196.t4 574.43
R6799 a_16812_n6196.n0 a_16812_n6196.t7 285.109
R6800 a_16812_n6196.n2 a_16812_n6196.n1 197.217
R6801 a_16812_n6196.n4 a_16812_n6196.n3 192.754
R6802 a_16812_n6196.n0 a_16812_n6196.t6 160.666
R6803 a_16812_n6196.n1 a_16812_n6196.t5 160.666
R6804 a_16812_n6196.n1 a_16812_n6196.n0 114.829
R6805 a_16812_n6196.n3 a_16812_n6196.t1 28.568
R6806 a_16812_n6196.n4 a_16812_n6196.t2 28.565
R6807 a_16812_n6196.t3 a_16812_n6196.n4 28.565
R6808 a_16812_n6196.n2 a_16812_n6196.t0 18.838
R6809 a_16812_n6196.n3 a_16812_n6196.n2 1.129
R6810 B[0].t12 B[0].t14 437.233
R6811 B[0].t0 B[0].t7 437.233
R6812 B[0].t4 B[0].t10 437.233
R6813 B[0].t5 B[0].t8 415.315
R6814 B[0].n2 B[0].t5 225.375
R6815 B[0].n5 B[0].t4 223.992
R6816 B[0].n5 B[0].t0 217.885
R6817 B[0].n2 B[0].t12 216.848
R6818 B[0].n1 B[0].t11 214.686
R6819 B[0].t14 B[0].n1 214.686
R6820 B[0].n3 B[0].t15 214.686
R6821 B[0].t7 B[0].n3 214.686
R6822 B[0].n4 B[0].t3 214.686
R6823 B[0].t10 B[0].n4 214.686
R6824 B[0].n0 B[0].t2 214.335
R6825 B[0].t8 B[0].n0 214.335
R6826 B[0].n1 B[0].t1 80.333
R6827 B[0].n0 B[0].t9 80.333
R6828 B[0].n3 B[0].t6 80.333
R6829 B[0].n4 B[0].t13 80.333
R6830 B[0].n6 B[0].n2 62.925
R6831 B[0].n6 B[0].n5 0.469
R6832 B[0] B[0].n6 0.446
R6833 a_114_n5080.n0 a_114_n5080.t9 214.335
R6834 a_114_n5080.t7 a_114_n5080.n0 214.335
R6835 a_114_n5080.n1 a_114_n5080.t7 143.851
R6836 a_114_n5080.n1 a_114_n5080.t10 135.658
R6837 a_114_n5080.n0 a_114_n5080.t8 80.333
R6838 a_114_n5080.n2 a_114_n5080.t4 28.565
R6839 a_114_n5080.n2 a_114_n5080.t5 28.565
R6840 a_114_n5080.n4 a_114_n5080.t6 28.565
R6841 a_114_n5080.n4 a_114_n5080.t2 28.565
R6842 a_114_n5080.t3 a_114_n5080.n7 28.565
R6843 a_114_n5080.n7 a_114_n5080.t1 28.565
R6844 a_114_n5080.n6 a_114_n5080.t0 9.714
R6845 a_114_n5080.n7 a_114_n5080.n6 1.003
R6846 a_114_n5080.n5 a_114_n5080.n3 0.833
R6847 a_114_n5080.n3 a_114_n5080.n2 0.653
R6848 a_114_n5080.n5 a_114_n5080.n4 0.653
R6849 a_114_n5080.n6 a_114_n5080.n5 0.341
R6850 a_114_n5080.n3 a_114_n5080.n1 0.032
R6851 a_351_n5717.t0 a_351_n5717.t1 17.4
R6852 a_17578_1029.n1 a_17578_1029.t5 318.922
R6853 a_17578_1029.n0 a_17578_1029.t7 273.935
R6854 a_17578_1029.n0 a_17578_1029.t4 273.935
R6855 a_17578_1029.n1 a_17578_1029.t6 269.116
R6856 a_17578_1029.n4 a_17578_1029.n3 193.227
R6857 a_17578_1029.t5 a_17578_1029.n0 179.142
R6858 a_17578_1029.n2 a_17578_1029.n1 106.999
R6859 a_17578_1029.n3 a_17578_1029.t1 28.568
R6860 a_17578_1029.t3 a_17578_1029.n4 28.565
R6861 a_17578_1029.n4 a_17578_1029.t2 28.565
R6862 a_17578_1029.n2 a_17578_1029.t0 18.149
R6863 a_17578_1029.n3 a_17578_1029.n2 3.726
R6864 a_11463_n6198.t0 a_11463_n6198.t1 380.209
R6865 a_117_958.n4 a_117_958.t9 214.335
R6866 a_117_958.t8 a_117_958.n4 214.335
R6867 a_117_958.n5 a_117_958.t8 143.851
R6868 a_117_958.n5 a_117_958.t10 135.658
R6869 a_117_958.n4 a_117_958.t7 80.333
R6870 a_117_958.n0 a_117_958.t4 28.565
R6871 a_117_958.n0 a_117_958.t6 28.565
R6872 a_117_958.n2 a_117_958.t0 28.565
R6873 a_117_958.n2 a_117_958.t5 28.565
R6874 a_117_958.t2 a_117_958.n7 28.565
R6875 a_117_958.n7 a_117_958.t1 28.565
R6876 a_117_958.n1 a_117_958.t3 9.714
R6877 a_117_958.n1 a_117_958.n0 1.003
R6878 a_117_958.n6 a_117_958.n3 0.833
R6879 a_117_958.n3 a_117_958.n2 0.653
R6880 a_117_958.n7 a_117_958.n6 0.653
R6881 a_117_958.n3 a_117_958.n1 0.341
R6882 a_117_958.n6 a_117_958.n5 0.032
R6883 a_4367_n4771.n2 a_4367_n4771.t6 318.922
R6884 a_4367_n4771.n1 a_4367_n4771.t5 273.935
R6885 a_4367_n4771.n1 a_4367_n4771.t7 273.935
R6886 a_4367_n4771.n2 a_4367_n4771.t4 269.116
R6887 a_4367_n4771.n4 a_4367_n4771.n0 193.227
R6888 a_4367_n4771.t6 a_4367_n4771.n1 179.142
R6889 a_4367_n4771.n3 a_4367_n4771.n2 106.999
R6890 a_4367_n4771.t3 a_4367_n4771.n4 28.568
R6891 a_4367_n4771.n0 a_4367_n4771.t1 28.565
R6892 a_4367_n4771.n0 a_4367_n4771.t2 28.565
R6893 a_4367_n4771.n3 a_4367_n4771.t0 18.149
R6894 a_4367_n4771.n4 a_4367_n4771.n3 3.726
R6895 a_4912_n6196.t0 a_4912_n6196.t1 380.209
R6896 a_5486_2565.t7 a_5486_2565.t6 800.071
R6897 a_5486_2565.n3 a_5486_2565.n2 672.951
R6898 a_5486_2565.n1 a_5486_2565.t4 285.109
R6899 a_5486_2565.n2 a_5486_2565.t7 193.602
R6900 a_5486_2565.n1 a_5486_2565.t5 160.666
R6901 a_5486_2565.n2 a_5486_2565.n1 91.507
R6902 a_5486_2565.n0 a_5486_2565.t1 28.57
R6903 a_5486_2565.t3 a_5486_2565.n4 28.565
R6904 a_5486_2565.n4 a_5486_2565.t2 28.565
R6905 a_5486_2565.n0 a_5486_2565.t0 17.638
R6906 a_5486_2565.n4 a_5486_2565.n3 0.69
R6907 a_5486_2565.n3 a_5486_2565.n0 0.6
R6908 a_30880_3466.t0 a_30880_3466.t1 380.209
R6909 a_11883_n2634.n0 a_11883_n2634.t5 14.282
R6910 a_11883_n2634.n0 a_11883_n2634.t0 14.282
R6911 a_11883_n2634.n1 a_11883_n2634.t3 14.282
R6912 a_11883_n2634.n1 a_11883_n2634.t4 14.282
R6913 a_11883_n2634.n3 a_11883_n2634.t1 14.282
R6914 a_11883_n2634.t2 a_11883_n2634.n3 14.282
R6915 a_11883_n2634.n3 a_11883_n2634.n2 2.546
R6916 a_11883_n2634.n2 a_11883_n2634.n1 2.367
R6917 a_11883_n2634.n2 a_11883_n2634.n0 0.001
R6918 a_23080_2727.t0 a_23080_2727.t1 17.4
R6919 a_10924_1097.n1 a_10924_1097.t6 318.922
R6920 a_10924_1097.n0 a_10924_1097.t7 273.935
R6921 a_10924_1097.n0 a_10924_1097.t5 273.935
R6922 a_10924_1097.n1 a_10924_1097.t4 269.116
R6923 a_10924_1097.n4 a_10924_1097.n3 193.227
R6924 a_10924_1097.t6 a_10924_1097.n0 179.142
R6925 a_10924_1097.n2 a_10924_1097.n1 106.999
R6926 a_10924_1097.n3 a_10924_1097.t2 28.568
R6927 a_10924_1097.n4 a_10924_1097.t1 28.565
R6928 a_10924_1097.t3 a_10924_1097.n4 28.565
R6929 a_10924_1097.n2 a_10924_1097.t0 18.149
R6930 a_10924_1097.n3 a_10924_1097.n2 3.726
R6931 a_5340_3148.n0 a_5340_3148.t5 14.282
R6932 a_5340_3148.n0 a_5340_3148.t3 14.282
R6933 a_5340_3148.n1 a_5340_3148.t1 14.282
R6934 a_5340_3148.n1 a_5340_3148.t0 14.282
R6935 a_5340_3148.t2 a_5340_3148.n3 14.282
R6936 a_5340_3148.n3 a_5340_3148.t4 14.282
R6937 a_5340_3148.n2 a_5340_3148.n0 2.546
R6938 a_5340_3148.n2 a_5340_3148.n1 2.367
R6939 a_5340_3148.n3 a_5340_3148.n2 0.001
R6940 a_18005_336.n3 a_18005_336.n1 267.767
R6941 a_18005_336.n7 a_18005_336.t9 16.058
R6942 a_18005_336.t2 a_18005_336.n9 16.058
R6943 a_18005_336.n2 a_18005_336.t4 14.282
R6944 a_18005_336.n2 a_18005_336.t6 14.282
R6945 a_18005_336.n1 a_18005_336.t3 14.282
R6946 a_18005_336.n1 a_18005_336.t5 14.282
R6947 a_18005_336.n4 a_18005_336.t8 14.282
R6948 a_18005_336.n4 a_18005_336.t7 14.282
R6949 a_18005_336.n6 a_18005_336.t11 14.282
R6950 a_18005_336.n6 a_18005_336.t10 14.282
R6951 a_18005_336.n0 a_18005_336.t1 14.282
R6952 a_18005_336.n0 a_18005_336.t0 14.282
R6953 a_18005_336.n5 a_18005_336.n4 1.511
R6954 a_18005_336.n7 a_18005_336.n6 0.999
R6955 a_18005_336.n9 a_18005_336.n0 0.999
R6956 a_18005_336.n5 a_18005_336.n3 0.669
R6957 a_18005_336.n8 a_18005_336.n7 0.575
R6958 a_18005_336.n8 a_18005_336.n5 0.227
R6959 a_18005_336.n9 a_18005_336.n8 0.2
R6960 a_18005_336.n3 a_18005_336.n2 0.001
R6961 a_19471_n4772.n2 a_19471_n4772.t6 318.922
R6962 a_19471_n4772.n1 a_19471_n4772.t4 273.935
R6963 a_19471_n4772.n1 a_19471_n4772.t7 273.935
R6964 a_19471_n4772.n2 a_19471_n4772.t5 269.116
R6965 a_19471_n4772.n4 a_19471_n4772.n0 193.227
R6966 a_19471_n4772.t6 a_19471_n4772.n1 179.142
R6967 a_19471_n4772.n3 a_19471_n4772.n2 106.999
R6968 a_19471_n4772.t3 a_19471_n4772.n4 28.568
R6969 a_19471_n4772.n0 a_19471_n4772.t1 28.565
R6970 a_19471_n4772.n0 a_19471_n4772.t2 28.565
R6971 a_19471_n4772.n3 a_19471_n4772.t0 18.149
R6972 a_19471_n4772.n4 a_19471_n4772.n3 3.726
R6973 B[3].n6 B[3].t1 5229.8
R6974 B[3].t7 B[3].t14 437.233
R6975 B[3].t3 B[3].t13 437.233
R6976 B[3].t1 B[3].t2 415.315
R6977 B[3].t15 B[3].t4 415.315
R6978 B[3].n4 B[3].t15 220.313
R6979 B[3].n5 B[3].t7 219.163
R6980 B[3].n4 B[3].t3 217.194
R6981 B[3].n1 B[3].t0 214.686
R6982 B[3].t14 B[3].n1 214.686
R6983 B[3].n3 B[3].t11 214.686
R6984 B[3].t13 B[3].n3 214.686
R6985 B[3].n0 B[3].t5 214.335
R6986 B[3].t2 B[3].n0 214.335
R6987 B[3].n2 B[3].t9 214.335
R6988 B[3].t4 B[3].n2 214.335
R6989 B[3].n0 B[3].t10 80.333
R6990 B[3].n1 B[3].t8 80.333
R6991 B[3].n2 B[3].t6 80.333
R6992 B[3].n3 B[3].t12 80.333
R6993 B[3].n6 B[3].n5 23.931
R6994 B[3].n5 B[3].n4 11.749
R6995 B[3] B[3].n6 3.368
R6996 a_16459_n6396.t0 a_16459_n6396.t1 17.4
R6997 a_3007_n2504.n0 a_3007_n2504.t9 214.335
R6998 a_3007_n2504.t7 a_3007_n2504.n0 214.335
R6999 a_3007_n2504.n1 a_3007_n2504.t7 143.851
R7000 a_3007_n2504.n1 a_3007_n2504.t10 135.658
R7001 a_3007_n2504.n0 a_3007_n2504.t8 80.333
R7002 a_3007_n2504.n2 a_3007_n2504.t5 28.565
R7003 a_3007_n2504.n2 a_3007_n2504.t6 28.565
R7004 a_3007_n2504.n4 a_3007_n2504.t4 28.565
R7005 a_3007_n2504.n4 a_3007_n2504.t2 28.565
R7006 a_3007_n2504.t3 a_3007_n2504.n7 28.565
R7007 a_3007_n2504.n7 a_3007_n2504.t1 28.565
R7008 a_3007_n2504.n6 a_3007_n2504.t0 9.714
R7009 a_3007_n2504.n7 a_3007_n2504.n6 1.003
R7010 a_3007_n2504.n5 a_3007_n2504.n3 0.833
R7011 a_3007_n2504.n3 a_3007_n2504.n2 0.653
R7012 a_3007_n2504.n5 a_3007_n2504.n4 0.653
R7013 a_3007_n2504.n6 a_3007_n2504.n5 0.341
R7014 a_3007_n2504.n3 a_3007_n2504.n1 0.032
R7015 a_31176_n3414.n1 a_31176_n3414.t7 318.922
R7016 a_31176_n3414.n0 a_31176_n3414.t6 274.739
R7017 a_31176_n3414.n0 a_31176_n3414.t4 274.739
R7018 a_31176_n3414.n1 a_31176_n3414.t5 269.116
R7019 a_31176_n3414.t7 a_31176_n3414.n0 179.946
R7020 a_31176_n3414.n2 a_31176_n3414.n1 107.263
R7021 a_31176_n3414.n3 a_31176_n3414.t1 29.444
R7022 a_31176_n3414.n4 a_31176_n3414.t2 28.565
R7023 a_31176_n3414.t3 a_31176_n3414.n4 28.565
R7024 a_31176_n3414.n2 a_31176_n3414.t0 18.145
R7025 a_31176_n3414.n3 a_31176_n3414.n2 2.878
R7026 a_31176_n3414.n4 a_31176_n3414.n3 0.764
R7027 Y[4].n4 Y[4].n2 157.665
R7028 Y[4] Y[4].n6 145.6
R7029 Y[4].n4 Y[4].n3 122.999
R7030 Y[4].n6 Y[4].n0 90.436
R7031 Y[4].n5 Y[4].n1 90.416
R7032 Y[4].n6 Y[4].n5 74.302
R7033 Y[4].n5 Y[4].n4 50.575
R7034 Y[4].n0 Y[4].t6 14.282
R7035 Y[4].n0 Y[4].t4 14.282
R7036 Y[4].n1 Y[4].t5 14.282
R7037 Y[4].n1 Y[4].t0 14.282
R7038 Y[4].n3 Y[4].t2 14.282
R7039 Y[4].n3 Y[4].t1 14.282
R7040 Y[4].n2 Y[4].t7 8.7
R7041 Y[4].n2 Y[4].t3 8.7
R7042 a_9801_2727.t0 a_9801_2727.t1 17.4
R7043 a_9810_n527.t0 a_9810_n527.t1 17.4
R7044 a_18420_n2633.t5 a_18420_n2633.n2 404.877
R7045 a_18420_n2633.n1 a_18420_n2633.t7 210.902
R7046 a_18420_n2633.n3 a_18420_n2633.t5 136.943
R7047 a_18420_n2633.n2 a_18420_n2633.n1 107.801
R7048 a_18420_n2633.n1 a_18420_n2633.t6 80.333
R7049 a_18420_n2633.n2 a_18420_n2633.t8 80.333
R7050 a_18420_n2633.n0 a_18420_n2633.t4 17.4
R7051 a_18420_n2633.n0 a_18420_n2633.t3 17.4
R7052 a_18420_n2633.n4 a_18420_n2633.t2 15.032
R7053 a_18420_n2633.t0 a_18420_n2633.n5 14.282
R7054 a_18420_n2633.n5 a_18420_n2633.t1 14.282
R7055 a_18420_n2633.n5 a_18420_n2633.n4 1.65
R7056 a_18420_n2633.n3 a_18420_n2633.n0 0.672
R7057 a_18420_n2633.n4 a_18420_n2633.n3 0.665
R7058 a_28877_2088.t0 a_28877_2088.t1 17.4
R7059 a_24748_n328.t0 a_24748_n328.t1 380.209
R7060 a_11757_n5492.n1 a_11757_n5492.t6 318.922
R7061 a_11757_n5492.n0 a_11757_n5492.t5 274.739
R7062 a_11757_n5492.n0 a_11757_n5492.t7 274.739
R7063 a_11757_n5492.n1 a_11757_n5492.t4 269.116
R7064 a_11757_n5492.t6 a_11757_n5492.n0 179.946
R7065 a_11757_n5492.n2 a_11757_n5492.n1 107.263
R7066 a_11757_n5492.n3 a_11757_n5492.t2 29.444
R7067 a_11757_n5492.t3 a_11757_n5492.n4 28.565
R7068 a_11757_n5492.n4 a_11757_n5492.t1 28.565
R7069 a_11757_n5492.n2 a_11757_n5492.t0 18.145
R7070 a_11757_n5492.n3 a_11757_n5492.n2 2.878
R7071 a_11757_n5492.n4 a_11757_n5492.n3 0.764
R7072 a_362_2906.t0 a_362_2906.t1 17.4
R7073 a_26101_1097.n1 a_26101_1097.t6 318.922
R7074 a_26101_1097.n0 a_26101_1097.t5 273.935
R7075 a_26101_1097.n0 a_26101_1097.t4 273.935
R7076 a_26101_1097.n1 a_26101_1097.t7 269.116
R7077 a_26101_1097.n4 a_26101_1097.n3 193.227
R7078 a_26101_1097.t6 a_26101_1097.n0 179.142
R7079 a_26101_1097.n2 a_26101_1097.n1 106.999
R7080 a_26101_1097.n3 a_26101_1097.t1 28.568
R7081 a_26101_1097.t3 a_26101_1097.n4 28.565
R7082 a_26101_1097.n4 a_26101_1097.t2 28.565
R7083 a_26101_1097.n2 a_26101_1097.t0 18.149
R7084 a_26101_1097.n3 a_26101_1097.n2 3.726
R7085 a_5156_n416.t0 a_5156_n416.t1 17.4
R7086 a_98_n2320.n0 a_98_n2320.t10 214.335
R7087 a_98_n2320.t8 a_98_n2320.n0 214.335
R7088 a_98_n2320.n1 a_98_n2320.t8 143.851
R7089 a_98_n2320.n1 a_98_n2320.t7 135.658
R7090 a_98_n2320.n0 a_98_n2320.t9 80.333
R7091 a_98_n2320.n2 a_98_n2320.t5 28.565
R7092 a_98_n2320.n2 a_98_n2320.t6 28.565
R7093 a_98_n2320.n4 a_98_n2320.t4 28.565
R7094 a_98_n2320.n4 a_98_n2320.t0 28.565
R7095 a_98_n2320.n7 a_98_n2320.t1 28.565
R7096 a_98_n2320.t2 a_98_n2320.n7 28.565
R7097 a_98_n2320.n6 a_98_n2320.t3 9.714
R7098 a_98_n2320.n7 a_98_n2320.n6 1.003
R7099 a_98_n2320.n5 a_98_n2320.n3 0.833
R7100 a_98_n2320.n3 a_98_n2320.n2 0.653
R7101 a_98_n2320.n5 a_98_n2320.n4 0.653
R7102 a_98_n2320.n6 a_98_n2320.n5 0.341
R7103 a_98_n2320.n3 a_98_n2320.n1 0.032
R7104 a_23442_n327.t5 a_23442_n327.t6 574.43
R7105 a_23442_n327.n1 a_23442_n327.t7 285.109
R7106 a_23442_n327.n3 a_23442_n327.n2 197.217
R7107 a_23442_n327.n4 a_23442_n327.n0 192.754
R7108 a_23442_n327.n1 a_23442_n327.t4 160.666
R7109 a_23442_n327.n2 a_23442_n327.t5 160.666
R7110 a_23442_n327.n2 a_23442_n327.n1 114.829
R7111 a_23442_n327.t3 a_23442_n327.n4 28.568
R7112 a_23442_n327.n0 a_23442_n327.t2 28.565
R7113 a_23442_n327.n0 a_23442_n327.t1 28.565
R7114 a_23442_n327.n3 a_23442_n327.t0 18.838
R7115 a_23442_n327.n4 a_23442_n327.n3 1.129
R7116 a_25168_3236.n0 a_25168_3236.t4 14.282
R7117 a_25168_3236.n0 a_25168_3236.t0 14.282
R7118 a_25168_3236.n1 a_25168_3236.t3 14.282
R7119 a_25168_3236.n1 a_25168_3236.t5 14.282
R7120 a_25168_3236.t2 a_25168_3236.n3 14.282
R7121 a_25168_3236.n3 a_25168_3236.t1 14.282
R7122 a_25168_3236.n3 a_25168_3236.n2 2.546
R7123 a_25168_3236.n2 a_25168_3236.n1 2.367
R7124 a_25168_3236.n2 a_25168_3236.n0 0.001
R7125 a_30337_n2695.n2 a_30337_n2695.t6 318.922
R7126 a_30337_n2695.n1 a_30337_n2695.t5 273.935
R7127 a_30337_n2695.n1 a_30337_n2695.t7 273.935
R7128 a_30337_n2695.n2 a_30337_n2695.t4 269.116
R7129 a_30337_n2695.n4 a_30337_n2695.n0 193.227
R7130 a_30337_n2695.t6 a_30337_n2695.n1 179.142
R7131 a_30337_n2695.n3 a_30337_n2695.n2 106.999
R7132 a_30337_n2695.t3 a_30337_n2695.n4 28.568
R7133 a_30337_n2695.n0 a_30337_n2695.t1 28.565
R7134 a_30337_n2695.n0 a_30337_n2695.t2 28.565
R7135 a_30337_n2695.n3 a_30337_n2695.t0 18.149
R7136 a_30337_n2695.n4 a_30337_n2695.n3 3.726
R7137 a_30882_n4120.t0 a_30882_n4120.t1 380.209
R7138 a_3597_n2941.t5 a_3597_n2941.t4 800.071
R7139 a_3597_n2941.n2 a_3597_n2941.n1 659.097
R7140 a_3597_n2941.n0 a_3597_n2941.t7 285.109
R7141 a_3597_n2941.n1 a_3597_n2941.t5 193.602
R7142 a_3597_n2941.n4 a_3597_n2941.n3 192.754
R7143 a_3597_n2941.n0 a_3597_n2941.t6 160.666
R7144 a_3597_n2941.n1 a_3597_n2941.n0 91.507
R7145 a_3597_n2941.n3 a_3597_n2941.t1 28.568
R7146 a_3597_n2941.n4 a_3597_n2941.t2 28.565
R7147 a_3597_n2941.t3 a_3597_n2941.n4 28.565
R7148 a_3597_n2941.n2 a_3597_n2941.t0 19.061
R7149 a_3597_n2941.n3 a_3597_n2941.n2 1.005
R7150 a_20229_4826.t0 a_20229_4826.t1 17.4
R7151 a_5478_n3215.t5 a_5478_n3215.t4 800.071
R7152 a_5478_n3215.n3 a_5478_n3215.n2 672.951
R7153 a_5478_n3215.n1 a_5478_n3215.t7 285.109
R7154 a_5478_n3215.n2 a_5478_n3215.t5 193.602
R7155 a_5478_n3215.n1 a_5478_n3215.t6 160.666
R7156 a_5478_n3215.n2 a_5478_n3215.n1 91.507
R7157 a_5478_n3215.t3 a_5478_n3215.n4 28.57
R7158 a_5478_n3215.n0 a_5478_n3215.t1 28.565
R7159 a_5478_n3215.n0 a_5478_n3215.t2 28.565
R7160 a_5478_n3215.n4 a_5478_n3215.t0 17.638
R7161 a_5478_n3215.n3 a_5478_n3215.n0 0.69
R7162 a_5478_n3215.n4 a_5478_n3215.n3 0.6
R7163 a_26184_n2628.t7 a_26184_n2628.n3 404.877
R7164 a_26184_n2628.n2 a_26184_n2628.t5 210.902
R7165 a_26184_n2628.n4 a_26184_n2628.t7 136.943
R7166 a_26184_n2628.n3 a_26184_n2628.n2 107.801
R7167 a_26184_n2628.n2 a_26184_n2628.t8 80.333
R7168 a_26184_n2628.n3 a_26184_n2628.t6 80.333
R7169 a_26184_n2628.n1 a_26184_n2628.t0 17.4
R7170 a_26184_n2628.n1 a_26184_n2628.t1 17.4
R7171 a_26184_n2628.t4 a_26184_n2628.n5 15.032
R7172 a_26184_n2628.n0 a_26184_n2628.t2 14.282
R7173 a_26184_n2628.n0 a_26184_n2628.t3 14.282
R7174 a_26184_n2628.n5 a_26184_n2628.n0 1.65
R7175 a_26184_n2628.n4 a_26184_n2628.n1 0.672
R7176 a_26184_n2628.n5 a_26184_n2628.n4 0.665
R7177 a_28948_n2865.t0 a_28948_n2865.t1 17.4
R7178 a_26310_3240.n0 a_26310_3240.t3 14.282
R7179 a_26310_3240.n0 a_26310_3240.t1 14.282
R7180 a_26310_3240.n1 a_26310_3240.t5 14.282
R7181 a_26310_3240.n1 a_26310_3240.t4 14.282
R7182 a_26310_3240.n3 a_26310_3240.t0 14.282
R7183 a_26310_3240.t2 a_26310_3240.n3 14.282
R7184 a_26310_3240.n3 a_26310_3240.n2 2.546
R7185 a_26310_3240.n2 a_26310_3240.n1 2.367
R7186 a_26310_3240.n2 a_26310_3240.n0 0.001
R7187 a_26638_n6196.t0 a_26638_n6196.t1 380.209
R7188 a_32483_4251.t0 a_32483_4251.t1 17.4
R7189 a_17573_n4772.n2 a_17573_n4772.t6 318.922
R7190 a_17573_n4772.n1 a_17573_n4772.t5 273.935
R7191 a_17573_n4772.n1 a_17573_n4772.t7 273.935
R7192 a_17573_n4772.n2 a_17573_n4772.t4 269.116
R7193 a_17573_n4772.n4 a_17573_n4772.n0 193.227
R7194 a_17573_n4772.t6 a_17573_n4772.n1 179.142
R7195 a_17573_n4772.n3 a_17573_n4772.n2 106.999
R7196 a_17573_n4772.t3 a_17573_n4772.n4 28.568
R7197 a_17573_n4772.n0 a_17573_n4772.t1 28.565
R7198 a_17573_n4772.n0 a_17573_n4772.t2 28.565
R7199 a_17573_n4772.n3 a_17573_n4772.t0 18.149
R7200 a_17573_n4772.n4 a_17573_n4772.n3 3.726
R7201 a_13603_n328.t0 a_13603_n328.t1 17.4
R7202 a_28715_n8143.n0 a_28715_n8143.t9 214.335
R7203 a_28715_n8143.t7 a_28715_n8143.n0 214.335
R7204 a_28715_n8143.n1 a_28715_n8143.t7 143.851
R7205 a_28715_n8143.n1 a_28715_n8143.t10 135.658
R7206 a_28715_n8143.n0 a_28715_n8143.t8 80.333
R7207 a_28715_n8143.n2 a_28715_n8143.t4 28.565
R7208 a_28715_n8143.n2 a_28715_n8143.t5 28.565
R7209 a_28715_n8143.n4 a_28715_n8143.t6 28.565
R7210 a_28715_n8143.n4 a_28715_n8143.t1 28.565
R7211 a_28715_n8143.n7 a_28715_n8143.t2 28.565
R7212 a_28715_n8143.t3 a_28715_n8143.n7 28.565
R7213 a_28715_n8143.n6 a_28715_n8143.t0 9.714
R7214 a_28715_n8143.n7 a_28715_n8143.n6 1.003
R7215 a_28715_n8143.n5 a_28715_n8143.n3 0.833
R7216 a_28715_n8143.n3 a_28715_n8143.n2 0.653
R7217 a_28715_n8143.n5 a_28715_n8143.n4 0.653
R7218 a_28715_n8143.n6 a_28715_n8143.n5 0.341
R7219 a_28715_n8143.n3 a_28715_n8143.n1 0.032
R7220 a_28952_n8780.t0 a_28952_n8780.t1 17.4
R7221 a_18118_n6197.t0 a_18118_n6197.t1 380.209
R7222 a_5148_n6196.t0 a_5148_n6196.t1 17.4
R7223 a_9795_n3143.t0 a_9795_n3143.t1 17.4
R7224 a_30337_800.n1 a_30337_800.t6 318.922
R7225 a_30337_800.n0 a_30337_800.t7 273.935
R7226 a_30337_800.n0 a_30337_800.t4 273.935
R7227 a_30337_800.n1 a_30337_800.t5 269.116
R7228 a_30337_800.n4 a_30337_800.n3 193.227
R7229 a_30337_800.t6 a_30337_800.n0 179.142
R7230 a_30337_800.n2 a_30337_800.n1 106.999
R7231 a_30337_800.n3 a_30337_800.t2 28.568
R7232 a_30337_800.t3 a_30337_800.n4 28.565
R7233 a_30337_800.n4 a_30337_800.t1 28.565
R7234 a_30337_800.n2 a_30337_800.t0 18.149
R7235 a_30337_800.n3 a_30337_800.n2 3.726
R7236 a_18538_n2633.n0 a_18538_n2633.t5 14.282
R7237 a_18538_n2633.n0 a_18538_n2633.t0 14.282
R7238 a_18538_n2633.n1 a_18538_n2633.t3 14.282
R7239 a_18538_n2633.n1 a_18538_n2633.t4 14.282
R7240 a_18538_n2633.n3 a_18538_n2633.t1 14.282
R7241 a_18538_n2633.t2 a_18538_n2633.n3 14.282
R7242 a_18538_n2633.n3 a_18538_n2633.n2 2.546
R7243 a_18538_n2633.n2 a_18538_n2633.n1 2.367
R7244 a_18538_n2633.n2 a_18538_n2633.n0 0.001
R7245 a_18354_n6197.t0 a_18354_n6197.t1 17.4
R7246 a_25042_378.n1 a_25042_378.t5 318.922
R7247 a_25042_378.n0 a_25042_378.t7 274.739
R7248 a_25042_378.n0 a_25042_378.t4 274.739
R7249 a_25042_378.n1 a_25042_378.t6 269.116
R7250 a_25042_378.t5 a_25042_378.n0 179.946
R7251 a_25042_378.n2 a_25042_378.n1 107.263
R7252 a_25042_378.n3 a_25042_378.t2 29.444
R7253 a_25042_378.t3 a_25042_378.n4 28.565
R7254 a_25042_378.n4 a_25042_378.t1 28.565
R7255 a_25042_378.n2 a_25042_378.t0 18.145
R7256 a_25042_378.n3 a_25042_378.n2 2.878
R7257 a_25042_378.n4 a_25042_378.n3 0.764
R7258 a_7104_n5490.n1 a_7104_n5490.t6 318.922
R7259 a_7104_n5490.n0 a_7104_n5490.t5 274.739
R7260 a_7104_n5490.n0 a_7104_n5490.t7 274.739
R7261 a_7104_n5490.n1 a_7104_n5490.t4 269.116
R7262 a_7104_n5490.t6 a_7104_n5490.n0 179.946
R7263 a_7104_n5490.n2 a_7104_n5490.n1 105.178
R7264 a_7104_n5490.n3 a_7104_n5490.t1 29.444
R7265 a_7104_n5490.n4 a_7104_n5490.t2 28.565
R7266 a_7104_n5490.t3 a_7104_n5490.n4 28.565
R7267 a_7104_n5490.n2 a_7104_n5490.t0 18.145
R7268 a_7104_n5490.n3 a_7104_n5490.n2 2.878
R7269 a_7104_n5490.n4 a_7104_n5490.n3 0.764
R7270 a_6818_n416.t0 a_6818_n416.t1 380.209
R7271 a_11469_n328.t0 a_11469_n328.t1 380.209
R7272 a_31118_n4120.t0 a_31118_n4120.t1 17.4
R7273 a_20252_n6197.t0 a_20252_n6197.t1 17.4
R7274 a_13661_378.n1 a_13661_378.t5 318.922
R7275 a_13661_378.n0 a_13661_378.t7 274.739
R7276 a_13661_378.n0 a_13661_378.t4 274.739
R7277 a_13661_378.n1 a_13661_378.t6 269.116
R7278 a_13661_378.t5 a_13661_378.n0 179.946
R7279 a_13661_378.n2 a_13661_378.n1 105.178
R7280 a_13661_378.n3 a_13661_378.t2 29.444
R7281 a_13661_378.n4 a_13661_378.t1 28.565
R7282 a_13661_378.t3 a_13661_378.n4 28.565
R7283 a_13661_378.n2 a_13661_378.t0 18.145
R7284 a_13661_378.n3 a_13661_378.n2 2.878
R7285 a_13661_378.n4 a_13661_378.n3 0.764
R7286 a_3244_n3141.t0 a_3244_n3141.t1 17.4
R7287 a_16464_n595.t0 a_16464_n595.t1 17.4
R7288 a_11699_n6198.t0 a_11699_n6198.t1 17.4
R7289 a_354_321.t0 a_354_321.t1 17.4
R7290 a_32485_n7683.t0 a_32485_n7683.t1 17.4
R7291 a_9809_n4793.t0 a_9809_n4793.t1 17.4
R7292 a_28877_n945.t0 a_28877_n945.t1 17.4
R7293 a_9804_n6397.t0 a_9804_n6397.t1 17.4
R7294 a_16455_2659.t0 a_16455_2659.t1 17.4
R7295 a_31116_3466.t0 a_31116_3466.t1 17.4
R7296 a_20257_n396.t0 a_20257_n396.t1 17.4
R7297 a_20264_n7831.t0 a_20264_n7831.t1 17.4
R7298 a_3261_n615.t0 a_3261_n615.t1 17.4
R7299 a_28882_4659.t0 a_28882_4659.t1 17.4
R7300 a_3258_n4791.t0 a_3258_n4791.t1 17.4
R7301 a_3253_n6395.t0 a_3253_n6395.t1 17.4
R7302 a_7061_n7824.t0 a_7061_n7824.t1 17.4
R7303 a_3266_989.t0 a_3266_989.t1 17.4
R7304 a_20021_n396.t0 a_20021_n396.t1 380.209
R7305 a_7026_4806.t0 a_7026_4806.t1 17.4
R7306 a_23089_n527.t0 a_23089_n527.t1 17.4
R7307 a_24740_n6196.t0 a_24740_n6196.t1 380.209
R7308 a_26874_n6196.t0 a_26874_n6196.t1 17.4
R7309 a_28945_n5935.t0 a_28945_n5935.t1 17.4
R7310 a_30882_n625.t0 a_30882_n625.t1 380.209
R7311 a_335_n2957.t0 a_335_n2957.t1 17.4
R7312 a_32485_n3335.t0 a_32485_n3335.t1 17.4
R7313 a_26646_n328.t0 a_26646_n328.t1 380.209
R7314 a_13615_n7819.t0 a_13615_n7819.t1 17.4
R7315 a_4920_n416.t0 a_4920_n416.t1 380.209
R7316 a_24984_n328.t0 a_24984_n328.t1 17.4
R7317 a_16464_n4792.t0 a_16464_n4792.t1 17.4
C0 A[2] B[2] 27.45fF
C1 A[3] B[3] 12.18fF
C2 B[1] B[0] 0.91fF
C3 VDD A[0] 7.69fF
C4 B[0] Y[6] 0.64fF
C5 A[0] Y[7] 0.05fF
C6 B[1] A[0] 1.78fF
C7 A[3] B[0] 3.66fF
C8 A[2] B[3] 1.27fF
C9 VDD Y[0] 1.01fF
C10 Y[0] Y[7] 0.00fF
C11 A[0] Y[6] 0.05fF
C12 VDD A[1] 3.51fF
C13 B[2] B[3] 1.54fF
C14 A[2] B[0] 5.07fF
C15 A[3] A[0] 1.09fF
C16 B[3] Y[5] 0.16fF
C17 Y[0] Y[6] 0.00fF
C18 B[2] B[0] 0.15fF
C19 B[1] A[1] 25.16fF
C20 VDD Y[2] 0.49fF
C21 A[2] A[0] 0.19fF
C22 A[3] A[1] 3.94fF
C23 B[3] B[0] 0.08fF
C24 VDD Y[7] 1.68fF
C25 B[2] A[0] 53.98fF
C26 A[0] Y[5] 0.14fF
C27 VDD B[1] 5.14fF
C28 B[3] A[0] 25.77fF
C29 A[2] A[1] 19.80fF
C30 VDD Y[6] 0.83fF
C31 Y[7] Y[6] 0.93fF
C32 VDD A[3] 3.19fF
C33 B[0] A[0] 58.43fF
C34 B[2] A[1] 1.69fF
C35 VDD Y[1] 0.49fF
C36 A[1] Y[5] 0.12fF
C37 B[1] A[3] 2.80fF
C38 VDD A[2] 2.67fF
C39 B[0] Y[0] 0.01fF
C40 VDD Y[4] 0.62fF
C41 B[3] A[1] 1.25fF
C42 B[1] A[2] 2.21fF
C43 VDD B[2] 8.32fF
C44 VDD Y[5] 1.26fF
C45 B[0] A[1] 1.35fF
C46 A[0] Y[0] 0.01fF
C47 B[2] Y[7] 0.13fF
C48 VDD B[3] 6.09fF
C49 B[1] B[2] 0.21fF
C50 A[3] A[2] 12.19fF
C51 B[2] Y[6] 0.08fF
C52 B[1] Y[5] 2.64fF
C53 VDD Y[3] 0.45fF
C54 A[0] A[1] 0.80fF
C55 VDD B[0] 2.62fF
C56 B[1] B[3] 27.63fF
C57 A[3] B[2] 18.53fF
C58 B[0] Y[7] 0.05fF
.ends

