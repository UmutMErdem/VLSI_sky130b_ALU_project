* NGSPICE file created from logic_unit_pex.ext - technology: sky130B

.subckt logic_unit B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] Y[0] Y[1] Y[2] Y[3]
+ Y[4] Y[5] Y[6] Y[7] VDD VSS opcode[0] opcode[1] A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7]
X0 VDD.t548 B[7].t0 a_20252_3694.t1 VDD.t547 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1 VDD.t1054 a_3891_1714.t4 a_3951_1740.t5 VDD.t1053 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2 a_3881_n3752.t3 A[1].t0 VDD.t739 VDD.t738 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 VSS.t154 A[0].t0 a_n25_n6671.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4 VDD.t326 A[7].t0 a_10615_3699.t2 VDD.t325 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 VDD.t714 opcode[0].t0 a_3392_1740.t2 VDD.t713 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6 a_12813_n7362.t11 a_12386_n6669.t4 a_12931_n7362.t7 VDD.t278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 a_3891_n1020.t2 a_4290_n3726.t8 VDD.t900 VDD.t899 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8 VDD.t546 B[7].t1 a_14881_n7360.t9 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X9 a_10852_3062.t0 A[7].t1 a_10615_3699.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10 VDD.t1216 a_3891_n1020.t4 a_3951_n994.t10 VDD.t1215 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 a_20054_n990.t0 opcode[1].t0 a_20290_n2323.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X12 a_4290_n3726.t6 a_2588_n7362.t8 a_3941_n3726.t8 VDD.t678 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X13 VDD.t763 a_747_1714.t4 a_807_1740.t11 VDD.t762 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X14 a_10217_n3722.t3 a_6725_n7362.t8 a_10566_n3722.t3 VDD.t404 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X15 VDD.t1059 opcode[1].t1 a_3392_n994.t2 VDD.t1058 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X16 a_21997_n6357.t2 A[7].t2 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X17 a_17916_3694.t5 A[5].t0 a_17798_3694.t1 VDD.t1036 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 a_7083_n990.t9 a_7023_n1016.t4 VDD.t414 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_10576_n990.t0 opcode[1].t2 a_10812_n2323.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X20 VDD.t902 A[5].t1 a_7669_3697.t3 VDD.t901 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X21 a_2588_n7362.t4 a_2043_n6669.t4 a_2588_n8094.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X22 VSS.t123 a_6725_n7362.t9 a_11038_n5055.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X23 a_7906_3060.t0 A[5].t2 a_7669_3697.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X24 a_7083_1744.t6 a_7023_1718.t4 VDD.t1074 VDD.t1073 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X25 VDD.t151 A[1].t1 a_3881_n3752.t2 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 VDD.t191 a_747_n1020.t4 a_807_n994.t11 VDD.t190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X27 Y[6].t2 a_20054_n990.t8 VDD.t403 VDD.t402 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 VDD.t166 a_10566_n3722.t8 a_10167_n1016.t2 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X29 VDD.t410 a_4290_n3726.t9 a_3891_n1020.t1 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X30 a_747_1714.t1 a_11952_3694.t5 VSS.t137 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X31 a_3951_1740.t6 a_3392_1740.t4 a_4300_1740.t4 VDD.t291 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X32 a_20579_n1475.t2 a_20054_1744.t8 VDD.t1048 VDD.t1047 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X33 a_15293_n7386.t2 B[7].t2 VDD.t544 VDD.t543 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X34 a_1382_n5059.t1 a_737_n3752.t4 VSS.t41 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X35 a_1156_1740.t5 a_897_3260.t4 a_807_1740.t4 VDD.t505 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X36 a_20526_n2323.t0 a_19146_n990.t4 a_20054_n990.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X37 VSS.t75 B[7].t3 a_20134_3694.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X38 a_10566_n3722.t2 a_6725_n7362.t10 a_10217_n3722.t2 VDD.t895 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 a_9668_n990.t2 opcode[1].t3 VDD.t1061 VDD.t1060 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X40 VSS.t144 opcode[1].t4 a_3392_n994.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X41 a_4951_n7390.t2 B[2].t0 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X42 a_3951_n994.t6 a_3392_n994.t4 a_4300_n994.t3 VDD.t457 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X43 a_22839_n3722.t7 a_21997_n6357.t4 VDD.t1031 VDD.t1030 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X44 a_9668_1744.t2 opcode[0].t1 VDD.t1148 VDD.t1147 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X45 a_1156_n994.t5 a_1681_n1479.t4 a_807_n994.t6 VDD.t589 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X46 a_2824_n8094.t0 A[1].t2 a_2588_n7362.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X47 VDD.t592 B[4].t0 a_16748_3696.t3 VDD.t591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X48 VSS.t68 a_14303_n1479.t4 a_14250_n2327.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X49 a_10167_n1016.t1 a_10566_n3722.t9 VDD.t168 VDD.t167 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X50 a_3891_n1020.t0 a_4290_n3726.t10 VDD.t412 VDD.t411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X51 a_13369_1714.t3 a_16630_3696.t5 VSS.t125 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X52 a_1146_n3726.t1 opcode[0].t2 a_1382_n5059.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X53 a_10227_n990.t2 opcode[1].t5 VDD.t1084 VDD.t1083 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X54 VSS.t142 a_20579_n1475.t4 a_20526_n2323.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X55 a_10227_1744.t5 opcode[0].t3 VDD.t1150 VDD.t1149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X56 Y[1].t3 a_4300_n994.t8 VSS.t165 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X57 a_15574_3694.t4 B[3].t0 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X58 VDD.t495 a_7432_n990.t8 Y[2].t2 VDD.t494 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X59 a_13238_3694.t2 A[1].t3 a_13120_3694.t0 VDD.t847 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X60 VDD.t368 a_7432_1744.t8 a_7957_n1475.t2 VDD.t367 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X61 VSS.t77 B[1].t0 a_2824_n8094.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X62 VDD.t560 B[1].t1 a_1755_3697.t6 VDD.t559 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 a_17158_n2327.t1 a_16513_n1020.t4 VSS.t27 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X64 VSS.t39 a_23723_n1475.t4 a_23670_n2323.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X65 Y[2].t1 a_7432_n990.t9 VDD.t520 VDD.t519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X66 a_7957_n1475.t1 a_7432_1744.t9 VDD.t370 VDD.t369 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X67 a_737_n3752.t3 A[0].t1 VSS.t153 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X68 VSS.t80 A[4].t0 a_8249_n6669.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X69 a_6221_3697.t2 B[4].t1 VDD.t594 VDD.t593 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X70 a_5291_3262.t2 a_4701_3699.t7 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X71 a_15293_n7386.t3 B[7].t4 VSS.t74 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X72 a_2470_n7362.t6 A[1].t4 VDD.t140 VDD.t139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X73 a_9757_3262.t2 a_9167_3699.t7 VDD.t604 VDD.t603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X74 VSS.t15 B[3].t1 a_15456_3694.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X75 VDD.t1086 opcode[1].t6 a_22290_n990.t2 VDD.t1085 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X76 VDD.t364 a_13120_3694.t5 a_3891_1714.t0 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X77 VDD.t581 a_15456_3694.t5 a_10167_1718.t2 VDD.t580 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X78 a_16014_1740.t2 opcode[0].t4 VDD.t240 VDD.t239 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X79 a_21997_n6357.t1 A[7].t3 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X80 a_4762_n5059.t1 a_3382_n3726.t4 a_4290_n3726.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X81 VDD.t242 opcode[0].t5 a_22290_1744.t2 VDD.t241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X82 a_10227_n990.t5 a_10167_n1016.t4 VDD.t733 VDD.t732 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X83 a_10227_1744.t8 a_10167_1718.t4 VDD.t586 VDD.t585 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X84 a_16014_n994.t2 opcode[1].t7 VDD.t1078 VDD.t1077 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X85 a_7013_n3748.t3 A[2].t0 VSS.t13 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X86 VDD.t244 opcode[0].t6 a_13429_1740.t2 VDD.t243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X87 a_7083_n990.t8 a_7023_n1016.t5 VDD.t416 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 a_13167_n8094.t1 A[6].t0 a_12931_n7362.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X89 a_7083_1744.t5 a_7023_1718.t5 VDD.t1076 VDD.t1075 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X90 VSS.t23 opcode[0].t7 a_16004_n3726.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X91 VDD.t162 opcode[0].t8 a_16004_n3726.t2 VDD.t161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X92 Y[6].t1 a_20054_n990.t9 VDD.t673 VDD.t672 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X93 a_807_1740.t7 a_248_1740.t4 a_1156_1740.t6 VDD.t937 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X94 VDD.t628 a_13778_1740.t8 a_14303_n1479.t0 VDD.t627 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X95 VSS.t150 a_8259_3260.t4 a_17394_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X96 VDD.t1080 opcode[1].t8 a_13429_n994.t5 VDD.t1079 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X97 VSS.t90 a_2588_n7362.t9 a_4762_n5059.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X98 VDD.t164 opcode[0].t9 a_248_1740.t2 VDD.t163 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X99 a_22849_n990.t6 a_22290_n990.t4 a_23198_n990.t3 VDD.t746 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X100 a_14881_n7360.t0 a_14454_n6667.t4 a_14999_n7360.t6 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X101 a_11038_n5055.t1 a_9658_n3722.t4 a_10566_n3722.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X102 a_20579_n1475.t1 a_20054_1744.t9 VDD.t1050 VDD.t1049 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X103 a_4825_n1479.t3 a_4300_1740.t8 VSS.t24 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X104 VSS.t133 a_5291_3262.t4 a_11048_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X105 a_13369_n1020.t3 a_13768_n3726.t8 VSS.t21 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X106 a_1156_1740.t4 a_897_3260.t5 a_807_1740.t5 VDD.t851 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X107 a_22849_1744.t9 a_22290_1744.t4 a_23198_1744.t5 VDD.t897 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X108 VDD.t652 B[5].t0 a_17916_3694.t0 VDD.t651 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X109 a_807_n994.t4 a_248_n994.t4 a_1156_n994.t1 VDD.t313 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X110 VDD.t805 a_13778_n994.t8 Y[4].t2 VDD.t804 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X111 VDD.t940 A[6].t1 a_19635_n3748.t2 VDD.t939 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X112 VDD.t122 A[2].t1 a_4112_n6671.t2 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X113 VDD.t1082 opcode[1].t9 a_248_n994.t2 VDD.t1081 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X114 VSS.t10 B[6].t0 a_13167_n8094.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X115 a_10167_n1016.t0 a_10566_n3722.t10 VDD.t170 VDD.t169 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X116 a_1156_n994.t4 a_1681_n1479.t5 a_807_n994.t7 VDD.t590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X117 a_402_n7364.t7 a_814_n7390.t4 a_520_n7364.t6 VDD.t812 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X118 a_16513_n1020.t2 a_16912_n3726.t8 VSS.t168 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X119 a_14406_3692.t5 A[2].t2 a_14288_3692.t3 VDD.t380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X120 a_6961_n8094.t1 A[3].t0 a_6725_n7362.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X121 VDD.t654 B[5].t1 a_11156_n7386.t2 VDD.t653 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X122 a_7422_n3722.t2 a_4657_n7364.t8 a_7073_n3722.t5 VDD.t723 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X123 a_20290_411.t1 a_19230_3112.t4 VSS.t109 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X124 a_3843_3262.t2 a_3253_3699.t7 VDD.t610 VDD.t609 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X125 a_14999_n7360.t5 a_14454_n6667.t5 a_14881_n7360.t1 VDD.t220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X126 VSS.t4 opcode[0].t10 a_238_n3726.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X127 VDD.t875 a_13369_1714.t4 a_13429_1740.t11 VDD.t874 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X128 a_19635_n3748.t1 A[6].t2 VDD.t624 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X129 a_12931_n8094.t0 a_13225_n7388.t4 VSS.t162 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X130 a_7083_n990.t10 a_7957_n1475.t4 a_7432_n990.t5 VDD.t565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X131 a_737_n3752.t2 A[0].t2 VDD.t681 VDD.t680 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X132 VSS.t172 opcode[1].t10 a_19146_n990.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X133 a_520_n7364.t5 a_814_n7390.t5 a_402_n7364.t6 VDD.t813 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X134 a_12070_3694.t4 A[0].t3 a_11952_3694.t1 VDD.t331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X135 a_11156_n7386.t1 B[5].t2 VDD.t771 VDD.t770 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X136 a_7073_n3722.t4 a_4657_n7364.t9 a_7422_n3722.t1 VDD.t724 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X137 a_7083_1744.t7 a_3843_3262.t4 a_7432_1744.t2 VDD.t477 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X138 VDD.t224 a_13369_n1020.t4 a_13429_n994.t0 VDD.t223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X139 a_13419_n3726.t6 opcode[0].t11 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X140 a_897_3260.t1 a_307_3697.t7 VDD.t646 VDD.t645 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X141 a_4701_3699.t6 A[3].t1 VDD.t959 VDD.t958 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X142 VSS.t173 opcode[1].t11 a_9668_n990.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X143 a_14881_n7360.t10 a_15293_n7386.t4 a_14999_n7360.t2 VDD.t891 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X144 a_19645_n1016.t2 a_20044_n3722.t8 VDD.t831 VDD.t830 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X145 VSS.t5 opcode[0].t12 a_22290_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X146 Y[0].t3 a_1156_n994.t8 VSS.t57 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X147 a_2588_n7362.t5 a_2043_n6669.t5 a_2470_n7362.t2 VDD.t1069 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X148 a_19695_n3722.t8 a_19136_n3722.t4 a_20044_n3722.t6 VDD.t760 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X149 a_6811_3260.t2 a_6221_3697.t7 VDD.t500 VDD.t499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X150 a_20252_3694.t0 A[7].t4 a_20134_3694.t3 VDD.t203 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X151 a_23188_n3722.t3 a_14999_n7360.t8 a_22839_n3722.t10 VDD.t838 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X152 VDD.t626 A[6].t3 a_12813_n7362.t5 VDD.t625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X153 VDD.t388 A[0].t4 a_737_n3752.t1 VDD.t387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X154 a_6607_n7362.t11 A[3].t2 VDD.t312 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X155 VSS.t78 B[1].t2 a_13120_3694.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X156 a_19705_n990.t11 a_19645_n1016.t4 VDD.t753 VDD.t752 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X157 a_7422_n3722.t0 a_4657_n7364.t10 a_7073_n3722.t3 VDD.t855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X158 Y[3].t3 a_10576_n990.t8 VSS.t175 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X159 a_19705_1744.t5 a_19230_3112.t5 VDD.t841 VDD.t840 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X160 a_2470_n7362.t1 a_2043_n6669.t6 a_2588_n7362.t6 VDD.t1070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X161 a_20044_n3722.t7 a_19136_n3722.t5 a_19695_n3722.t7 VDD.t761 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X162 a_22839_n3722.t11 a_14999_n7360.t9 a_23188_n3722.t2 VDD.t839 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X163 a_11101_n1475.t3 a_10576_1744.t8 VSS.t114 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X164 a_10227_n990.t4 a_10167_n1016.t5 VDD.t735 VDD.t734 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X165 VSS.t44 A[3].t3 a_6180_n6669.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X166 a_12813_n7362.t1 A[6].t4 VDD.t262 VDD.t261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X167 a_13778_1740.t2 a_6811_3260.t4 a_13429_1740.t4 VDD.t800 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X168 VDD.t1259 opcode[1].t12 a_6524_n990.t2 VDD.t1258 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X169 VDD.t246 a_7422_n3722.t8 a_7023_n1016.t0 VDD.t245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X170 a_10227_1744.t6 a_10167_1718.t5 VDD.t502 VDD.t501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X171 a_11205_3262.t2 a_10615_3699.t7 VDD.t1193 VDD.t1192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X172 a_807_1740.t2 opcode[0].t13 VDD.t302 VDD.t301 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X173 VDD.t304 opcode[0].t14 a_6524_1744.t2 VDD.t303 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X174 VDD.t809 A[3].t4 a_6607_n7362.t10 VDD.t808 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X175 a_16922_1740.t3 a_16014_1740.t4 a_16573_1740.t2 VDD.t450 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X176 a_13778_n994.t5 a_14303_n1479.t5 a_13429_n994.t9 VDD.t514 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X177 a_20054_n990.t5 a_20579_n1475.t5 a_19705_n990.t8 VDD.t1062 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X178 a_16922_1740.t7 a_8259_3260.t5 a_16573_1740.t10 VDD.t1126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X179 a_20054_1744.t2 a_9757_3262.t4 a_19705_1744.t11 VDD.t578 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X180 a_16912_n3726.t6 a_10862_n7360.t8 a_16563_n3726.t9 VDD.t853 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X181 VDD.t773 B[5].t3 a_17916_3694.t2 VDD.t772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X182 a_807_n994.t2 opcode[1].t13 VDD.t1100 VDD.t1099 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X183 a_8259_3260.t2 a_7669_3697.t7 VDD.t1067 VDD.t1066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X184 a_8794_n8094.t0 a_9088_n7388.t4 VSS.t55 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X185 a_14999_n7360.t4 a_14454_n6667.t6 a_14881_n7360.t2 VDD.t221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X186 a_2588_n7362.t3 a_2043_n6669.t7 a_2470_n7362.t0 VDD.t1068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X187 VSS.t43 opcode[0].t15 a_248_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X188 a_16922_n994.t3 a_16014_n994.t4 a_16573_n994.t1 VDD.t250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X189 a_23198_n990.t7 a_23723_n1475.t5 a_22849_n990.t9 VDD.t743 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X190 a_10862_n7360.t4 a_10317_n6667.t4 a_10744_n7360.t11 VDD.t881 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X191 VDD.t104 B[6].t1 a_12813_n7362.t0 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X192 a_16922_n994.t5 a_17447_n1479.t4 a_16573_n994.t6 VDD.t460 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X193 a_19084_3696.t5 A[6].t5 a_18966_3696.t4 VDD.t263 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X194 a_7073_n3722.t9 a_6514_n3722.t4 a_7422_n3722.t4 VDD.t185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X195 a_23198_1744.t6 a_11205_3262.t4 a_22849_1744.t10 VDD.t1155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X196 a_1392_n2327.t1 a_747_n1020.t5 VSS.t28 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X197 a_4825_n1479.t2 a_4300_1740.t9 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X198 VDD.t1238 a_16912_n3726.t9 a_16513_n1020.t3 VDD.t1237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X199 a_10576_n990.t6 a_9668_n990.t4 a_10227_n990.t8 VDD.t990 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X200 Y[2].t3 a_7432_n990.t10 VSS.t70 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X201 a_10576_1744.t2 a_9668_1744.t4 a_10227_1744.t0 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X202 a_17447_n1479.t3 a_16922_1740.t8 VSS.t99 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X203 VDD.t974 a_18966_3696.t5 a_19230_3112.t2 VDD.t973 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X204 VDD.t1102 opcode[1].t14 a_7083_n990.t2 VDD.t1101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X205 a_10227_n990.t11 a_11101_n1475.t4 a_10576_n990.t7 VDD.t1158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X206 Y[1].t2 a_4300_n994.t9 VDD.t702 VDD.t701 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X207 a_2470_n7362.t7 a_2882_n7388.t4 a_2588_n7362.t2 VDD.t725 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X208 a_7422_n3722.t3 opcode[0].t16 a_7658_n5055.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X209 a_16513_1714.t3 a_17798_3694.t5 VSS.t141 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X210 VDD.t919 opcode[0].t17 a_7083_1744.t2 VDD.t918 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X211 a_10227_1744.t11 a_5291_3262.t5 a_10576_1744.t7 VDD.t970 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X212 VDD.t205 A[7].t5 a_14454_n6667.t2 VDD.t204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X213 a_1755_3697.t3 A[1].t5 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X214 a_10744_n7360.t10 a_10317_n6667.t5 a_10862_n7360.t5 VDD.t1125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X215 VDD.t904 A[5].t3 a_10317_n6667.t2 VDD.t903 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X216 a_12070_3694.t3 A[0].t5 a_11952_3694.t3 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X217 a_797_n3726.t2 a_520_n7364.t8 a_1146_n3726.t4 VDD.t926 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X218 a_10157_n3748.t2 A[3].t5 VDD.t811 VDD.t810 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X219 a_814_n7390.t3 B[0].t0 VSS.t169 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X220 VSS.t124 opcode[0].t18 a_16014_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X221 a_1156_n994.t0 opcode[1].t15 a_1392_n2327.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X222 a_4701_3699.t5 A[3].t6 VDD.t479 VDD.t478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X223 VDD.t1010 opcode[0].t19 a_12870_1740.t2 VDD.t1009 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X224 a_23424_n5055.t1 a_21997_n6357.t5 VSS.t140 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X225 VDD.t1012 opcode[0].t20 a_22839_n3722.t4 VDD.t1011 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X226 VSS.t16 B[3].t2 a_4938_3062.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X227 a_7013_n3748.t2 A[2].t3 VDD.t382 VDD.t381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X228 a_13768_n3726.t2 opcode[0].t21 a_14004_n5059.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X229 VDD.t869 a_16630_3696.t6 a_13369_1714.t2 VDD.t868 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X230 a_8676_n7362.t8 A[4].t1 VDD.t573 VDD.t572 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X231 VDD.t398 A[6].t6 a_9167_3699.t1 VDD.t397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X232 VDD.t1104 opcode[1].t16 a_12870_n994.t2 VDD.t1103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X233 a_7894_n5055.t1 a_6514_n3722.t5 a_7422_n3722.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X234 a_10217_n3722.t7 a_10157_n3748.t4 VDD.t741 VDD.t740 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X235 a_9404_3062.t1 A[6].t7 a_9167_3699.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X236 VDD.t863 opcode[0].t22 a_16014_1740.t1 VDD.t862 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X237 a_21997_n6357.t3 A[7].t6 VSS.t31 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X238 a_16912_n3726.t0 opcode[0].t23 a_17148_n5059.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X239 a_1146_n3726.t5 a_520_n7364.t9 a_797_n3726.t1 VDD.t927 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X240 a_14999_n7360.t7 a_14454_n6667.t7 a_14999_n8092.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X241 a_12813_n7362.t4 A[6].t8 VDD.t620 VDD.t619 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X242 VSS.t2 B[2].t1 a_14288_3692.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X243 VSS.t60 a_2345_3260.t4 a_4772_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X244 a_13768_n3726.t5 a_8794_n7362.t8 a_13419_n3726.t9 VDD.t730 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X245 a_12931_n7362.t5 a_12386_n6669.t5 a_12813_n7362.t10 VDD.t279 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X246 a_23188_n3722.t5 opcode[0].t24 a_23424_n5055.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X247 VDD.t1106 opcode[1].t17 a_16014_n994.t1 VDD.t1105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X248 a_13359_n3752.t3 A[4].t2 VSS.t81 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X249 VDD.t1163 a_14288_3692.t5 a_7023_1718.t3 VDD.t1162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X250 a_14240_n5059.t0 a_12860_n3726.t4 a_13768_n3726.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X251 a_3843_3262.t3 a_3253_3699.t8 VSS.t91 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X252 VDD.t596 B[4].t2 a_8676_n7362.t5 VDD.t595 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X253 a_13778_1740.t3 a_6811_3260.t5 a_13429_1740.t5 VDD.t801 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X254 a_19146_n990.t2 opcode[1].t18 VDD.t1108 VDD.t1107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X255 a_4772_n2327.t0 a_3392_n994.t5 a_4300_n994.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X256 VDD.t656 a_3881_n3752.t4 a_3941_n3726.t11 VDD.t655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X257 VDD.t1094 B[5].t4 a_10744_n7360.t5 VDD.t1093 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X258 VSS.t116 a_4657_n7364.t11 a_7894_n5055.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X259 VDD.t1121 a_10157_n3748.t5 a_10217_n3722.t11 VDD.t1120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X260 VSS.t86 A[6].t9 a_12386_n6669.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X261 a_11205_3262.t1 a_10615_3699.t8 VDD.t622 VDD.t621 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X262 VDD.t472 opcode[0].t25 a_13429_1740.t1 VDD.t471 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X263 a_19146_1744.t2 opcode[0].t26 VDD.t474 VDD.t473 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X264 a_19705_n990.t5 opcode[1].t19 VDD.t1261 VDD.t1260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X265 a_17384_n5059.t0 a_16004_n3726.t4 a_16912_n3726.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X266 a_19705_1744.t2 opcode[0].t27 VDD.t476 VDD.t475 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X267 a_11048_411.t0 a_9668_1744.t5 a_10576_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X268 a_15235_n8092.t0 A[7].t7 a_14999_n7360.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X269 a_13778_n994.t4 a_14303_n1479.t6 a_13429_n994.t8 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X270 a_13419_n3726.t8 a_8794_n7362.t9 a_13768_n3726.t4 VDD.t330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X271 a_17394_407.t0 a_16014_1740.t5 a_16922_1740.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X272 a_12813_n7362.t8 a_13225_n7388.t5 a_12931_n7362.t3 VDD.t1166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X273 VDD.t90 a_20134_3694.t5 a_20398_3112.t2 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X274 VDD.t1263 opcode[1].t20 a_13429_n994.t4 VDD.t1262 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X275 a_3253_3699.t5 A[2].t4 VDD.t1172 VDD.t1171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X276 a_22849_n990.t3 opcode[1].t21 VDD.t1265 VDD.t1264 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X277 VDD.t437 opcode[0].t28 a_16573_1740.t5 VDD.t436 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X278 VSS.t47 B[2].t2 a_3490_3062.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X279 a_16630_3696.t0 A[4].t3 a_16748_3696.t0 VDD.t496 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X280 a_22849_1744.t4 opcode[0].t29 VDD.t439 VDD.t438 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X281 a_6725_n7362.t4 a_6180_n6669.t4 a_6607_n7362.t7 VDD.t905 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X282 a_8676_n7362.t4 B[4].t3 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X283 a_402_n7364.t11 A[0].t6 VDD.t608 VDD.t607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X284 VSS.t33 a_4825_n1479.t4 a_4772_n2327.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X285 VSS.t69 B[3].t3 a_6961_n8094.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X286 a_16563_n3726.t8 a_10862_n7360.t9 a_16912_n3726.t7 VDD.t854 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X287 a_10217_n3722.t8 a_10157_n3748.t6 VDD.t883 VDD.t882 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X288 a_1681_n1479.t2 a_1156_1740.t8 VDD.t815 VDD.t814 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X289 VDD.t358 B[2].t3 a_3253_3699.t2 VDD.t357 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X290 a_19084_3696.t2 B[6].t2 VDD.t843 VDD.t842 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X291 Y[7].t2 a_23198_n990.t8 VDD.t757 VDD.t756 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X292 a_11048_n2323.t0 a_9668_n990.t5 a_10576_n990.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X293 VDD.t1038 opcode[1].t22 a_16573_n994.t5 VDD.t1037 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X294 a_814_n7390.t1 B[0].t1 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X295 VSS.t113 a_10862_n7360.t10 a_17384_n5059.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X296 a_23723_n1475.t2 a_23198_1744.t8 VDD.t1255 VDD.t1254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X297 VDD.t1040 opcode[1].t23 a_10227_n990.t1 VDD.t1039 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X298 VSS.t73 B[7].t5 a_15235_n8092.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X299 a_14406_3692.t2 B[2].t4 VDD.t360 VDD.t359 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X300 a_4300_1740.t6 a_2345_3260.t5 a_3951_1740.t8 VDD.t791 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X301 a_3881_n3752.t1 A[1].t6 VDD.t1144 VDD.t1143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X302 Y[0].t2 a_1156_n994.t9 VDD.t443 VDD.t442 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X303 a_12931_n7362.t0 a_13225_n7388.t6 a_12813_n7362.t2 VDD.t453 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X304 VDD.t986 a_18966_3696.t6 a_19230_3112.t3 VDD.t985 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X305 VDD.t441 opcode[0].t30 a_10227_1744.t4 VDD.t440 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X306 a_238_n3726.t2 opcode[0].t31 VDD.t1160 VDD.t1159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X307 a_3941_n3726.t5 a_3382_n3726.t5 a_4290_n3726.t5 VDD.t587 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X308 a_5291_3262.t3 a_4701_3699.t8 VSS.t9 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X309 VSS.t158 opcode[0].t32 a_6514_n3722.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X310 a_18966_3696.t2 A[6].t10 VSS.t126 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X311 a_4300_n994.t4 a_4825_n1479.t5 a_3951_n994.t3 VDD.t253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X312 VDD.t180 B[4].t4 a_8676_n7362.t3 VDD.t179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X313 VDD.t211 A[0].t7 a_402_n7364.t10 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X314 a_15456_3694.t4 A[3].t7 a_15574_3694.t5 VDD.t480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X315 a_6725_n8094.t0 a_7019_n7388.t4 VSS.t96 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X316 VDD.t1056 A[0].t8 a_307_3697.t3 VDD.t1055 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X317 VSS.t159 opcode[0].t33 a_12870_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X318 a_2588_n8094.t1 a_2882_n7388.t5 VSS.t103 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X319 a_544_3060.t1 A[0].t9 a_307_3697.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X320 a_3881_n3752.t0 A[1].t7 VSS.t64 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X321 VDD.t1146 B[0].t2 a_814_n7390.t2 VDD.t1145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X322 a_1755_3697.t2 A[1].t8 VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X323 VSS.t110 B[6].t3 a_18966_3696.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X324 VDD.t498 A[4].t4 a_6221_3697.t5 VDD.t497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X325 a_12813_n7362.t3 a_13225_n7388.t7 a_12931_n7362.t1 VDD.t454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X326 a_6458_3060.t1 A[4].t5 a_6221_3697.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X327 a_22849_n990.t11 a_22789_n1016.t4 VDD.t890 VDD.t889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X328 VDD.t1233 opcode[0].t34 a_238_n3726.t1 VDD.t1232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X329 a_4290_n3726.t2 a_3382_n3726.t6 a_3941_n3726.t3 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X330 a_22849_1744.t1 a_20398_3112.t4 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X331 a_13359_n3752.t2 A[4].t6 VDD.t567 VDD.t566 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X332 a_1618_n5059.t1 a_238_n3726.t4 a_1146_n3726.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X333 a_402_n7364.t9 A[0].t10 VDD.t213 VDD.t212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X334 a_14004_n5059.t0 a_13359_n3752.t4 VSS.t19 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X335 a_19136_n3722.t2 opcode[0].t35 VDD.t1235 VDD.t1234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X336 a_4300_1740.t0 opcode[0].t36 a_4536_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X337 a_7957_n1475.t3 a_7432_1744.t10 VSS.t48 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X338 VDD.t516 B[3].t4 a_4701_3699.t4 VDD.t515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X339 a_20252_3694.t2 B[7].t6 VDD.t542 VDD.t541 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X340 a_747_n1020.t3 a_1146_n3726.t8 VDD.t992 VDD.t991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X341 VDD.t569 A[4].t7 a_8676_n7362.t7 VDD.t568 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X342 a_814_n7390.t0 B[0].t3 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X343 a_10615_3699.t1 A[7].t8 VDD.t980 VDD.t979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X344 a_3392_1740.t1 opcode[0].t37 VDD.t803 VDD.t802 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X345 a_13225_n7388.t2 B[6].t4 VDD.t1168 VDD.t1167 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X346 VSS.t100 opcode[0].t38 a_22280_n3722.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X347 VSS.t101 opcode[0].t39 a_6524_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X348 a_807_1740.t10 a_747_1714.t5 VDD.t765 VDD.t764 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X349 a_3941_n3726.t4 a_3382_n3726.t7 a_4290_n3726.t3 VDD.t430 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X350 a_3392_n994.t1 opcode[1].t24 VDD.t1042 VDD.t1041 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X351 VDD.t571 A[4].t8 a_13359_n3752.t1 VDD.t570 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X352 VSS.t18 a_520_n7364.t10 a_1618_n5059.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X353 a_16563_n3726.t5 a_16004_n3726.t5 a_16912_n3726.t4 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X354 a_7669_3697.t2 A[5].t4 VDD.t932 VDD.t931 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X355 VDD.t143 B[0].t4 a_402_n7364.t0 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X356 VDD.t664 opcode[0].t40 a_19136_n3722.t1 VDD.t663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X357 a_17158_407.t1 a_16513_1714.t4 VSS.t119 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X358 a_14250_407.t1 a_12870_1740.t4 a_13778_1740.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X359 a_807_n994.t10 a_747_n1020.t6 VDD.t193 VDD.t192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X360 VDD.t1240 opcode[1].t25 a_6524_n990.t1 VDD.t1239 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X361 Y[5].t3 a_16922_n994.t8 VSS.t151 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X362 VDD.t124 a_1146_n3726.t9 a_747_n1020.t0 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X363 a_8794_n7362.t2 a_9088_n7388.t5 a_8676_n7362.t2 VDD.t1212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X364 VDD.t666 opcode[0].t41 a_6524_1744.t1 VDD.t665 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X365 VDD.t1170 B[6].t5 a_13225_n7388.t1 VDD.t1169 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X366 VDD.t1096 B[5].t5 a_7669_3697.t4 VDD.t1095 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X367 VSS.t20 B[0].t5 a_11952_3694.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X368 VDD.t113 a_20134_3694.t6 a_20398_3112.t1 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X369 a_20134_3694.t0 A[7].t9 VSS.t136 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X370 VSS.t170 opcode[1].t26 a_248_n994.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X371 a_10862_n7360.t7 a_10317_n6667.t6 a_10862_n8092.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X372 VDD.t1242 opcode[1].t27 a_9668_n990.t1 VDD.t1241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X373 a_7669_3697.t6 B[5].t6 VDD.t1267 VDD.t1266 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X374 VSS.t115 a_897_3260.t6 a_1628_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X375 VDD.t518 B[3].t5 a_6607_n7362.t6 VDD.t517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X376 a_3951_1740.t9 a_3392_1740.t5 a_4300_1740.t3 VDD.t910 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X377 VDD.t668 opcode[0].t42 a_9668_1744.t1 VDD.t667 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X378 VDD.t799 a_16922_1740.t9 a_17447_n1479.t2 VDD.t798 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X379 a_19635_n3748.t3 A[6].t11 VSS.t127 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X380 a_23198_n990.t6 a_23723_n1475.t6 a_22849_n990.t8 VDD.t744 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X381 a_7073_n3722.t2 a_7013_n3748.t4 VDD.t1199 VDD.t1198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X382 a_747_n1020.t1 a_1146_n3726.t10 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X383 a_2345_3260.t3 a_1755_3697.t7 VSS.t166 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X384 a_7668_n2323.t1 a_7023_n1016.t6 VSS.t52 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X385 a_9088_n7388.t3 B[4].t5 VSS.t26 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X386 a_8676_n7362.t1 a_9088_n7388.t6 a_8794_n7362.t1 VDD.t1035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X387 a_23198_1744.t7 a_11205_3262.t5 a_22849_1744.t11 VDD.t1156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X388 VSS.t25 B[4].t6 a_16630_3696.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X389 a_3951_n994.t0 a_3392_n994.t6 a_4300_n994.t2 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X390 VDD.t1129 a_16922_n994.t9 Y[5].t2 VDD.t1128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X391 a_4300_1740.t7 a_2345_3260.t6 a_3951_1740.t11 VDD.t1057 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X392 a_10862_n7360.t6 a_10317_n6667.t7 a_10744_n7360.t9 VDD.t1127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X393 VDD.t1024 a_17798_3694.t6 a_16513_1714.t2 VDD.t1023 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X394 VDD.t600 B[3].t6 a_15574_3694.t3 VDD.t599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X395 a_4657_n7364.t1 a_4112_n6671.t4 a_4539_n7364.t8 VDD.t371 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X396 a_6607_n7362.t5 B[3].t7 VDD.t602 VDD.t601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X397 a_4112_n6671.t1 A[2].t5 VDD.t1174 VDD.t1173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X398 a_4300_n994.t6 a_4825_n1479.t6 a_3951_n994.t4 VDD.t392 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X399 a_9088_n7388.t2 B[4].t7 VDD.t173 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X400 VDD.t1201 a_7013_n3748.t5 a_7073_n3722.t1 VDD.t1200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X401 VDD.t27 B[0].t6 a_307_3697.t0 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X402 a_10576_1744.t4 opcode[0].t43 a_10812_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X403 a_7432_n990.t0 opcode[1].t28 a_7668_n2323.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X404 a_13238_3694.t3 B[1].t3 VDD.t554 VDD.t553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X405 Y[3].t2 a_10576_n990.t9 VDD.t1269 VDD.t1268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X406 VDD.t556 B[1].t4 a_1755_3697.t5 VDD.t555 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X407 VDD.t175 B[4].t8 a_6221_3697.t1 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X408 VDD.t583 a_15456_3694.t6 a_10167_1718.t1 VDD.t582 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X409 a_11101_n1475.t2 a_10576_1744.t9 VDD.t850 VDD.t849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X410 a_10744_n7360.t2 a_11156_n7386.t4 a_10862_n7360.t1 VDD.t396 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X411 VDD.t1208 opcode[0].t44 a_22280_n3722.t2 VDD.t1207 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X412 VDD.t459 a_16513_1714.t5 a_16573_1740.t7 VDD.t458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X413 a_12860_n3726.t2 opcode[0].t45 VDD.t1210 VDD.t1209 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X414 VDD.t132 a_4701_3699.t9 a_5291_3262.t1 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X415 a_23434_n2323.t0 a_22789_n1016.t5 VSS.t98 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X416 a_737_n3752.t0 A[0].t11 VDD.t288 VDD.t287 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X417 a_15456_3694.t2 A[3].t8 VSS.t49 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X418 a_22290_n990.t1 opcode[1].t29 VDD.t885 VDD.t884 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X419 a_10217_n3722.t9 a_9658_n3722.t5 a_10566_n3722.t5 VDD.t929 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X420 VDD.t708 opcode[0].t46 a_6514_n3722.t2 VDD.t707 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X421 a_3891_1714.t1 a_13120_3694.t6 VDD.t820 VDD.t819 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X422 a_10167_1718.t0 a_15456_3694.t7 VDD.t1250 VDD.t1249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X423 VDD.t710 opcode[0].t47 a_16014_1740.t0 VDD.t709 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X424 a_13778_n994.t1 opcode[1].t30 a_14014_n2327.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X425 VDD.t749 A[6].t12 a_12386_n6669.t1 VDD.t748 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X426 VDD.t489 B[4].t9 a_9088_n7388.t1 VDD.t488 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X427 a_22290_1744.t1 opcode[0].t48 VDD.t712 VDD.t711 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X428 a_4772_407.t0 a_3392_1740.t6 a_4300_1740.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X429 VDD.t182 a_16513_n1020.t5 a_16573_n994.t9 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X430 a_7904_n2323.t1 a_6524_n990.t4 a_7432_n990.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X431 a_14881_n7360.t5 A[7].t10 VDD.t1019 VDD.t1018 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X432 VDD.t976 opcode[1].t31 a_16014_n994.t0 VDD.t975 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X433 a_13429_1740.t0 opcode[0].t49 VDD.t234 VDD.t233 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X434 a_16922_n994.t4 opcode[1].t32 a_17158_n2327.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X435 a_10862_n7360.t2 a_11156_n7386.t5 a_10744_n7360.t1 VDD.t455 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X436 a_22280_n3722.t1 opcode[0].t50 VDD.t236 VDD.t235 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X437 VSS.t72 B[7].t7 a_10852_3062.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X438 VDD.t238 opcode[0].t51 a_12860_n3726.t1 VDD.t237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X439 VSS.t22 opcode[0].t52 a_12860_n3726.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X440 a_7023_n1016.t1 a_7422_n3722.t9 VDD.t248 VDD.t247 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X441 a_23198_n990.t0 opcode[1].t33 a_23434_n2323.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X442 a_14250_n2327.t0 a_12870_n994.t4 a_13778_n994.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X443 a_10566_n3722.t6 a_9658_n3722.t6 a_10217_n3722.t10 VDD.t930 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X444 a_248_1740.t1 opcode[0].t53 VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X445 a_1156_1740.t7 a_248_1740.t5 a_807_1740.t8 VDD.t938 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X446 a_14303_n1479.t1 a_13778_1740.t9 VDD.t630 VDD.t629 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X447 a_13429_n994.t3 opcode[1].t34 VDD.t775 VDD.t774 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X448 a_12386_n6669.t2 A[6].t13 VDD.t751 VDD.t750 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X449 VSS.t63 A[1].t9 a_2043_n6669.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X450 a_9088_n7388.t0 B[4].t10 VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X451 a_807_1740.t6 a_897_3260.t7 a_1156_1740.t3 VDD.t852 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X452 a_16573_1740.t1 a_16014_1740.t6 a_16922_1740.t2 VDD.t893 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X453 a_1681_n1479.t3 a_1156_1740.t9 VSS.t104 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X454 a_16922_1740.t4 opcode[0].t54 a_17158_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X455 VSS.t79 a_7957_n1475.t5 a_7904_n2323.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X456 a_6607_n7362.t8 a_7019_n7388.t5 a_6725_n7362.t7 VDD.t982 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X457 VDD.t612 A[1].t10 a_2470_n7362.t5 VDD.t611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X458 a_20398_3112.t3 a_20134_3694.t7 VSS.t12 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X459 a_1156_n994.t2 a_248_n994.t5 a_807_n994.t5 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X460 a_248_n994.t1 opcode[1].t35 VDD.t777 VDD.t776 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X461 Y[4].t1 a_13778_n994.t9 VDD.t807 VDD.t806 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X462 a_3253_3699.t4 A[2].t6 VDD.t390 VDD.t389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X463 a_22849_n990.t5 a_22290_n990.t5 a_23198_n990.t2 VDD.t747 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X464 a_17394_n2327.t0 a_16014_n994.t5 a_16922_n994.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X465 a_10744_n7360.t0 a_11156_n7386.t6 a_10862_n7360.t0 VDD.t456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X466 VDD.t33 opcode[0].t55 a_22280_n3722.t0 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X467 a_897_3260.t2 a_307_3697.t8 VSS.t128 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X468 a_807_n994.t3 a_1681_n1479.t6 a_1156_n994.t3 VDD.t300 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X469 a_16573_n994.t0 a_16014_n994.t6 a_16922_n994.t2 VDD.t316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X470 a_19695_n3722.t6 a_19136_n3722.t6 a_20044_n3722.t1 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X471 a_22849_1744.t8 a_22290_1744.t5 a_23198_1744.t4 VDD.t898 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X472 a_19645_n1016.t3 a_20044_n3722.t9 VSS.t108 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X473 a_10217_n3722.t0 a_9658_n3722.t7 a_10566_n3722.t0 VDD.t171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X474 VDD.t696 a_3253_3699.t9 a_3843_3262.t1 VDD.t695 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X475 VDD.t1205 A[6].t14 a_12386_n6669.t3 VDD.t1204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X476 a_3951_1740.t2 opcode[0].t56 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X477 a_6607_n7362.t9 A[3].t9 VDD.t379 VDD.t378 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X478 a_897_3260.t3 a_307_3697.t9 VDD.t936 VDD.t935 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X479 a_14406_3692.t4 A[2].t7 a_14288_3692.t2 VDD.t391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X480 VSS.t174 B[5].t7 a_17798_3694.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X481 a_6725_n7362.t1 a_7019_n7388.t6 a_6607_n7362.t1 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X482 a_2470_n7362.t4 A[1].t11 VDD.t1014 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X483 a_13429_1740.t10 a_13369_1714.t5 VDD.t877 VDD.t876 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X484 VSS.t58 a_3843_3262.t5 a_7904_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X485 a_2588_n7362.t0 a_2882_n7388.t6 a_2470_n7362.t3 VDD.t201 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X486 a_520_n7364.t0 a_n25_n6671.t4 a_402_n7364.t4 VDD.t928 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X487 a_22789_n1016.t3 a_23188_n3722.t8 VSS.t167 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X488 a_3951_n994.t11 opcode[1].t36 VDD.t779 VDD.t778 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X489 VSS.t120 a_17447_n1479.t5 a_17394_n2327.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X490 a_n25_n6671.t2 A[0].t12 VDD.t464 VDD.t463 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X491 a_7432_n990.t1 a_7957_n1475.t6 a_7083_n990.t3 VDD.t280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X492 VDD.t37 opcode[0].t57 a_19695_n3722.t2 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X493 VDD.t1026 a_17798_3694.t7 a_16513_1714.t1 VDD.t1025 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X494 VDD.t373 A[4].t9 a_8249_n6669.t2 VDD.t372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X495 a_7432_1744.t4 a_3843_3262.t6 a_7083_1744.t9 VDD.t956 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X496 a_13429_n994.t1 a_13369_n1020.t5 VDD.t226 VDD.t225 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X497 a_7422_n3722.t5 a_6514_n3722.t6 a_7073_n3722.t10 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X498 VDD.t1253 B[0].t7 a_307_3697.t6 VDD.t1252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X499 VSS.t160 a_6811_3260.t6 a_14250_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X500 a_7019_n7388.t3 B[3].t8 VSS.t83 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X501 a_6607_n7362.t0 a_7019_n7388.t7 a_6725_n7362.t0 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X502 a_11205_3262.t3 a_10615_3699.t9 VSS.t148 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X503 VDD.t273 B[2].t5 a_4539_n7364.t2 VDD.t272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X504 VDD.t718 a_1755_3697.t8 a_2345_3260.t2 VDD.t717 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X505 a_4536_407.t0 a_3891_1714.t5 VSS.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X506 a_19695_n3722.t1 opcode[0].t58 VDD.t295 VDD.t294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X507 a_8249_n6669.t1 A[4].t10 VDD.t375 VDD.t374 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X508 a_7023_1718.t1 a_14288_3692.t6 VDD.t1152 VDD.t1151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X509 a_3951_1740.t4 a_3891_1714.t6 VDD.t1134 VDD.t1133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X510 VDD.t297 opcode[0].t59 a_12860_n3726.t0 VDD.t296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X511 a_7019_n7388.t2 B[3].t9 VDD.t306 VDD.t305 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X512 a_1628_n2327.t0 a_248_n994.t6 a_1156_n994.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X513 a_14014_n2327.t1 a_13369_n1020.t6 VSS.t56 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X514 a_2882_n7388.t2 B[1].t5 VDD.t558 VDD.t557 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X515 a_22839_n3722.t3 opcode[0].t60 VDD.t299 VDD.t298 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X516 a_16912_n3726.t3 a_16004_n3726.t6 a_16563_n3726.t4 VDD.t251 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X517 VDD.t1116 A[2].t8 a_7013_n3748.t1 VDD.t1115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X518 a_3951_n994.t9 a_3891_n1020.t5 VDD.t1218 VDD.t1217 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X519 a_19705_n990.t10 a_19645_n1016.t5 VDD.t755 VDD.t754 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X520 VDD.t913 opcode[0].t61 a_13419_n3726.t5 VDD.t912 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X521 a_20054_n990.t6 a_20579_n1475.t6 a_19705_n990.t7 VDD.t1063 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X522 a_3941_n3726.t10 a_3881_n3752.t5 VDD.t1017 VDD.t1016 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X523 a_14999_n7360.t1 a_15293_n7386.t5 a_14881_n7360.t11 VDD.t892 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X524 a_19705_1744.t4 a_19230_3112.t6 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X525 a_4539_n7364.t1 B[2].t6 VDD.t275 VDD.t274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X526 a_16563_n3726.t10 a_16503_n3752.t4 VDD.t1046 VDD.t1045 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X527 VDD.t540 B[7].t8 a_10615_3699.t6 VDD.t539 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X528 a_20054_1744.t3 a_9757_3262.t5 a_19705_1744.t10 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X529 a_20054_n990.t2 a_19146_n990.t5 a_19705_n990.t2 VDD.t345 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X530 VDD.t915 opcode[0].t62 a_19695_n3722.t0 VDD.t914 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X531 a_13369_n1020.t2 a_13768_n3726.t9 VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X532 VDD.t917 opcode[0].t63 a_807_1740.t1 VDD.t916 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X533 VDD.t377 A[4].t11 a_8249_n6669.t0 VDD.t376 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X534 a_20054_1744.t7 a_19146_1744.t4 a_19705_1744.t8 VDD.t994 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X535 a_13778_1740.t0 opcode[0].t64 a_14014_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X536 a_19705_n990.t6 a_20579_n1475.t7 a_20054_n990.t7 VDD.t1064 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X537 VDD.t308 B[3].t10 a_7019_n7388.t1 VDD.t307 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X538 a_19705_1744.t9 a_9757_3262.t6 a_20054_1744.t5 VDD.t846 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X539 VSS.t42 a_1681_n1479.t7 a_1628_n2327.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X540 a_11098_n8092.t1 A[5].t5 a_10862_n7360.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X541 a_17916_3694.t1 B[5].t8 VDD.t662 VDD.t661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X542 VDD.t658 opcode[1].t37 a_807_n994.t1 VDD.t657 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X543 VDD.t550 B[1].t6 a_2882_n7388.t1 VDD.t549 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X544 VDD.t1008 opcode[0].t65 a_22839_n3722.t2 VDD.t1007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X545 a_7013_n3748.t0 A[2].t9 VDD.t1118 VDD.t1117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X546 VSS.t35 a_8794_n7362.t10 a_14240_n5059.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X547 VSS.t87 opcode[1].t38 a_6524_n990.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X548 VSS.t139 opcode[0].t66 a_19146_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X549 VDD.t277 B[2].t7 a_4539_n7364.t0 VDD.t276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X550 a_22789_n1016.t2 a_23188_n3722.t9 VDD.t1226 VDD.t1225 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X551 VDD.t1214 a_16503_n3752.t5 a_16563_n3726.t11 VDD.t1213 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X552 a_18966_3696.t1 A[6].t15 a_19084_3696.t4 VDD.t1206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X553 a_1628_407.t1 a_248_1740.t6 a_1156_1740.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X554 VSS.t157 a_11101_n1475.t5 a_11048_n2323.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X555 VDD.t1140 a_13768_n3726.t10 a_13369_n1020.t1 VDD.t1139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X556 a_8259_3260.t1 a_7669_3697.t8 VDD.t1088 VDD.t1087 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X557 a_10227_n990.t7 a_9668_n990.t6 a_10576_n990.t2 VDD.t435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X558 a_7019_n7388.t0 B[3].t11 VDD.t310 VDD.t309 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X559 a_10227_1744.t2 a_9668_1744.t6 a_10576_1744.t1 VDD.t693 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X560 VSS.t88 B[5].t9 a_11098_n8092.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X561 a_13768_n3726.t1 a_8794_n7362.t11 a_13419_n3726.t3 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X562 a_7083_n990.t11 a_6524_n990.t5 a_7432_n990.t7 VDD.t699 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X563 a_4825_n1479.t1 a_4300_1740.t10 VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X564 a_7083_1744.t3 a_6524_1744.t4 a_7432_1744.t1 VDD.t315 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X565 VDD.t857 opcode[0].t67 a_12870_1740.t1 VDD.t856 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X566 a_14303_n1479.t2 a_13778_1740.t10 VSS.t134 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X567 a_13429_1740.t9 a_13369_1714.t6 VDD.t524 VDD.t523 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X568 VDD.t1222 a_23188_n3722.t10 a_22789_n1016.t1 VDD.t1221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X569 a_11952_3694.t4 A[0].t13 a_12070_3694.t2 VDD.t727 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X570 a_20280_n5055.t1 a_19635_n3748.t4 VSS.t161 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X571 a_13369_n1020.t0 a_13768_n3726.t11 VDD.t1142 VDD.t1141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X572 VDD.t366 A[3].t10 a_4701_3699.t0 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X573 Y[1].t1 a_4300_n994.t10 VDD.t704 VDD.t703 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X574 a_12870_1740.t0 opcode[0].t68 VDD.t859 VDD.t858 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X575 VDD.t660 opcode[1].t39 a_12870_n994.t1 VDD.t659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X576 a_12813_n7362.t7 B[6].t6 VDD.t1131 VDD.t1130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X577 a_4938_3062.t1 A[3].t11 a_4701_3699.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X578 a_10812_411.t1 a_10167_1718.t6 VSS.t61 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X579 a_13429_n994.t6 a_13369_n1020.t7 VDD.t462 VDD.t461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X580 VSS.t97 opcode[1].t40 a_22290_n990.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X581 a_13369_1714.t1 a_16630_3696.t7 VDD.t871 VDD.t870 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X582 a_10862_n8092.t0 a_11156_n7386.t7 VSS.t117 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X583 a_12070_3694.t5 B[0].t8 VDD.t1203 VDD.t1202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X584 a_13225_n7388.t3 B[6].t7 VSS.t155 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X585 a_16513_n1020.t0 a_16912_n3726.t10 VDD.t1177 VDD.t1176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X586 a_9167_3699.t4 A[6].t16 VDD.t648 VDD.t647 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X587 a_12870_n994.t0 opcode[1].t41 VDD.t787 VDD.t786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X588 a_9757_3262.t1 a_9167_3699.t8 VDD.t606 VDD.t605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X589 a_20134_3694.t2 A[7].t11 a_20252_3694.t5 VDD.t1020 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X590 a_22789_n1016.t0 a_23188_n3722.t11 VDD.t1224 VDD.t1223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X591 a_14288_3692.t1 A[2].t10 VSS.t92 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X592 VDD.t1002 a_11952_3694.t6 a_747_1714.t2 VDD.t1001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X593 VDD.t616 A[3].t12 a_6180_n6669.t2 VDD.t615 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X594 VDD.t1183 B[6].t8 a_9167_3699.t6 VDD.t1182 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X595 VSS.t46 a_11205_3262.t6 a_23670_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X596 a_520_n7364.t3 a_n25_n6671.t5 a_520_n8096.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X597 a_6811_3260.t1 a_6221_3697.t8 VDD.t575 VDD.t574 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X598 a_13778_1740.t1 a_12870_1740.t5 a_13429_1740.t3 VDD.t790 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X599 VDD.t1092 A[1].t12 a_2043_n6669.t2 VDD.t1091 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X600 a_4657_n7364.t2 a_4112_n6671.t5 a_4657_n8096.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X601 VDD.t789 opcode[1].t42 a_19146_n990.t1 VDD.t788 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X602 VDD.t948 opcode[1].t43 a_19705_n990.t4 VDD.t947 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X603 a_13429_1740.t7 a_12870_1740.t6 a_13778_1740.t5 VDD.t987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X604 VDD.t861 opcode[0].t69 a_19146_1744.t1 VDD.t860 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X605 a_13778_n994.t6 a_12870_n994.t5 a_13429_n994.t10 VDD.t829 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X606 VDD.t54 opcode[0].t70 a_19705_1744.t1 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X607 a_10167_n1016.t3 a_10566_n3722.t11 VSS.t156 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X608 a_6180_n6669.t1 A[3].t13 VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X609 a_13225_n7388.t0 B[6].t9 VDD.t1185 VDD.t1184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X610 a_756_n8096.t1 A[0].t14 a_520_n7364.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X611 VDD.t56 opcode[0].t71 a_807_1740.t0 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X612 a_13429_n994.t2 a_12870_n994.t6 a_13778_n994.t0 VDD.t260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X613 a_11952_3694.t2 A[0].t15 VSS.t152 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X614 a_16573_1740.t0 a_16014_1740.t7 a_16922_1740.t1 VDD.t894 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X615 a_10744_n7360.t8 A[5].t6 VDD.t934 VDD.t933 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X616 a_4893_n8096.t1 A[2].t11 a_4657_n7364.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X617 a_23660_n5055.t1 a_22280_n3722.t4 a_23188_n3722.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X618 VDD.t817 a_1156_1740.t10 a_1681_n1479.t1 VDD.t816 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X619 VDD.t950 opcode[1].t44 a_807_n994.t0 VDD.t949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X620 a_3253_3699.t1 B[2].t8 VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X621 VDD.t384 B[6].t10 a_19084_3696.t1 VDD.t383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X622 a_16573_n994.t2 a_16014_n994.t7 a_16922_n994.t1 VDD.t317 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X623 a_13359_n3752.t0 A[4].t12 VDD.t965 VDD.t964 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X624 a_402_n7364.t1 B[0].t9 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X625 VDD.t58 opcode[0].t72 a_16573_1740.t4 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X626 a_23198_1744.t0 opcode[0].t73 a_23434_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X627 VDD.t406 opcode[0].t74 a_3382_n3726.t2 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X628 VDD.t136 A[3].t14 a_6180_n6669.t0 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X629 VDD.t445 a_1156_n994.t10 Y[0].t1 VDD.t444 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X630 a_797_n3726.t8 a_238_n3726.t5 a_1146_n3726.t7 VDD.t1236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X631 Y[7].t1 a_23198_n990.t9 VDD.t759 VDD.t758 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X632 a_4290_n3726.t7 a_2588_n7362.t10 a_3941_n3726.t7 VDD.t679 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X633 a_16503_n3752.t2 A[5].t7 VDD.t638 VDD.t637 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X634 VDD.t952 opcode[1].t45 a_16573_n994.t4 VDD.t951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X635 a_16748_3696.t2 B[4].t11 VDD.t493 VDD.t492 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X636 a_23723_n1475.t3 a_23198_1744.t9 VDD.t1257 VDD.t1256 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X637 a_7904_411.t1 a_6524_1744.t5 a_7432_1744.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X638 VSS.t65 B[2].t9 a_4893_n8096.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X639 a_9757_3262.t3 a_9167_3699.t9 VSS.t84 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X640 a_15574_3694.t0 A[3].t15 a_15456_3694.t0 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X641 a_307_3697.t2 A[0].t16 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X642 a_10217_n3722.t6 opcode[0].t75 VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X643 a_13120_3694.t1 A[1].t13 a_13238_3694.t1 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X644 VDD.t449 A[1].t14 a_1755_3697.t1 VDD.t448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X645 a_797_n3726.t11 a_737_n3752.t5 VDD.t284 VDD.t283 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X646 a_2470_n7362.t10 B[1].t7 VDD.t552 VDD.t551 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X647 a_1992_3060.t0 A[1].t15 a_1755_3697.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X648 a_1146_n3726.t2 a_238_n3726.t6 a_797_n3726.t7 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X649 VDD.t511 B[2].t10 a_4951_n7390.t1 VDD.t510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X650 a_3941_n3726.t6 a_2588_n7362.t11 a_4290_n3726.t1 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X651 a_14999_n8092.t0 a_15293_n7386.t6 VSS.t40 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X652 a_23723_n1475.t0 a_23198_1744.t10 VSS.t129 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X653 VSS.t76 B[1].t8 a_1992_3060.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X654 a_8794_n7362.t4 a_8249_n6669.t4 a_8794_n8094.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X655 a_4701_3699.t3 B[3].t12 VDD.t921 VDD.t920 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X656 VDD.t538 B[7].t9 a_20252_3694.t3 VDD.t537 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X657 VSS.t131 opcode[1].t46 a_12870_n994.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X658 VSS.t112 a_9757_3262.t7 a_20526_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X659 VDD.t386 B[6].t11 a_9167_3699.t0 VDD.t385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X660 VDD.t1004 a_11952_3694.t7 a_747_1714.t3 VDD.t1003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X661 a_1156_1740.t0 opcode[0].t76 a_1392_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X662 VDD.t286 a_737_n3752.t6 a_797_n3726.t10 VDD.t285 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X663 VDD.t1244 B[1].t9 a_2470_n7362.t9 VDD.t1243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X664 a_7073_n3722.t0 a_7013_n3748.t6 VDD.t828 VDD.t827 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X665 a_3951_1740.t3 a_3891_1714.t7 VDD.t698 VDD.t697 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X666 a_797_n3726.t6 a_238_n3726.t7 a_1146_n3726.t3 VDD.t199 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X667 VSS.t17 A[2].t12 a_4112_n6671.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X668 a_4951_n7390.t0 B[2].t11 VDD.t267 VDD.t266 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X669 a_19695_n3722.t11 a_19635_n3748.t5 VDD.t1165 VDD.t1164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X670 VSS.t132 opcode[1].t47 a_16014_n994.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X671 VDD.t1022 A[7].t12 a_14881_n7360.t4 VDD.t1021 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X672 a_10615_3699.t0 A[7].t13 VDD.t255 VDD.t254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X673 a_3951_n994.t8 a_3891_n1020.t6 VDD.t1220 VDD.t1219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X674 Y[4].t3 a_13778_n994.t10 VSS.t32 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X675 a_9030_n8094.t1 A[4].t13 a_8794_n7362.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X676 a_10744_n7360.t7 A[5].t8 VDD.t640 VDD.t639 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X677 a_807_1740.t9 a_747_1714.t6 VDD.t767 VDD.t766 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X678 VDD.t954 opcode[1].t48 a_19705_n990.t3 VDD.t953 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X679 Y[6].t3 a_20054_n990.t10 VSS.t89 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X680 a_17798_3694.t3 A[5].t9 a_17916_3694.t4 VDD.t641 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X681 a_20398_3112.t0 a_20134_3694.t8 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X682 VDD.t1044 a_7023_n1016.t7 a_7083_n990.t7 VDD.t1043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X683 a_797_n3726.t9 a_737_n3752.t7 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X684 a_7669_3697.t1 A[5].t10 VDD.t320 VDD.t319 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X685 VDD.t92 opcode[0].t77 a_19705_1744.t0 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X686 VDD.t1072 a_7023_1718.t6 a_7083_1744.t4 VDD.t1071 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X687 VDD.t484 a_19635_n3748.t6 a_19695_n3722.t10 VDD.t483 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X688 VSS.t130 B[5].t10 a_7906_3060.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X689 a_807_n994.t9 a_747_n1020.t7 VDD.t769 VDD.t768 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X690 a_14881_n7360.t3 A[7].t14 VDD.t257 VDD.t256 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X691 VDD.t675 a_20054_n990.t11 Y[6].t0 VDD.t674 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X692 a_17916_3694.t3 A[5].t11 a_17798_3694.t2 VDD.t321 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X693 Y[7].t3 a_23198_n990.t10 VSS.t135 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X694 VDD.t1052 a_20054_1744.t10 a_20579_n1475.t0 VDD.t1051 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X695 a_4300_1740.t2 a_3392_1740.t7 a_3951_1740.t10 VDD.t911 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X696 VDD.t323 A[5].t12 a_10744_n7360.t6 VDD.t322 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X697 a_4526_n5059.t1 a_3881_n3752.t6 VSS.t121 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X698 VDD.t94 opcode[0].t78 a_3941_n3726.t2 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X699 VDD.t781 opcode[1].t49 a_9668_n990.t0 VDD.t780 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X700 a_10157_n3748.t1 A[3].t16 VDD.t482 VDD.t481 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X701 a_3843_3262.t0 a_3253_3699.t10 VDD.t716 VDD.t715 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X702 VDD.t865 B[6].t12 a_19084_3696.t0 VDD.t864 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X703 VDD.t17 opcode[0].t79 a_9668_1744.t0 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X704 a_4300_n994.t1 a_3392_n994.t7 a_3951_n994.t1 VDD.t184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X705 a_23670_411.t1 a_22290_1744.t6 a_23198_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X706 a_19695_n3722.t9 a_19635_n3748.t7 VDD.t486 VDD.t485 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X707 a_3951_1740.t7 a_2345_3260.t7 a_4300_1740.t5 VDD.t487 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X708 VDD.t536 B[7].t10 a_14881_n7360.t8 VDD.t535 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X709 a_6811_3260.t3 a_6221_3697.t9 VSS.t82 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X710 a_7083_n990.t5 a_6524_n990.t6 a_7432_n990.t3 VDD.t289 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X711 a_8676_n7362.t6 A[4].t14 VDD.t967 VDD.t966 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X712 a_7083_1744.t11 a_6524_1744.t6 a_7432_1744.t7 VDD.t1157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X713 VDD.t783 opcode[1].t50 a_10227_n990.t0 VDD.t782 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X714 Y[3].t1 a_10576_n990.t10 VDD.t1271 VDD.t1270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X715 a_3951_n994.t5 a_4825_n1479.t7 a_4300_n994.t7 VDD.t393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X716 a_4290_n3726.t0 opcode[0].t80 a_4526_n5059.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X717 VDD.t19 opcode[0].t81 a_10227_1744.t3 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X718 a_11101_n1475.t1 a_10576_1744.t10 VDD.t795 VDD.t794 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X719 a_3941_n3726.t1 opcode[0].t82 VDD.t352 VDD.t351 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X720 VDD.t354 opcode[0].t83 a_10217_n3722.t5 VDD.t353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X721 VDD.t1246 B[1].t10 a_13238_3694.t5 VDD.t1245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X722 VDD.t1112 a_10576_n990.t11 Y[3].t0 VDD.t1111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X723 VSS.t30 B[0].t10 a_544_3060.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X724 a_1755_3697.t4 B[1].t11 VDD.t1248 VDD.t1247 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X725 a_20579_n1475.t3 a_20054_1744.t11 VSS.t146 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X726 a_12931_n7362.t4 a_12386_n6669.t6 a_12813_n7362.t9 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X727 VDD.t797 a_10576_1744.t11 a_11101_n1475.t0 VDD.t796 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X728 VDD.t195 B[1].t12 a_2470_n7362.t8 VDD.t194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X729 VDD.t826 a_22789_n1016.t6 a_22849_n990.t10 VDD.t825 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X730 a_20290_n2323.t1 a_19645_n1016.t6 VSS.t149 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X731 VSS.t66 B[4].t12 a_6458_3060.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X732 a_16573_1740.t11 a_16513_1714.t6 VDD.t1110 VDD.t1109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X733 a_2882_n7388.t3 B[1].t13 VSS.t29 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X734 a_2470_n7362.t11 a_2882_n7388.t7 a_2588_n7362.t7 VDD.t1132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X735 a_5291_3262.t0 a_4701_3699.t10 VDD.t134 VDD.t133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X736 VDD.t984 a_20398_3112.t5 a_22849_1744.t6 VDD.t983 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X737 a_402_n7364.t3 a_n25_n6671.t6 a_520_n7364.t2 VDD.t1211 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X738 VDD.t837 A[0].t17 a_n25_n6671.t1 VDD.t836 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X739 a_10566_n3722.t1 a_6725_n7362.t11 a_10217_n3722.t1 VDD.t896 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X740 VDD.t785 opcode[1].t51 a_22290_n990.t0 VDD.t784 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X741 VDD.t822 a_13120_3694.t7 a_3891_1714.t2 VDD.t821 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X742 VDD.t513 B[4].t13 a_6221_3697.t0 VDD.t512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X743 a_13120_3694.t2 A[1].t16 VSS.t62 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X744 VDD.t356 opcode[0].t84 a_22290_1744.t0 VDD.t355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X745 a_22849_n990.t0 a_22789_n1016.t7 VDD.t102 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X746 a_4539_n7364.t7 a_4112_n6671.t6 a_4657_n7364.t4 VDD.t249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X747 a_16573_n994.t8 a_16513_n1020.t6 VDD.t562 VDD.t561 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X748 VDD.t923 B[3].t13 a_6607_n7362.t4 VDD.t922 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X749 VDD.t130 A[2].t13 a_4112_n6671.t0 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X750 a_8259_3260.t3 a_7669_3697.t9 VSS.t145 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X751 a_22849_1744.t0 a_20398_3112.t6 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X752 a_13419_n3726.t2 a_13359_n3752.t5 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X753 VDD.t1138 a_9167_3699.t10 a_9757_3262.t0 VDD.t1137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X754 a_10167_1718.t3 a_15456_3694.t8 VSS.t171 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X755 a_19635_n3748.t0 A[6].t17 VDD.t650 VDD.t649 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X756 a_19695_n3722.t5 a_12931_n7362.t8 a_20044_n3722.t4 VDD.t1065 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X757 VDD.t737 a_10167_n1016.t6 a_10227_n990.t3 VDD.t736 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X758 a_11156_n7386.t0 B[5].t11 VDD.t946 VDD.t945 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X759 a_520_n7364.t1 a_n25_n6671.t7 a_402_n7364.t2 VDD.t671 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X760 a_807_1740.t3 a_248_1740.t7 a_1156_1740.t2 VDD.t324 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X761 VDD.t504 a_10167_1718.t7 a_10227_1744.t7 VDD.t503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X762 a_6725_n7362.t5 a_6180_n6669.t5 a_6725_n8094.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X763 VDD.t84 opcode[0].t85 a_248_1740.t0 VDD.t83 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X764 a_4657_n7364.t3 a_4112_n6671.t7 a_4539_n7364.t6 VDD.t878 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X765 a_22839_n3722.t6 a_21997_n6357.t6 VDD.t1033 VDD.t1032 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X766 a_6524_n990.t0 opcode[1].t52 VDD.t228 VDD.t227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X767 VDD.t29 a_13359_n3752.t6 a_13419_n3726.t0 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X768 a_807_n994.t8 a_248_n994.t7 a_1156_n994.t7 VDD.t726 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X769 a_6524_1744.t0 opcode[0].t86 VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X770 a_14303_n1479.t3 a_13778_1740.t11 VDD.t972 VDD.t971 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X771 VDD.t230 opcode[1].t53 a_248_n994.t0 VDD.t229 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X772 VDD.t1195 B[5].t12 a_7669_3697.t5 VDD.t1194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X773 a_23198_n990.t1 a_22290_n990.t6 a_22849_n990.t4 VDD.t584 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X774 VSS.t34 A[7].t15 a_14454_n6667.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X775 a_20044_n3722.t3 a_12931_n7362.t9 a_19695_n3722.t4 VDD.t1005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X776 VDD.t88 opcode[0].t87 a_6514_n3722.t1 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X777 a_23198_1744.t2 a_22290_1744.t7 a_22849_1744.t7 VDD.t588 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X778 VSS.t36 A[5].t13 a_10317_n6667.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X779 a_14881_n7360.t6 a_15293_n7386.t7 a_14999_n7360.t0 VDD.t282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X780 a_23434_411.t1 a_20398_3112.t7 VSS.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X781 Y[4].t0 a_13778_n994.t11 VDD.t218 VDD.t217 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X782 VDD.t11 opcode[0].t88 a_3951_1740.t1 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X783 a_17447_n1479.t1 a_16922_1740.t10 VDD.t907 VDD.t906 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X784 a_4539_n7364.t11 a_4951_n7390.t4 a_4657_n7364.t5 VDD.t742 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X785 VDD.t1098 B[0].t11 a_402_n7364.t8 VDD.t1097 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X786 a_23188_n3722.t1 a_14999_n7360.t10 a_22839_n3722.t9 VDD.t399 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X787 VDD.t13 opcode[0].t89 a_7073_n3722.t8 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X788 VDD.t395 a_307_3697.t10 a_897_3260.t0 VDD.t394 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X789 a_22849_n990.t7 a_23723_n1475.t7 a_23198_n990.t5 VDD.t745 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X790 a_23670_n2323.t0 a_22290_n990.t7 a_23198_n990.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X791 a_8794_n7362.t7 a_8249_n6669.t5 a_8676_n7362.t10 VDD.t1186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X792 VDD.t42 a_21997_n6357.t7 a_22839_n3722.t5 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X793 a_14288_3692.t4 A[2].t14 a_14406_3692.t3 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X794 a_17798_3694.t0 A[5].t14 VSS.t37 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X795 a_4657_n8096.t1 a_4951_n7390.t5 VSS.t95 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X796 a_13419_n3726.t1 a_13359_n3752.t7 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X797 VDD.t15 opcode[0].t90 a_9658_n3722.t2 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X798 a_22849_1744.t5 a_11205_3262.t7 a_23198_1744.t1 VDD.t338 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X799 VDD.t232 opcode[1].t54 a_3951_n994.t2 VDD.t231 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X800 Y[5].t1 a_16922_n994.t10 VDD.t207 VDD.t206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X801 a_2882_n7388.t0 B[1].t14 VDD.t197 VDD.t196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X802 a_7432_1744.t0 opcode[0].t91 a_7668_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X803 a_6514_n3722.t0 opcode[0].t92 VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X804 a_16513_1714.t0 a_17798_3694.t8 VDD.t1028 VDD.t1027 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X805 a_10576_n990.t3 a_11101_n1475.t6 a_10227_n990.t9 VDD.t792 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X806 a_16563_n3726.t6 a_16503_n3752.t6 VDD.t401 VDD.t400 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X807 a_307_3697.t5 B[0].t12 VDD.t1189 VDD.t1188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X808 VSS.t54 opcode[0].t93 a_3382_n3726.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X809 a_10576_1744.t6 a_5291_3262.t6 a_10227_1744.t9 VDD.t968 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X810 a_16503_n3752.t3 A[5].t15 VSS.t38 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X811 VDD.t348 opcode[0].t94 a_16004_n3726.t1 VDD.t347 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X812 VDD.t824 B[1].t15 a_13238_3694.t4 VDD.t823 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X813 a_7432_n990.t2 a_7957_n1475.t7 a_7083_n990.t4 VDD.t281 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X814 a_8676_n7362.t11 a_8249_n6669.t6 a_8794_n7362.t6 VDD.t1187 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X815 VDD.t1 A[0].t18 a_n25_n6671.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X816 VDD.t925 B[3].t14 a_15574_3694.t2 VDD.t924 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X817 a_10802_n5055.t1 a_10157_n3748.t7 VSS.t94 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X818 a_9658_n3722.t1 opcode[0].t95 VDD.t350 VDD.t349 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X819 a_7432_1744.t5 a_3843_3262.t7 a_7083_1744.t10 VDD.t957 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X820 a_16573_1740.t6 a_16513_1714.t7 VDD.t452 VDD.t451 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X821 a_2345_3260.t1 a_1755_3697.t9 VDD.t720 VDD.t719 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X822 a_3891_n1020.t3 a_4290_n3726.t11 VSS.t51 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X823 VDD.t577 a_6221_3697.t10 a_6811_3260.t0 VDD.t576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X824 VDD.t1154 a_14288_3692.t7 a_7023_1718.t2 VDD.t1153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X825 a_20526_411.t0 a_19146_1744.t5 a_20054_1744.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X826 a_16573_n994.t7 a_16513_n1020.t7 VDD.t564 VDD.t563 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X827 a_22839_n3722.t8 a_22280_n3722.t5 a_23188_n3722.t6 VDD.t329 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X828 a_1392_407.t1 a_747_1714.t7 VSS.t107 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X829 a_20044_n3722.t0 opcode[0].t96 a_20280_n5055.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X830 a_16004_n3726.t0 opcode[0].t97 VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X831 VDD.t534 B[7].t11 a_10615_3699.t5 VDD.t533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X832 VDD.t867 B[6].t13 a_12813_n7362.t6 VDD.t866 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X833 a_8794_n7362.t5 a_8249_n6669.t7 a_8676_n7362.t9 VDD.t1251 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X834 a_3891_1714.t3 a_13120_3694.t8 VSS.t105 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X835 VDD.t1124 a_19645_n1016.t7 a_19705_n990.t9 VDD.t1123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X836 VSS.t67 B[4].t14 a_9030_n8094.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X837 a_10566_n3722.t4 opcode[0].t98 a_10802_n5055.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X838 VDD.t82 opcode[0].t99 a_9658_n3722.t0 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X839 a_7073_n3722.t11 a_6514_n3722.t7 a_7422_n3722.t7 VDD.t1119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X840 VDD.t25 a_19230_3112.t7 a_19705_1744.t3 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X841 a_19705_n990.t1 a_19146_n990.t6 a_20054_n990.t3 VDD.t346 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X842 a_10615_3699.t4 B[7].t12 VDD.t532 VDD.t531 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X843 VDD.t632 A[5].t16 a_10317_n6667.t1 VDD.t631 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X844 a_15293_n7386.t1 B[7].t13 VDD.t530 VDD.t529 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X845 a_20044_n3722.t5 a_12931_n7362.t10 a_19695_n3722.t3 VDD.t1006 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X846 a_19705_1744.t6 a_19146_1744.t6 a_20054_1744.t4 VDD.t731 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X847 a_12931_n7362.t6 a_12386_n6669.t7 a_12931_n8094.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X848 a_23188_n3722.t0 a_22280_n3722.t6 a_22839_n3722.t0 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X849 a_13429_1740.t8 a_6811_3260.t7 a_13778_1740.t7 VDD.t1161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X850 a_20516_n5055.t1 a_19136_n3722.t7 a_20044_n3722.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X851 a_13419_n3726.t10 a_12860_n3726.t5 a_13768_n3726.t6 VDD.t1015 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X852 VDD.t729 a_10615_3699.t10 a_11205_3262.t0 VDD.t728 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X853 a_2043_n6669.t1 A[1].t17 VDD.t507 VDD.t506 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X854 a_7658_n5055.t0 a_7013_n3748.t7 VSS.t106 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X855 a_19645_n1016.t1 a_20044_n3722.t10 VDD.t833 VDD.t832 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X856 VDD.t7 opcode[0].t100 a_7073_n3722.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X857 a_16748_3696.t4 A[4].t15 a_16630_3696.t3 VDD.t960 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X858 VSS.t1 opcode[0].t101 a_3392_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X859 a_13429_n994.t7 a_14303_n1479.t7 a_13778_n994.t3 VDD.t362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X860 a_10157_n3748.t3 A[3].t17 VSS.t59 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X861 a_16573_1740.t9 a_8259_3260.t6 a_16922_1740.t6 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X862 VDD.t120 A[2].t15 a_3253_3699.t3 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X863 a_19084_3696.t3 A[6].t18 a_18966_3696.t3 VDD.t642 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X864 a_10317_n6667.t0 A[5].t17 VDD.t634 VDD.t633 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X865 a_16563_n3726.t3 a_16004_n3726.t7 a_16912_n3726.t2 VDD.t252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X866 VDD.t1090 a_7669_3697.t10 a_8259_3260.t0 VDD.t1089 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X867 VDD.t688 opcode[1].t55 a_22849_n990.t2 VDD.t687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X868 VDD.t528 B[7].t14 a_15293_n7386.t0 VDD.t527 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X869 a_3490_3062.t1 A[2].t16 a_3253_3699.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X870 VDD.t9 opcode[0].t102 a_3951_1740.t0 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X871 VDD.t422 opcode[0].t103 a_22849_1744.t3 VDD.t421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X872 a_22839_n3722.t1 a_22280_n3722.t7 a_23188_n3722.t4 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X873 a_16922_1740.t5 a_8259_3260.t7 a_16573_1740.t8 VDD.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X874 a_16573_n994.t10 a_17447_n1479.t6 a_16922_n994.t6 VDD.t993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X875 VSS.t138 a_12931_n7362.t11 a_20516_n5055.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X876 VDD.t424 opcode[0].t104 a_13419_n3726.t4 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X877 a_7432_n990.t4 a_6524_n990.t7 a_7083_n990.t6 VDD.t290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X878 VDD.t52 a_4300_1740.t11 a_4825_n1479.t0 VDD.t51 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X879 VDD.t690 opcode[1].t56 a_3951_n994.t7 VDD.t689 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X880 VDD.t96 A[1].t18 a_2043_n6669.t0 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X881 a_7432_1744.t3 a_6524_1744.t7 a_7083_1744.t8 VDD.t700 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X882 a_10227_n990.t6 a_9668_n990.t7 a_10576_n990.t5 VDD.t955 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X883 a_4536_n2327.t1 a_3891_n1020.t7 VSS.t122 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X884 VDD.t835 a_20044_n3722.t11 a_19645_n1016.t0 VDD.t834 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X885 a_7073_n3722.t6 opcode[0].t105 VDD.t426 VDD.t425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X886 VDD.t269 B[2].t12 a_14406_3692.t1 VDD.t268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X887 a_16922_n994.t7 a_17447_n1479.t7 a_16573_n994.t11 VDD.t1034 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X888 a_10227_1744.t1 a_9668_1744.t7 a_10576_1744.t0 VDD.t694 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X889 VSS.t50 a_14999_n7360.t11 a_23660_n5055.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X890 a_17148_n5059.t1 a_16503_n3752.t7 VSS.t102 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X891 a_19230_3112.t1 a_18966_3696.t7 VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X892 a_7083_n990.t1 opcode[1].t57 VDD.t692 VDD.t691 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X893 a_10576_n990.t4 a_11101_n1475.t7 a_10227_n990.t10 VDD.t793 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X894 VDD.t340 opcode[0].t106 a_16563_n3726.t2 VDD.t339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X895 VDD.t706 a_4300_n994.t11 Y[1].t0 VDD.t705 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X896 a_7083_1744.t1 opcode[0].t107 VDD.t342 VDD.t341 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X897 a_10576_1744.t5 a_5291_3262.t7 a_10227_1744.t10 VDD.t969 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X898 VDD.t887 B[0].t13 a_12070_3694.t1 VDD.t886 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X899 VDD.t873 a_16630_3696.t8 a_13369_1714.t0 VDD.t872 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X900 VDD.t63 opcode[1].t58 a_7083_n990.t0 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X901 Y[2].t0 a_7432_n990.t11 VDD.t522 VDD.t521 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X902 a_3382_n3726.t1 opcode[0].t108 VDD.t344 VDD.t343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X903 a_6725_n7362.t2 a_6180_n6669.t6 a_6607_n7362.t2 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X904 VDD.t598 B[3].t15 a_4701_3699.t2 VDD.t597 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X905 VDD.t74 opcode[0].t109 a_7083_1744.t0 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X906 a_7957_n1475.t0 a_7432_1744.t11 VDD.t265 VDD.t264 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X907 VDD.t636 A[5].t18 a_16503_n3752.t1 VDD.t635 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X908 a_4300_n994.t5 opcode[1].t59 a_4536_n2327.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X909 a_2345_3260.t0 a_1755_3697.t10 VDD.t722 VDD.t721 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X910 a_6221_3697.t4 A[4].t16 VDD.t962 VDD.t961 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X911 a_16563_n3726.t1 opcode[0].t110 VDD.t76 VDD.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X912 a_7023_n1016.t2 a_7422_n3722.t10 VDD.t1191 VDD.t1190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X913 a_9167_3699.t3 A[6].t19 VDD.t644 VDD.t643 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X914 VSS.t8 opcode[0].t111 a_19136_n3722.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X915 VSS.t111 B[6].t14 a_9404_3062.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X916 a_13429_1740.t6 a_12870_1740.t7 a_13778_1740.t4 VDD.t981 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X917 VDD.t3 opcode[0].t112 a_3382_n3726.t0 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X918 VSS.t0 opcode[0].t113 a_9658_n3722.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X919 a_7023_1718.t0 a_14288_3692.t8 VSS.t85 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X920 a_6607_n7362.t3 a_6180_n6669.t7 a_6725_n7362.t3 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X921 a_16503_n3752.t0 A[5].t19 VDD.t677 VDD.t676 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X922 a_13419_n3726.t11 a_12860_n3726.t6 a_13768_n3726.t7 VDD.t1122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X923 VDD.t5 opcode[0].t114 a_3392_1740.t0 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X924 a_19705_n990.t0 a_19146_n990.t7 a_20054_n990.t4 VDD.t818 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X925 a_16912_n3726.t5 a_10862_n7360.t11 a_16563_n3726.t7 VDD.t848 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X926 a_13429_n994.t11 a_12870_n994.t7 a_13778_n994.t7 VDD.t1029 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X927 a_747_n1020.t2 a_1146_n3726.t11 VSS.t14 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X928 a_19705_1744.t7 a_19146_1744.t7 a_20054_1744.t6 VDD.t888 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X929 VDD.t683 A[7].t16 a_14454_n6667.t1 VDD.t682 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X930 VDD.t418 opcode[0].t115 a_16563_n3726.t0 VDD.t417 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X931 VDD.t65 opcode[1].t60 a_19146_n990.t0 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X932 VSS.t53 opcode[0].t116 a_9668_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X933 VDD.t996 opcode[1].t61 a_3392_n994.t0 VDD.t995 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X934 VDD.t420 opcode[0].t117 a_19146_1744.t0 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X935 a_16513_n1020.t1 a_16912_n3726.t11 VDD.t1179 VDD.t1178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X936 a_14014_407.t1 a_13369_1714.t7 VSS.t71 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X937 VDD.t333 opcode[0].t118 a_238_n3726.t0 VDD.t332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X938 VDD.t335 opcode[0].t119 a_797_n3726.t5 VDD.t334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X939 a_13768_n3726.t3 a_12860_n3726.t7 a_13419_n3726.t7 VDD.t219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X940 a_1681_n1479.t0 a_1156_1740.t11 VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X941 VDD.t271 B[2].t13 a_3253_3699.t0 VDD.t270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X942 VDD.t998 opcode[1].t62 a_22849_n990.t1 VDD.t997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X943 a_14454_n6667.t0 A[7].t17 VDD.t685 VDD.t684 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X944 a_16573_1740.t3 opcode[0].t120 VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X945 a_4657_n7364.t7 a_4951_n7390.t6 a_4539_n7364.t10 VDD.t292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X946 a_4539_n7364.t5 A[2].t17 VDD.t1181 VDD.t1180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X947 a_16748_3696.t5 A[4].t17 a_16630_3696.t4 VDD.t963 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X948 VDD.t466 opcode[0].t121 a_22849_1744.t2 VDD.t465 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X949 Y[0].t0 a_1156_n994.t11 VDD.t447 VDD.t446 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X950 a_1146_n3726.t0 a_520_n7364.t11 a_797_n3726.t0 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X951 VDD.t215 A[3].t18 a_10157_n3748.t0 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X952 a_17447_n1479.t0 a_16922_1740.t11 VDD.t909 VDD.t908 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X953 VDD.t978 a_23198_n990.t11 Y[7].t0 VDD.t977 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X954 a_16630_3696.t1 A[4].t18 VSS.t118 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X955 a_16573_n994.t3 opcode[1].t63 VDD.t1000 VDD.t999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X956 VDD.t670 B[4].t15 a_16748_3696.t1 VDD.t669 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X957 VDD.t944 a_23198_1744.t11 a_23723_n1475.t1 VDD.t943 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X958 a_797_n3726.t4 opcode[0].t122 VDD.t468 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X959 VDD.t1114 B[2].t14 a_14406_3692.t0 VDD.t1113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X960 VSS.t7 B[0].t14 a_756_n8096.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X961 VDD.t470 opcode[0].t123 a_19136_n3722.t0 VDD.t469 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X962 Y[5].t0 a_16922_n994.t11 VDD.t209 VDD.t208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X963 VDD.t1197 B[5].t13 a_10744_n7360.t4 VDD.t1196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X964 a_13238_3694.t0 A[1].t19 a_13120_3694.t3 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X965 a_7668_411.t1 a_7023_1718.t7 VSS.t143 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X966 a_4951_n7390.t3 B[2].t15 VSS.t147 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X967 a_4539_n7364.t9 a_4951_n7390.t7 a_4657_n7364.t6 VDD.t293 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X968 VDD.t1229 A[2].t18 a_4539_n7364.t4 VDD.t1228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X969 a_15574_3694.t1 A[3].t19 a_15456_3694.t1 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X970 a_402_n7364.t5 a_814_n7390.t6 a_520_n7364.t4 VDD.t1175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X971 a_307_3697.t1 A[0].t19 VDD.t259 VDD.t258 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X972 a_7023_n1016.t3 a_7422_n3722.t11 VSS.t164 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X973 a_19230_3112.t0 a_18966_3696.t8 VSS.t11 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X974 VDD.t432 opcode[0].t124 a_797_n3726.t3 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X975 a_14881_n7360.t7 B[7].t15 VDD.t526 VDD.t525 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X976 a_520_n8096.t1 a_814_n7390.t7 VSS.t163 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X977 a_6221_3697.t3 A[4].t19 VDD.t880 VDD.t879 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X978 VDD.t187 B[0].t15 a_12070_3694.t0 VDD.t186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X979 a_20252_3694.t4 A[7].t18 a_20134_3694.t1 VDD.t686 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X980 a_3941_n3726.t9 a_3881_n3752.t7 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X981 a_10744_n7360.t3 B[5].t14 VDD.t328 VDD.t327 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X982 a_9167_3699.t5 B[6].t15 VDD.t845 VDD.t844 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X983 a_747_1714.t0 a_11952_3694.t8 VDD.t989 VDD.t988 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X984 VDD.t942 A[7].t19 a_21997_n6357.t0 VDD.t941 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X985 a_4539_n7364.t3 A[2].t19 VDD.t1231 VDD.t1230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X986 a_10812_n2323.t1 a_10167_n1016.t7 VSS.t93 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X987 a_8676_n7362.t0 a_9088_n7388.t7 a_8794_n7362.t0 VDD.t1227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X988 a_20054_1744.t1 opcode[0].t125 a_20290_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X989 VDD.t434 opcode[0].t126 a_3941_n3726.t0 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X990 a_11156_n7386.t3 B[5].t15 VSS.t45 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X991 VDD.t1136 opcode[0].t127 a_10217_n3722.t4 VDD.t1135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
R0 B[7].t9 B[7].t3 799.268
R1 B[7].n9 B[7].n1 648.503
R2 B[7].n7 B[7].n6 592.056
R3 B[7].t7 B[7].t11 415.315
R4 B[7].t13 B[7].n4 313.873
R5 B[7].n6 B[7].t5 294.986
R6 B[7].n0 B[7].t0 285.543
R7 B[7].n3 B[7].t10 272.288
R8 B[7].n8 B[7].t7 217.472
R9 B[7].n2 B[7].t8 214.335
R10 B[7].t11 B[7].n2 214.335
R11 B[7].n7 B[7].t14 204.68
R12 B[7].n1 B[7].t9 194.406
R13 B[7].n5 B[7].t13 190.152
R14 B[7].n5 B[7].t2 190.152
R15 B[7].n0 B[7].t6 160.666
R16 B[7].n3 B[7].t15 160.666
R17 B[7].n4 B[7].t1 160.666
R18 B[7].n6 B[7].t4 110.859
R19 B[7].n4 B[7].n3 96.129
R20 B[7].n1 B[7].n0 91.137
R21 B[7].n2 B[7].t12 80.333
R22 B[7].t14 B[7].n5 80.333
R23 B[7].n8 B[7].n7 61.581
R24 B[7] B[7].n9 33.418
R25 B[7].n9 B[7].n8 6.999
R26 a_20252_3694.n0 a_20252_3694.t3 14.282
R27 a_20252_3694.n0 a_20252_3694.t4 14.282
R28 a_20252_3694.n1 a_20252_3694.t1 14.282
R29 a_20252_3694.n1 a_20252_3694.t2 14.282
R30 a_20252_3694.n3 a_20252_3694.t5 14.282
R31 a_20252_3694.t0 a_20252_3694.n3 14.282
R32 a_20252_3694.n3 a_20252_3694.n2 2.554
R33 a_20252_3694.n2 a_20252_3694.n1 2.361
R34 a_20252_3694.n2 a_20252_3694.n0 0.001
R35 VDD.t851 VDD.t77 95474.9
R36 VDD.t1057 VDD.t47 95474.9
R37 VDD.t801 VDD.t629 95474.9
R38 VDD.t69 VDD.t908 95474.9
R39 VDD.t1155 VDD.t1254 95474.9
R40 VDD.t578 VDD.t1047 95474.9
R41 VDD.t969 VDD.t794 95474.9
R42 VDD.t957 VDD.t264 95474.9
R43 VDD.t590 VDD.t446 95474.9
R44 VDD.t392 VDD.t701 95474.9
R45 VDD.t361 VDD.t806 95474.9
R46 VDD.t1034 VDD.t208 95474.9
R47 VDD.t743 VDD.t756 95474.9
R48 VDD.t1062 VDD.t402 95474.9
R49 VDD.t793 VDD.t1270 95474.9
R50 VDD.t281 VDD.t521 95474.9
R51 VDD.t927 VDD.t991 95474.9
R52 VDD.t678 VDD.t899 95474.9
R53 VDD.t141 VDD.t157 95474.9
R54 VDD.t853 VDD.t1178 95474.9
R55 VDD.t399 VDD.t1225 95474.9
R56 VDD.t1005 VDD.t832 95474.9
R57 VDD.t895 VDD.t169 95474.9
R58 VDD.t855 VDD.t1190 95474.9
R59 VDD.n45 VDD.t872 77361
R60 VDD.n74 VDD.n73 604.435
R61 VDD.n5 VDD.n4 604.408
R62 VDD.n60 VDD.n59 600.509
R63 VDD.n88 VDD.n87 600.503
R64 VDD.n19 VDD.n18 600.482
R65 VDD.n46 VDD.n45 563.326
R66 VDD.t1243 VDD.t557 413.681
R67 VDD.t1093 VDD.t945 413.681
R68 VDD.t1097 VDD.t188 413.681
R69 VDD.t276 VDD.t20 413.681
R70 VDD.t922 VDD.t305 413.681
R71 VDD.t179 VDD.t172 413.681
R72 VDD.t866 VDD.t1167 413.681
R73 VDD.t545 VDD.t529 413.681
R74 VDD.t819 VDD.t363 406.159
R75 VDD.t1151 VDD.t1162 406.159
R76 VDD.n4 VDD.t821 404.97
R77 VDD.n18 VDD.t1153 404.97
R78 VDD.t870 VDD.t872 397.517
R79 VDD.t114 VDD.t112 397.517
R80 VDD.n87 VDD.t89 396.391
R81 VDD.t613 VDD.t985 396.113
R82 VDD.t1027 VDD.t1025 396.113
R83 VDD.n73 VDD.t973 394.999
R84 VDD.n59 VDD.t1023 394.999
R85 VDD.n44 VDD.t868 394.148
R86 VDD.t764 VDD.t163 382.217
R87 VDD.t1133 VDD.t713 382.217
R88 VDD.t876 VDD.t1009 382.217
R89 VDD.t1109 VDD.t862 382.217
R90 VDD.t154 VDD.t241 382.217
R91 VDD.t840 VDD.t419 382.217
R92 VDD.t585 VDD.t16 382.217
R93 VDD.t1073 VDD.t303 382.217
R94 VDD.t192 VDD.t1081 382.217
R95 VDD.t1217 VDD.t1058 382.217
R96 VDD.t225 VDD.t1103 382.217
R97 VDD.t561 VDD.t1105 382.217
R98 VDD.t889 VDD.t1085 382.217
R99 VDD.t752 VDD.t64 382.217
R100 VDD.t732 VDD.t780 382.217
R101 VDD.t413 VDD.t1258 382.217
R102 VDD.t283 VDD.t1232 382.217
R103 VDD.t107 VDD.t2 382.217
R104 VDD.t70 VDD.t237 382.217
R105 VDD.t1045 VDD.t161 382.217
R106 VDD.t1032 VDD.t32 382.217
R107 VDD.t1164 VDD.t663 382.217
R108 VDD.t740 VDD.t81 382.217
R109 VDD.t1198 VDD.t707 382.217
R110 VDD.t163 VDD.t159 345.987
R111 VDD.t159 VDD.t83 345.987
R112 VDD.t816 VDD.t814 345.987
R113 VDD.t77 VDD.t816 345.987
R114 VDD.t713 VDD.t802 345.987
R115 VDD.t802 VDD.t4 345.987
R116 VDD.t51 VDD.t49 345.987
R117 VDD.t47 VDD.t51 345.987
R118 VDD.t1009 VDD.t858 345.987
R119 VDD.t858 VDD.t856 345.987
R120 VDD.t627 VDD.t971 345.987
R121 VDD.t629 VDD.t627 345.987
R122 VDD.t862 VDD.t239 345.987
R123 VDD.t239 VDD.t709 345.987
R124 VDD.t798 VDD.t906 345.987
R125 VDD.t908 VDD.t798 345.987
R126 VDD.t241 VDD.t711 345.987
R127 VDD.t711 VDD.t355 345.987
R128 VDD.t943 VDD.t1256 345.987
R129 VDD.t1254 VDD.t943 345.987
R130 VDD.t419 VDD.t473 345.987
R131 VDD.t473 VDD.t860 345.987
R132 VDD.t1051 VDD.t1049 345.987
R133 VDD.t1047 VDD.t1051 345.987
R134 VDD.t16 VDD.t1147 345.987
R135 VDD.t1147 VDD.t667 345.987
R136 VDD.t796 VDD.t849 345.987
R137 VDD.t794 VDD.t796 345.987
R138 VDD.t303 VDD.t85 345.987
R139 VDD.t85 VDD.t665 345.987
R140 VDD.t367 VDD.t369 345.987
R141 VDD.t264 VDD.t367 345.987
R142 VDD.t95 VDD.t506 345.987
R143 VDD.t506 VDD.t1091 345.987
R144 VDD.t549 VDD.t196 345.987
R145 VDD.t557 VDD.t549 345.987
R146 VDD.t903 VDD.t633 345.987
R147 VDD.t633 VDD.t631 345.987
R148 VDD.t653 VDD.t770 345.987
R149 VDD.t945 VDD.t653 345.987
R150 VDD.t836 VDD.t463 345.987
R151 VDD.t463 VDD.t0 345.987
R152 VDD.t1145 VDD.t152 345.987
R153 VDD.t188 VDD.t1145 345.987
R154 VDD.t129 VDD.t1173 345.987
R155 VDD.t1173 VDD.t121 345.987
R156 VDD.t510 VDD.t266 345.987
R157 VDD.t20 VDD.t510 345.987
R158 VDD.t135 VDD.t617 345.987
R159 VDD.t617 VDD.t615 345.987
R160 VDD.t307 VDD.t309 345.987
R161 VDD.t305 VDD.t307 345.987
R162 VDD.t376 VDD.t374 345.987
R163 VDD.t374 VDD.t372 345.987
R164 VDD.t488 VDD.t490 345.987
R165 VDD.t172 VDD.t488 345.987
R166 VDD.t1204 VDD.t750 345.987
R167 VDD.t750 VDD.t748 345.987
R168 VDD.t1169 VDD.t1184 345.987
R169 VDD.t1167 VDD.t1169 345.987
R170 VDD.t204 VDD.t684 345.987
R171 VDD.t684 VDD.t682 345.987
R172 VDD.t527 VDD.t543 345.987
R173 VDD.t529 VDD.t527 345.987
R174 VDD.t1081 VDD.t776 345.987
R175 VDD.t776 VDD.t229 345.987
R176 VDD.t444 VDD.t442 345.987
R177 VDD.t446 VDD.t444 345.987
R178 VDD.t1058 VDD.t1041 345.987
R179 VDD.t1041 VDD.t995 345.987
R180 VDD.t705 VDD.t703 345.987
R181 VDD.t701 VDD.t705 345.987
R182 VDD.t1103 VDD.t786 345.987
R183 VDD.t786 VDD.t659 345.987
R184 VDD.t804 VDD.t217 345.987
R185 VDD.t806 VDD.t804 345.987
R186 VDD.t1105 VDD.t1077 345.987
R187 VDD.t1077 VDD.t975 345.987
R188 VDD.t1128 VDD.t206 345.987
R189 VDD.t208 VDD.t1128 345.987
R190 VDD.t1085 VDD.t884 345.987
R191 VDD.t884 VDD.t784 345.987
R192 VDD.t977 VDD.t758 345.987
R193 VDD.t756 VDD.t977 345.987
R194 VDD.t64 VDD.t1107 345.987
R195 VDD.t1107 VDD.t788 345.987
R196 VDD.t674 VDD.t672 345.987
R197 VDD.t402 VDD.t674 345.987
R198 VDD.t780 VDD.t1060 345.987
R199 VDD.t1060 VDD.t1241 345.987
R200 VDD.t1111 VDD.t1268 345.987
R201 VDD.t1270 VDD.t1111 345.987
R202 VDD.t1258 VDD.t227 345.987
R203 VDD.t227 VDD.t1239 345.987
R204 VDD.t494 VDD.t519 345.987
R205 VDD.t521 VDD.t494 345.987
R206 VDD.t1232 VDD.t1159 345.987
R207 VDD.t1159 VDD.t332 345.987
R208 VDD.t123 VDD.t125 345.987
R209 VDD.t991 VDD.t123 345.987
R210 VDD.t2 VDD.t343 345.987
R211 VDD.t343 VDD.t405 345.987
R212 VDD.t409 VDD.t411 345.987
R213 VDD.t899 VDD.t409 345.987
R214 VDD.t237 VDD.t1209 345.987
R215 VDD.t1209 VDD.t296 345.987
R216 VDD.t1139 VDD.t1141 345.987
R217 VDD.t157 VDD.t1139 345.987
R218 VDD.t161 VDD.t79 345.987
R219 VDD.t79 VDD.t347 345.987
R220 VDD.t1237 VDD.t1176 345.987
R221 VDD.t1178 VDD.t1237 345.987
R222 VDD.t32 VDD.t235 345.987
R223 VDD.t235 VDD.t1207 345.987
R224 VDD.t1221 VDD.t1223 345.987
R225 VDD.t1225 VDD.t1221 345.987
R226 VDD.t663 VDD.t1234 345.987
R227 VDD.t1234 VDD.t469 345.987
R228 VDD.t834 VDD.t830 345.987
R229 VDD.t832 VDD.t834 345.987
R230 VDD.t81 VDD.t349 345.987
R231 VDD.t349 VDD.t14 345.987
R232 VDD.t165 VDD.t167 345.987
R233 VDD.t169 VDD.t165 345.987
R234 VDD.t707 VDD.t427 345.987
R235 VDD.t427 VDD.t87 345.987
R236 VDD.t245 VDD.t247 345.987
R237 VDD.t1190 VDD.t245 345.987
R238 VDD.t1069 VDD.t95 312.28
R239 VDD.t881 VDD.t903 312.28
R240 VDD.t928 VDD.t836 312.28
R241 VDD.t371 VDD.t129 312.28
R242 VDD.t116 VDD.t135 312.28
R243 VDD.t1186 VDD.t376 312.28
R244 VDD.t40 VDD.t1204 312.28
R245 VDD.t221 VDD.t204 312.28
R246 VDD.t55 VDD.t505 276.597
R247 VDD.t8 VDD.t791 276.597
R248 VDD.t243 VDD.t800 276.597
R249 VDD.t57 VDD.t1126 276.597
R250 VDD.t465 VDD.t1156 276.597
R251 VDD.t91 VDD.t579 276.597
R252 VDD.t18 VDD.t968 276.597
R253 VDD.t73 VDD.t956 276.597
R254 VDD.t949 VDD.t589 276.597
R255 VDD.t689 VDD.t253 276.597
R256 VDD.t1079 VDD.t514 276.597
R257 VDD.t951 VDD.t460 276.597
R258 VDD.t997 VDD.t744 276.597
R259 VDD.t953 VDD.t1063 276.597
R260 VDD.t782 VDD.t792 276.597
R261 VDD.t62 VDD.t280 276.597
R262 VDD.t431 VDD.t138 276.597
R263 VDD.t433 VDD.t679 276.597
R264 VDD.t912 VDD.t730 276.597
R265 VDD.t417 VDD.t848 276.597
R266 VDD.t1007 VDD.t838 276.597
R267 VDD.t914 VDD.t1006 276.597
R268 VDD.t1135 VDD.t896 276.597
R269 VDD.t12 VDD.t723 276.597
R270 VDD.t324 VDD.t766 269.594
R271 VDD.t291 VDD.t697 269.594
R272 VDD.t981 VDD.t523 269.594
R273 VDD.t893 VDD.t451 269.594
R274 VDD.t897 VDD.t66 269.594
R275 VDD.t731 VDD.t22 269.594
R276 VDD.t693 VDD.t501 269.594
R277 VDD.t1157 VDD.t1075 269.594
R278 VDD.t726 VDD.t768 269.594
R279 VDD.t457 VDD.t1219 269.594
R280 VDD.t1029 VDD.t461 269.594
R281 VDD.t316 VDD.t563 269.594
R282 VDD.t746 VDD.t101 269.594
R283 VDD.t346 VDD.t754 269.594
R284 VDD.t435 VDD.t734 269.594
R285 VDD.t289 VDD.t415 269.594
R286 VDD.t1236 VDD.t110 269.594
R287 VDD.t587 VDD.t1016 269.594
R288 VDD.t1122 VDD.t59 269.594
R289 VDD.t222 VDD.t400 269.594
R290 VDD.t329 VDD.t1030 269.594
R291 VDD.t760 VDD.t485 269.594
R292 VDD.t929 VDD.t882 269.594
R293 VDD.t185 VDD.t827 269.594
R294 VDD.n329 VDD.n326 258.915
R295 VDD.n309 VDD.n306 258.915
R296 VDD.n249 VDD.n246 258.915
R297 VDD.n229 VDD.n226 258.915
R298 VDD.n190 VDD.n187 258.915
R299 VDD.n209 VDD.n206 258.915
R300 VDD.n269 VDD.n266 258.915
R301 VDD.n289 VDD.n286 258.915
R302 VDD.n488 VDD.n485 258.915
R303 VDD.n468 VDD.n465 258.915
R304 VDD.n408 VDD.n405 258.915
R305 VDD.n388 VDD.n385 258.915
R306 VDD.n349 VDD.n346 258.915
R307 VDD.n368 VDD.n365 258.915
R308 VDD.n428 VDD.n425 258.915
R309 VDD.n448 VDD.n445 258.915
R310 VDD.n647 VDD.n644 258.915
R311 VDD.n627 VDD.n624 258.915
R312 VDD.n567 VDD.n564 258.915
R313 VDD.n547 VDD.n544 258.915
R314 VDD.n508 VDD.n505 258.915
R315 VDD.n527 VDD.n524 258.915
R316 VDD.n587 VDD.n584 258.915
R317 VDD.n607 VDD.n604 258.915
R318 VDD.n332 VDD.n331 258.161
R319 VDD.n312 VDD.n311 258.161
R320 VDD.n252 VDD.n251 258.161
R321 VDD.n232 VDD.n231 258.161
R322 VDD.n193 VDD.n192 258.161
R323 VDD.n212 VDD.n211 258.161
R324 VDD.n272 VDD.n271 258.161
R325 VDD.n292 VDD.n291 258.161
R326 VDD.n491 VDD.n490 258.161
R327 VDD.n471 VDD.n470 258.161
R328 VDD.n411 VDD.n410 258.161
R329 VDD.n391 VDD.n390 258.161
R330 VDD.n352 VDD.n351 258.161
R331 VDD.n371 VDD.n370 258.161
R332 VDD.n431 VDD.n430 258.161
R333 VDD.n451 VDD.n450 258.161
R334 VDD.n650 VDD.n649 258.161
R335 VDD.n630 VDD.n629 258.161
R336 VDD.n570 VDD.n569 258.161
R337 VDD.n550 VDD.n549 258.161
R338 VDD.n511 VDD.n510 258.161
R339 VDD.n530 VDD.n529 258.161
R340 VDD.n590 VDD.n589 258.161
R341 VDD.n610 VDD.n609 258.161
R342 VDD.n1 VDD.n0 222.796
R343 VDD.n15 VDD.n14 222.796
R344 VDD.n29 VDD.n28 222.796
R345 VDD.n41 VDD.n40 222.796
R346 VDD.n70 VDD.n69 222.796
R347 VDD.n84 VDD.n83 222.796
R348 VDD.n56 VDD.n55 222.796
R349 VDD.n108 VDD.n107 222.796
R350 VDD.t394 VDD.t935 196.666
R351 VDD.t645 VDD.t394 196.666
R352 VDD.t1252 VDD.t645 196.666
R353 VDD.t1188 VDD.t1252 196.666
R354 VDD.t26 VDD.t1188 196.666
R355 VDD.t258 VDD.t1055 196.666
R356 VDD.t1055 VDD.t105 196.666
R357 VDD.t717 VDD.t721 196.666
R358 VDD.t719 VDD.t717 196.666
R359 VDD.t555 VDD.t719 196.666
R360 VDD.t1247 VDD.t555 196.666
R361 VDD.t559 VDD.t1247 196.666
R362 VDD.t148 VDD.t448 196.666
R363 VDD.t448 VDD.t144 196.666
R364 VDD.t576 VDD.t574 196.666
R365 VDD.t499 VDD.t576 196.666
R366 VDD.t512 VDD.t499 196.666
R367 VDD.t593 VDD.t512 196.666
R368 VDD.t174 VDD.t593 196.666
R369 VDD.t879 VDD.t497 196.666
R370 VDD.t497 VDD.t961 196.666
R371 VDD.t1089 VDD.t1087 196.666
R372 VDD.t1066 VDD.t1089 196.666
R373 VDD.t1194 VDD.t1066 196.666
R374 VDD.t1266 VDD.t1194 196.666
R375 VDD.t1095 VDD.t1266 196.666
R376 VDD.t319 VDD.t901 196.666
R377 VDD.t901 VDD.t931 196.666
R378 VDD.t728 VDD.t621 196.666
R379 VDD.t1192 VDD.t728 196.666
R380 VDD.t539 VDD.t1192 196.666
R381 VDD.t531 VDD.t539 196.666
R382 VDD.t533 VDD.t531 196.666
R383 VDD.t254 VDD.t325 196.666
R384 VDD.t325 VDD.t979 196.666
R385 VDD.t1137 VDD.t605 196.666
R386 VDD.t603 VDD.t1137 196.666
R387 VDD.t385 VDD.t603 196.666
R388 VDD.t844 VDD.t385 196.666
R389 VDD.t1182 VDD.t844 196.666
R390 VDD.t643 VDD.t397 196.666
R391 VDD.t397 VDD.t647 196.666
R392 VDD.t131 VDD.t98 196.666
R393 VDD.t133 VDD.t131 196.666
R394 VDD.t515 VDD.t133 196.666
R395 VDD.t920 VDD.t515 196.666
R396 VDD.t597 VDD.t920 196.666
R397 VDD.t478 VDD.t365 196.666
R398 VDD.t365 VDD.t958 196.666
R399 VDD.t695 VDD.t609 196.666
R400 VDD.t715 VDD.t695 196.666
R401 VDD.t357 VDD.t715 196.666
R402 VDD.t508 VDD.t357 196.666
R403 VDD.t270 VDD.t508 196.666
R404 VDD.t1171 VDD.t119 196.666
R405 VDD.t119 VDD.t389 196.666
R406 VDD.t1249 VDD.t580 191.952
R407 VDD.t1249 VDD.t582 191.952
R408 VDD.t988 VDD.t1003 190
R409 VDD.t988 VDD.t1001 190
R410 VDD.n334 VDD.n333 184.375
R411 VDD.n314 VDD.n313 184.375
R412 VDD.n254 VDD.n253 184.375
R413 VDD.n234 VDD.n233 184.375
R414 VDD.n195 VDD.n194 184.375
R415 VDD.n214 VDD.n213 184.375
R416 VDD.n274 VDD.n273 184.375
R417 VDD.n294 VDD.n293 184.375
R418 VDD.n493 VDD.n492 184.375
R419 VDD.n473 VDD.n472 184.375
R420 VDD.n413 VDD.n412 184.375
R421 VDD.n393 VDD.n392 184.375
R422 VDD.n354 VDD.n353 184.375
R423 VDD.n373 VDD.n372 184.375
R424 VDD.n433 VDD.n432 184.375
R425 VDD.n453 VDD.n452 184.375
R426 VDD.n652 VDD.n651 184.375
R427 VDD.n632 VDD.n631 184.375
R428 VDD.n572 VDD.n571 184.375
R429 VDD.n552 VDD.n551 184.375
R430 VDD.n513 VDD.n512 184.375
R431 VDD.n532 VDD.n531 184.375
R432 VDD.n592 VDD.n591 184.375
R433 VDD.n612 VDD.n611 184.375
R434 VDD.n325 VDD.n324 182.117
R435 VDD.n305 VDD.n304 182.117
R436 VDD.n245 VDD.n244 182.117
R437 VDD.n225 VDD.n224 182.117
R438 VDD.n186 VDD.n185 182.117
R439 VDD.n205 VDD.n204 182.117
R440 VDD.n265 VDD.n264 182.117
R441 VDD.n285 VDD.n284 182.117
R442 VDD.n484 VDD.n483 182.117
R443 VDD.n464 VDD.n463 182.117
R444 VDD.n404 VDD.n403 182.117
R445 VDD.n384 VDD.n383 182.117
R446 VDD.n345 VDD.n344 182.117
R447 VDD.n364 VDD.n363 182.117
R448 VDD.n424 VDD.n423 182.117
R449 VDD.n444 VDD.n443 182.117
R450 VDD.n643 VDD.n642 182.117
R451 VDD.n623 VDD.n622 182.117
R452 VDD.n563 VDD.n562 182.117
R453 VDD.n543 VDD.n542 182.117
R454 VDD.n504 VDD.n503 182.117
R455 VDD.n523 VDD.n522 182.117
R456 VDD.n583 VDD.n582 182.117
R457 VDD.n603 VDD.n602 182.117
R458 VDD.n864 VDD.t1143 174.172
R459 VDD.n870 VDD.t1117 173.061
R460 VDD.n900 VDD.t43 172.51
R461 VDD.n894 VDD.t623 172.51
R462 VDD.n888 VDD.t676 172.51
R463 VDD.n882 VDD.t964 172.51
R464 VDD.n876 VDD.t810 172.51
R465 VDD.n858 VDD.t287 172.51
R466 VDD.n863 VDD.t738 170.712
R467 VDD.n702 VDD.t194 170.677
R468 VDD.n802 VDD.t1196 170.677
R469 VDD.n677 VDD.t142 170.677
R470 VDD.n727 VDD.t272 170.677
R471 VDD.n752 VDD.t517 170.677
R472 VDD.n777 VDD.t595 170.677
R473 VDD.n827 VDD.t103 170.677
R474 VDD.n852 VDD.t535 170.677
R475 VDD.n869 VDD.t381 169.626
R476 VDD.n899 VDD.t45 169.088
R477 VDD.n893 VDD.t649 169.088
R478 VDD.n887 VDD.t637 169.088
R479 VDD.n881 VDD.t566 169.088
R480 VDD.n875 VDD.t481 169.088
R481 VDD.n857 VDD.t680 169.088
R482 VDD.n703 VDD.n702 151.379
R483 VDD.n803 VDD.n802 151.379
R484 VDD.n678 VDD.n677 151.379
R485 VDD.n728 VDD.n727 151.379
R486 VDD.n753 VDD.n752 151.379
R487 VDD.n778 VDD.n777 151.379
R488 VDD.n828 VDD.n827 151.379
R489 VDD.n853 VDD.n852 151.379
R490 VDD.t1245 VDD.t847 144.087
R491 VDD.t847 VDD.t109 144.087
R492 VDD.t109 VDD.t97 144.087
R493 VDD.t599 VDD.t216 144.087
R494 VDD.t216 VDD.t480 144.087
R495 VDD.t480 VDD.t137 144.087
R496 VDD.t669 VDD.t963 144.087
R497 VDD.t963 VDD.t496 144.087
R498 VDD.t496 VDD.t960 144.087
R499 VDD.t383 VDD.t263 144.087
R500 VDD.t263 VDD.t1206 144.087
R501 VDD.t1206 VDD.t642 144.087
R502 VDD.t886 VDD.t100 144.087
R503 VDD.t100 VDD.t727 144.087
R504 VDD.t727 VDD.t331 144.087
R505 VDD.t268 VDD.t391 143.717
R506 VDD.t391 VDD.t118 143.717
R507 VDD.t118 VDD.t380 143.717
R508 VDD.t537 VDD.t686 143.717
R509 VDD.t686 VDD.t1020 143.717
R510 VDD.t1020 VDD.t203 143.717
R511 VDD.t651 VDD.t321 143.717
R512 VDD.t321 VDD.t641 143.717
R513 VDD.t641 VDD.t1036 143.717
R514 VDD.n1 VDD.t1245 137.982
R515 VDD.n29 VDD.t599 137.982
R516 VDD.n41 VDD.t669 137.982
R517 VDD.n70 VDD.t383 137.982
R518 VDD.n107 VDD.t886 137.982
R519 VDD.t852 VDD.t851 137.714
R520 VDD.t505 VDD.t852 137.714
R521 VDD.t301 VDD.t55 137.714
R522 VDD.t938 VDD.t324 137.714
R523 VDD.t766 VDD.t762 137.714
R524 VDD.t762 VDD.t764 137.714
R525 VDD.t487 VDD.t1057 137.714
R526 VDD.t791 VDD.t487 137.714
R527 VDD.t34 VDD.t8 137.714
R528 VDD.t911 VDD.t291 137.714
R529 VDD.t697 VDD.t1053 137.714
R530 VDD.t1053 VDD.t1133 137.714
R531 VDD.t1161 VDD.t801 137.714
R532 VDD.t800 VDD.t1161 137.714
R533 VDD.t233 VDD.t243 137.714
R534 VDD.t790 VDD.t981 137.714
R535 VDD.t523 VDD.t874 137.714
R536 VDD.t874 VDD.t876 137.714
R537 VDD.t68 VDD.t69 137.714
R538 VDD.t1126 VDD.t68 137.714
R539 VDD.t336 VDD.t57 137.714
R540 VDD.t450 VDD.t893 137.714
R541 VDD.t451 VDD.t458 137.714
R542 VDD.t458 VDD.t1109 137.714
R543 VDD.t338 VDD.t1155 137.714
R544 VDD.t1156 VDD.t338 137.714
R545 VDD.t438 VDD.t465 137.714
R546 VDD.t588 VDD.t897 137.714
R547 VDD.t66 VDD.t983 137.714
R548 VDD.t983 VDD.t154 137.714
R549 VDD.t846 VDD.t578 137.714
R550 VDD.t579 VDD.t846 137.714
R551 VDD.t475 VDD.t91 137.714
R552 VDD.t994 VDD.t731 137.714
R553 VDD.t22 VDD.t24 137.714
R554 VDD.t24 VDD.t840 137.714
R555 VDD.t970 VDD.t969 137.714
R556 VDD.t968 VDD.t970 137.714
R557 VDD.t1149 VDD.t18 137.714
R558 VDD.t176 VDD.t693 137.714
R559 VDD.t501 VDD.t503 137.714
R560 VDD.t503 VDD.t585 137.714
R561 VDD.t477 VDD.t957 137.714
R562 VDD.t956 VDD.t477 137.714
R563 VDD.t341 VDD.t73 137.714
R564 VDD.t700 VDD.t1157 137.714
R565 VDD.t1075 VDD.t1071 137.714
R566 VDD.t1071 VDD.t1073 137.714
R567 VDD.t300 VDD.t590 137.714
R568 VDD.t589 VDD.t300 137.714
R569 VDD.t1099 VDD.t949 137.714
R570 VDD.t314 VDD.t726 137.714
R571 VDD.t768 VDD.t190 137.714
R572 VDD.t190 VDD.t192 137.714
R573 VDD.t393 VDD.t392 137.714
R574 VDD.t253 VDD.t393 137.714
R575 VDD.t778 VDD.t689 137.714
R576 VDD.t184 VDD.t457 137.714
R577 VDD.t1219 VDD.t1215 137.714
R578 VDD.t1215 VDD.t1217 137.714
R579 VDD.t362 VDD.t361 137.714
R580 VDD.t514 VDD.t362 137.714
R581 VDD.t774 VDD.t1079 137.714
R582 VDD.t829 VDD.t1029 137.714
R583 VDD.t461 VDD.t223 137.714
R584 VDD.t223 VDD.t225 137.714
R585 VDD.t993 VDD.t1034 137.714
R586 VDD.t460 VDD.t993 137.714
R587 VDD.t999 VDD.t951 137.714
R588 VDD.t250 VDD.t316 137.714
R589 VDD.t563 VDD.t181 137.714
R590 VDD.t181 VDD.t561 137.714
R591 VDD.t745 VDD.t743 137.714
R592 VDD.t744 VDD.t745 137.714
R593 VDD.t1264 VDD.t997 137.714
R594 VDD.t584 VDD.t746 137.714
R595 VDD.t101 VDD.t825 137.714
R596 VDD.t825 VDD.t889 137.714
R597 VDD.t1064 VDD.t1062 137.714
R598 VDD.t1063 VDD.t1064 137.714
R599 VDD.t1260 VDD.t953 137.714
R600 VDD.t345 VDD.t346 137.714
R601 VDD.t754 VDD.t1123 137.714
R602 VDD.t1123 VDD.t752 137.714
R603 VDD.t1158 VDD.t793 137.714
R604 VDD.t792 VDD.t1158 137.714
R605 VDD.t1083 VDD.t782 137.714
R606 VDD.t990 VDD.t435 137.714
R607 VDD.t734 VDD.t736 137.714
R608 VDD.t736 VDD.t732 137.714
R609 VDD.t565 VDD.t281 137.714
R610 VDD.t280 VDD.t565 137.714
R611 VDD.t691 VDD.t62 137.714
R612 VDD.t290 VDD.t289 137.714
R613 VDD.t415 VDD.t1043 137.714
R614 VDD.t1043 VDD.t413 137.714
R615 VDD.t926 VDD.t927 137.714
R616 VDD.t138 VDD.t926 137.714
R617 VDD.t467 VDD.t431 137.714
R618 VDD.t198 VDD.t1236 137.714
R619 VDD.t110 VDD.t285 137.714
R620 VDD.t285 VDD.t283 137.714
R621 VDD.t318 VDD.t678 137.714
R622 VDD.t679 VDD.t318 137.714
R623 VDD.t351 VDD.t433 137.714
R624 VDD.t429 VDD.t587 137.714
R625 VDD.t1016 VDD.t655 137.714
R626 VDD.t655 VDD.t107 137.714
R627 VDD.t330 VDD.t141 137.714
R628 VDD.t730 VDD.t330 137.714
R629 VDD.t38 VDD.t912 137.714
R630 VDD.t219 VDD.t1122 137.714
R631 VDD.t59 VDD.t28 137.714
R632 VDD.t28 VDD.t70 137.714
R633 VDD.t854 VDD.t853 137.714
R634 VDD.t848 VDD.t854 137.714
R635 VDD.t75 VDD.t417 137.714
R636 VDD.t251 VDD.t222 137.714
R637 VDD.t400 VDD.t1213 137.714
R638 VDD.t1213 VDD.t1045 137.714
R639 VDD.t839 VDD.t399 137.714
R640 VDD.t838 VDD.t839 137.714
R641 VDD.t298 VDD.t1007 137.714
R642 VDD.t31 VDD.t329 137.714
R643 VDD.t1030 VDD.t41 137.714
R644 VDD.t41 VDD.t1032 137.714
R645 VDD.t1065 VDD.t1005 137.714
R646 VDD.t1006 VDD.t1065 137.714
R647 VDD.t294 VDD.t914 137.714
R648 VDD.t761 VDD.t760 137.714
R649 VDD.t485 VDD.t483 137.714
R650 VDD.t483 VDD.t1164 137.714
R651 VDD.t404 VDD.t895 137.714
R652 VDD.t896 VDD.t404 137.714
R653 VDD.t407 VDD.t1135 137.714
R654 VDD.t930 VDD.t929 137.714
R655 VDD.t882 VDD.t1120 137.714
R656 VDD.t1120 VDD.t740 137.714
R657 VDD.t724 VDD.t855 137.714
R658 VDD.t723 VDD.t724 137.714
R659 VDD.t425 VDD.t12 137.714
R660 VDD.t202 VDD.t185 137.714
R661 VDD.t827 VDD.t1200 137.714
R662 VDD.t1200 VDD.t1198 137.714
R663 VDD.n15 VDD.t268 137.628
R664 VDD.n84 VDD.t537 137.628
R665 VDD.n56 VDD.t651 137.628
R666 VDD.n319 VDD.t938 136.641
R667 VDD.n299 VDD.t911 136.641
R668 VDD.n239 VDD.t790 136.641
R669 VDD.n219 VDD.t450 136.641
R670 VDD.n180 VDD.t588 136.641
R671 VDD.n199 VDD.t994 136.641
R672 VDD.n259 VDD.t176 136.641
R673 VDD.n279 VDD.t700 136.641
R674 VDD.n478 VDD.t314 136.641
R675 VDD.n458 VDD.t184 136.641
R676 VDD.n398 VDD.t829 136.641
R677 VDD.n378 VDD.t250 136.641
R678 VDD.n339 VDD.t584 136.641
R679 VDD.n358 VDD.t345 136.641
R680 VDD.n418 VDD.t990 136.641
R681 VDD.n438 VDD.t290 136.641
R682 VDD.n637 VDD.t198 136.641
R683 VDD.n617 VDD.t429 136.641
R684 VDD.n557 VDD.t219 136.641
R685 VDD.n537 VDD.t251 136.641
R686 VDD.n498 VDD.t31 136.641
R687 VDD.n517 VDD.t761 136.641
R688 VDD.n577 VDD.t930 136.641
R689 VDD.n597 VDD.t202 136.641
R690 VDD.n322 VDD.t301 120.208
R691 VDD.n302 VDD.t34 120.208
R692 VDD.n242 VDD.t233 120.208
R693 VDD.n222 VDD.t336 120.208
R694 VDD.n183 VDD.t438 120.208
R695 VDD.n202 VDD.t475 120.208
R696 VDD.n262 VDD.t1149 120.208
R697 VDD.n282 VDD.t341 120.208
R698 VDD.n481 VDD.t1099 120.208
R699 VDD.n461 VDD.t778 120.208
R700 VDD.n401 VDD.t774 120.208
R701 VDD.n381 VDD.t999 120.208
R702 VDD.n342 VDD.t1264 120.208
R703 VDD.n361 VDD.t1260 120.208
R704 VDD.n421 VDD.t1083 120.208
R705 VDD.n441 VDD.t691 120.208
R706 VDD.n640 VDD.t467 120.208
R707 VDD.n620 VDD.t351 120.208
R708 VDD.n560 VDD.t38 120.208
R709 VDD.n540 VDD.t75 120.208
R710 VDD.n501 VDD.t298 120.208
R711 VDD.n520 VDD.t294 120.208
R712 VDD.n580 VDD.t407 120.208
R713 VDD.n600 VDD.t425 120.208
R714 VDD.n702 VDD.n701 115.932
R715 VDD.n802 VDD.n801 115.932
R716 VDD.n677 VDD.n676 115.932
R717 VDD.n727 VDD.n726 115.932
R718 VDD.n752 VDD.n751 115.932
R719 VDD.n777 VDD.n776 115.932
R720 VDD.n827 VDD.n826 115.932
R721 VDD.n852 VDD.n851 115.932
R722 VDD.n328 VDD.n327 85.695
R723 VDD.n308 VDD.n307 85.695
R724 VDD.n248 VDD.n247 85.695
R725 VDD.n228 VDD.n227 85.695
R726 VDD.n189 VDD.n188 85.695
R727 VDD.n208 VDD.n207 85.695
R728 VDD.n268 VDD.n267 85.695
R729 VDD.n288 VDD.n287 85.695
R730 VDD.n487 VDD.n486 85.695
R731 VDD.n467 VDD.n466 85.695
R732 VDD.n407 VDD.n406 85.695
R733 VDD.n387 VDD.n386 85.695
R734 VDD.n348 VDD.n347 85.695
R735 VDD.n367 VDD.n366 85.695
R736 VDD.n427 VDD.n426 85.695
R737 VDD.n447 VDD.n446 85.695
R738 VDD.n646 VDD.n645 85.695
R739 VDD.n626 VDD.n625 85.695
R740 VDD.n566 VDD.n565 85.695
R741 VDD.n546 VDD.n545 85.695
R742 VDD.n507 VDD.n506 85.695
R743 VDD.n526 VDD.n525 85.695
R744 VDD.n586 VDD.n585 85.695
R745 VDD.n606 VDD.n605 85.695
R746 VDD.n2 VDD.t553 61.054
R747 VDD.n30 VDD.t127 61.054
R748 VDD.n42 VDD.t492 61.054
R749 VDD.n71 VDD.t842 61.054
R750 VDD.t1202 VDD.n106 61.054
R751 VDD.n16 VDD.t359 60.898
R752 VDD.n85 VDD.t541 60.898
R753 VDD.n57 VDD.t661 60.898
R754 VDD.t916 VDD.n321 58.354
R755 VDD.t10 VDD.n301 58.354
R756 VDD.t471 VDD.n241 58.354
R757 VDD.t436 VDD.n221 58.354
R758 VDD.t421 VDD.n182 58.354
R759 VDD.t53 VDD.n201 58.354
R760 VDD.t440 VDD.n261 58.354
R761 VDD.t918 VDD.n281 58.354
R762 VDD.t657 VDD.n480 58.354
R763 VDD.t231 VDD.n460 58.354
R764 VDD.t1262 VDD.n400 58.354
R765 VDD.t1037 VDD.n380 58.354
R766 VDD.t687 VDD.n341 58.354
R767 VDD.t947 VDD.n360 58.354
R768 VDD.t1039 VDD.n420 58.354
R769 VDD.t1101 VDD.n440 58.354
R770 VDD.t334 VDD.n639 58.354
R771 VDD.t93 VDD.n619 58.354
R772 VDD.t423 VDD.n559 58.354
R773 VDD.t339 VDD.n539 58.354
R774 VDD.t1011 VDD.n500 58.354
R775 VDD.t36 VDD.n519 58.354
R776 VDD.t353 VDD.n579 58.354
R777 VDD.t6 VDD.n599 58.354
R778 VDD.t725 VDD.t194 53.244
R779 VDD.t139 VDD.t1069 53.244
R780 VDD.t396 VDD.t1196 53.244
R781 VDD.t639 VDD.t881 53.244
R782 VDD.t812 VDD.t142 53.244
R783 VDD.t607 VDD.t928 53.244
R784 VDD.t742 VDD.t272 53.244
R785 VDD.t1180 VDD.t371 53.244
R786 VDD.t982 VDD.t517 53.244
R787 VDD.t311 VDD.t116 53.244
R788 VDD.t1227 VDD.t595 53.244
R789 VDD.t966 VDD.t1186 53.244
R790 VDD.t1166 VDD.t103 53.244
R791 VDD.t619 VDD.t40 53.244
R792 VDD.t891 VDD.t535 53.244
R793 VDD.t1018 VDD.t221 53.244
R794 VDD.t551 VDD.n697 44.17
R795 VDD.t194 VDD.n698 44.17
R796 VDD.n700 VDD.t611 44.17
R797 VDD.n699 VDD.t139 44.17
R798 VDD.t327 VDD.n797 44.17
R799 VDD.t1196 VDD.n798 44.17
R800 VDD.n800 VDD.t322 44.17
R801 VDD.n799 VDD.t639 44.17
R802 VDD.t146 VDD.n672 44.17
R803 VDD.t142 VDD.n673 44.17
R804 VDD.n675 VDD.t210 44.17
R805 VDD.n674 VDD.t607 44.17
R806 VDD.t274 VDD.n722 44.17
R807 VDD.t272 VDD.n723 44.17
R808 VDD.n725 VDD.t1228 44.17
R809 VDD.n724 VDD.t1180 44.17
R810 VDD.t601 VDD.n747 44.17
R811 VDD.t517 VDD.n748 44.17
R812 VDD.n750 VDD.t808 44.17
R813 VDD.n749 VDD.t311 44.17
R814 VDD.t177 VDD.n772 44.17
R815 VDD.t595 VDD.n773 44.17
R816 VDD.n775 VDD.t568 44.17
R817 VDD.n774 VDD.t966 44.17
R818 VDD.t1130 VDD.n822 44.17
R819 VDD.t103 VDD.n823 44.17
R820 VDD.n825 VDD.t625 44.17
R821 VDD.n824 VDD.t619 44.17
R822 VDD.t525 VDD.n847 44.17
R823 VDD.t535 VDD.n848 44.17
R824 VDD.n850 VDD.t1021 44.17
R825 VDD.n849 VDD.t1018 44.17
R826 VDD.n698 VDD.t551 41.273
R827 VDD.t1013 VDD.n700 41.273
R828 VDD.t611 VDD.n699 41.273
R829 VDD.n697 VDD.t1243 41.273
R830 VDD.n798 VDD.t327 41.273
R831 VDD.t933 VDD.n800 41.273
R832 VDD.t322 VDD.n799 41.273
R833 VDD.n797 VDD.t1093 41.273
R834 VDD.n673 VDD.t146 41.273
R835 VDD.t212 VDD.n675 41.273
R836 VDD.t210 VDD.n674 41.273
R837 VDD.n672 VDD.t1097 41.273
R838 VDD.n723 VDD.t274 41.273
R839 VDD.t1230 VDD.n725 41.273
R840 VDD.t1228 VDD.n724 41.273
R841 VDD.n722 VDD.t276 41.273
R842 VDD.n748 VDD.t601 41.273
R843 VDD.t378 VDD.n750 41.273
R844 VDD.t808 VDD.n749 41.273
R845 VDD.n747 VDD.t922 41.273
R846 VDD.n773 VDD.t177 41.273
R847 VDD.t572 VDD.n775 41.273
R848 VDD.t568 VDD.n774 41.273
R849 VDD.n772 VDD.t179 41.273
R850 VDD.n823 VDD.t1130 41.273
R851 VDD.t261 VDD.n825 41.273
R852 VDD.t625 VDD.n824 41.273
R853 VDD.n822 VDD.t866 41.273
R854 VDD.n848 VDD.t525 41.273
R855 VDD.t256 VDD.n850 41.273
R856 VDD.t1021 VDD.n849 41.273
R857 VDD.n847 VDD.t545 41.273
R858 VDD.n45 VDD.n44 41.219
R859 VDD.n6 VDD.n5 37.853
R860 VDD.n32 VDD.t1249 37.853
R861 VDD.n47 VDD.n46 37.853
R862 VDD.n75 VDD.n74 37.853
R863 VDD.t988 VDD.n104 37.853
R864 VDD.n20 VDD.n19 37.756
R865 VDD.n89 VDD.n88 37.756
R866 VDD.n61 VDD.n60 37.756
R867 VDD.n179 VDD.t106 30.163
R868 VDD.n171 VDD.t145 30.163
R869 VDD.n147 VDD.t962 30.163
R870 VDD.n139 VDD.t932 30.163
R871 VDD.n123 VDD.t980 30.163
R872 VDD.n131 VDD.t648 30.163
R873 VDD.n155 VDD.t959 30.163
R874 VDD.n163 VDD.t390 30.163
R875 VDD.n701 VDD.t725 29.891
R876 VDD.n801 VDD.t396 29.891
R877 VDD.n676 VDD.t812 29.891
R878 VDD.n726 VDD.t742 29.891
R879 VDD.n751 VDD.t982 29.891
R880 VDD.n776 VDD.t1227 29.891
R881 VDD.n826 VDD.t1166 29.891
R882 VDD.n851 VDD.t891 29.891
R883 VDD.n5 VDD.n3 29.305
R884 VDD.t1249 VDD.n31 29.305
R885 VDD.n46 VDD.n43 29.305
R886 VDD.n74 VDD.n72 29.305
R887 VDD.n105 VDD.t988 29.305
R888 VDD.n19 VDD.n17 29.23
R889 VDD.n88 VDD.n86 29.23
R890 VDD.n60 VDD.n58 29.23
R891 VDD.n903 VDD.t46 29.208
R892 VDD.n897 VDD.t650 29.208
R893 VDD.n891 VDD.t638 29.208
R894 VDD.n885 VDD.t567 29.208
R895 VDD.n879 VDD.t482 29.208
R896 VDD.n861 VDD.t681 29.208
R897 VDD.n873 VDD.t382 29.202
R898 VDD.n867 VDD.t739 29.191
R899 VDD.n684 VDD.t96 28.664
R900 VDD.n691 VDD.t558 28.664
R901 VDD.n784 VDD.t904 28.664
R902 VDD.n791 VDD.t946 28.664
R903 VDD.n659 VDD.t837 28.664
R904 VDD.n666 VDD.t189 28.664
R905 VDD.n709 VDD.t130 28.664
R906 VDD.n716 VDD.t21 28.664
R907 VDD.n734 VDD.t136 28.664
R908 VDD.n741 VDD.t306 28.664
R909 VDD.n759 VDD.t377 28.664
R910 VDD.n766 VDD.t173 28.664
R911 VDD.n809 VDD.t1205 28.664
R912 VDD.n816 VDD.t1168 28.664
R913 VDD.n834 VDD.t205 28.664
R914 VDD.n841 VDD.t530 28.664
R915 VDD.n9 VDD.t364 28.57
R916 VDD.n23 VDD.t1163 28.57
R917 VDD.n35 VDD.t581 28.57
R918 VDD.n50 VDD.t869 28.57
R919 VDD.n78 VDD.t986 28.57
R920 VDD.n92 VDD.t113 28.57
R921 VDD.n64 VDD.t1026 28.57
R922 VDD.n110 VDD.t1004 28.57
R923 VDD.n334 VDD.t78 28.568
R924 VDD.n314 VDD.t48 28.568
R925 VDD.n254 VDD.t630 28.568
R926 VDD.n234 VDD.t909 28.568
R927 VDD.n195 VDD.t1255 28.568
R928 VDD.n214 VDD.t1048 28.568
R929 VDD.n274 VDD.t795 28.568
R930 VDD.n294 VDD.t265 28.568
R931 VDD.n493 VDD.t447 28.568
R932 VDD.n473 VDD.t702 28.568
R933 VDD.n413 VDD.t807 28.568
R934 VDD.n393 VDD.t209 28.568
R935 VDD.n354 VDD.t757 28.568
R936 VDD.n373 VDD.t403 28.568
R937 VDD.n433 VDD.t1271 28.568
R938 VDD.n453 VDD.t522 28.568
R939 VDD.n652 VDD.t992 28.568
R940 VDD.n632 VDD.t900 28.568
R941 VDD.n572 VDD.t158 28.568
R942 VDD.n552 VDD.t1179 28.568
R943 VDD.n513 VDD.t1226 28.568
R944 VDD.n532 VDD.t833 28.568
R945 VDD.n592 VDD.t170 28.568
R946 VDD.n612 VDD.t1191 28.568
R947 VDD.n178 VDD.t259 28.565
R948 VDD.n178 VDD.t1056 28.565
R949 VDD.n173 VDD.t936 28.565
R950 VDD.n173 VDD.t395 28.565
R951 VDD.n174 VDD.t646 28.565
R952 VDD.n174 VDD.t1253 28.565
R953 VDD.n176 VDD.t1189 28.565
R954 VDD.n176 VDD.t27 28.565
R955 VDD.n170 VDD.t149 28.565
R956 VDD.n170 VDD.t449 28.565
R957 VDD.n165 VDD.t722 28.565
R958 VDD.n165 VDD.t718 28.565
R959 VDD.n166 VDD.t720 28.565
R960 VDD.n166 VDD.t556 28.565
R961 VDD.n168 VDD.t1248 28.565
R962 VDD.n168 VDD.t560 28.565
R963 VDD.n146 VDD.t880 28.565
R964 VDD.n146 VDD.t498 28.565
R965 VDD.n141 VDD.t575 28.565
R966 VDD.n141 VDD.t577 28.565
R967 VDD.n142 VDD.t500 28.565
R968 VDD.n142 VDD.t513 28.565
R969 VDD.n144 VDD.t594 28.565
R970 VDD.n144 VDD.t175 28.565
R971 VDD.n138 VDD.t320 28.565
R972 VDD.n138 VDD.t902 28.565
R973 VDD.n133 VDD.t1088 28.565
R974 VDD.n133 VDD.t1090 28.565
R975 VDD.n134 VDD.t1067 28.565
R976 VDD.n134 VDD.t1195 28.565
R977 VDD.n136 VDD.t1267 28.565
R978 VDD.n136 VDD.t1096 28.565
R979 VDD.n122 VDD.t255 28.565
R980 VDD.n122 VDD.t326 28.565
R981 VDD.n117 VDD.t622 28.565
R982 VDD.n117 VDD.t729 28.565
R983 VDD.n118 VDD.t1193 28.565
R984 VDD.n118 VDD.t540 28.565
R985 VDD.n120 VDD.t532 28.565
R986 VDD.n120 VDD.t534 28.565
R987 VDD.n130 VDD.t644 28.565
R988 VDD.n130 VDD.t398 28.565
R989 VDD.n125 VDD.t606 28.565
R990 VDD.n125 VDD.t1138 28.565
R991 VDD.n126 VDD.t604 28.565
R992 VDD.n126 VDD.t386 28.565
R993 VDD.n128 VDD.t845 28.565
R994 VDD.n128 VDD.t1183 28.565
R995 VDD.n154 VDD.t479 28.565
R996 VDD.n154 VDD.t366 28.565
R997 VDD.n149 VDD.t99 28.565
R998 VDD.n149 VDD.t132 28.565
R999 VDD.n150 VDD.t134 28.565
R1000 VDD.n150 VDD.t516 28.565
R1001 VDD.n152 VDD.t921 28.565
R1002 VDD.n152 VDD.t598 28.565
R1003 VDD.n162 VDD.t1172 28.565
R1004 VDD.n162 VDD.t120 28.565
R1005 VDD.n157 VDD.t610 28.565
R1006 VDD.n157 VDD.t696 28.565
R1007 VDD.n158 VDD.t716 28.565
R1008 VDD.n158 VDD.t358 28.565
R1009 VDD.n160 VDD.t509 28.565
R1010 VDD.n160 VDD.t271 28.565
R1011 VDD.n333 VDD.t815 28.565
R1012 VDD.n333 VDD.t817 28.565
R1013 VDD.n324 VDD.t160 28.565
R1014 VDD.n324 VDD.t84 28.565
R1015 VDD.n327 VDD.t164 28.565
R1016 VDD.n313 VDD.t50 28.565
R1017 VDD.n313 VDD.t52 28.565
R1018 VDD.n304 VDD.t803 28.565
R1019 VDD.n304 VDD.t5 28.565
R1020 VDD.n307 VDD.t714 28.565
R1021 VDD.n253 VDD.t972 28.565
R1022 VDD.n253 VDD.t628 28.565
R1023 VDD.n244 VDD.t859 28.565
R1024 VDD.n244 VDD.t857 28.565
R1025 VDD.n247 VDD.t1010 28.565
R1026 VDD.n233 VDD.t907 28.565
R1027 VDD.n233 VDD.t799 28.565
R1028 VDD.n224 VDD.t240 28.565
R1029 VDD.n224 VDD.t710 28.565
R1030 VDD.n227 VDD.t863 28.565
R1031 VDD.n194 VDD.t1257 28.565
R1032 VDD.n194 VDD.t944 28.565
R1033 VDD.n185 VDD.t712 28.565
R1034 VDD.n185 VDD.t356 28.565
R1035 VDD.n188 VDD.t242 28.565
R1036 VDD.n213 VDD.t1050 28.565
R1037 VDD.n213 VDD.t1052 28.565
R1038 VDD.n204 VDD.t474 28.565
R1039 VDD.n204 VDD.t861 28.565
R1040 VDD.n207 VDD.t420 28.565
R1041 VDD.n273 VDD.t850 28.565
R1042 VDD.n273 VDD.t797 28.565
R1043 VDD.n264 VDD.t1148 28.565
R1044 VDD.n264 VDD.t668 28.565
R1045 VDD.n267 VDD.t17 28.565
R1046 VDD.n293 VDD.t370 28.565
R1047 VDD.n293 VDD.t368 28.565
R1048 VDD.n284 VDD.t86 28.565
R1049 VDD.n284 VDD.t666 28.565
R1050 VDD.n287 VDD.t304 28.565
R1051 VDD.n685 VDD.t507 28.565
R1052 VDD.n685 VDD.t1092 28.565
R1053 VDD.n692 VDD.t197 28.565
R1054 VDD.n692 VDD.t550 28.565
R1055 VDD.n785 VDD.t634 28.565
R1056 VDD.n785 VDD.t632 28.565
R1057 VDD.n792 VDD.t771 28.565
R1058 VDD.n792 VDD.t654 28.565
R1059 VDD.n660 VDD.t464 28.565
R1060 VDD.n660 VDD.t1 28.565
R1061 VDD.n667 VDD.t153 28.565
R1062 VDD.n667 VDD.t1146 28.565
R1063 VDD.n710 VDD.t1174 28.565
R1064 VDD.n710 VDD.t122 28.565
R1065 VDD.n717 VDD.t267 28.565
R1066 VDD.n717 VDD.t511 28.565
R1067 VDD.n735 VDD.t618 28.565
R1068 VDD.n735 VDD.t616 28.565
R1069 VDD.n742 VDD.t310 28.565
R1070 VDD.n742 VDD.t308 28.565
R1071 VDD.n760 VDD.t375 28.565
R1072 VDD.n760 VDD.t373 28.565
R1073 VDD.n767 VDD.t491 28.565
R1074 VDD.n767 VDD.t489 28.565
R1075 VDD.n810 VDD.t751 28.565
R1076 VDD.n810 VDD.t749 28.565
R1077 VDD.n817 VDD.t1185 28.565
R1078 VDD.n817 VDD.t1170 28.565
R1079 VDD.n835 VDD.t685 28.565
R1080 VDD.n835 VDD.t683 28.565
R1081 VDD.n842 VDD.t544 28.565
R1082 VDD.n842 VDD.t528 28.565
R1083 VDD.n902 VDD.t44 28.565
R1084 VDD.n902 VDD.t942 28.565
R1085 VDD.n896 VDD.t624 28.565
R1086 VDD.n896 VDD.t940 28.565
R1087 VDD.n890 VDD.t677 28.565
R1088 VDD.n890 VDD.t636 28.565
R1089 VDD.n884 VDD.t965 28.565
R1090 VDD.n884 VDD.t571 28.565
R1091 VDD.n878 VDD.t811 28.565
R1092 VDD.n878 VDD.t215 28.565
R1093 VDD.n872 VDD.t1118 28.565
R1094 VDD.n872 VDD.t1116 28.565
R1095 VDD.n866 VDD.t1144 28.565
R1096 VDD.n866 VDD.t151 28.565
R1097 VDD.n860 VDD.t288 28.565
R1098 VDD.n860 VDD.t388 28.565
R1099 VDD.n492 VDD.t443 28.565
R1100 VDD.n492 VDD.t445 28.565
R1101 VDD.n483 VDD.t777 28.565
R1102 VDD.n483 VDD.t230 28.565
R1103 VDD.n486 VDD.t1082 28.565
R1104 VDD.n472 VDD.t704 28.565
R1105 VDD.n472 VDD.t706 28.565
R1106 VDD.n463 VDD.t1042 28.565
R1107 VDD.n463 VDD.t996 28.565
R1108 VDD.n466 VDD.t1059 28.565
R1109 VDD.n412 VDD.t218 28.565
R1110 VDD.n412 VDD.t805 28.565
R1111 VDD.n403 VDD.t787 28.565
R1112 VDD.n403 VDD.t660 28.565
R1113 VDD.n406 VDD.t1104 28.565
R1114 VDD.n392 VDD.t207 28.565
R1115 VDD.n392 VDD.t1129 28.565
R1116 VDD.n383 VDD.t1078 28.565
R1117 VDD.n383 VDD.t976 28.565
R1118 VDD.n386 VDD.t1106 28.565
R1119 VDD.n353 VDD.t759 28.565
R1120 VDD.n353 VDD.t978 28.565
R1121 VDD.n344 VDD.t885 28.565
R1122 VDD.n344 VDD.t785 28.565
R1123 VDD.n347 VDD.t1086 28.565
R1124 VDD.n372 VDD.t673 28.565
R1125 VDD.n372 VDD.t675 28.565
R1126 VDD.n363 VDD.t1108 28.565
R1127 VDD.n363 VDD.t789 28.565
R1128 VDD.n366 VDD.t65 28.565
R1129 VDD.n432 VDD.t1269 28.565
R1130 VDD.n432 VDD.t1112 28.565
R1131 VDD.n423 VDD.t1061 28.565
R1132 VDD.n423 VDD.t1242 28.565
R1133 VDD.n426 VDD.t781 28.565
R1134 VDD.n452 VDD.t520 28.565
R1135 VDD.n452 VDD.t495 28.565
R1136 VDD.n443 VDD.t228 28.565
R1137 VDD.n443 VDD.t1240 28.565
R1138 VDD.n446 VDD.t1259 28.565
R1139 VDD.n651 VDD.t126 28.565
R1140 VDD.n651 VDD.t124 28.565
R1141 VDD.n642 VDD.t1160 28.565
R1142 VDD.n642 VDD.t333 28.565
R1143 VDD.n645 VDD.t1233 28.565
R1144 VDD.n631 VDD.t412 28.565
R1145 VDD.n631 VDD.t410 28.565
R1146 VDD.n622 VDD.t344 28.565
R1147 VDD.n622 VDD.t406 28.565
R1148 VDD.n625 VDD.t3 28.565
R1149 VDD.n571 VDD.t1142 28.565
R1150 VDD.n571 VDD.t1140 28.565
R1151 VDD.n562 VDD.t1210 28.565
R1152 VDD.n562 VDD.t297 28.565
R1153 VDD.n565 VDD.t238 28.565
R1154 VDD.n551 VDD.t1177 28.565
R1155 VDD.n551 VDD.t1238 28.565
R1156 VDD.n542 VDD.t80 28.565
R1157 VDD.n542 VDD.t348 28.565
R1158 VDD.n545 VDD.t162 28.565
R1159 VDD.n512 VDD.t1224 28.565
R1160 VDD.n512 VDD.t1222 28.565
R1161 VDD.n503 VDD.t236 28.565
R1162 VDD.n503 VDD.t1208 28.565
R1163 VDD.n506 VDD.t33 28.565
R1164 VDD.n531 VDD.t831 28.565
R1165 VDD.n531 VDD.t835 28.565
R1166 VDD.n522 VDD.t1235 28.565
R1167 VDD.n522 VDD.t470 28.565
R1168 VDD.n525 VDD.t664 28.565
R1169 VDD.n591 VDD.t168 28.565
R1170 VDD.n591 VDD.t166 28.565
R1171 VDD.n582 VDD.t350 28.565
R1172 VDD.n582 VDD.t15 28.565
R1173 VDD.n585 VDD.t82 28.565
R1174 VDD.n611 VDD.t248 28.565
R1175 VDD.n611 VDD.t246 28.565
R1176 VDD.n602 VDD.t428 28.565
R1177 VDD.n602 VDD.t88 28.565
R1178 VDD.n605 VDD.t708 28.565
R1179 VDD.n8 VDD.t820 28.565
R1180 VDD.n8 VDD.t822 28.565
R1181 VDD.n22 VDD.t1152 28.565
R1182 VDD.n22 VDD.t1154 28.565
R1183 VDD.n34 VDD.t1250 28.565
R1184 VDD.n34 VDD.t583 28.565
R1185 VDD.n49 VDD.t871 28.565
R1186 VDD.n49 VDD.t873 28.565
R1187 VDD.n77 VDD.t614 28.565
R1188 VDD.n77 VDD.t974 28.565
R1189 VDD.n91 VDD.t115 28.565
R1190 VDD.n91 VDD.t90 28.565
R1191 VDD.n63 VDD.t1028 28.565
R1192 VDD.n63 VDD.t1024 28.565
R1193 VDD.n109 VDD.t989 28.565
R1194 VDD.n109 VDD.t1002 28.565
R1195 VDD.n172 VDD.t258 23.317
R1196 VDD.n164 VDD.t148 23.317
R1197 VDD.n140 VDD.t879 23.317
R1198 VDD.n132 VDD.t319 23.317
R1199 VDD.n116 VDD.t254 23.317
R1200 VDD.n124 VDD.t643 23.317
R1201 VDD.n148 VDD.t478 23.317
R1202 VDD.n156 VDD.t1171 23.317
R1203 VDD.n701 VDD.t1013 20.998
R1204 VDD.n801 VDD.t933 20.998
R1205 VDD.n676 VDD.t212 20.998
R1206 VDD.n726 VDD.t1230 20.998
R1207 VDD.n751 VDD.t378 20.998
R1208 VDD.n776 VDD.t572 20.998
R1209 VDD.n826 VDD.t261 20.998
R1210 VDD.n851 VDD.t256 20.998
R1211 VDD.n172 VDD.t26 20.183
R1212 VDD.n164 VDD.t559 20.183
R1213 VDD.n140 VDD.t174 20.183
R1214 VDD.n132 VDD.t1095 20.183
R1215 VDD.n116 VDD.t533 20.183
R1216 VDD.n124 VDD.t1182 20.183
R1217 VDD.n148 VDD.t597 20.183
R1218 VDD.n156 VDD.t270 20.183
R1219 VDD.n322 VDD.t916 17.506
R1220 VDD.n302 VDD.t10 17.506
R1221 VDD.n242 VDD.t471 17.506
R1222 VDD.n222 VDD.t436 17.506
R1223 VDD.n183 VDD.t421 17.506
R1224 VDD.n202 VDD.t53 17.506
R1225 VDD.n262 VDD.t440 17.506
R1226 VDD.n282 VDD.t918 17.506
R1227 VDD.n481 VDD.t657 17.506
R1228 VDD.n461 VDD.t231 17.506
R1229 VDD.n401 VDD.t1262 17.506
R1230 VDD.n381 VDD.t1037 17.506
R1231 VDD.n342 VDD.t687 17.506
R1232 VDD.n361 VDD.t947 17.506
R1233 VDD.n421 VDD.t1039 17.506
R1234 VDD.n441 VDD.t1101 17.506
R1235 VDD.n640 VDD.t334 17.506
R1236 VDD.n620 VDD.t93 17.506
R1237 VDD.n560 VDD.t423 17.506
R1238 VDD.n540 VDD.t339 17.506
R1239 VDD.n501 VDD.t1011 17.506
R1240 VDD.n520 VDD.t36 17.506
R1241 VDD.n580 VDD.t353 17.506
R1242 VDD.n600 VDD.t6 17.506
R1243 VDD.n684 VDD.t140 14.284
R1244 VDD.n691 VDD.t1244 14.284
R1245 VDD.n784 VDD.t640 14.284
R1246 VDD.n791 VDD.t1094 14.284
R1247 VDD.n659 VDD.t608 14.284
R1248 VDD.n666 VDD.t1098 14.284
R1249 VDD.n709 VDD.t1181 14.284
R1250 VDD.n716 VDD.t277 14.284
R1251 VDD.n734 VDD.t312 14.284
R1252 VDD.n741 VDD.t923 14.284
R1253 VDD.n759 VDD.t967 14.284
R1254 VDD.n766 VDD.t180 14.284
R1255 VDD.n809 VDD.t620 14.284
R1256 VDD.n816 VDD.t867 14.284
R1257 VDD.n834 VDD.t1019 14.284
R1258 VDD.n841 VDD.t546 14.284
R1259 VDD.n10 VDD.t824 14.284
R1260 VDD.n24 VDD.t1114 14.284
R1261 VDD.n36 VDD.t925 14.284
R1262 VDD.n51 VDD.t592 14.284
R1263 VDD.n79 VDD.t865 14.284
R1264 VDD.n93 VDD.t548 14.284
R1265 VDD.n65 VDD.t773 14.284
R1266 VDD.n111 VDD.t187 14.284
R1267 VDD.n332 VDD.t56 14.283
R1268 VDD.n312 VDD.t9 14.283
R1269 VDD.n252 VDD.t244 14.283
R1270 VDD.n232 VDD.t58 14.283
R1271 VDD.n193 VDD.t466 14.283
R1272 VDD.n212 VDD.t92 14.283
R1273 VDD.n272 VDD.t19 14.283
R1274 VDD.n292 VDD.t74 14.283
R1275 VDD.n491 VDD.t950 14.283
R1276 VDD.n471 VDD.t690 14.283
R1277 VDD.n411 VDD.t1080 14.283
R1278 VDD.n391 VDD.t952 14.283
R1279 VDD.n352 VDD.t998 14.283
R1280 VDD.n371 VDD.t954 14.283
R1281 VDD.n431 VDD.t783 14.283
R1282 VDD.n451 VDD.t63 14.283
R1283 VDD.n650 VDD.t432 14.283
R1284 VDD.n630 VDD.t434 14.283
R1285 VDD.n570 VDD.t913 14.283
R1286 VDD.n550 VDD.t418 14.283
R1287 VDD.n511 VDD.t1008 14.283
R1288 VDD.n530 VDD.t915 14.283
R1289 VDD.n590 VDD.t1136 14.283
R1290 VDD.n610 VDD.t13 14.283
R1291 VDD.n328 VDD.t765 14.283
R1292 VDD.n308 VDD.t1134 14.283
R1293 VDD.n248 VDD.t877 14.283
R1294 VDD.n228 VDD.t1110 14.283
R1295 VDD.n189 VDD.t155 14.283
R1296 VDD.n208 VDD.t841 14.283
R1297 VDD.n268 VDD.t586 14.283
R1298 VDD.n288 VDD.t1074 14.283
R1299 VDD.n487 VDD.t193 14.283
R1300 VDD.n467 VDD.t1218 14.283
R1301 VDD.n407 VDD.t226 14.283
R1302 VDD.n387 VDD.t562 14.283
R1303 VDD.n348 VDD.t890 14.283
R1304 VDD.n367 VDD.t753 14.283
R1305 VDD.n427 VDD.t733 14.283
R1306 VDD.n447 VDD.t414 14.283
R1307 VDD.n646 VDD.t284 14.283
R1308 VDD.n626 VDD.t108 14.283
R1309 VDD.n566 VDD.t71 14.283
R1310 VDD.n546 VDD.t1046 14.283
R1311 VDD.n507 VDD.t1033 14.283
R1312 VDD.n526 VDD.t1165 14.283
R1313 VDD.n586 VDD.t741 14.283
R1314 VDD.n606 VDD.t1199 14.283
R1315 VDD.n331 VDD.t302 14.282
R1316 VDD.n331 VDD.t917 14.282
R1317 VDD.n326 VDD.t767 14.282
R1318 VDD.n326 VDD.t763 14.282
R1319 VDD.n311 VDD.t35 14.282
R1320 VDD.n311 VDD.t11 14.282
R1321 VDD.n306 VDD.t698 14.282
R1322 VDD.n306 VDD.t1054 14.282
R1323 VDD.n251 VDD.t234 14.282
R1324 VDD.n251 VDD.t472 14.282
R1325 VDD.n246 VDD.t524 14.282
R1326 VDD.n246 VDD.t875 14.282
R1327 VDD.n231 VDD.t337 14.282
R1328 VDD.n231 VDD.t437 14.282
R1329 VDD.n226 VDD.t452 14.282
R1330 VDD.n226 VDD.t459 14.282
R1331 VDD.n192 VDD.t439 14.282
R1332 VDD.n192 VDD.t422 14.282
R1333 VDD.n187 VDD.t67 14.282
R1334 VDD.n187 VDD.t984 14.282
R1335 VDD.n211 VDD.t476 14.282
R1336 VDD.n211 VDD.t54 14.282
R1337 VDD.n206 VDD.t23 14.282
R1338 VDD.n206 VDD.t25 14.282
R1339 VDD.n271 VDD.t1150 14.282
R1340 VDD.n271 VDD.t441 14.282
R1341 VDD.n266 VDD.t502 14.282
R1342 VDD.n266 VDD.t504 14.282
R1343 VDD.n291 VDD.t342 14.282
R1344 VDD.n291 VDD.t919 14.282
R1345 VDD.n286 VDD.t1076 14.282
R1346 VDD.n286 VDD.t1072 14.282
R1347 VDD.n683 VDD.t1014 14.282
R1348 VDD.n683 VDD.t612 14.282
R1349 VDD.n690 VDD.t552 14.282
R1350 VDD.n690 VDD.t195 14.282
R1351 VDD.n783 VDD.t934 14.282
R1352 VDD.n783 VDD.t323 14.282
R1353 VDD.n790 VDD.t328 14.282
R1354 VDD.n790 VDD.t1197 14.282
R1355 VDD.n658 VDD.t213 14.282
R1356 VDD.n658 VDD.t211 14.282
R1357 VDD.n665 VDD.t147 14.282
R1358 VDD.n665 VDD.t143 14.282
R1359 VDD.n708 VDD.t1231 14.282
R1360 VDD.n708 VDD.t1229 14.282
R1361 VDD.n715 VDD.t275 14.282
R1362 VDD.n715 VDD.t273 14.282
R1363 VDD.n733 VDD.t379 14.282
R1364 VDD.n733 VDD.t809 14.282
R1365 VDD.n740 VDD.t602 14.282
R1366 VDD.n740 VDD.t518 14.282
R1367 VDD.n758 VDD.t573 14.282
R1368 VDD.n758 VDD.t569 14.282
R1369 VDD.n765 VDD.t178 14.282
R1370 VDD.n765 VDD.t596 14.282
R1371 VDD.n808 VDD.t262 14.282
R1372 VDD.n808 VDD.t626 14.282
R1373 VDD.n815 VDD.t1131 14.282
R1374 VDD.n815 VDD.t104 14.282
R1375 VDD.n833 VDD.t257 14.282
R1376 VDD.n833 VDD.t1022 14.282
R1377 VDD.n840 VDD.t526 14.282
R1378 VDD.n840 VDD.t536 14.282
R1379 VDD.n490 VDD.t1100 14.282
R1380 VDD.n490 VDD.t658 14.282
R1381 VDD.n485 VDD.t769 14.282
R1382 VDD.n485 VDD.t191 14.282
R1383 VDD.n470 VDD.t779 14.282
R1384 VDD.n470 VDD.t232 14.282
R1385 VDD.n465 VDD.t1220 14.282
R1386 VDD.n465 VDD.t1216 14.282
R1387 VDD.n410 VDD.t775 14.282
R1388 VDD.n410 VDD.t1263 14.282
R1389 VDD.n405 VDD.t462 14.282
R1390 VDD.n405 VDD.t224 14.282
R1391 VDD.n390 VDD.t1000 14.282
R1392 VDD.n390 VDD.t1038 14.282
R1393 VDD.n385 VDD.t564 14.282
R1394 VDD.n385 VDD.t182 14.282
R1395 VDD.n351 VDD.t1265 14.282
R1396 VDD.n351 VDD.t688 14.282
R1397 VDD.n346 VDD.t102 14.282
R1398 VDD.n346 VDD.t826 14.282
R1399 VDD.n370 VDD.t1261 14.282
R1400 VDD.n370 VDD.t948 14.282
R1401 VDD.n365 VDD.t755 14.282
R1402 VDD.n365 VDD.t1124 14.282
R1403 VDD.n430 VDD.t1084 14.282
R1404 VDD.n430 VDD.t1040 14.282
R1405 VDD.n425 VDD.t735 14.282
R1406 VDD.n425 VDD.t737 14.282
R1407 VDD.n450 VDD.t692 14.282
R1408 VDD.n450 VDD.t1102 14.282
R1409 VDD.n445 VDD.t416 14.282
R1410 VDD.n445 VDD.t1044 14.282
R1411 VDD.n649 VDD.t468 14.282
R1412 VDD.n649 VDD.t335 14.282
R1413 VDD.n644 VDD.t111 14.282
R1414 VDD.n644 VDD.t286 14.282
R1415 VDD.n629 VDD.t352 14.282
R1416 VDD.n629 VDD.t94 14.282
R1417 VDD.n624 VDD.t1017 14.282
R1418 VDD.n624 VDD.t656 14.282
R1419 VDD.n569 VDD.t39 14.282
R1420 VDD.n569 VDD.t424 14.282
R1421 VDD.n564 VDD.t60 14.282
R1422 VDD.n564 VDD.t29 14.282
R1423 VDD.n549 VDD.t76 14.282
R1424 VDD.n549 VDD.t340 14.282
R1425 VDD.n544 VDD.t401 14.282
R1426 VDD.n544 VDD.t1214 14.282
R1427 VDD.n510 VDD.t299 14.282
R1428 VDD.n510 VDD.t1012 14.282
R1429 VDD.n505 VDD.t1031 14.282
R1430 VDD.n505 VDD.t42 14.282
R1431 VDD.n529 VDD.t295 14.282
R1432 VDD.n529 VDD.t37 14.282
R1433 VDD.n524 VDD.t486 14.282
R1434 VDD.n524 VDD.t484 14.282
R1435 VDD.n589 VDD.t408 14.282
R1436 VDD.n589 VDD.t354 14.282
R1437 VDD.n584 VDD.t883 14.282
R1438 VDD.n584 VDD.t1121 14.282
R1439 VDD.n609 VDD.t426 14.282
R1440 VDD.n609 VDD.t7 14.282
R1441 VDD.n604 VDD.t828 14.282
R1442 VDD.n604 VDD.t1201 14.282
R1443 VDD.n11 VDD.t554 14.282
R1444 VDD.n11 VDD.t1246 14.282
R1445 VDD.n25 VDD.t360 14.282
R1446 VDD.n25 VDD.t269 14.282
R1447 VDD.n37 VDD.t128 14.282
R1448 VDD.n37 VDD.t600 14.282
R1449 VDD.n52 VDD.t493 14.282
R1450 VDD.n52 VDD.t670 14.282
R1451 VDD.n80 VDD.t843 14.282
R1452 VDD.n80 VDD.t384 14.282
R1453 VDD.n94 VDD.t542 14.282
R1454 VDD.n94 VDD.t538 14.282
R1455 VDD.n66 VDD.t662 14.282
R1456 VDD.n66 VDD.t652 14.282
R1457 VDD.n112 VDD.t1203 14.282
R1458 VDD.n112 VDD.t887 14.282
R1459 VDD.n6 VDD.t823 13.431
R1460 VDD.n32 VDD.t924 13.431
R1461 VDD.n47 VDD.t591 13.431
R1462 VDD.n75 VDD.t864 13.431
R1463 VDD.n104 VDD.t186 13.431
R1464 VDD.n20 VDD.t1113 13.397
R1465 VDD.n89 VDD.t547 13.397
R1466 VDD.n61 VDD.t772 13.397
R1467 VDD.n706 VDD.n688 9.03
R1468 VDD.n806 VDD.n788 9.03
R1469 VDD.n681 VDD.n663 9.03
R1470 VDD.n731 VDD.n713 9.03
R1471 VDD.n756 VDD.n738 9.03
R1472 VDD.n781 VDD.n763 9.03
R1473 VDD.n831 VDD.n813 9.03
R1474 VDD.n856 VDD.n838 9.03
R1475 VDD.n695 VDD.n682 9
R1476 VDD.n795 VDD.n782 9
R1477 VDD.n670 VDD.n657 9
R1478 VDD.n720 VDD.n707 9
R1479 VDD.n745 VDD.n732 9
R1480 VDD.n770 VDD.n757 9
R1481 VDD.n820 VDD.n807 9
R1482 VDD.n845 VDD.n832 9
R1483 VDD.n323 VDD.n322 6.626
R1484 VDD.n303 VDD.n302 6.626
R1485 VDD.n243 VDD.n242 6.626
R1486 VDD.n223 VDD.n222 6.626
R1487 VDD.n184 VDD.n183 6.626
R1488 VDD.n203 VDD.n202 6.626
R1489 VDD.n263 VDD.n262 6.626
R1490 VDD.n283 VDD.n282 6.626
R1491 VDD.n482 VDD.n481 6.626
R1492 VDD.n462 VDD.n461 6.626
R1493 VDD.n402 VDD.n401 6.626
R1494 VDD.n382 VDD.n381 6.626
R1495 VDD.n343 VDD.n342 6.626
R1496 VDD.n362 VDD.n361 6.626
R1497 VDD.n422 VDD.n421 6.626
R1498 VDD.n442 VDD.n441 6.626
R1499 VDD.n641 VDD.n640 6.626
R1500 VDD.n621 VDD.n620 6.626
R1501 VDD.n561 VDD.n560 6.626
R1502 VDD.n541 VDD.n540 6.626
R1503 VDD.n502 VDD.n501 6.626
R1504 VDD.n521 VDD.n520 6.626
R1505 VDD.n581 VDD.n580 6.626
R1506 VDD.n601 VDD.n600 6.626
R1507 VDD.n697 VDD.t1132 6.189
R1508 VDD.n698 VDD.t201 6.189
R1509 VDD.n700 VDD.t1068 6.189
R1510 VDD.n699 VDD.t1070 6.189
R1511 VDD.n797 VDD.t456 6.189
R1512 VDD.n798 VDD.t455 6.189
R1513 VDD.n800 VDD.t1127 6.189
R1514 VDD.n799 VDD.t1125 6.189
R1515 VDD.n672 VDD.t1175 6.189
R1516 VDD.n673 VDD.t813 6.189
R1517 VDD.n675 VDD.t671 6.189
R1518 VDD.n674 VDD.t1211 6.189
R1519 VDD.n722 VDD.t293 6.189
R1520 VDD.n723 VDD.t292 6.189
R1521 VDD.n725 VDD.t878 6.189
R1522 VDD.n724 VDD.t249 6.189
R1523 VDD.n747 VDD.t30 6.189
R1524 VDD.n748 VDD.t61 6.189
R1525 VDD.n750 VDD.t905 6.189
R1526 VDD.n749 VDD.t117 6.189
R1527 VDD.n772 VDD.t1035 6.189
R1528 VDD.n773 VDD.t1212 6.189
R1529 VDD.n775 VDD.t1251 6.189
R1530 VDD.n774 VDD.t1187 6.189
R1531 VDD.n822 VDD.t454 6.189
R1532 VDD.n823 VDD.t453 6.189
R1533 VDD.n825 VDD.t279 6.189
R1534 VDD.n824 VDD.t278 6.189
R1535 VDD.n847 VDD.t282 6.189
R1536 VDD.n848 VDD.t892 6.189
R1537 VDD.n850 VDD.t220 6.189
R1538 VDD.n849 VDD.t156 6.189
R1539 VDD.t553 VDD.n1 6.105
R1540 VDD.t127 VDD.n29 6.105
R1541 VDD.t492 VDD.n41 6.105
R1542 VDD.t842 VDD.n70 6.105
R1543 VDD.n107 VDD.t1202 6.105
R1544 VDD.t359 VDD.n15 6.089
R1545 VDD.t541 VDD.n84 6.089
R1546 VDD.t661 VDD.n56 6.089
R1547 VDD.n320 VDD.n319 6
R1548 VDD.n300 VDD.n299 6
R1549 VDD.n240 VDD.n239 6
R1550 VDD.n220 VDD.n219 6
R1551 VDD.n181 VDD.n180 6
R1552 VDD.n200 VDD.n199 6
R1553 VDD.n260 VDD.n259 6
R1554 VDD.n280 VDD.n279 6
R1555 VDD.n479 VDD.n478 6
R1556 VDD.n459 VDD.n458 6
R1557 VDD.n399 VDD.n398 6
R1558 VDD.n379 VDD.n378 6
R1559 VDD.n340 VDD.n339 6
R1560 VDD.n359 VDD.n358 6
R1561 VDD.n419 VDD.n418 6
R1562 VDD.n439 VDD.n438 6
R1563 VDD.n638 VDD.n637 6
R1564 VDD.n618 VDD.n617 6
R1565 VDD.n558 VDD.n557 6
R1566 VDD.n538 VDD.n537 6
R1567 VDD.n499 VDD.n498 6
R1568 VDD.n518 VDD.n517 6
R1569 VDD.n578 VDD.n577 6
R1570 VDD.n598 VDD.n597 6
R1571 VDD.n7 VDD.n6 5.506
R1572 VDD.n21 VDD.n20 5.506
R1573 VDD.n33 VDD.n32 5.506
R1574 VDD.n48 VDD.n47 5.506
R1575 VDD.n76 VDD.n75 5.506
R1576 VDD.n90 VDD.n89 5.506
R1577 VDD.n62 VDD.n61 5.506
R1578 VDD.n104 VDD.n103 5.506
R1579 VDD.n44 VDD.t870 3.368
R1580 VDD.n336 VDD.n330 2.572
R1581 VDD.n316 VDD.n310 2.572
R1582 VDD.n256 VDD.n250 2.572
R1583 VDD.n236 VDD.n230 2.572
R1584 VDD.n197 VDD.n191 2.572
R1585 VDD.n216 VDD.n210 2.572
R1586 VDD.n276 VDD.n270 2.572
R1587 VDD.n296 VDD.n290 2.572
R1588 VDD.n495 VDD.n489 2.572
R1589 VDD.n475 VDD.n469 2.572
R1590 VDD.n415 VDD.n409 2.572
R1591 VDD.n395 VDD.n389 2.572
R1592 VDD.n356 VDD.n350 2.572
R1593 VDD.n375 VDD.n369 2.572
R1594 VDD.n435 VDD.n429 2.572
R1595 VDD.n455 VDD.n449 2.572
R1596 VDD.n654 VDD.n648 2.572
R1597 VDD.n634 VDD.n628 2.572
R1598 VDD.n574 VDD.n568 2.572
R1599 VDD.n554 VDD.n548 2.572
R1600 VDD.n515 VDD.n509 2.572
R1601 VDD.n534 VDD.n528 2.572
R1602 VDD.n594 VDD.n588 2.572
R1603 VDD.n614 VDD.n608 2.572
R1604 VDD.n335 VDD.n334 2.54
R1605 VDD.n315 VDD.n314 2.54
R1606 VDD.n255 VDD.n254 2.54
R1607 VDD.n235 VDD.n234 2.54
R1608 VDD.n196 VDD.n195 2.54
R1609 VDD.n215 VDD.n214 2.54
R1610 VDD.n275 VDD.n274 2.54
R1611 VDD.n295 VDD.n294 2.54
R1612 VDD.n494 VDD.n493 2.54
R1613 VDD.n474 VDD.n473 2.54
R1614 VDD.n414 VDD.n413 2.54
R1615 VDD.n394 VDD.n393 2.54
R1616 VDD.n355 VDD.n354 2.54
R1617 VDD.n374 VDD.n373 2.54
R1618 VDD.n434 VDD.n433 2.54
R1619 VDD.n454 VDD.n453 2.54
R1620 VDD.n653 VDD.n652 2.54
R1621 VDD.n633 VDD.n632 2.54
R1622 VDD.n573 VDD.n572 2.54
R1623 VDD.n553 VDD.n552 2.54
R1624 VDD.n514 VDD.n513 2.54
R1625 VDD.n533 VDD.n532 2.54
R1626 VDD.n593 VDD.n592 2.54
R1627 VDD.n613 VDD.n612 2.54
R1628 VDD.n93 VDD.n92 2.521
R1629 VDD.n686 VDD.n685 2.451
R1630 VDD.n786 VDD.n785 2.451
R1631 VDD.n661 VDD.n660 2.451
R1632 VDD.n711 VDD.n710 2.451
R1633 VDD.n736 VDD.n735 2.451
R1634 VDD.n761 VDD.n760 2.451
R1635 VDD.n811 VDD.n810 2.451
R1636 VDD.n836 VDD.n835 2.451
R1637 VDD.n693 VDD.n692 2.449
R1638 VDD.n793 VDD.n792 2.449
R1639 VDD.n668 VDD.n667 2.449
R1640 VDD.n718 VDD.n717 2.449
R1641 VDD.n743 VDD.n742 2.449
R1642 VDD.n768 VDD.n767 2.449
R1643 VDD.n818 VDD.n817 2.449
R1644 VDD.n843 VDD.n842 2.449
R1645 VDD.n79 VDD.n78 2.225
R1646 VDD.n51 VDD.n50 2.221
R1647 VDD.n111 VDD.n110 2.221
R1648 VDD.n65 VDD.n64 2.218
R1649 VDD.n10 VDD.n9 2.199
R1650 VDD.n36 VDD.n35 2.199
R1651 VDD.n24 VDD.n23 2.192
R1652 VDD.n321 VDD.n320 1.929
R1653 VDD.n301 VDD.n300 1.929
R1654 VDD.n241 VDD.n240 1.929
R1655 VDD.n221 VDD.n220 1.929
R1656 VDD.n182 VDD.n181 1.929
R1657 VDD.n201 VDD.n200 1.929
R1658 VDD.n261 VDD.n260 1.929
R1659 VDD.n281 VDD.n280 1.929
R1660 VDD.n480 VDD.n479 1.929
R1661 VDD.n460 VDD.n459 1.929
R1662 VDD.n400 VDD.n399 1.929
R1663 VDD.n380 VDD.n379 1.929
R1664 VDD.n341 VDD.n340 1.929
R1665 VDD.n360 VDD.n359 1.929
R1666 VDD.n420 VDD.n419 1.929
R1667 VDD.n440 VDD.n439 1.929
R1668 VDD.n639 VDD.n638 1.929
R1669 VDD.n619 VDD.n618 1.929
R1670 VDD.n559 VDD.n558 1.929
R1671 VDD.n539 VDD.n538 1.929
R1672 VDD.n500 VDD.n499 1.929
R1673 VDD.n519 VDD.n518 1.929
R1674 VDD.n579 VDD.n578 1.929
R1675 VDD.n599 VDD.n598 1.929
R1676 VDD.n918 VDD.n682 1.738
R1677 VDD.n914 VDD.n782 1.738
R1678 VDD.n919 VDD.n657 1.738
R1679 VDD.n917 VDD.n707 1.738
R1680 VDD.n916 VDD.n732 1.738
R1681 VDD.n915 VDD.n757 1.738
R1682 VDD.n913 VDD.n807 1.738
R1683 VDD.n912 VDD.n832 1.738
R1684 VDD.n9 VDD.n8 1.651
R1685 VDD.n23 VDD.n22 1.651
R1686 VDD.n35 VDD.n34 1.651
R1687 VDD.n50 VDD.n49 1.607
R1688 VDD.n92 VDD.n91 1.607
R1689 VDD.n110 VDD.n109 1.607
R1690 VDD.n78 VDD.n77 1.599
R1691 VDD.n64 VDD.n63 1.599
R1692 VDD.n175 VDD.n173 1.564
R1693 VDD.n167 VDD.n165 1.564
R1694 VDD.n143 VDD.n141 1.564
R1695 VDD.n135 VDD.n133 1.564
R1696 VDD.n119 VDD.n117 1.564
R1697 VDD.n127 VDD.n125 1.564
R1698 VDD.n151 VDD.n149 1.564
R1699 VDD.n159 VDD.n157 1.564
R1700 VDD.n26 VDD.n24 1.161
R1701 VDD.n95 VDD.n93 1.161
R1702 VDD.n67 VDD.n65 1.161
R1703 VDD.n12 VDD.n10 1.154
R1704 VDD.n38 VDD.n36 1.154
R1705 VDD.n53 VDD.n51 1.154
R1706 VDD.n81 VDD.n79 1.154
R1707 VDD.n113 VDD.n111 1.154
R1708 VDD.n26 VDD.n25 1.107
R1709 VDD.n95 VDD.n94 1.107
R1710 VDD.n67 VDD.n66 1.107
R1711 VDD.n12 VDD.n11 1.1
R1712 VDD.n38 VDD.n37 1.1
R1713 VDD.n53 VDD.n52 1.1
R1714 VDD.n81 VDD.n80 1.1
R1715 VDD.n113 VDD.n112 1.1
R1716 VDD.n319 VDD.t937 1.057
R1717 VDD.n299 VDD.t910 1.057
R1718 VDD.n239 VDD.t987 1.057
R1719 VDD.n219 VDD.t894 1.057
R1720 VDD.n180 VDD.t898 1.057
R1721 VDD.n199 VDD.t888 1.057
R1722 VDD.n259 VDD.t694 1.057
R1723 VDD.n279 VDD.t315 1.057
R1724 VDD.n478 VDD.t313 1.057
R1725 VDD.n458 VDD.t183 1.057
R1726 VDD.n398 VDD.t260 1.057
R1727 VDD.n378 VDD.t317 1.057
R1728 VDD.n339 VDD.t747 1.057
R1729 VDD.n358 VDD.t818 1.057
R1730 VDD.n418 VDD.t955 1.057
R1731 VDD.n438 VDD.t699 1.057
R1732 VDD.n637 VDD.t199 1.057
R1733 VDD.n617 VDD.t430 1.057
R1734 VDD.n557 VDD.t1015 1.057
R1735 VDD.n537 VDD.t252 1.057
R1736 VDD.n498 VDD.t72 1.057
R1737 VDD.n517 VDD.t200 1.057
R1738 VDD.n577 VDD.t171 1.057
R1739 VDD.n597 VDD.t1119 1.057
R1740 VDD.n3 VDD.n2 1.008
R1741 VDD.n31 VDD.n30 1.008
R1742 VDD.n43 VDD.n42 1.008
R1743 VDD.n72 VDD.n71 1.008
R1744 VDD.n106 VDD.n105 1.008
R1745 VDD.n17 VDD.n16 1.006
R1746 VDD.n86 VDD.n85 1.006
R1747 VDD.n58 VDD.n57 1.006
R1748 VDD.n687 VDD.n683 0.922
R1749 VDD.n694 VDD.n690 0.922
R1750 VDD.n787 VDD.n783 0.922
R1751 VDD.n794 VDD.n790 0.922
R1752 VDD.n662 VDD.n658 0.922
R1753 VDD.n669 VDD.n665 0.922
R1754 VDD.n712 VDD.n708 0.922
R1755 VDD.n719 VDD.n715 0.922
R1756 VDD.n737 VDD.n733 0.922
R1757 VDD.n744 VDD.n740 0.922
R1758 VDD.n762 VDD.n758 0.922
R1759 VDD.n769 VDD.n765 0.922
R1760 VDD.n812 VDD.n808 0.922
R1761 VDD.n819 VDD.n815 0.922
R1762 VDD.n837 VDD.n833 0.922
R1763 VDD.n844 VDD.n840 0.922
R1764 VDD.n686 VDD.n684 0.921
R1765 VDD.n693 VDD.n691 0.921
R1766 VDD.n786 VDD.n784 0.921
R1767 VDD.n793 VDD.n791 0.921
R1768 VDD.n661 VDD.n659 0.921
R1769 VDD.n668 VDD.n666 0.921
R1770 VDD.n711 VDD.n709 0.921
R1771 VDD.n718 VDD.n716 0.921
R1772 VDD.n736 VDD.n734 0.921
R1773 VDD.n743 VDD.n741 0.921
R1774 VDD.n761 VDD.n759 0.921
R1775 VDD.n768 VDD.n766 0.921
R1776 VDD.n811 VDD.n809 0.921
R1777 VDD.n818 VDD.n816 0.921
R1778 VDD.n836 VDD.n834 0.921
R1779 VDD.n843 VDD.n841 0.921
R1780 VDD.n335 VDD.n332 0.863
R1781 VDD.n315 VDD.n312 0.863
R1782 VDD.n255 VDD.n252 0.863
R1783 VDD.n235 VDD.n232 0.863
R1784 VDD.n196 VDD.n193 0.863
R1785 VDD.n215 VDD.n212 0.863
R1786 VDD.n275 VDD.n272 0.863
R1787 VDD.n295 VDD.n292 0.863
R1788 VDD.n494 VDD.n491 0.863
R1789 VDD.n474 VDD.n471 0.863
R1790 VDD.n414 VDD.n411 0.863
R1791 VDD.n394 VDD.n391 0.863
R1792 VDD.n355 VDD.n352 0.863
R1793 VDD.n374 VDD.n371 0.863
R1794 VDD.n434 VDD.n431 0.863
R1795 VDD.n454 VDD.n451 0.863
R1796 VDD.n653 VDD.n650 0.863
R1797 VDD.n633 VDD.n630 0.863
R1798 VDD.n573 VDD.n570 0.863
R1799 VDD.n553 VDD.n550 0.863
R1800 VDD.n514 VDD.n511 0.863
R1801 VDD.n533 VDD.n530 0.863
R1802 VDD.n593 VDD.n590 0.863
R1803 VDD.n613 VDD.n610 0.863
R1804 VDD.n177 VDD.n175 0.85
R1805 VDD.n169 VDD.n167 0.85
R1806 VDD.n145 VDD.n143 0.85
R1807 VDD.n137 VDD.n135 0.85
R1808 VDD.n121 VDD.n119 0.85
R1809 VDD.n129 VDD.n127 0.85
R1810 VDD.n153 VDD.n151 0.85
R1811 VDD.n161 VDD.n159 0.85
R1812 VDD.n179 VDD.n178 0.747
R1813 VDD.n175 VDD.n174 0.747
R1814 VDD.n177 VDD.n176 0.747
R1815 VDD.n171 VDD.n170 0.747
R1816 VDD.n167 VDD.n166 0.747
R1817 VDD.n169 VDD.n168 0.747
R1818 VDD.n147 VDD.n146 0.747
R1819 VDD.n143 VDD.n142 0.747
R1820 VDD.n145 VDD.n144 0.747
R1821 VDD.n139 VDD.n138 0.747
R1822 VDD.n135 VDD.n134 0.747
R1823 VDD.n137 VDD.n136 0.747
R1824 VDD.n123 VDD.n122 0.747
R1825 VDD.n119 VDD.n118 0.747
R1826 VDD.n121 VDD.n120 0.747
R1827 VDD.n131 VDD.n130 0.747
R1828 VDD.n127 VDD.n126 0.747
R1829 VDD.n129 VDD.n128 0.747
R1830 VDD.n155 VDD.n154 0.747
R1831 VDD.n151 VDD.n150 0.747
R1832 VDD.n153 VDD.n152 0.747
R1833 VDD.n163 VDD.n162 0.747
R1834 VDD.n159 VDD.n158 0.747
R1835 VDD.n161 VDD.n160 0.747
R1836 VDD.n687 VDD.n686 0.686
R1837 VDD.n694 VDD.n693 0.686
R1838 VDD.n787 VDD.n786 0.686
R1839 VDD.n794 VDD.n793 0.686
R1840 VDD.n662 VDD.n661 0.686
R1841 VDD.n669 VDD.n668 0.686
R1842 VDD.n712 VDD.n711 0.686
R1843 VDD.n719 VDD.n718 0.686
R1844 VDD.n737 VDD.n736 0.686
R1845 VDD.n744 VDD.n743 0.686
R1846 VDD.n762 VDD.n761 0.686
R1847 VDD.n769 VDD.n768 0.686
R1848 VDD.n812 VDD.n811 0.686
R1849 VDD.n819 VDD.n818 0.686
R1850 VDD.n837 VDD.n836 0.686
R1851 VDD.n844 VDD.n843 0.686
R1852 VDD.n336 VDD.n335 0.646
R1853 VDD.n316 VDD.n315 0.646
R1854 VDD.n256 VDD.n255 0.646
R1855 VDD.n236 VDD.n235 0.646
R1856 VDD.n197 VDD.n196 0.646
R1857 VDD.n216 VDD.n215 0.646
R1858 VDD.n276 VDD.n275 0.646
R1859 VDD.n296 VDD.n295 0.646
R1860 VDD.n495 VDD.n494 0.646
R1861 VDD.n475 VDD.n474 0.646
R1862 VDD.n415 VDD.n414 0.646
R1863 VDD.n395 VDD.n394 0.646
R1864 VDD.n356 VDD.n355 0.646
R1865 VDD.n375 VDD.n374 0.646
R1866 VDD.n435 VDD.n434 0.646
R1867 VDD.n455 VDD.n454 0.646
R1868 VDD.n654 VDD.n653 0.646
R1869 VDD.n634 VDD.n633 0.646
R1870 VDD.n574 VDD.n573 0.646
R1871 VDD.n554 VDD.n553 0.646
R1872 VDD.n515 VDD.n514 0.646
R1873 VDD.n534 VDD.n533 0.646
R1874 VDD.n594 VDD.n593 0.646
R1875 VDD.n614 VDD.n613 0.646
R1876 VDD.n278 VDD.n258 0.643
R1877 VDD.n437 VDD.n417 0.643
R1878 VDD.n596 VDD.n576 0.643
R1879 VDD.n218 VDD.n198 0.638
R1880 VDD.n377 VDD.n357 0.638
R1881 VDD.n536 VDD.n516 0.638
R1882 VDD.n258 VDD.n238 0.631
R1883 VDD.n298 VDD.n278 0.631
R1884 VDD.n338 VDD.n318 0.631
R1885 VDD.n417 VDD.n397 0.631
R1886 VDD.n457 VDD.n437 0.631
R1887 VDD.n497 VDD.n477 0.631
R1888 VDD.n576 VDD.n556 0.631
R1889 VDD.n616 VDD.n596 0.631
R1890 VDD.n656 VDD.n636 0.631
R1891 VDD.n238 VDD.n218 0.629
R1892 VDD.n318 VDD.n298 0.629
R1893 VDD.n397 VDD.n377 0.629
R1894 VDD.n477 VDD.n457 0.629
R1895 VDD.n556 VDD.n536 0.629
R1896 VDD.n636 VDD.n616 0.629
R1897 VDD.n920 VDD.n919 0.573
R1898 VDD.n337 VDD.n320 0.465
R1899 VDD.n317 VDD.n300 0.465
R1900 VDD.n257 VDD.n240 0.465
R1901 VDD.n237 VDD.n220 0.465
R1902 VDD.n198 VDD.n181 0.465
R1903 VDD.n217 VDD.n200 0.465
R1904 VDD.n277 VDD.n260 0.465
R1905 VDD.n297 VDD.n280 0.465
R1906 VDD.n496 VDD.n479 0.465
R1907 VDD.n476 VDD.n459 0.465
R1908 VDD.n416 VDD.n399 0.465
R1909 VDD.n396 VDD.n379 0.465
R1910 VDD.n357 VDD.n340 0.465
R1911 VDD.n376 VDD.n359 0.465
R1912 VDD.n436 VDD.n419 0.465
R1913 VDD.n456 VDD.n439 0.465
R1914 VDD.n655 VDD.n638 0.465
R1915 VDD.n635 VDD.n618 0.465
R1916 VDD.n575 VDD.n558 0.465
R1917 VDD.n555 VDD.n538 0.465
R1918 VDD.n516 VDD.n499 0.465
R1919 VDD.n535 VDD.n518 0.465
R1920 VDD.n595 VDD.n578 0.465
R1921 VDD.n615 VDD.n598 0.465
R1922 VDD.n927 VDD.n926 0.452
R1923 VDD.n925 VDD.n924 0.446
R1924 VDD.n929 VDD.n928 0.446
R1925 VDD.n921 VDD.n920 0.444
R1926 VDD.n922 VDD.n921 0.431
R1927 VDD.n926 VDD.n925 0.431
R1928 VDD.n930 VDD.n929 0.431
R1929 VDD.n928 VDD.n927 0.431
R1930 VDD.n924 VDD.n923 0.431
R1931 VDD.n913 VDD.n912 0.398
R1932 VDD.n914 VDD.n913 0.398
R1933 VDD.n915 VDD.n914 0.398
R1934 VDD.n916 VDD.n915 0.398
R1935 VDD.n917 VDD.n916 0.398
R1936 VDD.n918 VDD.n917 0.398
R1937 VDD.n919 VDD.n918 0.398
R1938 VDD.n903 VDD.n902 0.386
R1939 VDD.n897 VDD.n896 0.386
R1940 VDD.n891 VDD.n890 0.386
R1941 VDD.n885 VDD.n884 0.386
R1942 VDD.n879 VDD.n878 0.386
R1943 VDD.n861 VDD.n860 0.386
R1944 VDD.n873 VDD.n872 0.38
R1945 VDD.n867 VDD.n866 0.369
R1946 VDD.n912 VDD.n911 0.308
R1947 VDD.n923 VDD.n922 0.291
R1948 VDD.n901 VDD.n900 0.285
R1949 VDD.n895 VDD.n894 0.285
R1950 VDD.n889 VDD.n888 0.285
R1951 VDD.n883 VDD.n882 0.285
R1952 VDD.n877 VDD.n876 0.285
R1953 VDD.n859 VDD.n858 0.285
R1954 VDD.n871 VDD.n870 0.285
R1955 VDD.n865 VDD.n864 0.285
R1956 VDD.n97 VDD.n96 0.283
R1957 VDD.n100 VDD.n99 0.281
R1958 VDD.n115 VDD.n102 0.28
R1959 VDD.n98 VDD.n97 0.28
R1960 VDD.n99 VDD.n98 0.28
R1961 VDD.n101 VDD.n100 0.28
R1962 VDD.n102 VDD.n101 0.28
R1963 VDD.n922 VDD.n338 0.262
R1964 VDD.t150 VDD.n863 0.244
R1965 VDD.t1115 VDD.n869 0.243
R1966 VDD.t941 VDD.n899 0.243
R1967 VDD.t939 VDD.n893 0.243
R1968 VDD.t635 VDD.n887 0.243
R1969 VDD.t570 VDD.n881 0.243
R1970 VDD.t214 VDD.n875 0.243
R1971 VDD.t387 VDD.n857 0.243
R1972 VDD.n921 VDD.n497 0.243
R1973 VDD.n13 VDD.n12 0.241
R1974 VDD.n27 VDD.n26 0.241
R1975 VDD.n39 VDD.n38 0.241
R1976 VDD.n54 VDD.n53 0.241
R1977 VDD.n82 VDD.n81 0.241
R1978 VDD.n96 VDD.n95 0.241
R1979 VDD.n68 VDD.n67 0.241
R1980 VDD.n114 VDD.n113 0.241
R1981 VDD.n920 VDD.n656 0.241
R1982 VDD.n923 VDD.n179 0.208
R1983 VDD.n924 VDD.n171 0.208
R1984 VDD.n927 VDD.n147 0.208
R1985 VDD.n928 VDD.n139 0.208
R1986 VDD.n930 VDD.n123 0.208
R1987 VDD.n929 VDD.n131 0.208
R1988 VDD.n926 VDD.n155 0.208
R1989 VDD.n925 VDD.n163 0.208
R1990 VDD.n923 VDD.n177 0.195
R1991 VDD.n924 VDD.n169 0.195
R1992 VDD.n927 VDD.n145 0.195
R1993 VDD.n928 VDD.n137 0.195
R1994 VDD.n930 VDD.n121 0.195
R1995 VDD.n929 VDD.n129 0.195
R1996 VDD.n926 VDD.n153 0.195
R1997 VDD.n925 VDD.n161 0.195
R1998 VDD VDD.n115 0.193
R1999 VDD.n688 VDD.n687 0.193
R2000 VDD.n788 VDD.n787 0.193
R2001 VDD.n663 VDD.n662 0.193
R2002 VDD.n713 VDD.n712 0.193
R2003 VDD.n738 VDD.n737 0.193
R2004 VDD.n763 VDD.n762 0.193
R2005 VDD.n813 VDD.n812 0.193
R2006 VDD.n838 VDD.n837 0.193
R2007 VDD.n695 VDD.n694 0.189
R2008 VDD.n795 VDD.n794 0.189
R2009 VDD.n670 VDD.n669 0.189
R2010 VDD.n720 VDD.n719 0.189
R2011 VDD.n745 VDD.n744 0.189
R2012 VDD.n770 VDD.n769 0.189
R2013 VDD.n820 VDD.n819 0.189
R2014 VDD.n845 VDD.n844 0.189
R2015 VDD.n905 VDD.n904 0.183
R2016 VDD.n909 VDD.n908 0.182
R2017 VDD.n13 VDD.n7 0.182
R2018 VDD.n27 VDD.n21 0.182
R2019 VDD.n39 VDD.n33 0.182
R2020 VDD.n54 VDD.n48 0.182
R2021 VDD.n82 VDD.n76 0.182
R2022 VDD.n96 VDD.n90 0.182
R2023 VDD.n68 VDD.n62 0.182
R2024 VDD.n114 VDD.n103 0.182
R2025 VDD.n906 VDD.n905 0.181
R2026 VDD.n907 VDD.n906 0.181
R2027 VDD.n908 VDD.n907 0.181
R2028 VDD.n910 VDD.n909 0.181
R2029 VDD.n911 VDD.n910 0.181
R2030 VDD.n4 VDD.t819 0.124
R2031 VDD.n18 VDD.t1151 0.124
R2032 VDD.n337 VDD.n336 0.12
R2033 VDD.n317 VDD.n316 0.12
R2034 VDD.n257 VDD.n256 0.12
R2035 VDD.n237 VDD.n236 0.12
R2036 VDD.n198 VDD.n197 0.12
R2037 VDD.n217 VDD.n216 0.12
R2038 VDD.n277 VDD.n276 0.12
R2039 VDD.n297 VDD.n296 0.12
R2040 VDD.n496 VDD.n495 0.12
R2041 VDD.n476 VDD.n475 0.12
R2042 VDD.n416 VDD.n415 0.12
R2043 VDD.n396 VDD.n395 0.12
R2044 VDD.n357 VDD.n356 0.12
R2045 VDD.n376 VDD.n375 0.12
R2046 VDD.n436 VDD.n435 0.12
R2047 VDD.n456 VDD.n455 0.12
R2048 VDD.n655 VDD.n654 0.12
R2049 VDD.n635 VDD.n634 0.12
R2050 VDD.n575 VDD.n574 0.12
R2051 VDD.n555 VDD.n554 0.12
R2052 VDD.n516 VDD.n515 0.12
R2053 VDD.n535 VDD.n534 0.12
R2054 VDD.n595 VDD.n594 0.12
R2055 VDD.n615 VDD.n614 0.12
R2056 VDD.n87 VDD.t114 0.106
R2057 VDD.n73 VDD.t613 0.101
R2058 VDD.n59 VDD.t1027 0.101
R2059 VDD.n330 VDD.n325 0.095
R2060 VDD.n310 VDD.n305 0.095
R2061 VDD.n250 VDD.n245 0.095
R2062 VDD.n230 VDD.n225 0.095
R2063 VDD.n191 VDD.n186 0.095
R2064 VDD.n210 VDD.n205 0.095
R2065 VDD.n270 VDD.n265 0.095
R2066 VDD.n290 VDD.n285 0.095
R2067 VDD.n489 VDD.n484 0.095
R2068 VDD.n469 VDD.n464 0.095
R2069 VDD.n409 VDD.n404 0.095
R2070 VDD.n389 VDD.n384 0.095
R2071 VDD.n350 VDD.n345 0.095
R2072 VDD.n369 VDD.n364 0.095
R2073 VDD.n429 VDD.n424 0.095
R2074 VDD.n449 VDD.n444 0.095
R2075 VDD.n648 VDD.n643 0.095
R2076 VDD.n628 VDD.n623 0.095
R2077 VDD.n568 VDD.n563 0.095
R2078 VDD.n548 VDD.n543 0.095
R2079 VDD.n509 VDD.n504 0.095
R2080 VDD.n528 VDD.n523 0.095
R2081 VDD.n588 VDD.n583 0.095
R2082 VDD.n608 VDD.n603 0.095
R2083 VDD VDD.n930 0.081
R2084 VDD.n904 VDD.n903 0.079
R2085 VDD.n898 VDD.n897 0.079
R2086 VDD.n892 VDD.n891 0.079
R2087 VDD.n886 VDD.n885 0.079
R2088 VDD.n880 VDD.n879 0.079
R2089 VDD.n874 VDD.n873 0.079
R2090 VDD.n868 VDD.n867 0.079
R2091 VDD.n862 VDD.n861 0.079
R2092 VDD.n7 VDD.n3 0.065
R2093 VDD.n21 VDD.n17 0.065
R2094 VDD.n33 VDD.n31 0.065
R2095 VDD.n48 VDD.n43 0.065
R2096 VDD.n76 VDD.n72 0.065
R2097 VDD.n90 VDD.n86 0.065
R2098 VDD.n62 VDD.n58 0.065
R2099 VDD.n105 VDD.n103 0.065
R2100 VDD.n689 VDD.n682 0.03
R2101 VDD.n789 VDD.n782 0.03
R2102 VDD.n664 VDD.n657 0.03
R2103 VDD.n714 VDD.n707 0.03
R2104 VDD.n739 VDD.n732 0.03
R2105 VDD.n764 VDD.n757 0.03
R2106 VDD.n814 VDD.n807 0.03
R2107 VDD.n839 VDD.n832 0.03
R2108 VDD.n931 VDD 0.028
R2109 VDD VDD.n931 0.028
R2110 VDD.n696 VDD.n695 0.021
R2111 VDD.n704 VDD.n688 0.021
R2112 VDD.n796 VDD.n795 0.021
R2113 VDD.n804 VDD.n788 0.021
R2114 VDD.n671 VDD.n670 0.021
R2115 VDD.n679 VDD.n663 0.021
R2116 VDD.n721 VDD.n720 0.021
R2117 VDD.n729 VDD.n713 0.021
R2118 VDD.n746 VDD.n745 0.021
R2119 VDD.n754 VDD.n738 0.021
R2120 VDD.n771 VDD.n770 0.021
R2121 VDD.n779 VDD.n763 0.021
R2122 VDD.n821 VDD.n820 0.021
R2123 VDD.n829 VDD.n813 0.021
R2124 VDD.n846 VDD.n845 0.021
R2125 VDD.n854 VDD.n838 0.021
R2126 VDD.n864 VDD.t150 0.021
R2127 VDD.n870 VDD.t1115 0.021
R2128 VDD.n900 VDD.t941 0.021
R2129 VDD.n894 VDD.t939 0.021
R2130 VDD.n888 VDD.t635 0.021
R2131 VDD.n882 VDD.t570 0.021
R2132 VDD.n876 VDD.t214 0.021
R2133 VDD.n858 VDD.t387 0.021
R2134 VDD.n931 VDD 0.014
R2135 VDD.n931 VDD 0.014
R2136 VDD.n338 VDD.n337 0.007
R2137 VDD.n318 VDD.n317 0.007
R2138 VDD.n258 VDD.n257 0.007
R2139 VDD.n238 VDD.n237 0.007
R2140 VDD.n218 VDD.n217 0.007
R2141 VDD.n278 VDD.n277 0.007
R2142 VDD.n298 VDD.n297 0.007
R2143 VDD.n497 VDD.n496 0.007
R2144 VDD.n477 VDD.n476 0.007
R2145 VDD.n417 VDD.n416 0.007
R2146 VDD.n397 VDD.n396 0.007
R2147 VDD.n377 VDD.n376 0.007
R2148 VDD.n437 VDD.n436 0.007
R2149 VDD.n457 VDD.n456 0.007
R2150 VDD.n656 VDD.n655 0.007
R2151 VDD.n636 VDD.n635 0.007
R2152 VDD.n576 VDD.n575 0.007
R2153 VDD.n556 VDD.n555 0.007
R2154 VDD.n536 VDD.n535 0.007
R2155 VDD.n596 VDD.n595 0.007
R2156 VDD.n616 VDD.n615 0.007
R2157 VDD.n100 VDD.n39 0.006
R2158 VDD.n115 VDD.n114 0.004
R2159 VDD.n102 VDD.n13 0.003
R2160 VDD.n101 VDD.n27 0.003
R2161 VDD.n99 VDD.n54 0.003
R2162 VDD.n97 VDD.n82 0.003
R2163 VDD.n327 VDD.n325 0.003
R2164 VDD.n307 VDD.n305 0.003
R2165 VDD.n247 VDD.n245 0.003
R2166 VDD.n227 VDD.n225 0.003
R2167 VDD.n188 VDD.n186 0.003
R2168 VDD.n207 VDD.n205 0.003
R2169 VDD.n267 VDD.n265 0.003
R2170 VDD.n287 VDD.n285 0.003
R2171 VDD.n486 VDD.n484 0.003
R2172 VDD.n466 VDD.n464 0.003
R2173 VDD.n406 VDD.n404 0.003
R2174 VDD.n386 VDD.n384 0.003
R2175 VDD.n347 VDD.n345 0.003
R2176 VDD.n366 VDD.n364 0.003
R2177 VDD.n426 VDD.n424 0.003
R2178 VDD.n446 VDD.n444 0.003
R2179 VDD.n645 VDD.n643 0.003
R2180 VDD.n625 VDD.n623 0.003
R2181 VDD.n565 VDD.n563 0.003
R2182 VDD.n545 VDD.n543 0.003
R2183 VDD.n506 VDD.n504 0.003
R2184 VDD.n525 VDD.n523 0.003
R2185 VDD.n585 VDD.n583 0.003
R2186 VDD.n605 VDD.n603 0.003
R2187 VDD.n901 VDD.n899 0.003
R2188 VDD.n895 VDD.n893 0.003
R2189 VDD.n889 VDD.n887 0.003
R2190 VDD.n883 VDD.n881 0.003
R2191 VDD.n877 VDD.n875 0.003
R2192 VDD.n859 VDD.n857 0.003
R2193 VDD.n871 VDD.n869 0.003
R2194 VDD.n865 VDD.n863 0.003
R2195 VDD.n704 VDD.n703 0.002
R2196 VDD.n804 VDD.n803 0.002
R2197 VDD.n679 VDD.n678 0.002
R2198 VDD.n729 VDD.n728 0.002
R2199 VDD.n754 VDD.n753 0.002
R2200 VDD.n779 VDD.n778 0.002
R2201 VDD.n829 VDD.n828 0.002
R2202 VDD.n854 VDD.n853 0.002
R2203 VDD.n705 VDD.n689 0.002
R2204 VDD.n805 VDD.n789 0.002
R2205 VDD.n680 VDD.n664 0.002
R2206 VDD.n730 VDD.n714 0.002
R2207 VDD.n755 VDD.n739 0.002
R2208 VDD.n780 VDD.n764 0.002
R2209 VDD.n830 VDD.n814 0.002
R2210 VDD.n855 VDD.n839 0.002
R2211 VDD.n705 VDD.n704 0.002
R2212 VDD.n805 VDD.n804 0.002
R2213 VDD.n680 VDD.n679 0.002
R2214 VDD.n730 VDD.n729 0.002
R2215 VDD.n755 VDD.n754 0.002
R2216 VDD.n780 VDD.n779 0.002
R2217 VDD.n830 VDD.n829 0.002
R2218 VDD.n855 VDD.n854 0.002
R2219 VDD.n98 VDD.n68 0.002
R2220 VDD.n323 VDD.n321 0.001
R2221 VDD.n303 VDD.n301 0.001
R2222 VDD.n243 VDD.n241 0.001
R2223 VDD.n223 VDD.n221 0.001
R2224 VDD.n184 VDD.n182 0.001
R2225 VDD.n203 VDD.n201 0.001
R2226 VDD.n263 VDD.n261 0.001
R2227 VDD.n283 VDD.n281 0.001
R2228 VDD.n696 VDD.n689 0.001
R2229 VDD.n796 VDD.n789 0.001
R2230 VDD.n671 VDD.n664 0.001
R2231 VDD.n721 VDD.n714 0.001
R2232 VDD.n746 VDD.n739 0.001
R2233 VDD.n771 VDD.n764 0.001
R2234 VDD.n821 VDD.n814 0.001
R2235 VDD.n846 VDD.n839 0.001
R2236 VDD.n482 VDD.n480 0.001
R2237 VDD.n462 VDD.n460 0.001
R2238 VDD.n402 VDD.n400 0.001
R2239 VDD.n382 VDD.n380 0.001
R2240 VDD.n343 VDD.n341 0.001
R2241 VDD.n362 VDD.n360 0.001
R2242 VDD.n422 VDD.n420 0.001
R2243 VDD.n442 VDD.n440 0.001
R2244 VDD.n641 VDD.n639 0.001
R2245 VDD.n621 VDD.n619 0.001
R2246 VDD.n561 VDD.n559 0.001
R2247 VDD.n541 VDD.n539 0.001
R2248 VDD.n502 VDD.n500 0.001
R2249 VDD.n521 VDD.n519 0.001
R2250 VDD.n581 VDD.n579 0.001
R2251 VDD.n601 VDD.n599 0.001
R2252 VDD.n2 VDD.n0 0.001
R2253 VDD.n16 VDD.n14 0.001
R2254 VDD.n30 VDD.n28 0.001
R2255 VDD.n42 VDD.n40 0.001
R2256 VDD.n71 VDD.n69 0.001
R2257 VDD.n85 VDD.n83 0.001
R2258 VDD.n57 VDD.n55 0.001
R2259 VDD.n108 VDD.n106 0.001
R2260 VDD.n706 VDD.n705 0.001
R2261 VDD.n806 VDD.n805 0.001
R2262 VDD.n681 VDD.n680 0.001
R2263 VDD.n731 VDD.n730 0.001
R2264 VDD.n756 VDD.n755 0.001
R2265 VDD.n781 VDD.n780 0.001
R2266 VDD.n831 VDD.n830 0.001
R2267 VDD.n856 VDD.n855 0.001
R2268 VDD.n329 VDD.n328 0.001
R2269 VDD.n309 VDD.n308 0.001
R2270 VDD.n249 VDD.n248 0.001
R2271 VDD.n229 VDD.n228 0.001
R2272 VDD.n190 VDD.n189 0.001
R2273 VDD.n209 VDD.n208 0.001
R2274 VDD.n269 VDD.n268 0.001
R2275 VDD.n289 VDD.n288 0.001
R2276 VDD.n488 VDD.n487 0.001
R2277 VDD.n468 VDD.n467 0.001
R2278 VDD.n408 VDD.n407 0.001
R2279 VDD.n388 VDD.n387 0.001
R2280 VDD.n349 VDD.n348 0.001
R2281 VDD.n368 VDD.n367 0.001
R2282 VDD.n428 VDD.n427 0.001
R2283 VDD.n448 VDD.n447 0.001
R2284 VDD.n647 VDD.n646 0.001
R2285 VDD.n627 VDD.n626 0.001
R2286 VDD.n567 VDD.n566 0.001
R2287 VDD.n547 VDD.n546 0.001
R2288 VDD.n508 VDD.n507 0.001
R2289 VDD.n527 VDD.n526 0.001
R2290 VDD.n587 VDD.n586 0.001
R2291 VDD.n607 VDD.n606 0.001
R2292 VDD.n923 VDD.n172 0.001
R2293 VDD.n924 VDD.n164 0.001
R2294 VDD.n927 VDD.n140 0.001
R2295 VDD.n928 VDD.n132 0.001
R2296 VDD.n930 VDD.n116 0.001
R2297 VDD.n929 VDD.n124 0.001
R2298 VDD.n926 VDD.n148 0.001
R2299 VDD.n925 VDD.n156 0.001
R2300 VDD.n918 VDD.n706 0.001
R2301 VDD.n914 VDD.n806 0.001
R2302 VDD.n919 VDD.n681 0.001
R2303 VDD.n917 VDD.n731 0.001
R2304 VDD.n916 VDD.n756 0.001
R2305 VDD.n915 VDD.n781 0.001
R2306 VDD.n913 VDD.n831 0.001
R2307 VDD.n912 VDD.n856 0.001
R2308 VDD.n703 VDD.n696 0.001
R2309 VDD.n803 VDD.n796 0.001
R2310 VDD.n678 VDD.n671 0.001
R2311 VDD.n728 VDD.n721 0.001
R2312 VDD.n753 VDD.n746 0.001
R2313 VDD.n778 VDD.n771 0.001
R2314 VDD.n828 VDD.n821 0.001
R2315 VDD.n853 VDD.n846 0.001
R2316 VDD.n337 VDD.n323 0.001
R2317 VDD.n330 VDD.n329 0.001
R2318 VDD.n317 VDD.n303 0.001
R2319 VDD.n310 VDD.n309 0.001
R2320 VDD.n257 VDD.n243 0.001
R2321 VDD.n250 VDD.n249 0.001
R2322 VDD.n237 VDD.n223 0.001
R2323 VDD.n230 VDD.n229 0.001
R2324 VDD.n198 VDD.n184 0.001
R2325 VDD.n191 VDD.n190 0.001
R2326 VDD.n217 VDD.n203 0.001
R2327 VDD.n210 VDD.n209 0.001
R2328 VDD.n277 VDD.n263 0.001
R2329 VDD.n270 VDD.n269 0.001
R2330 VDD.n297 VDD.n283 0.001
R2331 VDD.n290 VDD.n289 0.001
R2332 VDD.n904 VDD.n901 0.001
R2333 VDD.n905 VDD.n898 0.001
R2334 VDD.n898 VDD.n895 0.001
R2335 VDD.n906 VDD.n892 0.001
R2336 VDD.n892 VDD.n889 0.001
R2337 VDD.n907 VDD.n886 0.001
R2338 VDD.n886 VDD.n883 0.001
R2339 VDD.n908 VDD.n880 0.001
R2340 VDD.n880 VDD.n877 0.001
R2341 VDD.n909 VDD.n874 0.001
R2342 VDD.n874 VDD.n871 0.001
R2343 VDD.n910 VDD.n868 0.001
R2344 VDD.n868 VDD.n865 0.001
R2345 VDD.n911 VDD.n862 0.001
R2346 VDD.n862 VDD.n859 0.001
R2347 VDD.n496 VDD.n482 0.001
R2348 VDD.n489 VDD.n488 0.001
R2349 VDD.n476 VDD.n462 0.001
R2350 VDD.n469 VDD.n468 0.001
R2351 VDD.n416 VDD.n402 0.001
R2352 VDD.n409 VDD.n408 0.001
R2353 VDD.n396 VDD.n382 0.001
R2354 VDD.n389 VDD.n388 0.001
R2355 VDD.n357 VDD.n343 0.001
R2356 VDD.n350 VDD.n349 0.001
R2357 VDD.n376 VDD.n362 0.001
R2358 VDD.n369 VDD.n368 0.001
R2359 VDD.n436 VDD.n422 0.001
R2360 VDD.n429 VDD.n428 0.001
R2361 VDD.n456 VDD.n442 0.001
R2362 VDD.n449 VDD.n448 0.001
R2363 VDD.n655 VDD.n641 0.001
R2364 VDD.n648 VDD.n647 0.001
R2365 VDD.n635 VDD.n621 0.001
R2366 VDD.n628 VDD.n627 0.001
R2367 VDD.n575 VDD.n561 0.001
R2368 VDD.n568 VDD.n567 0.001
R2369 VDD.n555 VDD.n541 0.001
R2370 VDD.n548 VDD.n547 0.001
R2371 VDD.n516 VDD.n502 0.001
R2372 VDD.n509 VDD.n508 0.001
R2373 VDD.n535 VDD.n521 0.001
R2374 VDD.n528 VDD.n527 0.001
R2375 VDD.n595 VDD.n581 0.001
R2376 VDD.n588 VDD.n587 0.001
R2377 VDD.n615 VDD.n601 0.001
R2378 VDD.n608 VDD.n607 0.001
R2379 VDD.n13 VDD.n0 0.001
R2380 VDD.n27 VDD.n14 0.001
R2381 VDD.n39 VDD.n28 0.001
R2382 VDD.n54 VDD.n40 0.001
R2383 VDD.n82 VDD.n69 0.001
R2384 VDD.n96 VDD.n83 0.001
R2385 VDD.n68 VDD.n55 0.001
R2386 VDD.n114 VDD.n108 0.001
R2387 a_3891_1714.n0 a_3891_1714.t1 28.565
R2388 a_3891_1714.t0 a_3891_1714.n0 28.565
R2389 a_3891_1714.n0 a_3891_1714.n4 112.943
R2390 a_3891_1714.n4 a_3891_1714.n2 2880.87
R2391 a_3891_1714.n2 a_3891_1714.t5 408.211
R2392 a_3891_1714.n2 a_3891_1714.t4 990.34
R2393 a_3891_1714.t4 a_3891_1714.n3 160.666
R2394 a_3891_1714.n3 a_3891_1714.t7 286.438
R2395 a_3891_1714.n3 a_3891_1714.t6 286.438
R2396 a_3891_1714.n4 a_3891_1714.n1 112.94
R2397 a_3891_1714.n1 a_3891_1714.t2 28.568
R2398 a_3891_1714.n1 a_3891_1714.t3 17.64
R2399 a_3951_1740.n1 a_3951_1740.n0 167.433
R2400 a_3951_1740.n5 a_3951_1740.n4 167.433
R2401 a_3951_1740.n1 a_3951_1740.t8 104.259
R2402 a_3951_1740.n5 a_3951_1740.t3 104.259
R2403 a_3951_1740.n7 a_3951_1740.n2 89.977
R2404 a_3951_1740.n6 a_3951_1740.n3 89.977
R2405 a_3951_1740.n9 a_3951_1740.n8 89.977
R2406 a_3951_1740.n8 a_3951_1740.n1 77.784
R2407 a_3951_1740.n8 a_3951_1740.n7 77.456
R2408 a_3951_1740.n7 a_3951_1740.n6 77.456
R2409 a_3951_1740.n6 a_3951_1740.n5 75.815
R2410 a_3951_1740.n0 a_3951_1740.t11 14.282
R2411 a_3951_1740.n0 a_3951_1740.t7 14.282
R2412 a_3951_1740.n2 a_3951_1740.t1 14.282
R2413 a_3951_1740.n2 a_3951_1740.t9 14.282
R2414 a_3951_1740.n3 a_3951_1740.t10 14.282
R2415 a_3951_1740.n3 a_3951_1740.t6 14.282
R2416 a_3951_1740.n4 a_3951_1740.t5 14.282
R2417 a_3951_1740.n4 a_3951_1740.t4 14.282
R2418 a_3951_1740.t0 a_3951_1740.n9 14.282
R2419 a_3951_1740.n9 a_3951_1740.t2 14.282
R2420 A[1].n8 A[1].n7 3623.78
R2421 A[1].t19 A[1].t16 575.234
R2422 A[1].t15 A[1].t8 437.233
R2423 A[1].n5 A[1].n4 412.11
R2424 A[1].n1 A[1].t4 394.151
R2425 A[1].n4 A[1].t2 294.653
R2426 A[1].n9 A[1].t3 284.688
R2427 A[1].n0 A[1].t11 269.523
R2428 A[1].t4 A[1].n0 269.523
R2429 A[1].n5 A[1].n3 224.13
R2430 A[1].n12 A[1].t15 220.332
R2431 A[1].n11 A[1].t5 214.686
R2432 A[1].t8 A[1].n11 214.686
R2433 A[1].n2 A[1].t12 198.043
R2434 A[1].n6 A[1].t6 190.121
R2435 A[1].n6 A[1].t0 190.121
R2436 A[1].n12 A[1].n10 183.203
R2437 A[1].n9 A[1].t13 160.666
R2438 A[1].n10 A[1].t19 160.666
R2439 A[1].n0 A[1].t10 160.666
R2440 A[1].n8 A[1].n5 140.87
R2441 A[1].n7 A[1].t7 137.369
R2442 A[1].n10 A[1].n9 115.593
R2443 A[1].n6 A[1].t1 112.466
R2444 A[1].n4 A[1].t9 111.663
R2445 A[1].n3 A[1].n1 97.816
R2446 A[1].n2 A[1].t17 93.989
R2447 A[1].n11 A[1].t14 80.333
R2448 A[1].n1 A[1].t18 80.333
R2449 A[1].n7 A[1].n6 61.856
R2450 A[1].n13 A[1].n12 26.822
R2451 A[1].n13 A[1].n8 8.399
R2452 A[1].n3 A[1].n2 6.615
R2453 A[1] A[1].n13 3.227
R2454 a_3881_n3752.t3 a_3881_n3752.n0 28.565
R2455 a_3881_n3752.n0 a_3881_n3752.t2 28.565
R2456 a_3881_n3752.n0 a_3881_n3752.n1 192.754
R2457 a_3881_n3752.n1 a_3881_n3752.t1 28.568
R2458 a_3881_n3752.n1 a_3881_n3752.n2 0.478
R2459 a_3881_n3752.n2 a_3881_n3752.n3 44.147
R2460 a_3881_n3752.n3 a_3881_n3752.t6 408.211
R2461 a_3881_n3752.n3 a_3881_n3752.t4 990.34
R2462 a_3881_n3752.t4 a_3881_n3752.n4 160.666
R2463 a_3881_n3752.n4 a_3881_n3752.t5 286.438
R2464 a_3881_n3752.n4 a_3881_n3752.t7 286.438
R2465 a_3881_n3752.n2 a_3881_n3752.t0 18.09
R2466 A[0].n8 A[0].n7 4142.82
R2467 A[0].t3 A[0].t15 576.841
R2468 A[0].t9 A[0].t19 437.233
R2469 A[0].n5 A[0].n4 412.11
R2470 A[0].n1 A[0].t6 394.151
R2471 A[0].n4 A[0].t14 294.653
R2472 A[0].n10 A[0].t5 284.688
R2473 A[0].n0 A[0].t10 269.523
R2474 A[0].t6 A[0].n0 269.523
R2475 A[0].n5 A[0].n3 224.13
R2476 A[0].n13 A[0].t9 217.073
R2477 A[0].n12 A[0].t16 214.686
R2478 A[0].t19 A[0].n12 214.686
R2479 A[0].n2 A[0].t18 198.043
R2480 A[0].n13 A[0].n11 185.87
R2481 A[0].n6 A[0].t11 185.301
R2482 A[0].n6 A[0].t2 185.301
R2483 A[0].n0 A[0].t7 160.666
R2484 A[0].n10 A[0].t13 160.666
R2485 A[0].n11 A[0].t3 160.666
R2486 A[0].n7 A[0].t1 140.583
R2487 A[0].n9 A[0].n5 138.409
R2488 A[0].n11 A[0].n10 115.593
R2489 A[0].n4 A[0].t0 111.663
R2490 A[0].n6 A[0].t4 107.646
R2491 A[0].n3 A[0].n1 97.816
R2492 A[0].n2 A[0].t12 93.989
R2493 A[0].n1 A[0].t17 80.333
R2494 A[0].n12 A[0].t8 80.333
R2495 A[0].n7 A[0].n6 61.856
R2496 A[0].n14 A[0].n13 6.821
R2497 A[0].n3 A[0].n2 6.615
R2498 A[0] A[0].n15 4.756
R2499 A[0].n9 A[0].n8 0.198
R2500 A[0].n15 A[0].n14 0.038
R2501 A[0].n14 A[0].n9 0.004
R2502 a_n25_n6671.n1 a_n25_n6671.t6 318.922
R2503 a_n25_n6671.n0 a_n25_n6671.t4 273.935
R2504 a_n25_n6671.n0 a_n25_n6671.t7 273.935
R2505 a_n25_n6671.n1 a_n25_n6671.t5 269.116
R2506 a_n25_n6671.n4 a_n25_n6671.n3 193.227
R2507 a_n25_n6671.t6 a_n25_n6671.n0 179.142
R2508 a_n25_n6671.n2 a_n25_n6671.n1 106.999
R2509 a_n25_n6671.n3 a_n25_n6671.t0 28.568
R2510 a_n25_n6671.n4 a_n25_n6671.t1 28.565
R2511 a_n25_n6671.t2 a_n25_n6671.n4 28.565
R2512 a_n25_n6671.n2 a_n25_n6671.t3 18.149
R2513 a_n25_n6671.n3 a_n25_n6671.n2 3.726
R2514 VSS.n89 VSS.t29 20.763
R2515 VSS.n79 VSS.t83 20.763
R2516 VSS.n119 VSS.t147 20.763
R2517 VSS.n98 VSS.t169 20.763
R2518 VSS.n127 VSS.t26 20.763
R2519 VSS.n61 VSS.t45 20.763
R2520 VSS.n143 VSS.t155 20.763
R2521 VSS.n52 VSS.t74 20.763
R2522 VSS.n138 VSS.t36 20.676
R2523 VSS.n146 VSS.t86 20.676
R2524 VSS.n110 VSS.t63 20.675
R2525 VSS.n123 VSS.t44 20.675
R2526 VSS.n121 VSS.t17 20.675
R2527 VSS.n100 VSS.t154 20.675
R2528 VSS.n128 VSS.t80 20.675
R2529 VSS.n156 VSS.t34 20.675
R2530 VSS.n154 VSS.t92 18.459
R2531 VSS.n40 VSS.t136 18.459
R2532 VSS.n17 VSS.t126 18.459
R2533 VSS.n50 VSS.t49 18.459
R2534 VSS.n145 VSS.t62 18.459
R2535 VSS.n140 VSS.t152 18.452
R2536 VSS.n1 VSS.t118 18.452
R2537 VSS.n44 VSS.t37 18.452
R2538 VSS.n108 VSS.t166 18.178
R2539 VSS.n124 VSS.t145 18.178
R2540 VSS.n137 VSS.t148 18.178
R2541 VSS.n129 VSS.t84 18.178
R2542 VSS.n111 VSS.t91 18.178
R2543 VSS.n120 VSS.t9 18.178
R2544 VSS.n122 VSS.t82 18.178
R2545 VSS.n99 VSS.t128 18.178
R2546 VSS.n28 VSS.t31 17.972
R2547 VSS.n29 VSS.t127 17.97
R2548 VSS VSS.t64 17.97
R2549 VSS.n41 VSS.t38 17.961
R2550 VSS.n42 VSS.t59 17.959
R2551 VSS.n41 VSS.t81 17.959
R2552 VSS VSS.t153 17.959
R2553 VSS VSS.t13 17.959
R2554 VSS.n93 VSS.t4 17.509
R2555 VSS.n80 VSS.t54 17.509
R2556 VSS.n75 VSS.t158 17.509
R2557 VSS.n65 VSS.t0 17.509
R2558 VSS.n56 VSS.t22 17.509
R2559 VSS.n36 VSS.t8 17.509
R2560 VSS.n18 VSS.t100 17.509
R2561 VSS.n114 VSS.t144 17.509
R2562 VSS.n131 VSS.t173 17.509
R2563 VSS.n72 VSS.t87 17.509
R2564 VSS.n53 VSS.t131 17.509
R2565 VSS.n21 VSS.t97 17.509
R2566 VSS.n33 VSS.t172 17.509
R2567 VSS.n90 VSS.t170 17.509
R2568 VSS.n69 VSS.t101 17.509
R2569 VSS.n62 VSS.t53 17.509
R2570 VSS.n147 VSS.t159 17.509
R2571 VSS.n101 VSS.t43 17.509
R2572 VSS.n84 VSS.t1 17.509
R2573 VSS.n24 VSS.t5 17.509
R2574 VSS.n30 VSS.t139 17.509
R2575 VSS.n4 VSS.t23 17.509
R2576 VSS.n9 VSS.t132 17.509
R2577 VSS.n157 VSS.t124 17.509
R2578 VSS.n94 VSS.t14 17.505
R2579 VSS.n81 VSS.t51 17.505
R2580 VSS.n76 VSS.t164 17.505
R2581 VSS.n66 VSS.t156 17.505
R2582 VSS.n57 VSS.t21 17.505
R2583 VSS.n37 VSS.t108 17.505
R2584 VSS.n19 VSS.t167 17.505
R2585 VSS.n115 VSS.t165 17.505
R2586 VSS.n132 VSS.t175 17.505
R2587 VSS.n73 VSS.t70 17.505
R2588 VSS.n54 VSS.t32 17.505
R2589 VSS.n22 VSS.t135 17.505
R2590 VSS.n34 VSS.t89 17.505
R2591 VSS.n91 VSS.t57 17.505
R2592 VSS.n70 VSS.t48 17.505
R2593 VSS.n63 VSS.t114 17.505
R2594 VSS.n148 VSS.t134 17.505
R2595 VSS.n102 VSS.t104 17.505
R2596 VSS.n85 VSS.t24 17.505
R2597 VSS.n25 VSS.t129 17.505
R2598 VSS.n31 VSS.t146 17.505
R2599 VSS.n5 VSS.t168 17.505
R2600 VSS.n10 VSS.t151 17.505
R2601 VSS.n158 VSS.t99 17.505
R2602 VSS.n139 VSS.t137 17.4
R2603 VSS.n139 VSS.t20 17.4
R2604 VSS.n153 VSS.t85 17.4
R2605 VSS.n153 VSS.t2 17.4
R2606 VSS.n39 VSS.t12 17.4
R2607 VSS.n39 VSS.t75 17.4
R2608 VSS.n16 VSS.t11 17.4
R2609 VSS.n16 VSS.t110 17.4
R2610 VSS.n49 VSS.t171 17.4
R2611 VSS.n49 VSS.t15 17.4
R2612 VSS.n144 VSS.t105 17.4
R2613 VSS.n144 VSS.t78 17.4
R2614 VSS.n0 VSS.t125 17.4
R2615 VSS.n0 VSS.t25 17.4
R2616 VSS.n43 VSS.t141 17.4
R2617 VSS.n43 VSS.t174 17.4
R2618 VSS.n108 VSS.t76 9.319
R2619 VSS.n124 VSS.t130 9.319
R2620 VSS.n137 VSS.t72 9.319
R2621 VSS.n129 VSS.t111 9.319
R2622 VSS.n111 VSS.t47 9.319
R2623 VSS.n120 VSS.t16 9.319
R2624 VSS.n122 VSS.t66 9.319
R2625 VSS.n99 VSS.t30 9.319
R2626 VSS.n94 VSS.t18 8.702
R2627 VSS.n93 VSS.t41 8.702
R2628 VSS.n81 VSS.t90 8.702
R2629 VSS.n80 VSS.t121 8.702
R2630 VSS.n76 VSS.t116 8.702
R2631 VSS.n75 VSS.t106 8.702
R2632 VSS.n66 VSS.t123 8.702
R2633 VSS.n65 VSS.t94 8.702
R2634 VSS.n57 VSS.t35 8.702
R2635 VSS.n56 VSS.t19 8.702
R2636 VSS.n37 VSS.t138 8.702
R2637 VSS.n36 VSS.t161 8.702
R2638 VSS.n19 VSS.t50 8.702
R2639 VSS.n18 VSS.t140 8.702
R2640 VSS.n115 VSS.t33 8.702
R2641 VSS.n114 VSS.t122 8.702
R2642 VSS.n132 VSS.t157 8.702
R2643 VSS.n131 VSS.t93 8.702
R2644 VSS.n73 VSS.t79 8.702
R2645 VSS.n72 VSS.t52 8.702
R2646 VSS.n54 VSS.t68 8.702
R2647 VSS.n53 VSS.t56 8.702
R2648 VSS.n22 VSS.t39 8.702
R2649 VSS.n21 VSS.t98 8.702
R2650 VSS.n34 VSS.t142 8.702
R2651 VSS.n33 VSS.t149 8.702
R2652 VSS.n91 VSS.t42 8.702
R2653 VSS.n90 VSS.t28 8.702
R2654 VSS.n70 VSS.t58 8.702
R2655 VSS.n69 VSS.t143 8.702
R2656 VSS.n63 VSS.t133 8.702
R2657 VSS.n62 VSS.t61 8.702
R2658 VSS.n148 VSS.t160 8.702
R2659 VSS.n147 VSS.t71 8.702
R2660 VSS.n102 VSS.t115 8.702
R2661 VSS.n101 VSS.t107 8.702
R2662 VSS.n85 VSS.t60 8.702
R2663 VSS.n84 VSS.t6 8.702
R2664 VSS.n25 VSS.t46 8.702
R2665 VSS.n24 VSS.t3 8.702
R2666 VSS.n31 VSS.t112 8.702
R2667 VSS.n30 VSS.t109 8.702
R2668 VSS.n5 VSS.t113 8.702
R2669 VSS.n4 VSS.t102 8.702
R2670 VSS.n10 VSS.t120 8.702
R2671 VSS.n9 VSS.t27 8.702
R2672 VSS.n158 VSS.t150 8.702
R2673 VSS.n157 VSS.t119 8.702
R2674 VSS.n88 VSS.t103 8.7
R2675 VSS.n88 VSS.t77 8.7
R2676 VSS.n78 VSS.t96 8.7
R2677 VSS.n78 VSS.t69 8.7
R2678 VSS.n118 VSS.t95 8.7
R2679 VSS.n118 VSS.t65 8.7
R2680 VSS.n97 VSS.t163 8.7
R2681 VSS.n97 VSS.t7 8.7
R2682 VSS.n126 VSS.t55 8.7
R2683 VSS.n126 VSS.t67 8.7
R2684 VSS.n60 VSS.t117 8.7
R2685 VSS.n60 VSS.t88 8.7
R2686 VSS.n142 VSS.t162 8.7
R2687 VSS.n142 VSS.t10 8.7
R2688 VSS.n51 VSS.t40 8.7
R2689 VSS.n51 VSS.t73 8.7
R2690 VSS.n95 VSS.n93 2.025
R2691 VSS.n82 VSS.n80 2.025
R2692 VSS.n77 VSS.n75 2.025
R2693 VSS.n67 VSS.n65 2.025
R2694 VSS.n58 VSS.n56 2.025
R2695 VSS.n38 VSS.n36 2.025
R2696 VSS.n20 VSS.n18 2.025
R2697 VSS.n116 VSS.n114 2.025
R2698 VSS.n133 VSS.n131 2.025
R2699 VSS.n74 VSS.n72 2.025
R2700 VSS.n55 VSS.n53 2.025
R2701 VSS.n23 VSS.n21 2.025
R2702 VSS.n35 VSS.n33 2.025
R2703 VSS.n92 VSS.n90 2.025
R2704 VSS.n71 VSS.n69 2.025
R2705 VSS.n64 VSS.n62 2.025
R2706 VSS.n149 VSS.n147 2.025
R2707 VSS.n103 VSS.n101 2.025
R2708 VSS.n86 VSS.n84 2.025
R2709 VSS.n26 VSS.n24 2.025
R2710 VSS.n32 VSS.n30 2.025
R2711 VSS.n6 VSS.n4 2.025
R2712 VSS.n11 VSS.n9 2.025
R2713 VSS.n159 VSS.n157 2.025
R2714 VSS.n95 VSS.n94 1.953
R2715 VSS.n82 VSS.n81 1.953
R2716 VSS.n77 VSS.n76 1.953
R2717 VSS.n67 VSS.n66 1.953
R2718 VSS.n58 VSS.n57 1.953
R2719 VSS.n38 VSS.n37 1.953
R2720 VSS.n20 VSS.n19 1.953
R2721 VSS.n116 VSS.n115 1.953
R2722 VSS.n133 VSS.n132 1.953
R2723 VSS.n74 VSS.n73 1.953
R2724 VSS.n55 VSS.n54 1.953
R2725 VSS.n23 VSS.n22 1.953
R2726 VSS.n35 VSS.n34 1.953
R2727 VSS.n92 VSS.n91 1.953
R2728 VSS.n71 VSS.n70 1.953
R2729 VSS.n64 VSS.n63 1.953
R2730 VSS.n149 VSS.n148 1.953
R2731 VSS.n103 VSS.n102 1.953
R2732 VSS.n86 VSS.n85 1.953
R2733 VSS.n26 VSS.n25 1.953
R2734 VSS.n32 VSS.n31 1.953
R2735 VSS.n6 VSS.n5 1.953
R2736 VSS.n11 VSS.n10 1.953
R2737 VSS.n159 VSS.n158 1.953
R2738 VSS.n89 VSS.n88 0.948
R2739 VSS.n79 VSS.n78 0.948
R2740 VSS.n119 VSS.n118 0.948
R2741 VSS.n98 VSS.n97 0.948
R2742 VSS.n127 VSS.n126 0.948
R2743 VSS.n61 VSS.n60 0.948
R2744 VSS.n143 VSS.n142 0.948
R2745 VSS.n52 VSS.n51 0.948
R2746 VSS.n154 VSS.n153 0.533
R2747 VSS.n40 VSS.n39 0.533
R2748 VSS.n17 VSS.n16 0.533
R2749 VSS.n50 VSS.n49 0.533
R2750 VSS.n145 VSS.n144 0.533
R2751 VSS.n140 VSS.n139 0.526
R2752 VSS.n1 VSS.n0 0.526
R2753 VSS.n44 VSS.n43 0.526
R2754 VSS.n109 VSS.n108 0.309
R2755 VSS.n125 VSS.n124 0.309
R2756 VSS.n138 VSS.n137 0.309
R2757 VSS.n130 VSS.n129 0.309
R2758 VSS.n112 VSS.n111 0.309
R2759 VSS.n121 VSS.n120 0.309
R2760 VSS.n123 VSS.n122 0.309
R2761 VSS.n100 VSS.n99 0.309
R2762 VSS.n110 VSS.n89 0.197
R2763 VSS.n123 VSS.n79 0.197
R2764 VSS.n100 VSS.n98 0.197
R2765 VSS.n138 VSS.n61 0.197
R2766 VSS.n146 VSS.n143 0.197
R2767 VSS.n156 VSS.n52 0.197
R2768 VSS.n128 VSS.n127 0.196
R2769 VSS.n121 VSS.n119 0.196
R2770 VSS.n156 VSS.n50 0.176
R2771 VSS.n141 VSS.n140 0.174
R2772 VSS.n146 VSS.n145 0.173
R2773 VSS.n155 VSS.n154 0.172
R2774 VSS.n41 VSS.n40 0.172
R2775 VSS.n42 VSS.n17 0.172
R2776 VSS.n2 VSS.n1 0.17
R2777 VSS.n45 VSS.n44 0.17
R2778 VSS.n27 VSS.n20 0.103
R2779 VSS.n41 VSS.n38 0.101
R2780 VSS.n41 VSS.n32 0.099
R2781 VSS.n136 VSS.n64 0.099
R2782 VSS.n134 VSS.n133 0.099
R2783 VSS.n27 VSS.n23 0.098
R2784 VSS.n41 VSS.n35 0.098
R2785 VSS.n125 VSS.n74 0.098
R2786 VSS.n125 VSS.n71 0.098
R2787 VSS.n27 VSS.n26 0.098
R2788 VSS.n125 VSS.n77 0.098
R2789 VSS.n152 VSS.n55 0.098
R2790 VSS.n106 VSS.n92 0.098
R2791 VSS.n150 VSS.n149 0.098
R2792 VSS.n104 VSS.n103 0.098
R2793 VSS.n87 VSS.n86 0.097
R2794 VSS.n117 VSS.n116 0.097
R2795 VSS.n83 VSS.n82 0.097
R2796 VSS.n96 VSS.n95 0.097
R2797 VSS.n68 VSS.n67 0.097
R2798 VSS.n59 VSS.n58 0.097
R2799 VSS.n7 VSS.n6 0.095
R2800 VSS.n12 VSS.n11 0.095
R2801 VSS.n160 VSS.n159 0.095
R2802 VSS VSS.n48 0.019
R2803 VSS VSS.n47 0.019
R2804 VSS VSS.n15 0.019
R2805 VSS.n105 VSS.n96 0.006
R2806 VSS.n135 VSS.n68 0.006
R2807 VSS.n151 VSS.n59 0.006
R2808 VSS.n117 VSS.n113 0.003
R2809 VSS.n28 VSS.n27 0.003
R2810 VSS.n123 VSS.n121 0.003
R2811 VSS.n138 VSS.n136 0.002
R2812 VSS.n155 VSS.n152 0.002
R2813 VSS.n107 VSS.n106 0.002
R2814 VSS VSS.n2 0.002
R2815 VSS VSS.n45 0.002
R2816 VSS.n42 VSS.n41 0.002
R2817 VSS VSS.n156 0.002
R2818 VSS.n146 VSS.n141 0.002
R2819 VSS.n135 VSS.n130 0.002
R2820 VSS.n8 VSS.n7 0.001
R2821 VSS.n13 VSS.n12 0.001
R2822 VSS.n161 VSS.n160 0.001
R2823 VSS.n29 VSS.n28 0.001
R2824 VSS.n41 VSS.n29 0.001
R2825 VSS VSS.n42 0.001
R2826 VSS.n156 VSS.n155 0.001
R2827 VSS.n151 VSS.n146 0.001
R2828 VSS.n141 VSS.n138 0.001
R2829 VSS.n130 VSS.n128 0.001
R2830 VSS.n128 VSS.n125 0.001
R2831 VSS.n125 VSS.n123 0.001
R2832 VSS.n113 VSS.n112 0.001
R2833 VSS.n112 VSS.n110 0.001
R2834 VSS.n110 VSS.n109 0.001
R2835 VSS.n109 VSS.n107 0.001
R2836 VSS.n105 VSS.n100 0.001
R2837 VSS.n121 VSS.n87 0.001
R2838 VSS.n121 VSS.n117 0.001
R2839 VSS.n121 VSS.n83 0.001
R2840 VSS.n151 VSS.n150 0.001
R2841 VSS.n105 VSS.n104 0.001
R2842 VSS.n152 VSS.n151 0.001
R2843 VSS.n106 VSS.n105 0.001
R2844 VSS VSS.n3 0.001
R2845 VSS VSS.n14 0.001
R2846 VSS VSS.n46 0.001
R2847 VSS VSS.n8 0.001
R2848 VSS VSS.n13 0.001
R2849 VSS.n161 VSS 0.001
R2850 VSS.n135 VSS.n134 0.001
R2851 VSS.n136 VSS.n135 0.001
R2852 A[7].n8 A[7].n7 2070.12
R2853 A[7].t4 A[7].t9 573.627
R2854 A[7].t1 A[7].t13 437.233
R2855 A[7].n5 A[7].n4 412.11
R2856 A[7].n1 A[7].t10 394.151
R2857 A[7].n4 A[7].t7 294.653
R2858 A[7].n9 A[7].t18 285.543
R2859 A[7].n0 A[7].t14 269.523
R2860 A[7].t10 A[7].n0 269.523
R2861 A[7].n5 A[7].n3 224.13
R2862 A[7].n12 A[7].t1 223.33
R2863 A[7].n11 A[7].t8 214.686
R2864 A[7].t13 A[7].n11 214.686
R2865 A[7].n2 A[7].t16 198.043
R2866 A[7].n6 A[7].t2 185.301
R2867 A[7].n6 A[7].t3 185.301
R2868 A[7].n12 A[7].n10 181.056
R2869 A[7].n9 A[7].t11 160.666
R2870 A[7].n10 A[7].t4 160.666
R2871 A[7].n0 A[7].t12 160.666
R2872 A[7].n8 A[7].n5 142.556
R2873 A[7].n7 A[7].t6 137.369
R2874 A[7].n10 A[7].n9 114.089
R2875 A[7].n4 A[7].t15 111.663
R2876 A[7].n6 A[7].t19 107.646
R2877 A[7].n3 A[7].n1 97.816
R2878 A[7].n2 A[7].t17 93.989
R2879 A[7].n11 A[7].t0 80.333
R2880 A[7].n1 A[7].t5 80.333
R2881 A[7].n7 A[7].n6 61.856
R2882 A[7].n13 A[7].n12 42.073
R2883 A[7].n13 A[7].n8 32.163
R2884 A[7].n3 A[7].n2 6.615
R2885 A[7] A[7].n13 0.637
R2886 a_10615_3699.n0 a_10615_3699.t8 214.335
R2887 a_10615_3699.t7 a_10615_3699.n0 214.335
R2888 a_10615_3699.n1 a_10615_3699.t7 143.851
R2889 a_10615_3699.n1 a_10615_3699.t9 135.658
R2890 a_10615_3699.n0 a_10615_3699.t10 80.333
R2891 a_10615_3699.n2 a_10615_3699.t6 28.565
R2892 a_10615_3699.n2 a_10615_3699.t4 28.565
R2893 a_10615_3699.n4 a_10615_3699.t5 28.565
R2894 a_10615_3699.n4 a_10615_3699.t0 28.565
R2895 a_10615_3699.t2 a_10615_3699.n7 28.565
R2896 a_10615_3699.n7 a_10615_3699.t1 28.565
R2897 a_10615_3699.n6 a_10615_3699.t3 9.714
R2898 a_10615_3699.n7 a_10615_3699.n6 1.003
R2899 a_10615_3699.n5 a_10615_3699.n3 0.833
R2900 a_10615_3699.n3 a_10615_3699.n2 0.653
R2901 a_10615_3699.n5 a_10615_3699.n4 0.653
R2902 a_10615_3699.n6 a_10615_3699.n5 0.341
R2903 a_10615_3699.n3 a_10615_3699.n1 0.032
R2904 opcode[0].n45 opcode[0].t10 1374.12
R2905 opcode[0].n41 opcode[0].t93 1374.12
R2906 opcode[0].n37 opcode[0].t32 1374.12
R2907 opcode[0].n33 opcode[0].t113 1374.12
R2908 opcode[0].n29 opcode[0].t52 1374.12
R2909 opcode[0].n25 opcode[0].t7 1374.12
R2910 opcode[0].n21 opcode[0].t111 1374.12
R2911 opcode[0].n17 opcode[0].t38 1374.12
R2912 opcode[0].n48 opcode[0].t15 1374.12
R2913 opcode[0].n90 opcode[0].t101 1374.12
R2914 opcode[0].n86 opcode[0].t39 1374.12
R2915 opcode[0].n82 opcode[0].t116 1374.12
R2916 opcode[0].n78 opcode[0].t33 1374.12
R2917 opcode[0].n74 opcode[0].t18 1374.12
R2918 opcode[0].n70 opcode[0].t66 1374.12
R2919 opcode[0].n66 opcode[0].t12 1374.12
R2920 opcode[0].n1 opcode[0].t122 623.291
R2921 opcode[0].n3 opcode[0].t82 623.291
R2922 opcode[0].n5 opcode[0].t105 623.291
R2923 opcode[0].n7 opcode[0].t75 623.291
R2924 opcode[0].n9 opcode[0].t11 623.291
R2925 opcode[0].n11 opcode[0].t110 623.291
R2926 opcode[0].n13 opcode[0].t58 623.291
R2927 opcode[0].n15 opcode[0].t60 623.291
R2928 opcode[0].n50 opcode[0].t13 623.291
R2929 opcode[0].n52 opcode[0].t56 623.291
R2930 opcode[0].n54 opcode[0].t107 623.291
R2931 opcode[0].n56 opcode[0].t3 623.291
R2932 opcode[0].n58 opcode[0].t49 623.291
R2933 opcode[0].n60 opcode[0].t120 623.291
R2934 opcode[0].n62 opcode[0].t27 623.291
R2935 opcode[0].n64 opcode[0].t29 623.291
R2936 opcode[0].n1 opcode[0].t2 610.283
R2937 opcode[0].n3 opcode[0].t80 610.283
R2938 opcode[0].n5 opcode[0].t16 610.283
R2939 opcode[0].n7 opcode[0].t98 610.283
R2940 opcode[0].n9 opcode[0].t21 610.283
R2941 opcode[0].n11 opcode[0].t23 610.283
R2942 opcode[0].n13 opcode[0].t96 610.283
R2943 opcode[0].n15 opcode[0].t24 610.283
R2944 opcode[0].n50 opcode[0].t76 610.283
R2945 opcode[0].n52 opcode[0].t36 610.283
R2946 opcode[0].n54 opcode[0].t91 610.283
R2947 opcode[0].n56 opcode[0].t43 610.283
R2948 opcode[0].n58 opcode[0].t64 610.283
R2949 opcode[0].n60 opcode[0].t54 610.283
R2950 opcode[0].n62 opcode[0].t125 610.283
R2951 opcode[0].n64 opcode[0].t73 610.283
R2952 opcode[0].n45 opcode[0].t118 326.034
R2953 opcode[0].n41 opcode[0].t74 326.034
R2954 opcode[0].n37 opcode[0].t87 326.034
R2955 opcode[0].n33 opcode[0].t90 326.034
R2956 opcode[0].n29 opcode[0].t59 326.034
R2957 opcode[0].n25 opcode[0].t94 326.034
R2958 opcode[0].n21 opcode[0].t123 326.034
R2959 opcode[0].n17 opcode[0].t44 326.034
R2960 opcode[0].n48 opcode[0].t85 326.034
R2961 opcode[0].n90 opcode[0].t114 326.034
R2962 opcode[0].n86 opcode[0].t41 326.034
R2963 opcode[0].n82 opcode[0].t42 326.034
R2964 opcode[0].n78 opcode[0].t67 326.034
R2965 opcode[0].n74 opcode[0].t47 326.034
R2966 opcode[0].n70 opcode[0].t69 326.034
R2967 opcode[0].n66 opcode[0].t84 326.034
R2968 opcode[0].n0 opcode[0].t119 286.438
R2969 opcode[0].n0 opcode[0].t124 286.438
R2970 opcode[0].n2 opcode[0].t78 286.438
R2971 opcode[0].n2 opcode[0].t126 286.438
R2972 opcode[0].n4 opcode[0].t100 286.438
R2973 opcode[0].n4 opcode[0].t89 286.438
R2974 opcode[0].n6 opcode[0].t83 286.438
R2975 opcode[0].n6 opcode[0].t127 286.438
R2976 opcode[0].n8 opcode[0].t104 286.438
R2977 opcode[0].n8 opcode[0].t61 286.438
R2978 opcode[0].n10 opcode[0].t106 286.438
R2979 opcode[0].n10 opcode[0].t115 286.438
R2980 opcode[0].n12 opcode[0].t57 286.438
R2981 opcode[0].n12 opcode[0].t62 286.438
R2982 opcode[0].n14 opcode[0].t20 286.438
R2983 opcode[0].n14 opcode[0].t65 286.438
R2984 opcode[0].n49 opcode[0].t63 286.438
R2985 opcode[0].n49 opcode[0].t71 286.438
R2986 opcode[0].n51 opcode[0].t88 286.438
R2987 opcode[0].n51 opcode[0].t102 286.438
R2988 opcode[0].n53 opcode[0].t17 286.438
R2989 opcode[0].n53 opcode[0].t109 286.438
R2990 opcode[0].n55 opcode[0].t30 286.438
R2991 opcode[0].n55 opcode[0].t81 286.438
R2992 opcode[0].n57 opcode[0].t25 286.438
R2993 opcode[0].n57 opcode[0].t6 286.438
R2994 opcode[0].n59 opcode[0].t28 286.438
R2995 opcode[0].n59 opcode[0].t72 286.438
R2996 opcode[0].n61 opcode[0].t70 286.438
R2997 opcode[0].n61 opcode[0].t77 286.438
R2998 opcode[0].n63 opcode[0].t103 286.438
R2999 opcode[0].n63 opcode[0].t121 286.438
R3000 opcode[0].n44 opcode[0].t34 206.421
R3001 opcode[0].t118 opcode[0].n44 206.421
R3002 opcode[0].n40 opcode[0].t112 206.421
R3003 opcode[0].t74 opcode[0].n40 206.421
R3004 opcode[0].n36 opcode[0].t46 206.421
R3005 opcode[0].t87 opcode[0].n36 206.421
R3006 opcode[0].n32 opcode[0].t99 206.421
R3007 opcode[0].t90 opcode[0].n32 206.421
R3008 opcode[0].n28 opcode[0].t51 206.421
R3009 opcode[0].t59 opcode[0].n28 206.421
R3010 opcode[0].n24 opcode[0].t8 206.421
R3011 opcode[0].t94 opcode[0].n24 206.421
R3012 opcode[0].n20 opcode[0].t40 206.421
R3013 opcode[0].t123 opcode[0].n20 206.421
R3014 opcode[0].n16 opcode[0].t55 206.421
R3015 opcode[0].t44 opcode[0].n16 206.421
R3016 opcode[0].n47 opcode[0].t9 206.421
R3017 opcode[0].t85 opcode[0].n47 206.421
R3018 opcode[0].n89 opcode[0].t0 206.421
R3019 opcode[0].t114 opcode[0].n89 206.421
R3020 opcode[0].n85 opcode[0].t14 206.421
R3021 opcode[0].t41 opcode[0].n85 206.421
R3022 opcode[0].n81 opcode[0].t79 206.421
R3023 opcode[0].t42 opcode[0].n81 206.421
R3024 opcode[0].n77 opcode[0].t19 206.421
R3025 opcode[0].t67 opcode[0].n77 206.421
R3026 opcode[0].n73 opcode[0].t22 206.421
R3027 opcode[0].t47 opcode[0].n73 206.421
R3028 opcode[0].n69 opcode[0].t117 206.421
R3029 opcode[0].t69 opcode[0].n69 206.421
R3030 opcode[0].n65 opcode[0].t5 206.421
R3031 opcode[0].t84 opcode[0].n65 206.421
R3032 opcode[0].t122 opcode[0].n0 160.666
R3033 opcode[0].t82 opcode[0].n2 160.666
R3034 opcode[0].t105 opcode[0].n4 160.666
R3035 opcode[0].t75 opcode[0].n6 160.666
R3036 opcode[0].t11 opcode[0].n8 160.666
R3037 opcode[0].t110 opcode[0].n10 160.666
R3038 opcode[0].t58 opcode[0].n12 160.666
R3039 opcode[0].t60 opcode[0].n14 160.666
R3040 opcode[0].t13 opcode[0].n49 160.666
R3041 opcode[0].t56 opcode[0].n51 160.666
R3042 opcode[0].t107 opcode[0].n53 160.666
R3043 opcode[0].t3 opcode[0].n55 160.666
R3044 opcode[0].t49 opcode[0].n57 160.666
R3045 opcode[0].t120 opcode[0].n59 160.666
R3046 opcode[0].t27 opcode[0].n61 160.666
R3047 opcode[0].t29 opcode[0].n63 160.666
R3048 opcode[0].n44 opcode[0].t31 80.333
R3049 opcode[0].n40 opcode[0].t108 80.333
R3050 opcode[0].n36 opcode[0].t92 80.333
R3051 opcode[0].n32 opcode[0].t95 80.333
R3052 opcode[0].n28 opcode[0].t45 80.333
R3053 opcode[0].n24 opcode[0].t97 80.333
R3054 opcode[0].n20 opcode[0].t35 80.333
R3055 opcode[0].n16 opcode[0].t50 80.333
R3056 opcode[0].n47 opcode[0].t53 80.333
R3057 opcode[0].n89 opcode[0].t37 80.333
R3058 opcode[0].n85 opcode[0].t86 80.333
R3059 opcode[0].n81 opcode[0].t1 80.333
R3060 opcode[0].n77 opcode[0].t68 80.333
R3061 opcode[0].n73 opcode[0].t4 80.333
R3062 opcode[0].n69 opcode[0].t26 80.333
R3063 opcode[0].n65 opcode[0].t48 80.333
R3064 opcode[0].n94 opcode[0].n93 4.767
R3065 opcode[0].n94 opcode[0].n46 3.908
R3066 opcode[0].n80 opcode[0].n79 3.144
R3067 opcode[0].n31 opcode[0].n30 3.103
R3068 opcode[0].n76 opcode[0].n75 3.06
R3069 opcode[0].n92 opcode[0].n91 3.06
R3070 opcode[0].n68 opcode[0].n67 3.038
R3071 opcode[0].n84 opcode[0].n83 3.038
R3072 opcode[0].n72 opcode[0].n71 3.023
R3073 opcode[0].n88 opcode[0].n87 3.023
R3074 opcode[0].n27 opcode[0].n26 3.022
R3075 opcode[0].n43 opcode[0].n42 3.022
R3076 opcode[0].n19 opcode[0].n18 2.998
R3077 opcode[0].n35 opcode[0].n34 2.998
R3078 opcode[0] opcode[0].n94 2.993
R3079 opcode[0].n23 opcode[0].n22 2.985
R3080 opcode[0].n39 opcode[0].n38 2.985
R3081 opcode[0].n75 opcode[0].n72 1.616
R3082 opcode[0].n79 opcode[0].n76 1.616
R3083 opcode[0].n91 opcode[0].n88 1.616
R3084 opcode[0].n93 opcode[0].n92 1.616
R3085 opcode[0].n26 opcode[0].n23 1.597
R3086 opcode[0].n30 opcode[0].n27 1.597
R3087 opcode[0].n42 opcode[0].n39 1.597
R3088 opcode[0].n46 opcode[0].n43 1.597
R3089 opcode[0].n67 opcode[0].n64 1.544
R3090 opcode[0].n71 opcode[0].n68 1.543
R3091 opcode[0].n83 opcode[0].n80 1.543
R3092 opcode[0].n87 opcode[0].n84 1.543
R3093 opcode[0].n18 opcode[0].n15 1.526
R3094 opcode[0].n22 opcode[0].n19 1.525
R3095 opcode[0].n34 opcode[0].n31 1.525
R3096 opcode[0].n38 opcode[0].n35 1.525
R3097 opcode[0].n93 opcode[0].n48 0.003
R3098 opcode[0].n38 opcode[0].n37 0.003
R3099 opcode[0].n34 opcode[0].n33 0.003
R3100 opcode[0].n22 opcode[0].n21 0.003
R3101 opcode[0].n18 opcode[0].n17 0.003
R3102 opcode[0].n87 opcode[0].n86 0.003
R3103 opcode[0].n83 opcode[0].n82 0.003
R3104 opcode[0].n71 opcode[0].n70 0.003
R3105 opcode[0].n67 opcode[0].n66 0.003
R3106 opcode[0].n46 opcode[0].n45 0.003
R3107 opcode[0].n42 opcode[0].n41 0.003
R3108 opcode[0].n30 opcode[0].n29 0.003
R3109 opcode[0].n26 opcode[0].n25 0.003
R3110 opcode[0].n91 opcode[0].n90 0.003
R3111 opcode[0].n79 opcode[0].n78 0.003
R3112 opcode[0].n75 opcode[0].n74 0.003
R3113 opcode[0].n35 opcode[0].n5 0.001
R3114 opcode[0].n31 opcode[0].n7 0.001
R3115 opcode[0].n19 opcode[0].n13 0.001
R3116 opcode[0].n84 opcode[0].n54 0.001
R3117 opcode[0].n80 opcode[0].n56 0.001
R3118 opcode[0].n68 opcode[0].n62 0.001
R3119 opcode[0].n43 opcode[0].n1 0.001
R3120 opcode[0].n39 opcode[0].n3 0.001
R3121 opcode[0].n27 opcode[0].n9 0.001
R3122 opcode[0].n23 opcode[0].n11 0.001
R3123 opcode[0].n92 opcode[0].n50 0.001
R3124 opcode[0].n88 opcode[0].n52 0.001
R3125 opcode[0].n76 opcode[0].n58 0.001
R3126 opcode[0].n72 opcode[0].n60 0.001
R3127 a_3392_1740.n2 a_3392_1740.t7 448.382
R3128 a_3392_1740.n1 a_3392_1740.t4 286.438
R3129 a_3392_1740.n1 a_3392_1740.t5 286.438
R3130 a_3392_1740.n0 a_3392_1740.t6 247.69
R3131 a_3392_1740.n4 a_3392_1740.n3 182.117
R3132 a_3392_1740.t7 a_3392_1740.n1 160.666
R3133 a_3392_1740.n3 a_3392_1740.t0 28.568
R3134 a_3392_1740.t2 a_3392_1740.n4 28.565
R3135 a_3392_1740.n4 a_3392_1740.t1 28.565
R3136 a_3392_1740.n0 a_3392_1740.t3 18.127
R3137 a_3392_1740.n2 a_3392_1740.n0 4.039
R3138 a_3392_1740.n3 a_3392_1740.n2 0.937
R3139 a_12386_n6669.n2 a_12386_n6669.t4 318.922
R3140 a_12386_n6669.n1 a_12386_n6669.t6 273.935
R3141 a_12386_n6669.n1 a_12386_n6669.t5 273.935
R3142 a_12386_n6669.n2 a_12386_n6669.t7 269.116
R3143 a_12386_n6669.n4 a_12386_n6669.n0 193.227
R3144 a_12386_n6669.t4 a_12386_n6669.n1 179.142
R3145 a_12386_n6669.n3 a_12386_n6669.n2 106.999
R3146 a_12386_n6669.t1 a_12386_n6669.n4 28.568
R3147 a_12386_n6669.n0 a_12386_n6669.t3 28.565
R3148 a_12386_n6669.n0 a_12386_n6669.t2 28.565
R3149 a_12386_n6669.n3 a_12386_n6669.t0 18.149
R3150 a_12386_n6669.n4 a_12386_n6669.n3 3.726
R3151 a_12931_n7362.n7 a_12931_n7362.n1 1831.95
R3152 a_12931_n7362.n1 a_12931_n7362.t8 867.497
R3153 a_12931_n7362.n1 a_12931_n7362.t11 615.911
R3154 a_12931_n7362.n0 a_12931_n7362.t10 286.438
R3155 a_12931_n7362.n0 a_12931_n7362.t9 286.438
R3156 a_12931_n7362.t8 a_12931_n7362.n0 160.666
R3157 a_12931_n7362.n5 a_12931_n7362.n3 157.665
R3158 a_12931_n7362.n5 a_12931_n7362.n4 122.999
R3159 a_12931_n7362.n8 a_12931_n7362.n7 90.436
R3160 a_12931_n7362.n6 a_12931_n7362.n2 90.416
R3161 a_12931_n7362.n7 a_12931_n7362.n6 74.302
R3162 a_12931_n7362.n6 a_12931_n7362.n5 50.575
R3163 a_12931_n7362.n2 a_12931_n7362.t3 14.282
R3164 a_12931_n7362.n2 a_12931_n7362.t5 14.282
R3165 a_12931_n7362.n4 a_12931_n7362.t7 14.282
R3166 a_12931_n7362.n4 a_12931_n7362.t4 14.282
R3167 a_12931_n7362.n8 a_12931_n7362.t1 14.282
R3168 a_12931_n7362.t0 a_12931_n7362.n8 14.282
R3169 a_12931_n7362.n3 a_12931_n7362.t2 8.7
R3170 a_12931_n7362.n3 a_12931_n7362.t6 8.7
R3171 a_12813_n7362.n8 a_12813_n7362.n0 267.767
R3172 a_12813_n7362.n4 a_12813_n7362.t9 16.058
R3173 a_12813_n7362.n2 a_12813_n7362.t3 16.058
R3174 a_12813_n7362.n3 a_12813_n7362.t10 14.282
R3175 a_12813_n7362.n3 a_12813_n7362.t11 14.282
R3176 a_12813_n7362.n1 a_12813_n7362.t2 14.282
R3177 a_12813_n7362.n1 a_12813_n7362.t8 14.282
R3178 a_12813_n7362.n6 a_12813_n7362.t5 14.282
R3179 a_12813_n7362.n6 a_12813_n7362.t4 14.282
R3180 a_12813_n7362.n0 a_12813_n7362.t6 14.282
R3181 a_12813_n7362.n0 a_12813_n7362.t7 14.282
R3182 a_12813_n7362.t0 a_12813_n7362.n9 14.282
R3183 a_12813_n7362.n9 a_12813_n7362.t1 14.282
R3184 a_12813_n7362.n7 a_12813_n7362.n6 1.511
R3185 a_12813_n7362.n4 a_12813_n7362.n3 0.999
R3186 a_12813_n7362.n2 a_12813_n7362.n1 0.999
R3187 a_12813_n7362.n8 a_12813_n7362.n7 0.669
R3188 a_12813_n7362.n5 a_12813_n7362.n4 0.575
R3189 a_12813_n7362.n7 a_12813_n7362.n5 0.227
R3190 a_12813_n7362.n5 a_12813_n7362.n2 0.2
R3191 a_12813_n7362.n9 a_12813_n7362.n8 0.001
R3192 a_4290_n3726.n2 a_4290_n3726.t11 1527.4
R3193 a_4290_n3726.t11 a_4290_n3726.n1 657.379
R3194 a_4290_n3726.n4 a_4290_n3726.n3 258.161
R3195 a_4290_n3726.n7 a_4290_n3726.n6 258.161
R3196 a_4290_n3726.n0 a_4290_n3726.t8 206.421
R3197 a_4290_n3726.t10 a_4290_n3726.n0 206.421
R3198 a_4290_n3726.n2 a_4290_n3726.t10 200.029
R3199 a_4290_n3726.n5 a_4290_n3726.n2 97.614
R3200 a_4290_n3726.n0 a_4290_n3726.t9 80.333
R3201 a_4290_n3726.n4 a_4290_n3726.t5 14.283
R3202 a_4290_n3726.n6 a_4290_n3726.t6 14.283
R3203 a_4290_n3726.n3 a_4290_n3726.t3 14.282
R3204 a_4290_n3726.n3 a_4290_n3726.t2 14.282
R3205 a_4290_n3726.t1 a_4290_n3726.n7 14.282
R3206 a_4290_n3726.n7 a_4290_n3726.t7 14.282
R3207 a_4290_n3726.n1 a_4290_n3726.t4 8.7
R3208 a_4290_n3726.n1 a_4290_n3726.t0 8.7
R3209 a_4290_n3726.n5 a_4290_n3726.n4 4.366
R3210 a_4290_n3726.n6 a_4290_n3726.n5 0.852
R3211 a_3891_n1020.t2 a_3891_n1020.n0 28.565
R3212 a_3891_n1020.n0 a_3891_n1020.t1 28.565
R3213 a_3891_n1020.n0 a_3891_n1020.n1 185.55
R3214 a_3891_n1020.n1 a_3891_n1020.t0 28.568
R3215 a_3891_n1020.n1 a_3891_n1020.n4 1.537
R3216 a_3891_n1020.n4 a_3891_n1020.t3 21.473
R3217 a_3891_n1020.n4 a_3891_n1020.n2 13.979
R3218 a_3891_n1020.n2 a_3891_n1020.t7 408.211
R3219 a_3891_n1020.n2 a_3891_n1020.t4 990.34
R3220 a_3891_n1020.t4 a_3891_n1020.n3 160.666
R3221 a_3891_n1020.n3 a_3891_n1020.t6 286.438
R3222 a_3891_n1020.n3 a_3891_n1020.t5 286.438
R3223 a_14881_n7360.n2 a_14881_n7360.n0 267.767
R3224 a_14881_n7360.n8 a_14881_n7360.t2 16.058
R3225 a_14881_n7360.n6 a_14881_n7360.t6 16.058
R3226 a_14881_n7360.n1 a_14881_n7360.t8 14.282
R3227 a_14881_n7360.n1 a_14881_n7360.t3 14.282
R3228 a_14881_n7360.n0 a_14881_n7360.t9 14.282
R3229 a_14881_n7360.n0 a_14881_n7360.t7 14.282
R3230 a_14881_n7360.n3 a_14881_n7360.t4 14.282
R3231 a_14881_n7360.n3 a_14881_n7360.t5 14.282
R3232 a_14881_n7360.n5 a_14881_n7360.t11 14.282
R3233 a_14881_n7360.n5 a_14881_n7360.t10 14.282
R3234 a_14881_n7360.n9 a_14881_n7360.t1 14.282
R3235 a_14881_n7360.t0 a_14881_n7360.n9 14.282
R3236 a_14881_n7360.n4 a_14881_n7360.n3 1.511
R3237 a_14881_n7360.n6 a_14881_n7360.n5 0.999
R3238 a_14881_n7360.n9 a_14881_n7360.n8 0.999
R3239 a_14881_n7360.n4 a_14881_n7360.n2 0.669
R3240 a_14881_n7360.n8 a_14881_n7360.n7 0.575
R3241 a_14881_n7360.n7 a_14881_n7360.n4 0.227
R3242 a_14881_n7360.n7 a_14881_n7360.n6 0.2
R3243 a_14881_n7360.n2 a_14881_n7360.n1 0.001
R3244 a_10852_3062.t0 a_10852_3062.t1 17.4
R3245 a_3951_n994.n2 a_3951_n994.n1 167.433
R3246 a_3951_n994.n6 a_3951_n994.n5 167.433
R3247 a_3951_n994.n2 a_3951_n994.t3 104.259
R3248 a_3951_n994.n6 a_3951_n994.t8 104.259
R3249 a_3951_n994.n3 a_3951_n994.n0 89.977
R3250 a_3951_n994.n7 a_3951_n994.n4 89.977
R3251 a_3951_n994.n9 a_3951_n994.n8 89.977
R3252 a_3951_n994.n3 a_3951_n994.n2 77.784
R3253 a_3951_n994.n8 a_3951_n994.n3 77.456
R3254 a_3951_n994.n8 a_3951_n994.n7 77.456
R3255 a_3951_n994.n7 a_3951_n994.n6 75.815
R3256 a_3951_n994.n1 a_3951_n994.t4 14.282
R3257 a_3951_n994.n1 a_3951_n994.t5 14.282
R3258 a_3951_n994.n0 a_3951_n994.t7 14.282
R3259 a_3951_n994.n0 a_3951_n994.t11 14.282
R3260 a_3951_n994.n4 a_3951_n994.t1 14.282
R3261 a_3951_n994.n4 a_3951_n994.t6 14.282
R3262 a_3951_n994.n5 a_3951_n994.t10 14.282
R3263 a_3951_n994.n5 a_3951_n994.t9 14.282
R3264 a_3951_n994.n9 a_3951_n994.t2 14.282
R3265 a_3951_n994.t0 a_3951_n994.n9 14.282
R3266 opcode[1].n1 opcode[1].t26 1374.12
R3267 opcode[1].n42 opcode[1].t4 1374.12
R3268 opcode[1].n38 opcode[1].t38 1374.12
R3269 opcode[1].n34 opcode[1].t11 1374.12
R3270 opcode[1].n30 opcode[1].t46 1374.12
R3271 opcode[1].n26 opcode[1].t47 1374.12
R3272 opcode[1].n22 opcode[1].t10 1374.12
R3273 opcode[1].n18 opcode[1].t40 1374.12
R3274 opcode[1].n3 opcode[1].t13 623.291
R3275 opcode[1].n5 opcode[1].t36 623.291
R3276 opcode[1].n7 opcode[1].t57 623.291
R3277 opcode[1].n9 opcode[1].t5 623.291
R3278 opcode[1].n11 opcode[1].t34 623.291
R3279 opcode[1].n24 opcode[1].t63 623.291
R3280 opcode[1].n14 opcode[1].t19 623.291
R3281 opcode[1].n16 opcode[1].t21 623.291
R3282 opcode[1].n3 opcode[1].t15 610.283
R3283 opcode[1].n5 opcode[1].t59 610.283
R3284 opcode[1].n7 opcode[1].t28 610.283
R3285 opcode[1].n9 opcode[1].t2 610.283
R3286 opcode[1].n11 opcode[1].t30 610.283
R3287 opcode[1].n24 opcode[1].t32 610.283
R3288 opcode[1].n14 opcode[1].t0 610.283
R3289 opcode[1].n16 opcode[1].t33 610.283
R3290 opcode[1].n1 opcode[1].t53 326.034
R3291 opcode[1].n42 opcode[1].t61 326.034
R3292 opcode[1].n38 opcode[1].t25 326.034
R3293 opcode[1].n34 opcode[1].t27 326.034
R3294 opcode[1].n30 opcode[1].t39 326.034
R3295 opcode[1].n26 opcode[1].t31 326.034
R3296 opcode[1].n22 opcode[1].t42 326.034
R3297 opcode[1].n18 opcode[1].t51 326.034
R3298 opcode[1].n2 opcode[1].t37 286.438
R3299 opcode[1].n2 opcode[1].t44 286.438
R3300 opcode[1].n4 opcode[1].t54 286.438
R3301 opcode[1].n4 opcode[1].t56 286.438
R3302 opcode[1].n6 opcode[1].t14 286.438
R3303 opcode[1].n6 opcode[1].t58 286.438
R3304 opcode[1].n8 opcode[1].t23 286.438
R3305 opcode[1].n8 opcode[1].t50 286.438
R3306 opcode[1].n10 opcode[1].t20 286.438
R3307 opcode[1].n10 opcode[1].t8 286.438
R3308 opcode[1].n12 opcode[1].t22 286.438
R3309 opcode[1].n12 opcode[1].t45 286.438
R3310 opcode[1].n13 opcode[1].t43 286.438
R3311 opcode[1].n13 opcode[1].t48 286.438
R3312 opcode[1].n15 opcode[1].t55 286.438
R3313 opcode[1].n15 opcode[1].t62 286.438
R3314 opcode[1].n0 opcode[1].t9 206.421
R3315 opcode[1].t53 opcode[1].n0 206.421
R3316 opcode[1].n41 opcode[1].t1 206.421
R3317 opcode[1].t61 opcode[1].n41 206.421
R3318 opcode[1].n37 opcode[1].t12 206.421
R3319 opcode[1].t25 opcode[1].n37 206.421
R3320 opcode[1].n33 opcode[1].t49 206.421
R3321 opcode[1].t27 opcode[1].n33 206.421
R3322 opcode[1].n29 opcode[1].t16 206.421
R3323 opcode[1].t39 opcode[1].n29 206.421
R3324 opcode[1].n25 opcode[1].t17 206.421
R3325 opcode[1].t31 opcode[1].n25 206.421
R3326 opcode[1].n21 opcode[1].t60 206.421
R3327 opcode[1].t42 opcode[1].n21 206.421
R3328 opcode[1].n17 opcode[1].t6 206.421
R3329 opcode[1].t51 opcode[1].n17 206.421
R3330 opcode[1].t13 opcode[1].n2 160.666
R3331 opcode[1].t36 opcode[1].n4 160.666
R3332 opcode[1].t57 opcode[1].n6 160.666
R3333 opcode[1].t5 opcode[1].n8 160.666
R3334 opcode[1].t34 opcode[1].n10 160.666
R3335 opcode[1].t63 opcode[1].n12 160.666
R3336 opcode[1].t19 opcode[1].n13 160.666
R3337 opcode[1].t21 opcode[1].n15 160.666
R3338 opcode[1].n0 opcode[1].t35 80.333
R3339 opcode[1].n41 opcode[1].t24 80.333
R3340 opcode[1].n37 opcode[1].t52 80.333
R3341 opcode[1].n33 opcode[1].t3 80.333
R3342 opcode[1].n29 opcode[1].t41 80.333
R3343 opcode[1].n25 opcode[1].t7 80.333
R3344 opcode[1].n21 opcode[1].t18 80.333
R3345 opcode[1].n17 opcode[1].t29 80.333
R3346 opcode[1] opcode[1].n45 4.374
R3347 opcode[1].n32 opcode[1].n31 3.313
R3348 opcode[1].n28 opcode[1].n27 3.118
R3349 opcode[1].n20 opcode[1].n19 3.09
R3350 opcode[1].n36 opcode[1].n35 3.06
R3351 opcode[1].n44 opcode[1].n43 3.06
R3352 opcode[1].n40 opcode[1].n39 3.037
R3353 opcode[1].n24 opcode[1].n23 2.948
R3354 opcode[1].n39 opcode[1].n36 1.618
R3355 opcode[1].n19 opcode[1].n16 1.617
R3356 opcode[1].n23 opcode[1].n20 1.616
R3357 opcode[1].n31 opcode[1].n28 1.616
R3358 opcode[1].n35 opcode[1].n32 1.616
R3359 opcode[1].n43 opcode[1].n40 1.616
R3360 opcode[1].n45 opcode[1].n44 1.616
R3361 opcode[1].n27 opcode[1].n24 1.613
R3362 opcode[1].n45 opcode[1].n1 0.003
R3363 opcode[1].n43 opcode[1].n42 0.003
R3364 opcode[1].n35 opcode[1].n34 0.003
R3365 opcode[1].n31 opcode[1].n30 0.003
R3366 opcode[1].n27 opcode[1].n26 0.003
R3367 opcode[1].n23 opcode[1].n22 0.003
R3368 opcode[1].n19 opcode[1].n18 0.003
R3369 opcode[1].n39 opcode[1].n38 0.003
R3370 opcode[1].n44 opcode[1].n3 0.001
R3371 opcode[1].n40 opcode[1].n5 0.001
R3372 opcode[1].n36 opcode[1].n7 0.001
R3373 opcode[1].n32 opcode[1].n9 0.001
R3374 opcode[1].n28 opcode[1].n11 0.001
R3375 opcode[1].n20 opcode[1].n14 0.001
R3376 a_20290_n2323.t0 a_20290_n2323.t1 17.4
R3377 a_20054_n990.n4 a_20054_n990.t10 1527.4
R3378 a_20054_n990.t10 a_20054_n990.n3 657.379
R3379 a_20054_n990.n1 a_20054_n990.n0 258.161
R3380 a_20054_n990.n7 a_20054_n990.n6 258.161
R3381 a_20054_n990.n2 a_20054_n990.t8 206.421
R3382 a_20054_n990.t9 a_20054_n990.n2 206.421
R3383 a_20054_n990.n4 a_20054_n990.t9 200.029
R3384 a_20054_n990.n5 a_20054_n990.n4 97.614
R3385 a_20054_n990.n2 a_20054_n990.t11 80.333
R3386 a_20054_n990.n6 a_20054_n990.t3 14.283
R3387 a_20054_n990.n1 a_20054_n990.t5 14.283
R3388 a_20054_n990.n0 a_20054_n990.t7 14.282
R3389 a_20054_n990.n0 a_20054_n990.t6 14.282
R3390 a_20054_n990.n7 a_20054_n990.t4 14.282
R3391 a_20054_n990.t2 a_20054_n990.n7 14.282
R3392 a_20054_n990.n3 a_20054_n990.t1 8.7
R3393 a_20054_n990.n3 a_20054_n990.t0 8.7
R3394 a_20054_n990.n6 a_20054_n990.n5 4.366
R3395 a_20054_n990.n5 a_20054_n990.n1 0.852
R3396 a_2588_n7362.n7 a_2588_n7362.n1 1100.3
R3397 a_2588_n7362.n1 a_2588_n7362.t11 867.497
R3398 a_2588_n7362.n1 a_2588_n7362.t9 615.911
R3399 a_2588_n7362.n0 a_2588_n7362.t10 286.438
R3400 a_2588_n7362.n0 a_2588_n7362.t8 286.438
R3401 a_2588_n7362.t11 a_2588_n7362.n0 160.666
R3402 a_2588_n7362.n5 a_2588_n7362.n3 157.665
R3403 a_2588_n7362.n5 a_2588_n7362.n4 122.999
R3404 a_2588_n7362.n8 a_2588_n7362.n7 90.436
R3405 a_2588_n7362.n6 a_2588_n7362.n2 90.416
R3406 a_2588_n7362.n7 a_2588_n7362.n6 74.302
R3407 a_2588_n7362.n6 a_2588_n7362.n5 50.575
R3408 a_2588_n7362.n2 a_2588_n7362.t2 14.282
R3409 a_2588_n7362.n2 a_2588_n7362.t3 14.282
R3410 a_2588_n7362.n4 a_2588_n7362.t6 14.282
R3411 a_2588_n7362.n4 a_2588_n7362.t5 14.282
R3412 a_2588_n7362.n8 a_2588_n7362.t7 14.282
R3413 a_2588_n7362.t0 a_2588_n7362.n8 14.282
R3414 a_2588_n7362.n3 a_2588_n7362.t1 8.7
R3415 a_2588_n7362.n3 a_2588_n7362.t4 8.7
R3416 a_3941_n3726.n3 a_3941_n3726.n2 167.433
R3417 a_3941_n3726.n7 a_3941_n3726.n6 167.433
R3418 a_3941_n3726.n3 a_3941_n3726.t7 104.259
R3419 a_3941_n3726.n7 a_3941_n3726.t10 104.259
R3420 a_3941_n3726.n4 a_3941_n3726.n1 89.977
R3421 a_3941_n3726.n5 a_3941_n3726.n0 89.977
R3422 a_3941_n3726.n9 a_3941_n3726.n8 89.977
R3423 a_3941_n3726.n4 a_3941_n3726.n3 77.784
R3424 a_3941_n3726.n5 a_3941_n3726.n4 77.456
R3425 a_3941_n3726.n8 a_3941_n3726.n5 77.456
R3426 a_3941_n3726.n8 a_3941_n3726.n7 75.815
R3427 a_3941_n3726.n2 a_3941_n3726.t8 14.282
R3428 a_3941_n3726.n2 a_3941_n3726.t6 14.282
R3429 a_3941_n3726.n1 a_3941_n3726.t0 14.282
R3430 a_3941_n3726.n1 a_3941_n3726.t1 14.282
R3431 a_3941_n3726.n0 a_3941_n3726.t2 14.282
R3432 a_3941_n3726.n0 a_3941_n3726.t4 14.282
R3433 a_3941_n3726.n6 a_3941_n3726.t11 14.282
R3434 a_3941_n3726.n6 a_3941_n3726.t9 14.282
R3435 a_3941_n3726.t3 a_3941_n3726.n9 14.282
R3436 a_3941_n3726.n9 a_3941_n3726.t5 14.282
R3437 a_747_1714.t0 a_747_1714.n0 28.565
R3438 a_747_1714.n0 a_747_1714.t3 28.565
R3439 a_747_1714.n0 a_747_1714.n2 114.449
R3440 a_747_1714.n2 a_747_1714.n3 3288.22
R3441 a_747_1714.n3 a_747_1714.t7 408.211
R3442 a_747_1714.n3 a_747_1714.t4 990.34
R3443 a_747_1714.t4 a_747_1714.n4 160.666
R3444 a_747_1714.n4 a_747_1714.t6 286.438
R3445 a_747_1714.n4 a_747_1714.t5 286.438
R3446 a_747_1714.n2 a_747_1714.n1 99.011
R3447 a_747_1714.n1 a_747_1714.t2 28.568
R3448 a_747_1714.n1 a_747_1714.t1 17.641
R3449 a_807_1740.n3 a_807_1740.n2 167.433
R3450 a_807_1740.n7 a_807_1740.n6 167.433
R3451 a_807_1740.n3 a_807_1740.t4 104.259
R3452 a_807_1740.n7 a_807_1740.t9 104.259
R3453 a_807_1740.n4 a_807_1740.n1 89.977
R3454 a_807_1740.n5 a_807_1740.n0 89.977
R3455 a_807_1740.n9 a_807_1740.n8 89.977
R3456 a_807_1740.n4 a_807_1740.n3 77.784
R3457 a_807_1740.n5 a_807_1740.n4 77.456
R3458 a_807_1740.n8 a_807_1740.n5 77.456
R3459 a_807_1740.n8 a_807_1740.n7 75.815
R3460 a_807_1740.n2 a_807_1740.t5 14.282
R3461 a_807_1740.n2 a_807_1740.t6 14.282
R3462 a_807_1740.n1 a_807_1740.t0 14.282
R3463 a_807_1740.n1 a_807_1740.t2 14.282
R3464 a_807_1740.n0 a_807_1740.t1 14.282
R3465 a_807_1740.n0 a_807_1740.t7 14.282
R3466 a_807_1740.n6 a_807_1740.t11 14.282
R3467 a_807_1740.n6 a_807_1740.t10 14.282
R3468 a_807_1740.n9 a_807_1740.t8 14.282
R3469 a_807_1740.t3 a_807_1740.n9 14.282
R3470 a_6725_n7362.n7 a_6725_n7362.n1 1161.06
R3471 a_6725_n7362.n1 a_6725_n7362.t8 867.497
R3472 a_6725_n7362.n1 a_6725_n7362.t9 615.911
R3473 a_6725_n7362.n0 a_6725_n7362.t11 286.438
R3474 a_6725_n7362.n0 a_6725_n7362.t10 286.438
R3475 a_6725_n7362.t8 a_6725_n7362.n0 160.666
R3476 a_6725_n7362.n5 a_6725_n7362.n3 157.665
R3477 a_6725_n7362.n5 a_6725_n7362.n4 122.999
R3478 a_6725_n7362.n8 a_6725_n7362.n7 90.436
R3479 a_6725_n7362.n6 a_6725_n7362.n2 90.416
R3480 a_6725_n7362.n7 a_6725_n7362.n6 74.302
R3481 a_6725_n7362.n6 a_6725_n7362.n5 50.575
R3482 a_6725_n7362.n2 a_6725_n7362.t7 14.282
R3483 a_6725_n7362.n2 a_6725_n7362.t4 14.282
R3484 a_6725_n7362.n4 a_6725_n7362.t3 14.282
R3485 a_6725_n7362.n4 a_6725_n7362.t2 14.282
R3486 a_6725_n7362.t0 a_6725_n7362.n8 14.282
R3487 a_6725_n7362.n8 a_6725_n7362.t1 14.282
R3488 a_6725_n7362.n3 a_6725_n7362.t6 8.7
R3489 a_6725_n7362.n3 a_6725_n7362.t5 8.7
R3490 a_10566_n3722.n4 a_10566_n3722.t11 1527.4
R3491 a_10566_n3722.t11 a_10566_n3722.n3 657.379
R3492 a_10566_n3722.n1 a_10566_n3722.n0 258.161
R3493 a_10566_n3722.n7 a_10566_n3722.n6 258.161
R3494 a_10566_n3722.n2 a_10566_n3722.t10 206.421
R3495 a_10566_n3722.t9 a_10566_n3722.n2 206.421
R3496 a_10566_n3722.n4 a_10566_n3722.t9 200.029
R3497 a_10566_n3722.n5 a_10566_n3722.n4 97.614
R3498 a_10566_n3722.n2 a_10566_n3722.t8 80.333
R3499 a_10566_n3722.n6 a_10566_n3722.t5 14.283
R3500 a_10566_n3722.n1 a_10566_n3722.t2 14.283
R3501 a_10566_n3722.n0 a_10566_n3722.t3 14.282
R3502 a_10566_n3722.n0 a_10566_n3722.t1 14.282
R3503 a_10566_n3722.t0 a_10566_n3722.n7 14.282
R3504 a_10566_n3722.n7 a_10566_n3722.t6 14.282
R3505 a_10566_n3722.n3 a_10566_n3722.t7 8.7
R3506 a_10566_n3722.n3 a_10566_n3722.t4 8.7
R3507 a_10566_n3722.n6 a_10566_n3722.n5 4.366
R3508 a_10566_n3722.n5 a_10566_n3722.n1 0.852
R3509 a_10217_n3722.n2 a_10217_n3722.n1 167.433
R3510 a_10217_n3722.n6 a_10217_n3722.n5 167.433
R3511 a_10217_n3722.n2 a_10217_n3722.t1 104.259
R3512 a_10217_n3722.n6 a_10217_n3722.t8 104.259
R3513 a_10217_n3722.n3 a_10217_n3722.n0 89.977
R3514 a_10217_n3722.n7 a_10217_n3722.n4 89.977
R3515 a_10217_n3722.n9 a_10217_n3722.n8 89.977
R3516 a_10217_n3722.n3 a_10217_n3722.n2 77.784
R3517 a_10217_n3722.n8 a_10217_n3722.n3 77.456
R3518 a_10217_n3722.n8 a_10217_n3722.n7 77.456
R3519 a_10217_n3722.n7 a_10217_n3722.n6 75.815
R3520 a_10217_n3722.n1 a_10217_n3722.t2 14.282
R3521 a_10217_n3722.n1 a_10217_n3722.t3 14.282
R3522 a_10217_n3722.n0 a_10217_n3722.t4 14.282
R3523 a_10217_n3722.n0 a_10217_n3722.t6 14.282
R3524 a_10217_n3722.n4 a_10217_n3722.t10 14.282
R3525 a_10217_n3722.n4 a_10217_n3722.t9 14.282
R3526 a_10217_n3722.n5 a_10217_n3722.t11 14.282
R3527 a_10217_n3722.n5 a_10217_n3722.t7 14.282
R3528 a_10217_n3722.n9 a_10217_n3722.t5 14.282
R3529 a_10217_n3722.t0 a_10217_n3722.n9 14.282
R3530 a_3392_n994.n2 a_3392_n994.t7 448.382
R3531 a_3392_n994.n1 a_3392_n994.t4 286.438
R3532 a_3392_n994.n1 a_3392_n994.t6 286.438
R3533 a_3392_n994.n0 a_3392_n994.t5 247.69
R3534 a_3392_n994.n4 a_3392_n994.n3 182.117
R3535 a_3392_n994.t7 a_3392_n994.n1 160.666
R3536 a_3392_n994.n3 a_3392_n994.t0 28.568
R3537 a_3392_n994.t2 a_3392_n994.n4 28.565
R3538 a_3392_n994.n4 a_3392_n994.t1 28.565
R3539 a_3392_n994.n0 a_3392_n994.t3 18.127
R3540 a_3392_n994.n2 a_3392_n994.n0 4.039
R3541 a_3392_n994.n3 a_3392_n994.n2 0.937
R3542 a_21997_n6357.t2 a_21997_n6357.n0 28.568
R3543 a_21997_n6357.n0 a_21997_n6357.n4 197.272
R3544 a_21997_n6357.n4 a_21997_n6357.t1 28.565
R3545 a_21997_n6357.n4 a_21997_n6357.t0 28.565
R3546 a_21997_n6357.n0 a_21997_n6357.n1 0.459
R3547 a_21997_n6357.n1 a_21997_n6357.n2 6.445
R3548 a_21997_n6357.n2 a_21997_n6357.t5 408.211
R3549 a_21997_n6357.n2 a_21997_n6357.t7 990.34
R3550 a_21997_n6357.t7 a_21997_n6357.n3 160.666
R3551 a_21997_n6357.n3 a_21997_n6357.t4 286.438
R3552 a_21997_n6357.n3 a_21997_n6357.t6 286.438
R3553 a_21997_n6357.n1 a_21997_n6357.t3 18.092
R3554 A[5].n12 A[5].n5 2643.33
R3555 A[5].t0 A[5].t14 575.234
R3556 A[5].t2 A[5].t10 437.233
R3557 A[5].n11 A[5].n10 412.11
R3558 A[5].n7 A[5].t8 394.151
R3559 A[5].n10 A[5].t5 294.653
R3560 A[5].n0 A[5].t11 285.543
R3561 A[5].n6 A[5].t6 269.523
R3562 A[5].t8 A[5].n6 269.523
R3563 A[5].n11 A[5].n9 224.13
R3564 A[5].n3 A[5].t2 222.157
R3565 A[5].n2 A[5].t4 214.686
R3566 A[5].t10 A[5].n2 214.686
R3567 A[5].n8 A[5].t16 198.043
R3568 A[5].n4 A[5].t19 185.301
R3569 A[5].n4 A[5].t7 185.301
R3570 A[5].n3 A[5].n1 181.495
R3571 A[5].n0 A[5].t9 160.666
R3572 A[5].n1 A[5].t0 160.666
R3573 A[5].n6 A[5].t12 160.666
R3574 A[5].n12 A[5].n11 142.204
R3575 A[5].n5 A[5].t15 140.583
R3576 A[5].n1 A[5].n0 114.089
R3577 A[5].n10 A[5].t13 111.663
R3578 A[5].n4 A[5].t18 107.646
R3579 A[5].n9 A[5].n7 97.816
R3580 A[5].n8 A[5].t17 93.989
R3581 A[5].n2 A[5].t1 80.333
R3582 A[5].n7 A[5].t3 80.333
R3583 A[5].n5 A[5].n4 61.856
R3584 A[5].n13 A[5].n3 40.051
R3585 A[5].n13 A[5].n12 27.336
R3586 A[5].n9 A[5].n8 6.615
R3587 A[5] A[5].n13 1.546
R3588 a_17798_3694.t5 a_17798_3694.n3 405.372
R3589 a_17798_3694.n2 a_17798_3694.t7 207.38
R3590 a_17798_3694.n4 a_17798_3694.t5 138.55
R3591 a_17798_3694.n3 a_17798_3694.n2 112.003
R3592 a_17798_3694.n2 a_17798_3694.t8 80.333
R3593 a_17798_3694.n3 a_17798_3694.t6 80.333
R3594 a_17798_3694.n1 a_17798_3694.t4 17.4
R3595 a_17798_3694.n1 a_17798_3694.t0 17.4
R3596 a_17798_3694.t1 a_17798_3694.n5 15.029
R3597 a_17798_3694.n0 a_17798_3694.t2 14.282
R3598 a_17798_3694.n0 a_17798_3694.t3 14.282
R3599 a_17798_3694.n5 a_17798_3694.n0 1.647
R3600 a_17798_3694.n4 a_17798_3694.n1 0.679
R3601 a_17798_3694.n5 a_17798_3694.n4 0.665
R3602 a_17916_3694.n0 a_17916_3694.t4 14.282
R3603 a_17916_3694.n0 a_17916_3694.t5 14.282
R3604 a_17916_3694.n1 a_17916_3694.t2 14.282
R3605 a_17916_3694.n1 a_17916_3694.t1 14.282
R3606 a_17916_3694.t0 a_17916_3694.n3 14.282
R3607 a_17916_3694.n3 a_17916_3694.t3 14.282
R3608 a_17916_3694.n2 a_17916_3694.n0 2.554
R3609 a_17916_3694.n2 a_17916_3694.n1 2.361
R3610 a_17916_3694.n3 a_17916_3694.n2 0.001
R3611 a_7023_n1016.n0 a_7023_n1016.t2 28.565
R3612 a_7023_n1016.t0 a_7023_n1016.n0 28.565
R3613 a_7023_n1016.n0 a_7023_n1016.n1 185.55
R3614 a_7023_n1016.n1 a_7023_n1016.t1 28.568
R3615 a_7023_n1016.n1 a_7023_n1016.n4 1.537
R3616 a_7023_n1016.n4 a_7023_n1016.t3 21.497
R3617 a_7023_n1016.n4 a_7023_n1016.n2 12.948
R3618 a_7023_n1016.n2 a_7023_n1016.t6 408.211
R3619 a_7023_n1016.n2 a_7023_n1016.t7 990.34
R3620 a_7023_n1016.t7 a_7023_n1016.n3 160.666
R3621 a_7023_n1016.n3 a_7023_n1016.t5 286.438
R3622 a_7023_n1016.n3 a_7023_n1016.t4 286.438
R3623 a_7083_n990.n9 a_7083_n990.n0 167.433
R3624 a_7083_n990.n5 a_7083_n990.n4 167.433
R3625 a_7083_n990.n5 a_7083_n990.t8 104.259
R3626 a_7083_n990.t3 a_7083_n990.n9 104.259
R3627 a_7083_n990.n8 a_7083_n990.n1 89.977
R3628 a_7083_n990.n7 a_7083_n990.n2 89.977
R3629 a_7083_n990.n6 a_7083_n990.n3 89.977
R3630 a_7083_n990.n9 a_7083_n990.n8 77.784
R3631 a_7083_n990.n8 a_7083_n990.n7 77.456
R3632 a_7083_n990.n7 a_7083_n990.n6 77.456
R3633 a_7083_n990.n6 a_7083_n990.n5 75.815
R3634 a_7083_n990.n0 a_7083_n990.t4 14.282
R3635 a_7083_n990.n0 a_7083_n990.t10 14.282
R3636 a_7083_n990.n1 a_7083_n990.t0 14.282
R3637 a_7083_n990.n1 a_7083_n990.t1 14.282
R3638 a_7083_n990.n2 a_7083_n990.t2 14.282
R3639 a_7083_n990.n2 a_7083_n990.t11 14.282
R3640 a_7083_n990.n3 a_7083_n990.t6 14.282
R3641 a_7083_n990.n3 a_7083_n990.t5 14.282
R3642 a_7083_n990.n4 a_7083_n990.t7 14.282
R3643 a_7083_n990.n4 a_7083_n990.t9 14.282
R3644 a_10812_n2323.t0 a_10812_n2323.t1 17.4
R3645 a_10576_n990.n5 a_10576_n990.t8 1527.4
R3646 a_10576_n990.t8 a_10576_n990.n4 657.379
R3647 a_10576_n990.n7 a_10576_n990.n0 258.161
R3648 a_10576_n990.n2 a_10576_n990.n1 258.161
R3649 a_10576_n990.n3 a_10576_n990.t10 206.421
R3650 a_10576_n990.t9 a_10576_n990.n3 206.421
R3651 a_10576_n990.n5 a_10576_n990.t9 200.029
R3652 a_10576_n990.n6 a_10576_n990.n5 97.614
R3653 a_10576_n990.n3 a_10576_n990.t11 80.333
R3654 a_10576_n990.n2 a_10576_n990.t4 14.283
R3655 a_10576_n990.t2 a_10576_n990.n7 14.283
R3656 a_10576_n990.n0 a_10576_n990.t5 14.282
R3657 a_10576_n990.n0 a_10576_n990.t6 14.282
R3658 a_10576_n990.n1 a_10576_n990.t7 14.282
R3659 a_10576_n990.n1 a_10576_n990.t3 14.282
R3660 a_10576_n990.n4 a_10576_n990.t1 8.7
R3661 a_10576_n990.n4 a_10576_n990.t0 8.7
R3662 a_10576_n990.n7 a_10576_n990.n6 4.366
R3663 a_10576_n990.n6 a_10576_n990.n2 0.852
R3664 a_7669_3697.n2 a_7669_3697.t8 214.335
R3665 a_7669_3697.t7 a_7669_3697.n2 214.335
R3666 a_7669_3697.n3 a_7669_3697.t7 143.851
R3667 a_7669_3697.n3 a_7669_3697.t9 135.658
R3668 a_7669_3697.n2 a_7669_3697.t10 80.333
R3669 a_7669_3697.n4 a_7669_3697.t5 28.565
R3670 a_7669_3697.n4 a_7669_3697.t6 28.565
R3671 a_7669_3697.n0 a_7669_3697.t3 28.565
R3672 a_7669_3697.n0 a_7669_3697.t2 28.565
R3673 a_7669_3697.t4 a_7669_3697.n7 28.565
R3674 a_7669_3697.n7 a_7669_3697.t1 28.565
R3675 a_7669_3697.n1 a_7669_3697.t0 9.714
R3676 a_7669_3697.n1 a_7669_3697.n0 1.003
R3677 a_7669_3697.n6 a_7669_3697.n5 0.833
R3678 a_7669_3697.n5 a_7669_3697.n4 0.653
R3679 a_7669_3697.n7 a_7669_3697.n6 0.653
R3680 a_7669_3697.n6 a_7669_3697.n1 0.341
R3681 a_7669_3697.n5 a_7669_3697.n3 0.032
R3682 a_2043_n6669.n2 a_2043_n6669.t6 318.922
R3683 a_2043_n6669.n1 a_2043_n6669.t5 273.935
R3684 a_2043_n6669.n1 a_2043_n6669.t7 273.935
R3685 a_2043_n6669.n2 a_2043_n6669.t4 269.116
R3686 a_2043_n6669.n4 a_2043_n6669.n0 193.227
R3687 a_2043_n6669.t6 a_2043_n6669.n1 179.142
R3688 a_2043_n6669.n3 a_2043_n6669.n2 106.999
R3689 a_2043_n6669.t2 a_2043_n6669.n4 28.568
R3690 a_2043_n6669.n0 a_2043_n6669.t0 28.565
R3691 a_2043_n6669.n0 a_2043_n6669.t1 28.565
R3692 a_2043_n6669.n3 a_2043_n6669.t3 18.149
R3693 a_2043_n6669.n4 a_2043_n6669.n3 3.726
R3694 a_2588_n8094.t0 a_2588_n8094.t1 380.209
R3695 a_11038_n5055.t0 a_11038_n5055.t1 17.4
R3696 a_7906_3060.t0 a_7906_3060.t1 17.4
R3697 a_7023_1718.t1 a_7023_1718.n0 28.565
R3698 a_7023_1718.n0 a_7023_1718.t3 28.565
R3699 a_7023_1718.n0 a_7023_1718.n2 116.875
R3700 a_7023_1718.n2 a_7023_1718.n3 2682.43
R3701 a_7023_1718.n3 a_7023_1718.t7 408.211
R3702 a_7023_1718.n3 a_7023_1718.t6 990.34
R3703 a_7023_1718.t6 a_7023_1718.n4 160.666
R3704 a_7023_1718.n4 a_7023_1718.t5 286.438
R3705 a_7023_1718.n4 a_7023_1718.t4 286.438
R3706 a_7023_1718.n2 a_7023_1718.n1 99.45
R3707 a_7023_1718.n1 a_7023_1718.t2 28.568
R3708 a_7023_1718.n1 a_7023_1718.t0 17.64
R3709 a_7083_1744.n2 a_7083_1744.n1 167.433
R3710 a_7083_1744.n6 a_7083_1744.n5 167.433
R3711 a_7083_1744.n2 a_7083_1744.t9 104.259
R3712 a_7083_1744.n6 a_7083_1744.t5 104.259
R3713 a_7083_1744.n3 a_7083_1744.n0 89.977
R3714 a_7083_1744.n7 a_7083_1744.n4 89.977
R3715 a_7083_1744.n9 a_7083_1744.n8 89.977
R3716 a_7083_1744.n3 a_7083_1744.n2 77.784
R3717 a_7083_1744.n8 a_7083_1744.n3 77.456
R3718 a_7083_1744.n8 a_7083_1744.n7 77.456
R3719 a_7083_1744.n7 a_7083_1744.n6 75.815
R3720 a_7083_1744.n1 a_7083_1744.t10 14.282
R3721 a_7083_1744.n1 a_7083_1744.t7 14.282
R3722 a_7083_1744.n0 a_7083_1744.t0 14.282
R3723 a_7083_1744.n0 a_7083_1744.t1 14.282
R3724 a_7083_1744.n4 a_7083_1744.t8 14.282
R3725 a_7083_1744.n4 a_7083_1744.t11 14.282
R3726 a_7083_1744.n5 a_7083_1744.t4 14.282
R3727 a_7083_1744.n5 a_7083_1744.t6 14.282
R3728 a_7083_1744.n9 a_7083_1744.t2 14.282
R3729 a_7083_1744.t3 a_7083_1744.n9 14.282
R3730 a_747_n1020.n0 a_747_n1020.t3 28.565
R3731 a_747_n1020.t0 a_747_n1020.n0 28.565
R3732 a_747_n1020.n0 a_747_n1020.n1 185.55
R3733 a_747_n1020.n1 a_747_n1020.t1 28.568
R3734 a_747_n1020.n1 a_747_n1020.n4 2.677
R3735 a_747_n1020.n4 a_747_n1020.t2 21.468
R3736 a_747_n1020.n4 a_747_n1020.n2 12.581
R3737 a_747_n1020.n2 a_747_n1020.t5 408.211
R3738 a_747_n1020.n2 a_747_n1020.t4 990.34
R3739 a_747_n1020.t4 a_747_n1020.n3 160.666
R3740 a_747_n1020.n3 a_747_n1020.t7 286.438
R3741 a_747_n1020.n3 a_747_n1020.t6 286.438
R3742 a_807_n994.n4 a_807_n994.n3 167.433
R3743 a_807_n994.n9 a_807_n994.n8 167.433
R3744 a_807_n994.n8 a_807_n994.t6 104.259
R3745 a_807_n994.n4 a_807_n994.t9 104.259
R3746 a_807_n994.n7 a_807_n994.n0 89.977
R3747 a_807_n994.n6 a_807_n994.n1 89.977
R3748 a_807_n994.n5 a_807_n994.n2 89.977
R3749 a_807_n994.n8 a_807_n994.n7 77.784
R3750 a_807_n994.n7 a_807_n994.n6 77.456
R3751 a_807_n994.n6 a_807_n994.n5 77.456
R3752 a_807_n994.n5 a_807_n994.n4 75.815
R3753 a_807_n994.n0 a_807_n994.t0 14.282
R3754 a_807_n994.n0 a_807_n994.t2 14.282
R3755 a_807_n994.n1 a_807_n994.t1 14.282
R3756 a_807_n994.n1 a_807_n994.t4 14.282
R3757 a_807_n994.n2 a_807_n994.t5 14.282
R3758 a_807_n994.n2 a_807_n994.t8 14.282
R3759 a_807_n994.n3 a_807_n994.t11 14.282
R3760 a_807_n994.n3 a_807_n994.t10 14.282
R3761 a_807_n994.n9 a_807_n994.t7 14.282
R3762 a_807_n994.t3 a_807_n994.n9 14.282
R3763 Y[6].n1 Y[6].n0 185.55
R3764 Y[6].n1 Y[6].t1 28.568
R3765 Y[6].n0 Y[6].t0 28.565
R3766 Y[6].n0 Y[6].t2 28.565
R3767 Y[6].n2 Y[6].t3 21.373
R3768 Y[6] Y[6].n2 5.31
R3769 Y[6].n2 Y[6].n1 1.637
R3770 a_10167_n1016.n0 a_10167_n1016.t0 28.565
R3771 a_10167_n1016.t2 a_10167_n1016.n0 28.565
R3772 a_10167_n1016.n0 a_10167_n1016.n1 185.55
R3773 a_10167_n1016.n1 a_10167_n1016.t1 28.568
R3774 a_10167_n1016.n1 a_10167_n1016.n4 1.537
R3775 a_10167_n1016.n4 a_10167_n1016.t3 21.473
R3776 a_10167_n1016.n4 a_10167_n1016.n2 12.306
R3777 a_10167_n1016.n2 a_10167_n1016.t7 408.211
R3778 a_10167_n1016.n2 a_10167_n1016.t6 990.34
R3779 a_10167_n1016.t6 a_10167_n1016.n3 160.666
R3780 a_10167_n1016.n3 a_10167_n1016.t5 286.438
R3781 a_10167_n1016.n3 a_10167_n1016.t4 286.438
R3782 a_11952_3694.t5 a_11952_3694.n3 406.221
R3783 a_11952_3694.n2 a_11952_3694.t7 190.962
R3784 a_11952_3694.n4 a_11952_3694.t5 138.55
R3785 a_11952_3694.n3 a_11952_3694.n2 111.349
R3786 a_11952_3694.n2 a_11952_3694.t8 80.333
R3787 a_11952_3694.n3 a_11952_3694.t6 80.333
R3788 a_11952_3694.n1 a_11952_3694.t0 17.4
R3789 a_11952_3694.n1 a_11952_3694.t2 17.4
R3790 a_11952_3694.t1 a_11952_3694.n5 15.036
R3791 a_11952_3694.n0 a_11952_3694.t3 14.282
R3792 a_11952_3694.n0 a_11952_3694.t4 14.282
R3793 a_11952_3694.n5 a_11952_3694.n0 1.654
R3794 a_11952_3694.n4 a_11952_3694.n1 0.679
R3795 a_11952_3694.n5 a_11952_3694.n4 0.665
R3796 a_4300_1740.n2 a_4300_1740.t8 1527.4
R3797 a_4300_1740.t8 a_4300_1740.n1 657.379
R3798 a_4300_1740.n4 a_4300_1740.n3 258.161
R3799 a_4300_1740.n7 a_4300_1740.n6 258.161
R3800 a_4300_1740.n0 a_4300_1740.t9 206.421
R3801 a_4300_1740.t10 a_4300_1740.n0 206.421
R3802 a_4300_1740.n2 a_4300_1740.t10 200.029
R3803 a_4300_1740.n5 a_4300_1740.n2 97.614
R3804 a_4300_1740.n0 a_4300_1740.t11 80.333
R3805 a_4300_1740.n4 a_4300_1740.t4 14.283
R3806 a_4300_1740.n6 a_4300_1740.t7 14.283
R3807 a_4300_1740.n3 a_4300_1740.t3 14.282
R3808 a_4300_1740.n3 a_4300_1740.t2 14.282
R3809 a_4300_1740.t5 a_4300_1740.n7 14.282
R3810 a_4300_1740.n7 a_4300_1740.t6 14.282
R3811 a_4300_1740.n1 a_4300_1740.t1 8.7
R3812 a_4300_1740.n1 a_4300_1740.t0 8.7
R3813 a_4300_1740.n5 a_4300_1740.n4 4.366
R3814 a_4300_1740.n6 a_4300_1740.n5 0.852
R3815 a_20054_1744.n3 a_20054_1744.t11 1527.4
R3816 a_20054_1744.t11 a_20054_1744.n2 657.379
R3817 a_20054_1744.n5 a_20054_1744.n4 258.161
R3818 a_20054_1744.n7 a_20054_1744.n0 258.161
R3819 a_20054_1744.n1 a_20054_1744.t8 206.421
R3820 a_20054_1744.t9 a_20054_1744.n1 206.421
R3821 a_20054_1744.n3 a_20054_1744.t9 200.029
R3822 a_20054_1744.n6 a_20054_1744.n3 97.614
R3823 a_20054_1744.n1 a_20054_1744.t10 80.333
R3824 a_20054_1744.n5 a_20054_1744.t4 14.283
R3825 a_20054_1744.t2 a_20054_1744.n7 14.283
R3826 a_20054_1744.n4 a_20054_1744.t6 14.282
R3827 a_20054_1744.n4 a_20054_1744.t7 14.282
R3828 a_20054_1744.n0 a_20054_1744.t5 14.282
R3829 a_20054_1744.n0 a_20054_1744.t3 14.282
R3830 a_20054_1744.n2 a_20054_1744.t0 8.7
R3831 a_20054_1744.n2 a_20054_1744.t1 8.7
R3832 a_20054_1744.n6 a_20054_1744.n5 4.366
R3833 a_20054_1744.n7 a_20054_1744.n6 0.852
R3834 a_20579_n1475.t2 a_20579_n1475.n0 28.565
R3835 a_20579_n1475.n0 a_20579_n1475.t0 28.565
R3836 a_20579_n1475.n0 a_20579_n1475.n1 185.55
R3837 a_20579_n1475.n1 a_20579_n1475.t1 28.568
R3838 a_20579_n1475.n1 a_20579_n1475.n4 1.638
R3839 a_20579_n1475.n4 a_20579_n1475.t3 21.373
R3840 a_20579_n1475.n4 a_20579_n1475.n2 25.354
R3841 a_20579_n1475.n2 a_20579_n1475.t4 615.911
R3842 a_20579_n1475.n2 a_20579_n1475.t7 867.497
R3843 a_20579_n1475.t7 a_20579_n1475.n3 160.666
R3844 a_20579_n1475.n3 a_20579_n1475.t5 286.438
R3845 a_20579_n1475.n3 a_20579_n1475.t6 286.438
R3846 a_15293_n7386.n1 a_15293_n7386.t5 318.922
R3847 a_15293_n7386.n0 a_15293_n7386.t4 274.739
R3848 a_15293_n7386.n0 a_15293_n7386.t7 274.739
R3849 a_15293_n7386.n1 a_15293_n7386.t6 269.116
R3850 a_15293_n7386.t5 a_15293_n7386.n0 179.946
R3851 a_15293_n7386.n2 a_15293_n7386.n1 107.263
R3852 a_15293_n7386.t2 a_15293_n7386.n4 29.444
R3853 a_15293_n7386.n3 a_15293_n7386.t0 28.565
R3854 a_15293_n7386.n3 a_15293_n7386.t1 28.565
R3855 a_15293_n7386.n2 a_15293_n7386.t3 18.145
R3856 a_15293_n7386.n4 a_15293_n7386.n2 2.878
R3857 a_15293_n7386.n4 a_15293_n7386.n3 0.764
R3858 a_737_n3752.t2 a_737_n3752.n0 28.565
R3859 a_737_n3752.n0 a_737_n3752.t1 28.565
R3860 a_737_n3752.n0 a_737_n3752.n1 197.272
R3861 a_737_n3752.n1 a_737_n3752.t0 28.568
R3862 a_737_n3752.n1 a_737_n3752.n4 0.52
R3863 a_737_n3752.n4 a_737_n3752.t3 18.144
R3864 a_737_n3752.n4 a_737_n3752.n2 50.286
R3865 a_737_n3752.n2 a_737_n3752.t4 408.211
R3866 a_737_n3752.n2 a_737_n3752.t6 990.34
R3867 a_737_n3752.t6 a_737_n3752.n3 160.666
R3868 a_737_n3752.n3 a_737_n3752.t7 286.438
R3869 a_737_n3752.n3 a_737_n3752.t5 286.438
R3870 a_1382_n5059.t0 a_1382_n5059.t1 17.4
R3871 a_897_3260.n0 a_897_3260.t1 28.565
R3872 a_897_3260.t0 a_897_3260.n0 28.565
R3873 a_897_3260.n0 a_897_3260.n1 192.754
R3874 a_897_3260.n1 a_897_3260.t3 28.568
R3875 a_897_3260.n1 a_897_3260.n2 1.312
R3876 a_897_3260.n2 a_897_3260.n3 20.23
R3877 a_897_3260.n3 a_897_3260.t6 615.911
R3878 a_897_3260.n3 a_897_3260.t7 867.497
R3879 a_897_3260.t7 a_897_3260.n4 160.666
R3880 a_897_3260.n4 a_897_3260.t5 286.438
R3881 a_897_3260.n4 a_897_3260.t4 286.438
R3882 a_897_3260.n2 a_897_3260.t2 18.713
R3883 a_1156_1740.n5 a_1156_1740.t9 1527.4
R3884 a_1156_1740.t9 a_1156_1740.n4 657.379
R3885 a_1156_1740.n7 a_1156_1740.n0 258.161
R3886 a_1156_1740.n2 a_1156_1740.n1 258.161
R3887 a_1156_1740.n3 a_1156_1740.t11 206.421
R3888 a_1156_1740.t8 a_1156_1740.n3 206.421
R3889 a_1156_1740.n5 a_1156_1740.t8 200.029
R3890 a_1156_1740.n6 a_1156_1740.n5 97.614
R3891 a_1156_1740.n3 a_1156_1740.t10 80.333
R3892 a_1156_1740.n2 a_1156_1740.t4 14.283
R3893 a_1156_1740.t2 a_1156_1740.n7 14.283
R3894 a_1156_1740.n0 a_1156_1740.t6 14.282
R3895 a_1156_1740.n0 a_1156_1740.t7 14.282
R3896 a_1156_1740.n1 a_1156_1740.t3 14.282
R3897 a_1156_1740.n1 a_1156_1740.t5 14.282
R3898 a_1156_1740.n4 a_1156_1740.t1 8.7
R3899 a_1156_1740.n4 a_1156_1740.t0 8.7
R3900 a_1156_1740.n7 a_1156_1740.n6 4.366
R3901 a_1156_1740.n6 a_1156_1740.n2 0.852
R3902 a_19146_n990.n2 a_19146_n990.t5 448.382
R3903 a_19146_n990.n1 a_19146_n990.t6 286.438
R3904 a_19146_n990.n1 a_19146_n990.t7 286.438
R3905 a_19146_n990.n0 a_19146_n990.t4 247.69
R3906 a_19146_n990.n4 a_19146_n990.n3 182.117
R3907 a_19146_n990.t5 a_19146_n990.n1 160.666
R3908 a_19146_n990.n3 a_19146_n990.t1 28.568
R3909 a_19146_n990.n4 a_19146_n990.t0 28.565
R3910 a_19146_n990.t2 a_19146_n990.n4 28.565
R3911 a_19146_n990.n0 a_19146_n990.t3 18.127
R3912 a_19146_n990.n2 a_19146_n990.n0 4.039
R3913 a_19146_n990.n3 a_19146_n990.n2 0.937
R3914 a_20526_n2323.t0 a_20526_n2323.t1 17.4
R3915 a_20134_3694.t7 a_20134_3694.n3 406.651
R3916 a_20134_3694.n2 a_20134_3694.t6 207.856
R3917 a_20134_3694.n4 a_20134_3694.t7 136.943
R3918 a_20134_3694.n3 a_20134_3694.n2 111.349
R3919 a_20134_3694.n2 a_20134_3694.t8 80.333
R3920 a_20134_3694.n3 a_20134_3694.t5 80.333
R3921 a_20134_3694.n1 a_20134_3694.t4 17.4
R3922 a_20134_3694.n1 a_20134_3694.t0 17.4
R3923 a_20134_3694.t3 a_20134_3694.n5 15.029
R3924 a_20134_3694.n0 a_20134_3694.t1 14.282
R3925 a_20134_3694.n0 a_20134_3694.t2 14.282
R3926 a_20134_3694.n5 a_20134_3694.n0 1.647
R3927 a_20134_3694.n4 a_20134_3694.n1 0.672
R3928 a_20134_3694.n5 a_20134_3694.n4 0.665
R3929 a_9668_n990.n2 a_9668_n990.t4 448.382
R3930 a_9668_n990.n1 a_9668_n990.t6 286.438
R3931 a_9668_n990.n1 a_9668_n990.t7 286.438
R3932 a_9668_n990.n0 a_9668_n990.t5 247.69
R3933 a_9668_n990.n4 a_9668_n990.n3 182.117
R3934 a_9668_n990.t4 a_9668_n990.n1 160.666
R3935 a_9668_n990.n3 a_9668_n990.t1 28.568
R3936 a_9668_n990.n4 a_9668_n990.t0 28.565
R3937 a_9668_n990.t2 a_9668_n990.n4 28.565
R3938 a_9668_n990.n0 a_9668_n990.t3 18.127
R3939 a_9668_n990.n2 a_9668_n990.n0 4.039
R3940 a_9668_n990.n3 a_9668_n990.n2 0.937
R3941 B[2].t12 B[2].t1 799.268
R3942 B[2].n9 B[2].n8 650.893
R3943 B[2].n5 B[2].n4 592.056
R3944 B[2].t2 B[2].t13 415.315
R3945 B[2].t0 B[2].n2 313.873
R3946 B[2].n4 B[2].t9 294.986
R3947 B[2].n7 B[2].t14 285.543
R3948 B[2].n1 B[2].t5 272.288
R3949 B[2].n6 B[2].t2 217.526
R3950 B[2].n0 B[2].t3 214.335
R3951 B[2].t13 B[2].n0 214.335
R3952 B[2].n5 B[2].t10 204.68
R3953 B[2].n8 B[2].t12 194.406
R3954 B[2].n3 B[2].t0 190.152
R3955 B[2].n3 B[2].t11 190.152
R3956 B[2].n1 B[2].t6 160.666
R3957 B[2].n2 B[2].t7 160.666
R3958 B[2].n7 B[2].t4 160.666
R3959 B[2].n4 B[2].t15 110.859
R3960 B[2].n2 B[2].n1 96.129
R3961 B[2].n8 B[2].n7 91.137
R3962 B[2].n0 B[2].t8 80.333
R3963 B[2].t10 B[2].n3 80.333
R3964 B[2].n6 B[2].n5 50.415
R3965 B[2] B[2].n9 9.498
R3966 B[2].n9 B[2].n6 4.527
R3967 a_4951_n7390.n1 a_4951_n7390.t6 318.922
R3968 a_4951_n7390.n0 a_4951_n7390.t4 274.739
R3969 a_4951_n7390.n0 a_4951_n7390.t7 274.739
R3970 a_4951_n7390.n1 a_4951_n7390.t5 269.116
R3971 a_4951_n7390.t6 a_4951_n7390.n0 179.946
R3972 a_4951_n7390.n2 a_4951_n7390.n1 107.263
R3973 a_4951_n7390.n3 a_4951_n7390.t0 29.444
R3974 a_4951_n7390.n4 a_4951_n7390.t1 28.565
R3975 a_4951_n7390.t2 a_4951_n7390.n4 28.565
R3976 a_4951_n7390.n2 a_4951_n7390.t3 18.145
R3977 a_4951_n7390.n3 a_4951_n7390.n2 2.878
R3978 a_4951_n7390.n4 a_4951_n7390.n3 0.764
R3979 a_4300_n994.n2 a_4300_n994.t8 1527.4
R3980 a_4300_n994.t8 a_4300_n994.n1 657.379
R3981 a_4300_n994.n4 a_4300_n994.n3 258.161
R3982 a_4300_n994.n7 a_4300_n994.n6 258.161
R3983 a_4300_n994.n0 a_4300_n994.t9 206.421
R3984 a_4300_n994.t10 a_4300_n994.n0 206.421
R3985 a_4300_n994.n2 a_4300_n994.t10 200.029
R3986 a_4300_n994.n5 a_4300_n994.n2 97.614
R3987 a_4300_n994.n0 a_4300_n994.t11 80.333
R3988 a_4300_n994.n4 a_4300_n994.t3 14.283
R3989 a_4300_n994.n6 a_4300_n994.t6 14.283
R3990 a_4300_n994.n3 a_4300_n994.t2 14.282
R3991 a_4300_n994.n3 a_4300_n994.t1 14.282
R3992 a_4300_n994.n7 a_4300_n994.t7 14.282
R3993 a_4300_n994.t4 a_4300_n994.n7 14.282
R3994 a_4300_n994.n1 a_4300_n994.t0 8.7
R3995 a_4300_n994.n1 a_4300_n994.t5 8.7
R3996 a_4300_n994.n5 a_4300_n994.n4 4.366
R3997 a_4300_n994.n6 a_4300_n994.n5 0.852
R3998 a_22839_n3722.n3 a_22839_n3722.n2 167.433
R3999 a_22839_n3722.n7 a_22839_n3722.n6 167.433
R4000 a_22839_n3722.n3 a_22839_n3722.t10 104.259
R4001 a_22839_n3722.n7 a_22839_n3722.t7 104.259
R4002 a_22839_n3722.n4 a_22839_n3722.n1 89.977
R4003 a_22839_n3722.n5 a_22839_n3722.n0 89.977
R4004 a_22839_n3722.n9 a_22839_n3722.n8 89.977
R4005 a_22839_n3722.n4 a_22839_n3722.n3 77.784
R4006 a_22839_n3722.n5 a_22839_n3722.n4 77.456
R4007 a_22839_n3722.n8 a_22839_n3722.n5 77.456
R4008 a_22839_n3722.n8 a_22839_n3722.n7 75.815
R4009 a_22839_n3722.n2 a_22839_n3722.t9 14.282
R4010 a_22839_n3722.n2 a_22839_n3722.t11 14.282
R4011 a_22839_n3722.n1 a_22839_n3722.t2 14.282
R4012 a_22839_n3722.n1 a_22839_n3722.t3 14.282
R4013 a_22839_n3722.n0 a_22839_n3722.t4 14.282
R4014 a_22839_n3722.n0 a_22839_n3722.t1 14.282
R4015 a_22839_n3722.n6 a_22839_n3722.t5 14.282
R4016 a_22839_n3722.n6 a_22839_n3722.t6 14.282
R4017 a_22839_n3722.t0 a_22839_n3722.n9 14.282
R4018 a_22839_n3722.n9 a_22839_n3722.t8 14.282
R4019 a_9668_1744.n2 a_9668_1744.t4 448.382
R4020 a_9668_1744.n1 a_9668_1744.t6 286.438
R4021 a_9668_1744.n1 a_9668_1744.t7 286.438
R4022 a_9668_1744.n0 a_9668_1744.t5 247.69
R4023 a_9668_1744.n4 a_9668_1744.n3 182.117
R4024 a_9668_1744.t4 a_9668_1744.n1 160.666
R4025 a_9668_1744.n3 a_9668_1744.t1 28.568
R4026 a_9668_1744.n4 a_9668_1744.t0 28.565
R4027 a_9668_1744.t2 a_9668_1744.n4 28.565
R4028 a_9668_1744.n0 a_9668_1744.t3 18.127
R4029 a_9668_1744.n2 a_9668_1744.n0 4.039
R4030 a_9668_1744.n3 a_9668_1744.n2 0.937
R4031 a_1681_n1479.t2 a_1681_n1479.n0 28.568
R4032 a_1681_n1479.n0 a_1681_n1479.n4 185.55
R4033 a_1681_n1479.n4 a_1681_n1479.t0 28.565
R4034 a_1681_n1479.n4 a_1681_n1479.t1 28.565
R4035 a_1681_n1479.n0 a_1681_n1479.n3 1.637
R4036 a_1681_n1479.n3 a_1681_n1479.t3 21.373
R4037 a_1681_n1479.n3 a_1681_n1479.n1 26.067
R4038 a_1681_n1479.n1 a_1681_n1479.t7 615.911
R4039 a_1681_n1479.n1 a_1681_n1479.t6 867.497
R4040 a_1681_n1479.t6 a_1681_n1479.n2 160.666
R4041 a_1681_n1479.n2 a_1681_n1479.t5 286.438
R4042 a_1681_n1479.n2 a_1681_n1479.t4 286.438
R4043 a_1156_n994.n4 a_1156_n994.t8 1527.4
R4044 a_1156_n994.t8 a_1156_n994.n3 657.379
R4045 a_1156_n994.n1 a_1156_n994.n0 258.161
R4046 a_1156_n994.n7 a_1156_n994.n6 258.161
R4047 a_1156_n994.n2 a_1156_n994.t11 206.421
R4048 a_1156_n994.t9 a_1156_n994.n2 206.421
R4049 a_1156_n994.n4 a_1156_n994.t9 200.029
R4050 a_1156_n994.n5 a_1156_n994.n4 97.614
R4051 a_1156_n994.n2 a_1156_n994.t10 80.333
R4052 a_1156_n994.n6 a_1156_n994.t7 14.283
R4053 a_1156_n994.n1 a_1156_n994.t4 14.283
R4054 a_1156_n994.n0 a_1156_n994.t3 14.282
R4055 a_1156_n994.n0 a_1156_n994.t5 14.282
R4056 a_1156_n994.t1 a_1156_n994.n7 14.282
R4057 a_1156_n994.n7 a_1156_n994.t2 14.282
R4058 a_1156_n994.n3 a_1156_n994.t6 8.7
R4059 a_1156_n994.n3 a_1156_n994.t0 8.7
R4060 a_1156_n994.n6 a_1156_n994.n5 4.366
R4061 a_1156_n994.n5 a_1156_n994.n1 0.852
R4062 a_2824_n8094.t0 a_2824_n8094.t1 17.4
R4063 B[4].t15 B[4].t6 802.481
R4064 B[4].n9 B[4].n8 650.497
R4065 B[4].n4 B[4].n3 592.056
R4066 B[4].t12 B[4].t8 415.315
R4067 B[4].t7 B[4].n1 313.873
R4068 B[4].n3 B[4].t14 294.986
R4069 B[4].n7 B[4].t0 284.688
R4070 B[4].n0 B[4].t2 272.288
R4071 B[4].n6 B[4].t12 217.534
R4072 B[4].n5 B[4].t13 214.335
R4073 B[4].t8 B[4].n5 214.335
R4074 B[4].n4 B[4].t9 204.68
R4075 B[4].n8 B[4].t15 192.799
R4076 B[4].n2 B[4].t7 190.152
R4077 B[4].n2 B[4].t10 190.152
R4078 B[4].n7 B[4].t11 160.666
R4079 B[4].n0 B[4].t3 160.666
R4080 B[4].n1 B[4].t4 160.666
R4081 B[4].n3 B[4].t5 110.859
R4082 B[4].n1 B[4].n0 96.129
R4083 B[4].n8 B[4].n7 91.889
R4084 B[4].n5 B[4].t1 80.333
R4085 B[4].t9 B[4].n2 80.333
R4086 B[4].n6 B[4].n4 50.196
R4087 B[4] B[4].n9 15.176
R4088 B[4].n9 B[4].n6 5.535
R4089 a_16748_3696.n0 a_16748_3696.t1 14.282
R4090 a_16748_3696.n0 a_16748_3696.t5 14.282
R4091 a_16748_3696.n1 a_16748_3696.t3 14.282
R4092 a_16748_3696.n1 a_16748_3696.t2 14.282
R4093 a_16748_3696.t0 a_16748_3696.n3 14.282
R4094 a_16748_3696.n3 a_16748_3696.t4 14.282
R4095 a_16748_3696.n3 a_16748_3696.n2 2.538
R4096 a_16748_3696.n2 a_16748_3696.n1 2.375
R4097 a_16748_3696.n2 a_16748_3696.n0 0.001
R4098 a_14303_n1479.n0 a_14303_n1479.t1 28.565
R4099 a_14303_n1479.t0 a_14303_n1479.n0 28.565
R4100 a_14303_n1479.n0 a_14303_n1479.n1 185.55
R4101 a_14303_n1479.n1 a_14303_n1479.t3 28.568
R4102 a_14303_n1479.n1 a_14303_n1479.n4 1.637
R4103 a_14303_n1479.n4 a_14303_n1479.t2 21.373
R4104 a_14303_n1479.n4 a_14303_n1479.n2 25.444
R4105 a_14303_n1479.n2 a_14303_n1479.t4 615.911
R4106 a_14303_n1479.n2 a_14303_n1479.t7 867.497
R4107 a_14303_n1479.t7 a_14303_n1479.n3 160.666
R4108 a_14303_n1479.n3 a_14303_n1479.t6 286.438
R4109 a_14303_n1479.n3 a_14303_n1479.t5 286.438
R4110 a_14250_n2327.t0 a_14250_n2327.t1 17.4
R4111 a_16630_3696.t5 a_16630_3696.n2 403.87
R4112 a_16630_3696.n1 a_16630_3696.t6 191.682
R4113 a_16630_3696.n3 a_16630_3696.t5 138.55
R4114 a_16630_3696.n2 a_16630_3696.n1 111.349
R4115 a_16630_3696.n1 a_16630_3696.t7 80.333
R4116 a_16630_3696.n2 a_16630_3696.t8 80.333
R4117 a_16630_3696.n0 a_16630_3696.t2 17.4
R4118 a_16630_3696.n0 a_16630_3696.t1 17.4
R4119 a_16630_3696.n4 a_16630_3696.t3 15.036
R4120 a_16630_3696.n5 a_16630_3696.t4 14.282
R4121 a_16630_3696.t0 a_16630_3696.n5 14.282
R4122 a_16630_3696.n5 a_16630_3696.n4 1.654
R4123 a_16630_3696.n3 a_16630_3696.n0 0.679
R4124 a_16630_3696.n4 a_16630_3696.n3 0.665
R4125 a_13369_1714.n0 a_13369_1714.t1 28.565
R4126 a_13369_1714.t2 a_13369_1714.n0 28.565
R4127 a_13369_1714.n0 a_13369_1714.n2 97.476
R4128 a_13369_1714.n2 a_13369_1714.n3 940.604
R4129 a_13369_1714.n3 a_13369_1714.t7 408.211
R4130 a_13369_1714.n3 a_13369_1714.t4 990.34
R4131 a_13369_1714.t4 a_13369_1714.n4 160.666
R4132 a_13369_1714.n4 a_13369_1714.t6 286.438
R4133 a_13369_1714.n4 a_13369_1714.t5 286.438
R4134 a_13369_1714.n2 a_13369_1714.n1 109.176
R4135 a_13369_1714.n1 a_13369_1714.t0 28.568
R4136 a_13369_1714.n1 a_13369_1714.t3 17.638
R4137 a_1146_n3726.n2 a_1146_n3726.t11 1527.4
R4138 a_1146_n3726.t11 a_1146_n3726.n1 657.379
R4139 a_1146_n3726.n4 a_1146_n3726.n3 258.161
R4140 a_1146_n3726.n7 a_1146_n3726.n6 258.161
R4141 a_1146_n3726.n0 a_1146_n3726.t8 206.421
R4142 a_1146_n3726.t10 a_1146_n3726.n0 206.421
R4143 a_1146_n3726.n2 a_1146_n3726.t10 200.029
R4144 a_1146_n3726.n5 a_1146_n3726.n2 97.614
R4145 a_1146_n3726.n0 a_1146_n3726.t9 80.333
R4146 a_1146_n3726.n4 a_1146_n3726.t7 14.283
R4147 a_1146_n3726.n6 a_1146_n3726.t5 14.283
R4148 a_1146_n3726.n3 a_1146_n3726.t3 14.282
R4149 a_1146_n3726.n3 a_1146_n3726.t2 14.282
R4150 a_1146_n3726.n7 a_1146_n3726.t4 14.282
R4151 a_1146_n3726.t0 a_1146_n3726.n7 14.282
R4152 a_1146_n3726.n1 a_1146_n3726.t6 8.7
R4153 a_1146_n3726.n1 a_1146_n3726.t1 8.7
R4154 a_1146_n3726.n5 a_1146_n3726.n4 4.366
R4155 a_1146_n3726.n6 a_1146_n3726.n5 0.852
R4156 a_10227_n990.n9 a_10227_n990.n0 167.433
R4157 a_10227_n990.n5 a_10227_n990.n4 167.433
R4158 a_10227_n990.n5 a_10227_n990.t4 104.259
R4159 a_10227_n990.t9 a_10227_n990.n9 104.259
R4160 a_10227_n990.n8 a_10227_n990.n1 89.977
R4161 a_10227_n990.n7 a_10227_n990.n2 89.977
R4162 a_10227_n990.n6 a_10227_n990.n3 89.977
R4163 a_10227_n990.n9 a_10227_n990.n8 77.784
R4164 a_10227_n990.n8 a_10227_n990.n7 77.456
R4165 a_10227_n990.n7 a_10227_n990.n6 77.456
R4166 a_10227_n990.n6 a_10227_n990.n5 75.815
R4167 a_10227_n990.n0 a_10227_n990.t10 14.282
R4168 a_10227_n990.n0 a_10227_n990.t11 14.282
R4169 a_10227_n990.n1 a_10227_n990.t0 14.282
R4170 a_10227_n990.n1 a_10227_n990.t2 14.282
R4171 a_10227_n990.n2 a_10227_n990.t1 14.282
R4172 a_10227_n990.n2 a_10227_n990.t6 14.282
R4173 a_10227_n990.n3 a_10227_n990.t8 14.282
R4174 a_10227_n990.n3 a_10227_n990.t7 14.282
R4175 a_10227_n990.n4 a_10227_n990.t3 14.282
R4176 a_10227_n990.n4 a_10227_n990.t5 14.282
R4177 a_10227_1744.n3 a_10227_1744.n2 167.433
R4178 a_10227_1744.n7 a_10227_1744.n6 167.433
R4179 a_10227_1744.n3 a_10227_1744.t9 104.259
R4180 a_10227_1744.n7 a_10227_1744.t6 104.259
R4181 a_10227_1744.n4 a_10227_1744.n1 89.977
R4182 a_10227_1744.n5 a_10227_1744.n0 89.977
R4183 a_10227_1744.n9 a_10227_1744.n8 89.977
R4184 a_10227_1744.n4 a_10227_1744.n3 77.784
R4185 a_10227_1744.n5 a_10227_1744.n4 77.456
R4186 a_10227_1744.n8 a_10227_1744.n5 77.456
R4187 a_10227_1744.n8 a_10227_1744.n7 75.815
R4188 a_10227_1744.n2 a_10227_1744.t10 14.282
R4189 a_10227_1744.n2 a_10227_1744.t11 14.282
R4190 a_10227_1744.n1 a_10227_1744.t3 14.282
R4191 a_10227_1744.n1 a_10227_1744.t5 14.282
R4192 a_10227_1744.n0 a_10227_1744.t4 14.282
R4193 a_10227_1744.n0 a_10227_1744.t1 14.282
R4194 a_10227_1744.n6 a_10227_1744.t7 14.282
R4195 a_10227_1744.n6 a_10227_1744.t8 14.282
R4196 a_10227_1744.t0 a_10227_1744.n9 14.282
R4197 a_10227_1744.n9 a_10227_1744.t2 14.282
R4198 Y[1].n1 Y[1].n0 185.55
R4199 Y[1] Y[1].n2 29.697
R4200 Y[1].n1 Y[1].t1 28.568
R4201 Y[1].n0 Y[1].t0 28.565
R4202 Y[1].n0 Y[1].t2 28.565
R4203 Y[1].n2 Y[1].t3 21.879
R4204 Y[1].n2 Y[1].n1 1.625
R4205 B[3].t6 B[3].t1 800.875
R4206 B[3].n9 B[3].n8 650.874
R4207 B[3].n5 B[3].n4 592.056
R4208 B[3].t2 B[3].t15 415.315
R4209 B[3].t9 B[3].n2 313.873
R4210 B[3].n4 B[3].t3 294.986
R4211 B[3].n7 B[3].t14 284.688
R4212 B[3].n1 B[3].t5 272.288
R4213 B[3].n6 B[3].t2 217.532
R4214 B[3].n0 B[3].t4 214.335
R4215 B[3].t15 B[3].n0 214.335
R4216 B[3].n5 B[3].t10 204.68
R4217 B[3].n8 B[3].t6 192.799
R4218 B[3].n3 B[3].t9 190.152
R4219 B[3].n3 B[3].t11 190.152
R4220 B[3].n1 B[3].t7 160.666
R4221 B[3].n2 B[3].t13 160.666
R4222 B[3].n7 B[3].t0 160.666
R4223 B[3].n4 B[3].t8 110.859
R4224 B[3].n2 B[3].n1 96.129
R4225 B[3].n8 B[3].n7 91.889
R4226 B[3].n0 B[3].t12 80.333
R4227 B[3].t10 B[3].n3 80.333
R4228 B[3].n6 B[3].n5 50.557
R4229 B[3] B[3].n9 13.739
R4230 B[3].n9 B[3].n6 4.969
R4231 a_15574_3694.n0 a_15574_3694.t3 14.282
R4232 a_15574_3694.n0 a_15574_3694.t1 14.282
R4233 a_15574_3694.n1 a_15574_3694.t2 14.282
R4234 a_15574_3694.n1 a_15574_3694.t4 14.282
R4235 a_15574_3694.n3 a_15574_3694.t5 14.282
R4236 a_15574_3694.t0 a_15574_3694.n3 14.282
R4237 a_15574_3694.n3 a_15574_3694.n2 2.538
R4238 a_15574_3694.n2 a_15574_3694.n1 2.375
R4239 a_15574_3694.n2 a_15574_3694.n0 0.001
R4240 a_7432_n990.n2 a_7432_n990.t10 1527.4
R4241 a_7432_n990.t10 a_7432_n990.n1 657.379
R4242 a_7432_n990.n4 a_7432_n990.n3 258.161
R4243 a_7432_n990.n7 a_7432_n990.n6 258.161
R4244 a_7432_n990.n0 a_7432_n990.t11 206.421
R4245 a_7432_n990.t9 a_7432_n990.n0 206.421
R4246 a_7432_n990.n2 a_7432_n990.t9 200.029
R4247 a_7432_n990.n5 a_7432_n990.n2 97.614
R4248 a_7432_n990.n0 a_7432_n990.t8 80.333
R4249 a_7432_n990.n4 a_7432_n990.t3 14.283
R4250 a_7432_n990.n6 a_7432_n990.t2 14.283
R4251 a_7432_n990.n3 a_7432_n990.t7 14.282
R4252 a_7432_n990.n3 a_7432_n990.t4 14.282
R4253 a_7432_n990.n7 a_7432_n990.t5 14.282
R4254 a_7432_n990.t1 a_7432_n990.n7 14.282
R4255 a_7432_n990.n1 a_7432_n990.t6 8.7
R4256 a_7432_n990.n1 a_7432_n990.t0 8.7
R4257 a_7432_n990.n5 a_7432_n990.n4 4.366
R4258 a_7432_n990.n6 a_7432_n990.n5 0.852
R4259 Y[2].n1 Y[2].n0 185.55
R4260 Y[2].n1 Y[2].t1 28.568
R4261 Y[2].n0 Y[2].t2 28.565
R4262 Y[2].n0 Y[2].t0 28.565
R4263 Y[2] Y[2].n2 24.297
R4264 Y[2].n2 Y[2].t3 21.373
R4265 Y[2].n2 Y[2].n1 1.637
R4266 a_13120_3694.t8 a_13120_3694.n2 404.877
R4267 a_13120_3694.n1 a_13120_3694.t5 210.902
R4268 a_13120_3694.n3 a_13120_3694.t8 136.943
R4269 a_13120_3694.n2 a_13120_3694.n1 107.801
R4270 a_13120_3694.n1 a_13120_3694.t6 80.333
R4271 a_13120_3694.n2 a_13120_3694.t7 80.333
R4272 a_13120_3694.n0 a_13120_3694.t4 17.4
R4273 a_13120_3694.n0 a_13120_3694.t2 17.4
R4274 a_13120_3694.n4 a_13120_3694.t3 15.036
R4275 a_13120_3694.t0 a_13120_3694.n5 14.282
R4276 a_13120_3694.n5 a_13120_3694.t1 14.282
R4277 a_13120_3694.n5 a_13120_3694.n4 1.654
R4278 a_13120_3694.n3 a_13120_3694.n0 0.672
R4279 a_13120_3694.n4 a_13120_3694.n3 0.665
R4280 a_13238_3694.n1 a_13238_3694.t5 14.282
R4281 a_13238_3694.n1 a_13238_3694.t2 14.282
R4282 a_13238_3694.n0 a_13238_3694.t1 14.282
R4283 a_13238_3694.n0 a_13238_3694.t0 14.282
R4284 a_13238_3694.n3 a_13238_3694.t4 14.282
R4285 a_13238_3694.t3 a_13238_3694.n3 14.282
R4286 a_13238_3694.n2 a_13238_3694.n0 2.538
R4287 a_13238_3694.n3 a_13238_3694.n2 2.375
R4288 a_13238_3694.n2 a_13238_3694.n1 0.001
R4289 a_7432_1744.n4 a_7432_1744.t10 1527.4
R4290 a_7432_1744.t10 a_7432_1744.n3 657.379
R4291 a_7432_1744.n1 a_7432_1744.n0 258.161
R4292 a_7432_1744.n7 a_7432_1744.n6 258.161
R4293 a_7432_1744.n2 a_7432_1744.t11 206.421
R4294 a_7432_1744.t9 a_7432_1744.n2 206.421
R4295 a_7432_1744.n4 a_7432_1744.t9 200.029
R4296 a_7432_1744.n5 a_7432_1744.n4 97.614
R4297 a_7432_1744.n2 a_7432_1744.t8 80.333
R4298 a_7432_1744.n6 a_7432_1744.t7 14.283
R4299 a_7432_1744.n1 a_7432_1744.t5 14.283
R4300 a_7432_1744.n0 a_7432_1744.t2 14.282
R4301 a_7432_1744.n0 a_7432_1744.t4 14.282
R4302 a_7432_1744.t1 a_7432_1744.n7 14.282
R4303 a_7432_1744.n7 a_7432_1744.t3 14.282
R4304 a_7432_1744.n3 a_7432_1744.t6 8.7
R4305 a_7432_1744.n3 a_7432_1744.t0 8.7
R4306 a_7432_1744.n6 a_7432_1744.n5 4.366
R4307 a_7432_1744.n5 a_7432_1744.n1 0.852
R4308 a_7957_n1475.n0 a_7957_n1475.t0 28.565
R4309 a_7957_n1475.t2 a_7957_n1475.n0 28.565
R4310 a_7957_n1475.n0 a_7957_n1475.n1 185.55
R4311 a_7957_n1475.n1 a_7957_n1475.t1 28.568
R4312 a_7957_n1475.n1 a_7957_n1475.n4 1.638
R4313 a_7957_n1475.n4 a_7957_n1475.t3 21.373
R4314 a_7957_n1475.n4 a_7957_n1475.n2 26.1
R4315 a_7957_n1475.n2 a_7957_n1475.t5 615.911
R4316 a_7957_n1475.n2 a_7957_n1475.t4 867.497
R4317 a_7957_n1475.t4 a_7957_n1475.n3 160.666
R4318 a_7957_n1475.n3 a_7957_n1475.t7 286.438
R4319 a_7957_n1475.n3 a_7957_n1475.t6 286.438
R4320 B[1].t10 B[1].t2 800.875
R4321 B[1].n9 B[1].n1 654.791
R4322 B[1].n7 B[1].n6 592.056
R4323 B[1].t8 B[1].t1 415.315
R4324 B[1].t5 B[1].n4 313.873
R4325 B[1].n6 B[1].t0 294.986
R4326 B[1].n0 B[1].t15 284.688
R4327 B[1].n3 B[1].t12 272.288
R4328 B[1].n8 B[1].t8 217.528
R4329 B[1].n2 B[1].t4 214.335
R4330 B[1].t1 B[1].n2 214.335
R4331 B[1].n7 B[1].t6 204.68
R4332 B[1].n1 B[1].t10 192.799
R4333 B[1].n5 B[1].t5 190.152
R4334 B[1].n5 B[1].t14 190.152
R4335 B[1].n3 B[1].t7 160.666
R4336 B[1].n4 B[1].t9 160.666
R4337 B[1].n0 B[1].t3 160.666
R4338 B[1].n6 B[1].t13 110.859
R4339 B[1].n4 B[1].n3 96.129
R4340 B[1].n1 B[1].n0 91.889
R4341 B[1].n2 B[1].t11 80.333
R4342 B[1].t6 B[1].n5 80.333
R4343 B[1].n8 B[1].n7 49.906
R4344 B[1] B[1].n9 8.858
R4345 B[1].n9 B[1].n8 0.369
R4346 a_1755_3697.n0 a_1755_3697.t10 214.335
R4347 a_1755_3697.t9 a_1755_3697.n0 214.335
R4348 a_1755_3697.n1 a_1755_3697.t9 143.851
R4349 a_1755_3697.n1 a_1755_3697.t7 135.658
R4350 a_1755_3697.n0 a_1755_3697.t8 80.333
R4351 a_1755_3697.n2 a_1755_3697.t5 28.565
R4352 a_1755_3697.n2 a_1755_3697.t4 28.565
R4353 a_1755_3697.n4 a_1755_3697.t6 28.565
R4354 a_1755_3697.n4 a_1755_3697.t2 28.565
R4355 a_1755_3697.n7 a_1755_3697.t1 28.565
R4356 a_1755_3697.t3 a_1755_3697.n7 28.565
R4357 a_1755_3697.n6 a_1755_3697.t0 9.714
R4358 a_1755_3697.n7 a_1755_3697.n6 1.003
R4359 a_1755_3697.n5 a_1755_3697.n3 0.833
R4360 a_1755_3697.n3 a_1755_3697.n2 0.653
R4361 a_1755_3697.n5 a_1755_3697.n4 0.653
R4362 a_1755_3697.n6 a_1755_3697.n5 0.341
R4363 a_1755_3697.n3 a_1755_3697.n1 0.032
R4364 a_16513_n1020.t0 a_16513_n1020.n0 28.568
R4365 a_16513_n1020.n0 a_16513_n1020.n4 185.55
R4366 a_16513_n1020.n4 a_16513_n1020.t1 28.565
R4367 a_16513_n1020.n4 a_16513_n1020.t3 28.565
R4368 a_16513_n1020.n0 a_16513_n1020.n3 1.537
R4369 a_16513_n1020.n3 a_16513_n1020.t2 21.473
R4370 a_16513_n1020.n3 a_16513_n1020.n1 12.48
R4371 a_16513_n1020.n1 a_16513_n1020.t4 408.211
R4372 a_16513_n1020.n1 a_16513_n1020.t5 990.34
R4373 a_16513_n1020.t5 a_16513_n1020.n2 160.666
R4374 a_16513_n1020.n2 a_16513_n1020.t7 286.438
R4375 a_16513_n1020.n2 a_16513_n1020.t6 286.438
R4376 a_17158_n2327.t0 a_17158_n2327.t1 17.4
R4377 a_23723_n1475.n0 a_23723_n1475.t2 28.565
R4378 a_23723_n1475.t1 a_23723_n1475.n0 28.565
R4379 a_23723_n1475.n0 a_23723_n1475.n1 185.55
R4380 a_23723_n1475.n1 a_23723_n1475.t3 28.568
R4381 a_23723_n1475.n1 a_23723_n1475.n4 1.637
R4382 a_23723_n1475.n4 a_23723_n1475.t0 21.373
R4383 a_23723_n1475.n4 a_23723_n1475.n2 25.539
R4384 a_23723_n1475.n2 a_23723_n1475.t4 615.911
R4385 a_23723_n1475.n2 a_23723_n1475.t7 867.497
R4386 a_23723_n1475.t7 a_23723_n1475.n3 160.666
R4387 a_23723_n1475.n3 a_23723_n1475.t5 286.438
R4388 a_23723_n1475.n3 a_23723_n1475.t6 286.438
R4389 a_23670_n2323.t0 a_23670_n2323.t1 17.4
R4390 A[4].n8 A[4].n7 2886.86
R4391 A[4].t15 A[4].t18 576.841
R4392 A[4].t5 A[4].t19 437.233
R4393 A[4].n5 A[4].n4 412.11
R4394 A[4].n1 A[4].t14 394.151
R4395 A[4].n4 A[4].t13 294.653
R4396 A[4].n9 A[4].t17 284.688
R4397 A[4].n0 A[4].t1 269.523
R4398 A[4].t14 A[4].n0 269.523
R4399 A[4].n5 A[4].n3 224.13
R4400 A[4].n12 A[4].t5 221.772
R4401 A[4].n11 A[4].t16 214.686
R4402 A[4].t19 A[4].n11 214.686
R4403 A[4].n2 A[4].t9 198.043
R4404 A[4].n6 A[4].t12 185.301
R4405 A[4].n6 A[4].t6 185.301
R4406 A[4].n12 A[4].n10 182.459
R4407 A[4].n9 A[4].t3 160.666
R4408 A[4].n10 A[4].t15 160.666
R4409 A[4].n0 A[4].t7 160.666
R4410 A[4].n8 A[4].n5 141.986
R4411 A[4].n7 A[4].t2 140.583
R4412 A[4].n10 A[4].n9 115.593
R4413 A[4].n4 A[4].t0 111.663
R4414 A[4].n6 A[4].t8 107.646
R4415 A[4].n3 A[4].n1 97.816
R4416 A[4].n2 A[4].t10 93.989
R4417 A[4].n11 A[4].t4 80.333
R4418 A[4].n1 A[4].t11 80.333
R4419 A[4].n7 A[4].n6 61.856
R4420 A[4].n13 A[4].n12 33.949
R4421 A[4].n13 A[4].n8 19.007
R4422 A[4].n3 A[4].n2 6.615
R4423 A[4] A[4].n13 1.898
R4424 a_8249_n6669.n2 a_8249_n6669.t6 318.922
R4425 a_8249_n6669.n1 a_8249_n6669.t5 273.935
R4426 a_8249_n6669.n1 a_8249_n6669.t7 273.935
R4427 a_8249_n6669.n2 a_8249_n6669.t4 269.116
R4428 a_8249_n6669.n4 a_8249_n6669.n0 193.227
R4429 a_8249_n6669.t6 a_8249_n6669.n1 179.142
R4430 a_8249_n6669.n3 a_8249_n6669.n2 106.999
R4431 a_8249_n6669.t2 a_8249_n6669.n4 28.568
R4432 a_8249_n6669.n0 a_8249_n6669.t0 28.565
R4433 a_8249_n6669.n0 a_8249_n6669.t1 28.565
R4434 a_8249_n6669.n3 a_8249_n6669.t3 18.149
R4435 a_8249_n6669.n4 a_8249_n6669.n3 3.726
R4436 a_6221_3697.n4 a_6221_3697.t8 214.335
R4437 a_6221_3697.t7 a_6221_3697.n4 214.335
R4438 a_6221_3697.n5 a_6221_3697.t7 143.851
R4439 a_6221_3697.n5 a_6221_3697.t9 135.658
R4440 a_6221_3697.n4 a_6221_3697.t10 80.333
R4441 a_6221_3697.n0 a_6221_3697.t5 28.565
R4442 a_6221_3697.n0 a_6221_3697.t4 28.565
R4443 a_6221_3697.n2 a_6221_3697.t1 28.565
R4444 a_6221_3697.n2 a_6221_3697.t3 28.565
R4445 a_6221_3697.n7 a_6221_3697.t0 28.565
R4446 a_6221_3697.t2 a_6221_3697.n7 28.565
R4447 a_6221_3697.n1 a_6221_3697.t6 9.714
R4448 a_6221_3697.n1 a_6221_3697.n0 1.003
R4449 a_6221_3697.n6 a_6221_3697.n3 0.833
R4450 a_6221_3697.n3 a_6221_3697.n2 0.653
R4451 a_6221_3697.n7 a_6221_3697.n6 0.653
R4452 a_6221_3697.n3 a_6221_3697.n1 0.341
R4453 a_6221_3697.n6 a_6221_3697.n5 0.032
R4454 a_4701_3699.n0 a_4701_3699.t7 214.335
R4455 a_4701_3699.t10 a_4701_3699.n0 214.335
R4456 a_4701_3699.n1 a_4701_3699.t10 143.851
R4457 a_4701_3699.n1 a_4701_3699.t8 135.658
R4458 a_4701_3699.n0 a_4701_3699.t9 80.333
R4459 a_4701_3699.n2 a_4701_3699.t4 28.565
R4460 a_4701_3699.n2 a_4701_3699.t3 28.565
R4461 a_4701_3699.n4 a_4701_3699.t2 28.565
R4462 a_4701_3699.n4 a_4701_3699.t5 28.565
R4463 a_4701_3699.t0 a_4701_3699.n7 28.565
R4464 a_4701_3699.n7 a_4701_3699.t6 28.565
R4465 a_4701_3699.n6 a_4701_3699.t1 9.714
R4466 a_4701_3699.n7 a_4701_3699.n6 1.003
R4467 a_4701_3699.n5 a_4701_3699.n3 0.833
R4468 a_4701_3699.n3 a_4701_3699.n2 0.653
R4469 a_4701_3699.n5 a_4701_3699.n4 0.653
R4470 a_4701_3699.n6 a_4701_3699.n5 0.341
R4471 a_4701_3699.n3 a_4701_3699.n1 0.032
R4472 a_5291_3262.t2 a_5291_3262.n0 28.568
R4473 a_5291_3262.n0 a_5291_3262.n4 192.754
R4474 a_5291_3262.n4 a_5291_3262.t0 28.565
R4475 a_5291_3262.n4 a_5291_3262.t1 28.565
R4476 a_5291_3262.n0 a_5291_3262.n1 1.123
R4477 a_5291_3262.n1 a_5291_3262.n2 25.17
R4478 a_5291_3262.n2 a_5291_3262.t4 615.911
R4479 a_5291_3262.n2 a_5291_3262.t5 867.497
R4480 a_5291_3262.t5 a_5291_3262.n3 160.666
R4481 a_5291_3262.n3 a_5291_3262.t7 286.438
R4482 a_5291_3262.n3 a_5291_3262.t6 286.438
R4483 a_5291_3262.n1 a_5291_3262.t3 18.726
R4484 a_2470_n7362.n2 a_2470_n7362.n0 267.767
R4485 a_2470_n7362.n6 a_2470_n7362.t2 16.058
R4486 a_2470_n7362.n8 a_2470_n7362.t11 16.058
R4487 a_2470_n7362.n1 a_2470_n7362.t8 14.282
R4488 a_2470_n7362.n1 a_2470_n7362.t4 14.282
R4489 a_2470_n7362.n0 a_2470_n7362.t9 14.282
R4490 a_2470_n7362.n0 a_2470_n7362.t10 14.282
R4491 a_2470_n7362.n3 a_2470_n7362.t5 14.282
R4492 a_2470_n7362.n3 a_2470_n7362.t6 14.282
R4493 a_2470_n7362.n5 a_2470_n7362.t0 14.282
R4494 a_2470_n7362.n5 a_2470_n7362.t1 14.282
R4495 a_2470_n7362.t3 a_2470_n7362.n9 14.282
R4496 a_2470_n7362.n9 a_2470_n7362.t7 14.282
R4497 a_2470_n7362.n4 a_2470_n7362.n3 1.511
R4498 a_2470_n7362.n6 a_2470_n7362.n5 0.999
R4499 a_2470_n7362.n9 a_2470_n7362.n8 0.999
R4500 a_2470_n7362.n4 a_2470_n7362.n2 0.669
R4501 a_2470_n7362.n7 a_2470_n7362.n6 0.575
R4502 a_2470_n7362.n7 a_2470_n7362.n4 0.227
R4503 a_2470_n7362.n8 a_2470_n7362.n7 0.2
R4504 a_2470_n7362.n2 a_2470_n7362.n1 0.001
R4505 a_9167_3699.n4 a_9167_3699.t8 214.335
R4506 a_9167_3699.t7 a_9167_3699.n4 214.335
R4507 a_9167_3699.n5 a_9167_3699.t7 143.851
R4508 a_9167_3699.n5 a_9167_3699.t9 135.658
R4509 a_9167_3699.n4 a_9167_3699.t10 80.333
R4510 a_9167_3699.n0 a_9167_3699.t1 28.565
R4511 a_9167_3699.n0 a_9167_3699.t4 28.565
R4512 a_9167_3699.n2 a_9167_3699.t6 28.565
R4513 a_9167_3699.n2 a_9167_3699.t3 28.565
R4514 a_9167_3699.t0 a_9167_3699.n7 28.565
R4515 a_9167_3699.n7 a_9167_3699.t5 28.565
R4516 a_9167_3699.n1 a_9167_3699.t2 9.714
R4517 a_9167_3699.n1 a_9167_3699.n0 1.003
R4518 a_9167_3699.n6 a_9167_3699.n3 0.833
R4519 a_9167_3699.n3 a_9167_3699.n2 0.653
R4520 a_9167_3699.n7 a_9167_3699.n6 0.653
R4521 a_9167_3699.n3 a_9167_3699.n1 0.341
R4522 a_9167_3699.n6 a_9167_3699.n5 0.032
R4523 a_9757_3262.t2 a_9757_3262.n0 28.565
R4524 a_9757_3262.n0 a_9757_3262.t0 28.565
R4525 a_9757_3262.n0 a_9757_3262.n1 192.754
R4526 a_9757_3262.n1 a_9757_3262.t1 28.568
R4527 a_9757_3262.n1 a_9757_3262.n2 1.123
R4528 a_9757_3262.n2 a_9757_3262.n3 36.155
R4529 a_9757_3262.n3 a_9757_3262.t7 615.911
R4530 a_9757_3262.n3 a_9757_3262.t6 867.497
R4531 a_9757_3262.t6 a_9757_3262.n4 160.666
R4532 a_9757_3262.n4 a_9757_3262.t4 286.438
R4533 a_9757_3262.n4 a_9757_3262.t5 286.438
R4534 a_9757_3262.n2 a_9757_3262.t3 18.726
R4535 a_15456_3694.t8 a_15456_3694.n3 406.053
R4536 a_15456_3694.n2 a_15456_3694.t5 187.473
R4537 a_15456_3694.n4 a_15456_3694.t8 136.943
R4538 a_15456_3694.n3 a_15456_3694.n2 107.801
R4539 a_15456_3694.n2 a_15456_3694.t7 80.333
R4540 a_15456_3694.n3 a_15456_3694.t6 80.333
R4541 a_15456_3694.n1 a_15456_3694.t3 17.4
R4542 a_15456_3694.n1 a_15456_3694.t2 17.4
R4543 a_15456_3694.t0 a_15456_3694.n5 15.036
R4544 a_15456_3694.n0 a_15456_3694.t1 14.282
R4545 a_15456_3694.n0 a_15456_3694.t4 14.282
R4546 a_15456_3694.n5 a_15456_3694.n0 1.654
R4547 a_15456_3694.n4 a_15456_3694.n1 0.672
R4548 a_15456_3694.n5 a_15456_3694.n4 0.665
R4549 a_22290_n990.n2 a_22290_n990.t6 448.382
R4550 a_22290_n990.n1 a_22290_n990.t4 286.438
R4551 a_22290_n990.n1 a_22290_n990.t5 286.438
R4552 a_22290_n990.n0 a_22290_n990.t7 247.69
R4553 a_22290_n990.n4 a_22290_n990.n3 182.117
R4554 a_22290_n990.t6 a_22290_n990.n1 160.666
R4555 a_22290_n990.n3 a_22290_n990.t0 28.568
R4556 a_22290_n990.t2 a_22290_n990.n4 28.565
R4557 a_22290_n990.n4 a_22290_n990.t1 28.565
R4558 a_22290_n990.n0 a_22290_n990.t3 18.127
R4559 a_22290_n990.n2 a_22290_n990.n0 4.039
R4560 a_22290_n990.n3 a_22290_n990.n2 0.937
R4561 a_10167_1718.n0 a_10167_1718.t0 28.565
R4562 a_10167_1718.t2 a_10167_1718.n0 28.565
R4563 a_10167_1718.n0 a_10167_1718.n3 97.131
R4564 a_10167_1718.n3 a_10167_1718.n4 95.622
R4565 a_10167_1718.n4 a_10167_1718.t1 28.568
R4566 a_10167_1718.n4 a_10167_1718.t3 17.641
R4567 a_10167_1718.n3 a_10167_1718.n1 1642.26
R4568 a_10167_1718.n1 a_10167_1718.t6 408.211
R4569 a_10167_1718.n1 a_10167_1718.t7 990.34
R4570 a_10167_1718.t7 a_10167_1718.n2 160.666
R4571 a_10167_1718.n2 a_10167_1718.t5 286.438
R4572 a_10167_1718.n2 a_10167_1718.t4 286.438
R4573 a_16014_1740.n2 a_16014_1740.t4 448.382
R4574 a_16014_1740.n1 a_16014_1740.t6 286.438
R4575 a_16014_1740.n1 a_16014_1740.t7 286.438
R4576 a_16014_1740.n0 a_16014_1740.t5 247.69
R4577 a_16014_1740.n4 a_16014_1740.n3 182.117
R4578 a_16014_1740.t4 a_16014_1740.n1 160.666
R4579 a_16014_1740.n3 a_16014_1740.t0 28.568
R4580 a_16014_1740.n4 a_16014_1740.t1 28.565
R4581 a_16014_1740.t2 a_16014_1740.n4 28.565
R4582 a_16014_1740.n0 a_16014_1740.t3 18.127
R4583 a_16014_1740.n2 a_16014_1740.n0 4.039
R4584 a_16014_1740.n3 a_16014_1740.n2 0.937
R4585 a_3382_n3726.n3 a_3382_n3726.t6 448.382
R4586 a_3382_n3726.n2 a_3382_n3726.t5 286.438
R4587 a_3382_n3726.n2 a_3382_n3726.t7 286.438
R4588 a_3382_n3726.n1 a_3382_n3726.t4 247.69
R4589 a_3382_n3726.n4 a_3382_n3726.n0 182.117
R4590 a_3382_n3726.t6 a_3382_n3726.n2 160.666
R4591 a_3382_n3726.t2 a_3382_n3726.n4 28.568
R4592 a_3382_n3726.n0 a_3382_n3726.t0 28.565
R4593 a_3382_n3726.n0 a_3382_n3726.t1 28.565
R4594 a_3382_n3726.n1 a_3382_n3726.t3 18.127
R4595 a_3382_n3726.n3 a_3382_n3726.n1 4.039
R4596 a_3382_n3726.n4 a_3382_n3726.n3 0.937
R4597 a_4762_n5059.t0 a_4762_n5059.t1 17.4
R4598 a_22290_1744.n2 a_22290_1744.t7 448.382
R4599 a_22290_1744.n1 a_22290_1744.t4 286.438
R4600 a_22290_1744.n1 a_22290_1744.t5 286.438
R4601 a_22290_1744.n0 a_22290_1744.t6 247.69
R4602 a_22290_1744.n4 a_22290_1744.n3 182.117
R4603 a_22290_1744.t7 a_22290_1744.n1 160.666
R4604 a_22290_1744.n3 a_22290_1744.t0 28.568
R4605 a_22290_1744.t2 a_22290_1744.n4 28.565
R4606 a_22290_1744.n4 a_22290_1744.t1 28.565
R4607 a_22290_1744.n0 a_22290_1744.t3 18.127
R4608 a_22290_1744.n2 a_22290_1744.n0 4.039
R4609 a_22290_1744.n3 a_22290_1744.n2 0.937
R4610 a_16014_n994.n2 a_16014_n994.t4 448.382
R4611 a_16014_n994.n1 a_16014_n994.t6 286.438
R4612 a_16014_n994.n1 a_16014_n994.t7 286.438
R4613 a_16014_n994.n0 a_16014_n994.t5 247.69
R4614 a_16014_n994.n4 a_16014_n994.n3 182.117
R4615 a_16014_n994.t4 a_16014_n994.n1 160.666
R4616 a_16014_n994.n3 a_16014_n994.t0 28.568
R4617 a_16014_n994.n4 a_16014_n994.t1 28.565
R4618 a_16014_n994.t2 a_16014_n994.n4 28.565
R4619 a_16014_n994.n0 a_16014_n994.t3 18.127
R4620 a_16014_n994.n2 a_16014_n994.n0 4.039
R4621 a_16014_n994.n3 a_16014_n994.n2 0.937
R4622 A[2].n12 A[2].n5 3389.41
R4623 A[2].t2 A[2].t10 573.627
R4624 A[2].t16 A[2].t4 437.233
R4625 A[2].n11 A[2].n10 412.11
R4626 A[2].n7 A[2].t17 394.151
R4627 A[2].n10 A[2].t11 294.653
R4628 A[2].n0 A[2].t7 285.543
R4629 A[2].n6 A[2].t19 269.523
R4630 A[2].t17 A[2].n6 269.523
R4631 A[2].n11 A[2].n9 224.13
R4632 A[2].n3 A[2].t16 220.881
R4633 A[2].n2 A[2].t6 214.686
R4634 A[2].t4 A[2].n2 214.686
R4635 A[2].n8 A[2].t1 198.043
R4636 A[2].n4 A[2].t9 186.908
R4637 A[2].n4 A[2].t3 186.908
R4638 A[2].n3 A[2].n1 182.197
R4639 A[2].n0 A[2].t14 160.666
R4640 A[2].n1 A[2].t2 160.666
R4641 A[2].n6 A[2].t18 160.666
R4642 A[2].n12 A[2].n11 141.535
R4643 A[2].n5 A[2].t0 140.583
R4644 A[2].n1 A[2].n0 114.089
R4645 A[2].n10 A[2].t12 111.663
R4646 A[2].n4 A[2].t8 109.253
R4647 A[2].n9 A[2].n7 97.816
R4648 A[2].n8 A[2].t5 93.989
R4649 A[2].n2 A[2].t15 80.333
R4650 A[2].n7 A[2].t13 80.333
R4651 A[2].n5 A[2].n4 61.856
R4652 A[2].n13 A[2].n3 31.383
R4653 A[2].n13 A[2].n12 11.764
R4654 A[2].n9 A[2].n8 6.615
R4655 A[2] A[2].n13 2.713
R4656 a_7013_n3748.t2 a_7013_n3748.n0 28.565
R4657 a_7013_n3748.n0 a_7013_n3748.t1 28.565
R4658 a_7013_n3748.n0 a_7013_n3748.n1 195.766
R4659 a_7013_n3748.n1 a_7013_n3748.t0 28.568
R4660 a_7013_n3748.n1 a_7013_n3748.n2 0.462
R4661 a_7013_n3748.n2 a_7013_n3748.n3 38.314
R4662 a_7013_n3748.n3 a_7013_n3748.t7 408.211
R4663 a_7013_n3748.n3 a_7013_n3748.t5 990.34
R4664 a_7013_n3748.t5 a_7013_n3748.n4 160.666
R4665 a_7013_n3748.n4 a_7013_n3748.t6 286.438
R4666 a_7013_n3748.n4 a_7013_n3748.t4 286.438
R4667 a_7013_n3748.n2 a_7013_n3748.t3 18.111
R4668 a_13429_1740.n3 a_13429_1740.n2 167.433
R4669 a_13429_1740.n7 a_13429_1740.n6 167.433
R4670 a_13429_1740.n3 a_13429_1740.t4 104.259
R4671 a_13429_1740.n7 a_13429_1740.t9 104.259
R4672 a_13429_1740.n4 a_13429_1740.n1 89.977
R4673 a_13429_1740.n5 a_13429_1740.n0 89.977
R4674 a_13429_1740.n9 a_13429_1740.n8 89.977
R4675 a_13429_1740.n4 a_13429_1740.n3 77.784
R4676 a_13429_1740.n5 a_13429_1740.n4 77.456
R4677 a_13429_1740.n8 a_13429_1740.n5 77.456
R4678 a_13429_1740.n8 a_13429_1740.n7 75.815
R4679 a_13429_1740.n2 a_13429_1740.t5 14.282
R4680 a_13429_1740.n2 a_13429_1740.t8 14.282
R4681 a_13429_1740.n1 a_13429_1740.t2 14.282
R4682 a_13429_1740.n1 a_13429_1740.t0 14.282
R4683 a_13429_1740.n0 a_13429_1740.t1 14.282
R4684 a_13429_1740.n0 a_13429_1740.t7 14.282
R4685 a_13429_1740.n6 a_13429_1740.t11 14.282
R4686 a_13429_1740.n6 a_13429_1740.t10 14.282
R4687 a_13429_1740.t3 a_13429_1740.n9 14.282
R4688 a_13429_1740.n9 a_13429_1740.t6 14.282
R4689 A[6].n8 A[6].n7 2321.13
R4690 A[6].t18 A[6].t10 575.234
R4691 A[6].t7 A[6].t19 437.233
R4692 A[6].n5 A[6].n4 412.11
R4693 A[6].n1 A[6].t8 394.151
R4694 A[6].n4 A[6].t0 294.653
R4695 A[6].n9 A[6].t5 284.688
R4696 A[6].n0 A[6].t4 269.523
R4697 A[6].t8 A[6].n0 269.523
R4698 A[6].n5 A[6].n3 224.13
R4699 A[6].n12 A[6].t7 222.529
R4700 A[6].n11 A[6].t16 214.686
R4701 A[6].t19 A[6].n11 214.686
R4702 A[6].n2 A[6].t12 198.043
R4703 A[6].n6 A[6].t2 185.301
R4704 A[6].n6 A[6].t17 185.301
R4705 A[6].n12 A[6].n10 181.968
R4706 A[6].n0 A[6].t3 160.666
R4707 A[6].n9 A[6].t15 160.666
R4708 A[6].n10 A[6].t18 160.666
R4709 A[6].n8 A[6].n5 142.366
R4710 A[6].n7 A[6].t11 137.369
R4711 A[6].n10 A[6].n9 115.593
R4712 A[6].n4 A[6].t9 111.663
R4713 A[6].n6 A[6].t1 107.646
R4714 A[6].n3 A[6].n1 97.816
R4715 A[6].n2 A[6].t13 93.989
R4716 A[6].n1 A[6].t14 80.333
R4717 A[6].n11 A[6].t6 80.333
R4718 A[6].n7 A[6].n6 61.856
R4719 A[6].n13 A[6].n12 38.951
R4720 A[6].n13 A[6].n8 31.43
R4721 A[6].n3 A[6].n2 6.615
R4722 A[6] A[6].n13 1.096
R4723 a_13167_n8094.t0 a_13167_n8094.t1 17.4
R4724 a_16004_n3726.n2 a_16004_n3726.t6 448.382
R4725 a_16004_n3726.n1 a_16004_n3726.t5 286.438
R4726 a_16004_n3726.n1 a_16004_n3726.t7 286.438
R4727 a_16004_n3726.n0 a_16004_n3726.t4 247.69
R4728 a_16004_n3726.n4 a_16004_n3726.n3 182.117
R4729 a_16004_n3726.t6 a_16004_n3726.n1 160.666
R4730 a_16004_n3726.n3 a_16004_n3726.t1 28.568
R4731 a_16004_n3726.t2 a_16004_n3726.n4 28.565
R4732 a_16004_n3726.n4 a_16004_n3726.t0 28.565
R4733 a_16004_n3726.n0 a_16004_n3726.t3 18.127
R4734 a_16004_n3726.n2 a_16004_n3726.n0 4.039
R4735 a_16004_n3726.n3 a_16004_n3726.n2 0.937
R4736 a_248_1740.n2 a_248_1740.t5 448.382
R4737 a_248_1740.n1 a_248_1740.t7 286.438
R4738 a_248_1740.n1 a_248_1740.t4 286.438
R4739 a_248_1740.n0 a_248_1740.t6 247.69
R4740 a_248_1740.n4 a_248_1740.n3 182.117
R4741 a_248_1740.t5 a_248_1740.n1 160.666
R4742 a_248_1740.n3 a_248_1740.t0 28.568
R4743 a_248_1740.t2 a_248_1740.n4 28.565
R4744 a_248_1740.n4 a_248_1740.t1 28.565
R4745 a_248_1740.n0 a_248_1740.t3 18.127
R4746 a_248_1740.n2 a_248_1740.n0 4.039
R4747 a_248_1740.n3 a_248_1740.n2 0.937
R4748 a_13778_1740.n4 a_13778_1740.t10 1527.4
R4749 a_13778_1740.t10 a_13778_1740.n3 657.379
R4750 a_13778_1740.n1 a_13778_1740.n0 258.161
R4751 a_13778_1740.n7 a_13778_1740.n6 258.161
R4752 a_13778_1740.n2 a_13778_1740.t9 206.421
R4753 a_13778_1740.t11 a_13778_1740.n2 206.421
R4754 a_13778_1740.n4 a_13778_1740.t11 200.029
R4755 a_13778_1740.n5 a_13778_1740.n4 97.614
R4756 a_13778_1740.n2 a_13778_1740.t8 80.333
R4757 a_13778_1740.n6 a_13778_1740.t4 14.283
R4758 a_13778_1740.n1 a_13778_1740.t3 14.283
R4759 a_13778_1740.n0 a_13778_1740.t7 14.282
R4760 a_13778_1740.n0 a_13778_1740.t2 14.282
R4761 a_13778_1740.n7 a_13778_1740.t5 14.282
R4762 a_13778_1740.t1 a_13778_1740.n7 14.282
R4763 a_13778_1740.n3 a_13778_1740.t6 8.7
R4764 a_13778_1740.n3 a_13778_1740.t0 8.7
R4765 a_13778_1740.n6 a_13778_1740.n5 4.366
R4766 a_13778_1740.n5 a_13778_1740.n1 0.852
R4767 a_8259_3260.t2 a_8259_3260.n0 28.565
R4768 a_8259_3260.n0 a_8259_3260.t0 28.565
R4769 a_8259_3260.n0 a_8259_3260.n1 192.754
R4770 a_8259_3260.n1 a_8259_3260.t1 28.568
R4771 a_8259_3260.n1 a_8259_3260.n2 1.123
R4772 a_8259_3260.n2 a_8259_3260.n3 31.172
R4773 a_8259_3260.n3 a_8259_3260.t4 615.911
R4774 a_8259_3260.n3 a_8259_3260.t6 867.497
R4775 a_8259_3260.t6 a_8259_3260.n4 160.666
R4776 a_8259_3260.n4 a_8259_3260.t7 286.438
R4777 a_8259_3260.n4 a_8259_3260.t5 286.438
R4778 a_8259_3260.n2 a_8259_3260.t3 18.726
R4779 a_17394_407.t0 a_17394_407.t1 17.4
R4780 a_13429_n994.n4 a_13429_n994.n3 167.433
R4781 a_13429_n994.n9 a_13429_n994.n8 167.433
R4782 a_13429_n994.n4 a_13429_n994.t9 104.259
R4783 a_13429_n994.n8 a_13429_n994.t6 104.259
R4784 a_13429_n994.n5 a_13429_n994.n2 89.977
R4785 a_13429_n994.n6 a_13429_n994.n1 89.977
R4786 a_13429_n994.n7 a_13429_n994.n0 89.977
R4787 a_13429_n994.n5 a_13429_n994.n4 77.784
R4788 a_13429_n994.n6 a_13429_n994.n5 77.456
R4789 a_13429_n994.n7 a_13429_n994.n6 77.456
R4790 a_13429_n994.n8 a_13429_n994.n7 75.815
R4791 a_13429_n994.n3 a_13429_n994.t8 14.282
R4792 a_13429_n994.n3 a_13429_n994.t7 14.282
R4793 a_13429_n994.n2 a_13429_n994.t5 14.282
R4794 a_13429_n994.n2 a_13429_n994.t3 14.282
R4795 a_13429_n994.n1 a_13429_n994.t4 14.282
R4796 a_13429_n994.n1 a_13429_n994.t2 14.282
R4797 a_13429_n994.n0 a_13429_n994.t10 14.282
R4798 a_13429_n994.n0 a_13429_n994.t11 14.282
R4799 a_13429_n994.t0 a_13429_n994.n9 14.282
R4800 a_13429_n994.n9 a_13429_n994.t1 14.282
R4801 a_23198_n990.n4 a_23198_n990.t10 1527.4
R4802 a_23198_n990.t10 a_23198_n990.n3 657.379
R4803 a_23198_n990.n1 a_23198_n990.n0 258.161
R4804 a_23198_n990.n7 a_23198_n990.n6 258.161
R4805 a_23198_n990.n2 a_23198_n990.t8 206.421
R4806 a_23198_n990.t9 a_23198_n990.n2 206.421
R4807 a_23198_n990.n4 a_23198_n990.t9 200.029
R4808 a_23198_n990.n5 a_23198_n990.n4 97.614
R4809 a_23198_n990.n2 a_23198_n990.t11 80.333
R4810 a_23198_n990.n6 a_23198_n990.t3 14.283
R4811 a_23198_n990.n1 a_23198_n990.t7 14.283
R4812 a_23198_n990.n0 a_23198_n990.t5 14.282
R4813 a_23198_n990.n0 a_23198_n990.t6 14.282
R4814 a_23198_n990.n7 a_23198_n990.t2 14.282
R4815 a_23198_n990.t1 a_23198_n990.n7 14.282
R4816 a_23198_n990.n3 a_23198_n990.t4 8.7
R4817 a_23198_n990.n3 a_23198_n990.t0 8.7
R4818 a_23198_n990.n6 a_23198_n990.n5 4.366
R4819 a_23198_n990.n5 a_23198_n990.n1 0.852
R4820 a_22849_n990.n4 a_22849_n990.n3 167.433
R4821 a_22849_n990.n9 a_22849_n990.n8 167.433
R4822 a_22849_n990.n4 a_22849_n990.t8 104.259
R4823 a_22849_n990.t0 a_22849_n990.n9 104.259
R4824 a_22849_n990.n5 a_22849_n990.n2 89.977
R4825 a_22849_n990.n6 a_22849_n990.n1 89.977
R4826 a_22849_n990.n7 a_22849_n990.n0 89.977
R4827 a_22849_n990.n5 a_22849_n990.n4 77.784
R4828 a_22849_n990.n6 a_22849_n990.n5 77.456
R4829 a_22849_n990.n7 a_22849_n990.n6 77.456
R4830 a_22849_n990.n9 a_22849_n990.n7 75.815
R4831 a_22849_n990.n3 a_22849_n990.t9 14.282
R4832 a_22849_n990.n3 a_22849_n990.t7 14.282
R4833 a_22849_n990.n2 a_22849_n990.t1 14.282
R4834 a_22849_n990.n2 a_22849_n990.t3 14.282
R4835 a_22849_n990.n1 a_22849_n990.t2 14.282
R4836 a_22849_n990.n1 a_22849_n990.t5 14.282
R4837 a_22849_n990.n0 a_22849_n990.t4 14.282
R4838 a_22849_n990.n0 a_22849_n990.t6 14.282
R4839 a_22849_n990.n8 a_22849_n990.t10 14.282
R4840 a_22849_n990.n8 a_22849_n990.t11 14.282
R4841 a_14454_n6667.n1 a_14454_n6667.t4 318.922
R4842 a_14454_n6667.n0 a_14454_n6667.t6 273.935
R4843 a_14454_n6667.n0 a_14454_n6667.t5 273.935
R4844 a_14454_n6667.n1 a_14454_n6667.t7 269.116
R4845 a_14454_n6667.n4 a_14454_n6667.n3 193.227
R4846 a_14454_n6667.t4 a_14454_n6667.n0 179.142
R4847 a_14454_n6667.n2 a_14454_n6667.n1 106.999
R4848 a_14454_n6667.n3 a_14454_n6667.t1 28.568
R4849 a_14454_n6667.t2 a_14454_n6667.n4 28.565
R4850 a_14454_n6667.n4 a_14454_n6667.t0 28.565
R4851 a_14454_n6667.n2 a_14454_n6667.t3 18.149
R4852 a_14454_n6667.n3 a_14454_n6667.n2 3.726
R4853 a_14999_n7360.n3 a_14999_n7360.n2 2044.44
R4854 a_14999_n7360.n2 a_14999_n7360.t9 867.497
R4855 a_14999_n7360.n2 a_14999_n7360.t11 615.911
R4856 a_14999_n7360.n1 a_14999_n7360.t8 286.438
R4857 a_14999_n7360.n1 a_14999_n7360.t10 286.438
R4858 a_14999_n7360.t9 a_14999_n7360.n1 160.666
R4859 a_14999_n7360.n6 a_14999_n7360.n4 157.665
R4860 a_14999_n7360.n6 a_14999_n7360.n5 122.999
R4861 a_14999_n7360.n3 a_14999_n7360.n0 90.436
R4862 a_14999_n7360.n8 a_14999_n7360.n7 90.416
R4863 a_14999_n7360.n7 a_14999_n7360.n3 74.302
R4864 a_14999_n7360.n7 a_14999_n7360.n6 50.575
R4865 a_14999_n7360.n0 a_14999_n7360.t0 14.282
R4866 a_14999_n7360.n0 a_14999_n7360.t1 14.282
R4867 a_14999_n7360.n5 a_14999_n7360.t6 14.282
R4868 a_14999_n7360.n5 a_14999_n7360.t4 14.282
R4869 a_14999_n7360.t2 a_14999_n7360.n8 14.282
R4870 a_14999_n7360.n8 a_14999_n7360.t5 14.282
R4871 a_14999_n7360.n4 a_14999_n7360.t3 8.7
R4872 a_14999_n7360.n4 a_14999_n7360.t7 8.7
R4873 a_9658_n3722.n3 a_9658_n3722.t6 448.382
R4874 a_9658_n3722.n2 a_9658_n3722.t5 286.438
R4875 a_9658_n3722.n2 a_9658_n3722.t7 286.438
R4876 a_9658_n3722.n1 a_9658_n3722.t4 247.69
R4877 a_9658_n3722.n4 a_9658_n3722.n0 182.117
R4878 a_9658_n3722.t6 a_9658_n3722.n2 160.666
R4879 a_9658_n3722.t2 a_9658_n3722.n4 28.568
R4880 a_9658_n3722.n0 a_9658_n3722.t0 28.565
R4881 a_9658_n3722.n0 a_9658_n3722.t1 28.565
R4882 a_9658_n3722.n1 a_9658_n3722.t3 18.127
R4883 a_9658_n3722.n3 a_9658_n3722.n1 4.039
R4884 a_9658_n3722.n4 a_9658_n3722.n3 0.937
R4885 a_4825_n1479.t2 a_4825_n1479.n0 28.565
R4886 a_4825_n1479.n0 a_4825_n1479.t0 28.565
R4887 a_4825_n1479.n0 a_4825_n1479.n1 185.55
R4888 a_4825_n1479.n1 a_4825_n1479.t1 28.568
R4889 a_4825_n1479.n1 a_4825_n1479.n4 1.637
R4890 a_4825_n1479.n4 a_4825_n1479.t3 21.373
R4891 a_4825_n1479.n4 a_4825_n1479.n2 26.016
R4892 a_4825_n1479.n2 a_4825_n1479.t4 615.911
R4893 a_4825_n1479.n2 a_4825_n1479.t7 867.497
R4894 a_4825_n1479.t7 a_4825_n1479.n3 160.666
R4895 a_4825_n1479.n3 a_4825_n1479.t6 286.438
R4896 a_4825_n1479.n3 a_4825_n1479.t5 286.438
R4897 a_11048_411.t0 a_11048_411.t1 17.4
R4898 a_13768_n3726.n3 a_13768_n3726.t8 1527.4
R4899 a_13768_n3726.t8 a_13768_n3726.n2 657.379
R4900 a_13768_n3726.n5 a_13768_n3726.n4 258.161
R4901 a_13768_n3726.n7 a_13768_n3726.n0 258.161
R4902 a_13768_n3726.n1 a_13768_n3726.t9 206.421
R4903 a_13768_n3726.t11 a_13768_n3726.n1 206.421
R4904 a_13768_n3726.n3 a_13768_n3726.t11 200.029
R4905 a_13768_n3726.n6 a_13768_n3726.n3 97.614
R4906 a_13768_n3726.n1 a_13768_n3726.t10 80.333
R4907 a_13768_n3726.n5 a_13768_n3726.t7 14.283
R4908 a_13768_n3726.t1 a_13768_n3726.n7 14.283
R4909 a_13768_n3726.n4 a_13768_n3726.t6 14.282
R4910 a_13768_n3726.n4 a_13768_n3726.t3 14.282
R4911 a_13768_n3726.n0 a_13768_n3726.t4 14.282
R4912 a_13768_n3726.n0 a_13768_n3726.t5 14.282
R4913 a_13768_n3726.n2 a_13768_n3726.t0 8.7
R4914 a_13768_n3726.n2 a_13768_n3726.t2 8.7
R4915 a_13768_n3726.n6 a_13768_n3726.n5 4.366
R4916 a_13768_n3726.n7 a_13768_n3726.n6 0.852
R4917 a_13369_n1020.t2 a_13369_n1020.n0 28.565
R4918 a_13369_n1020.n0 a_13369_n1020.t1 28.565
R4919 a_13369_n1020.n1 a_13369_n1020.n2 0.002
R4920 a_13369_n1020.n0 a_13369_n1020.n1 185.55
R4921 a_13369_n1020.n1 a_13369_n1020.t0 28.568
R4922 a_13369_n1020.n2 a_13369_n1020.t3 23.43
R4923 a_13369_n1020.n2 a_13369_n1020.n3 11.505
R4924 a_13369_n1020.n3 a_13369_n1020.t6 408.211
R4925 a_13369_n1020.n3 a_13369_n1020.t4 990.34
R4926 a_13369_n1020.t4 a_13369_n1020.n4 160.666
R4927 a_13369_n1020.n4 a_13369_n1020.t7 286.438
R4928 a_13369_n1020.n4 a_13369_n1020.t5 286.438
R4929 a_23198_1744.n2 a_23198_1744.t10 1527.4
R4930 a_23198_1744.t10 a_23198_1744.n1 657.379
R4931 a_23198_1744.n4 a_23198_1744.n3 258.161
R4932 a_23198_1744.n7 a_23198_1744.n6 258.161
R4933 a_23198_1744.n0 a_23198_1744.t8 206.421
R4934 a_23198_1744.t9 a_23198_1744.n0 206.421
R4935 a_23198_1744.n2 a_23198_1744.t9 200.029
R4936 a_23198_1744.n5 a_23198_1744.n2 97.614
R4937 a_23198_1744.n0 a_23198_1744.t11 80.333
R4938 a_23198_1744.n4 a_23198_1744.t5 14.283
R4939 a_23198_1744.n6 a_23198_1744.t6 14.283
R4940 a_23198_1744.n3 a_23198_1744.t4 14.282
R4941 a_23198_1744.n3 a_23198_1744.t2 14.282
R4942 a_23198_1744.t1 a_23198_1744.n7 14.282
R4943 a_23198_1744.n7 a_23198_1744.t7 14.282
R4944 a_23198_1744.n1 a_23198_1744.t3 8.7
R4945 a_23198_1744.n1 a_23198_1744.t0 8.7
R4946 a_23198_1744.n5 a_23198_1744.n4 4.366
R4947 a_23198_1744.n6 a_23198_1744.n5 0.852
R4948 a_22849_1744.n4 a_22849_1744.n3 167.433
R4949 a_22849_1744.n9 a_22849_1744.n8 167.433
R4950 a_22849_1744.n4 a_22849_1744.t11 104.259
R4951 a_22849_1744.t0 a_22849_1744.n9 104.259
R4952 a_22849_1744.n5 a_22849_1744.n2 89.977
R4953 a_22849_1744.n6 a_22849_1744.n1 89.977
R4954 a_22849_1744.n7 a_22849_1744.n0 89.977
R4955 a_22849_1744.n5 a_22849_1744.n4 77.784
R4956 a_22849_1744.n6 a_22849_1744.n5 77.456
R4957 a_22849_1744.n7 a_22849_1744.n6 77.456
R4958 a_22849_1744.n9 a_22849_1744.n7 75.815
R4959 a_22849_1744.n3 a_22849_1744.t10 14.282
R4960 a_22849_1744.n3 a_22849_1744.t5 14.282
R4961 a_22849_1744.n2 a_22849_1744.t2 14.282
R4962 a_22849_1744.n2 a_22849_1744.t4 14.282
R4963 a_22849_1744.n1 a_22849_1744.t3 14.282
R4964 a_22849_1744.n1 a_22849_1744.t8 14.282
R4965 a_22849_1744.n0 a_22849_1744.t7 14.282
R4966 a_22849_1744.n0 a_22849_1744.t9 14.282
R4967 a_22849_1744.n8 a_22849_1744.t6 14.282
R4968 a_22849_1744.n8 a_22849_1744.t1 14.282
R4969 B[5].t0 B[5].t7 800.874
R4970 B[5].n9 B[5].n8 649.333
R4971 B[5].n5 B[5].n4 592.056
R4972 B[5].t10 B[5].t5 415.315
R4973 B[5].t11 B[5].n2 313.873
R4974 B[5].n4 B[5].t9 294.986
R4975 B[5].n7 B[5].t3 285.543
R4976 B[5].n1 B[5].t13 272.288
R4977 B[5].n6 B[5].t10 217.527
R4978 B[5].n0 B[5].t12 214.335
R4979 B[5].t5 B[5].n0 214.335
R4980 B[5].n5 B[5].t1 204.68
R4981 B[5].n8 B[5].t0 194.406
R4982 B[5].n3 B[5].t11 190.152
R4983 B[5].n3 B[5].t2 190.152
R4984 B[5].n1 B[5].t14 160.666
R4985 B[5].n2 B[5].t4 160.666
R4986 B[5].n7 B[5].t8 160.666
R4987 B[5].n4 B[5].t15 110.859
R4988 B[5].n2 B[5].n1 96.129
R4989 B[5].n8 B[5].n7 91.137
R4990 B[5].n0 B[5].t6 80.333
R4991 B[5].t1 B[5].n3 80.333
R4992 B[5].n6 B[5].n5 51.127
R4993 B[5] B[5].n9 18.713
R4994 B[5].n9 B[5].n6 5.864
R4995 a_248_n994.n2 a_248_n994.t5 448.382
R4996 a_248_n994.n1 a_248_n994.t7 286.438
R4997 a_248_n994.n1 a_248_n994.t4 286.438
R4998 a_248_n994.n0 a_248_n994.t6 247.69
R4999 a_248_n994.n4 a_248_n994.n3 182.117
R5000 a_248_n994.t5 a_248_n994.n1 160.666
R5001 a_248_n994.n3 a_248_n994.t0 28.568
R5002 a_248_n994.t2 a_248_n994.n4 28.565
R5003 a_248_n994.n4 a_248_n994.t1 28.565
R5004 a_248_n994.n0 a_248_n994.t3 18.127
R5005 a_248_n994.n2 a_248_n994.n0 4.039
R5006 a_248_n994.n3 a_248_n994.n2 0.937
R5007 a_13778_n994.n4 a_13778_n994.t10 1527.4
R5008 a_13778_n994.t10 a_13778_n994.n3 657.379
R5009 a_13778_n994.n1 a_13778_n994.n0 258.161
R5010 a_13778_n994.n7 a_13778_n994.n6 258.161
R5011 a_13778_n994.n2 a_13778_n994.t9 206.421
R5012 a_13778_n994.t11 a_13778_n994.n2 206.421
R5013 a_13778_n994.n4 a_13778_n994.t11 200.029
R5014 a_13778_n994.n5 a_13778_n994.n4 97.614
R5015 a_13778_n994.n2 a_13778_n994.t8 80.333
R5016 a_13778_n994.n6 a_13778_n994.t7 14.283
R5017 a_13778_n994.n1 a_13778_n994.t4 14.283
R5018 a_13778_n994.n0 a_13778_n994.t3 14.282
R5019 a_13778_n994.n0 a_13778_n994.t5 14.282
R5020 a_13778_n994.t0 a_13778_n994.n7 14.282
R5021 a_13778_n994.n7 a_13778_n994.t6 14.282
R5022 a_13778_n994.n3 a_13778_n994.t2 8.7
R5023 a_13778_n994.n3 a_13778_n994.t1 8.7
R5024 a_13778_n994.n6 a_13778_n994.n5 4.366
R5025 a_13778_n994.n5 a_13778_n994.n1 0.852
R5026 Y[4].n1 Y[4].n0 185.55
R5027 Y[4].n1 Y[4].t0 28.568
R5028 Y[4].n0 Y[4].t2 28.565
R5029 Y[4].n0 Y[4].t1 28.565
R5030 Y[4].n2 Y[4].t3 21.559
R5031 Y[4] Y[4].n2 13.933
R5032 Y[4].n2 Y[4].n1 1.603
R5033 a_19635_n3748.n0 a_19635_n3748.t0 28.565
R5034 a_19635_n3748.t2 a_19635_n3748.n0 28.565
R5035 a_19635_n3748.n0 a_19635_n3748.n1 197.272
R5036 a_19635_n3748.n1 a_19635_n3748.t1 28.568
R5037 a_19635_n3748.n1 a_19635_n3748.n2 0.467
R5038 a_19635_n3748.n2 a_19635_n3748.n3 13.505
R5039 a_19635_n3748.n3 a_19635_n3748.t4 408.211
R5040 a_19635_n3748.n3 a_19635_n3748.t6 990.34
R5041 a_19635_n3748.t6 a_19635_n3748.n4 160.666
R5042 a_19635_n3748.n4 a_19635_n3748.t7 286.438
R5043 a_19635_n3748.n4 a_19635_n3748.t5 286.438
R5044 a_19635_n3748.n2 a_19635_n3748.t3 18.085
R5045 a_4112_n6671.n2 a_4112_n6671.t6 318.922
R5046 a_4112_n6671.n1 a_4112_n6671.t4 273.935
R5047 a_4112_n6671.n1 a_4112_n6671.t7 273.935
R5048 a_4112_n6671.n2 a_4112_n6671.t5 269.116
R5049 a_4112_n6671.n4 a_4112_n6671.n0 193.227
R5050 a_4112_n6671.t6 a_4112_n6671.n1 179.142
R5051 a_4112_n6671.n3 a_4112_n6671.n2 106.999
R5052 a_4112_n6671.t2 a_4112_n6671.n4 28.568
R5053 a_4112_n6671.n0 a_4112_n6671.t0 28.565
R5054 a_4112_n6671.n0 a_4112_n6671.t1 28.565
R5055 a_4112_n6671.n3 a_4112_n6671.t3 18.149
R5056 a_4112_n6671.n4 a_4112_n6671.n3 3.726
R5057 B[6].t10 B[6].t3 800.875
R5058 B[6].n9 B[6].n8 648.993
R5059 B[6].n4 B[6].n3 592.056
R5060 B[6].t14 B[6].t8 415.315
R5061 B[6].t4 B[6].n1 313.873
R5062 B[6].n3 B[6].t0 294.986
R5063 B[6].n7 B[6].t12 284.688
R5064 B[6].n0 B[6].t1 272.288
R5065 B[6].n6 B[6].t14 217.532
R5066 B[6].n5 B[6].t11 214.335
R5067 B[6].t8 B[6].n5 214.335
R5068 B[6].n4 B[6].t5 204.68
R5069 B[6].n8 B[6].t10 192.799
R5070 B[6].n2 B[6].t4 190.152
R5071 B[6].n2 B[6].t9 190.152
R5072 B[6].n0 B[6].t6 160.666
R5073 B[6].n1 B[6].t13 160.666
R5074 B[6].n7 B[6].t2 160.666
R5075 B[6].n3 B[6].t7 110.859
R5076 B[6].n1 B[6].n0 96.129
R5077 B[6].n8 B[6].n7 91.889
R5078 B[6].n5 B[6].t15 80.333
R5079 B[6].t5 B[6].n2 80.333
R5080 B[6].n6 B[6].n4 51.824
R5081 B[6] B[6].n9 21.809
R5082 B[6].n9 B[6].n6 6.378
R5083 a_814_n7390.n1 a_814_n7390.t5 318.922
R5084 a_814_n7390.n0 a_814_n7390.t4 274.739
R5085 a_814_n7390.n0 a_814_n7390.t6 274.739
R5086 a_814_n7390.n1 a_814_n7390.t7 269.116
R5087 a_814_n7390.t5 a_814_n7390.n0 179.946
R5088 a_814_n7390.n2 a_814_n7390.n1 107.263
R5089 a_814_n7390.t0 a_814_n7390.n4 29.444
R5090 a_814_n7390.n3 a_814_n7390.t2 28.565
R5091 a_814_n7390.n3 a_814_n7390.t1 28.565
R5092 a_814_n7390.n2 a_814_n7390.t3 18.145
R5093 a_814_n7390.n4 a_814_n7390.n2 2.878
R5094 a_814_n7390.n4 a_814_n7390.n3 0.764
R5095 a_520_n7364.n5 a_520_n7364.n4 1297.25
R5096 a_520_n7364.n4 a_520_n7364.t8 867.497
R5097 a_520_n7364.n4 a_520_n7364.t10 615.911
R5098 a_520_n7364.n3 a_520_n7364.t11 286.438
R5099 a_520_n7364.n3 a_520_n7364.t9 286.438
R5100 a_520_n7364.t8 a_520_n7364.n3 160.666
R5101 a_520_n7364.n7 a_520_n7364.n0 157.665
R5102 a_520_n7364.n8 a_520_n7364.n7 122.999
R5103 a_520_n7364.n5 a_520_n7364.n2 90.436
R5104 a_520_n7364.n6 a_520_n7364.n1 90.416
R5105 a_520_n7364.n6 a_520_n7364.n5 74.302
R5106 a_520_n7364.n7 a_520_n7364.n6 50.575
R5107 a_520_n7364.n2 a_520_n7364.t4 14.282
R5108 a_520_n7364.n2 a_520_n7364.t5 14.282
R5109 a_520_n7364.n1 a_520_n7364.t6 14.282
R5110 a_520_n7364.n1 a_520_n7364.t1 14.282
R5111 a_520_n7364.n8 a_520_n7364.t2 14.282
R5112 a_520_n7364.t0 a_520_n7364.n8 14.282
R5113 a_520_n7364.n0 a_520_n7364.t7 8.7
R5114 a_520_n7364.n0 a_520_n7364.t3 8.7
R5115 a_402_n7364.n8 a_402_n7364.n0 267.767
R5116 a_402_n7364.n4 a_402_n7364.t4 16.058
R5117 a_402_n7364.n2 a_402_n7364.t5 16.058
R5118 a_402_n7364.n3 a_402_n7364.t2 14.282
R5119 a_402_n7364.n3 a_402_n7364.t3 14.282
R5120 a_402_n7364.n1 a_402_n7364.t6 14.282
R5121 a_402_n7364.n1 a_402_n7364.t7 14.282
R5122 a_402_n7364.n6 a_402_n7364.t10 14.282
R5123 a_402_n7364.n6 a_402_n7364.t11 14.282
R5124 a_402_n7364.n0 a_402_n7364.t8 14.282
R5125 a_402_n7364.n0 a_402_n7364.t1 14.282
R5126 a_402_n7364.t0 a_402_n7364.n9 14.282
R5127 a_402_n7364.n9 a_402_n7364.t9 14.282
R5128 a_402_n7364.n7 a_402_n7364.n6 1.511
R5129 a_402_n7364.n4 a_402_n7364.n3 0.999
R5130 a_402_n7364.n2 a_402_n7364.n1 0.999
R5131 a_402_n7364.n8 a_402_n7364.n7 0.669
R5132 a_402_n7364.n5 a_402_n7364.n4 0.575
R5133 a_402_n7364.n7 a_402_n7364.n5 0.227
R5134 a_402_n7364.n5 a_402_n7364.n2 0.2
R5135 a_402_n7364.n9 a_402_n7364.n8 0.001
R5136 a_16912_n3726.n4 a_16912_n3726.t8 1527.4
R5137 a_16912_n3726.t8 a_16912_n3726.n3 657.379
R5138 a_16912_n3726.n1 a_16912_n3726.n0 258.161
R5139 a_16912_n3726.n7 a_16912_n3726.n6 258.161
R5140 a_16912_n3726.n2 a_16912_n3726.t11 206.421
R5141 a_16912_n3726.t10 a_16912_n3726.n2 206.421
R5142 a_16912_n3726.n4 a_16912_n3726.t10 200.029
R5143 a_16912_n3726.n5 a_16912_n3726.n4 97.614
R5144 a_16912_n3726.n2 a_16912_n3726.t9 80.333
R5145 a_16912_n3726.n6 a_16912_n3726.t4 14.283
R5146 a_16912_n3726.n1 a_16912_n3726.t6 14.283
R5147 a_16912_n3726.n0 a_16912_n3726.t7 14.282
R5148 a_16912_n3726.n0 a_16912_n3726.t5 14.282
R5149 a_16912_n3726.t2 a_16912_n3726.n7 14.282
R5150 a_16912_n3726.n7 a_16912_n3726.t3 14.282
R5151 a_16912_n3726.n3 a_16912_n3726.t1 8.7
R5152 a_16912_n3726.n3 a_16912_n3726.t0 8.7
R5153 a_16912_n3726.n6 a_16912_n3726.n5 4.366
R5154 a_16912_n3726.n5 a_16912_n3726.n1 0.852
R5155 a_14288_3692.t8 a_14288_3692.n2 404.877
R5156 a_14288_3692.n1 a_14288_3692.t5 210.902
R5157 a_14288_3692.n3 a_14288_3692.t8 136.943
R5158 a_14288_3692.n2 a_14288_3692.n1 107.801
R5159 a_14288_3692.n1 a_14288_3692.t6 80.333
R5160 a_14288_3692.n2 a_14288_3692.t7 80.333
R5161 a_14288_3692.n0 a_14288_3692.t0 17.4
R5162 a_14288_3692.n0 a_14288_3692.t1 17.4
R5163 a_14288_3692.n4 a_14288_3692.t3 15.029
R5164 a_14288_3692.t2 a_14288_3692.n5 14.282
R5165 a_14288_3692.n5 a_14288_3692.t4 14.282
R5166 a_14288_3692.n5 a_14288_3692.n4 1.647
R5167 a_14288_3692.n3 a_14288_3692.n0 0.672
R5168 a_14288_3692.n4 a_14288_3692.n3 0.665
R5169 a_14406_3692.n1 a_14406_3692.t1 14.282
R5170 a_14406_3692.n1 a_14406_3692.t4 14.282
R5171 a_14406_3692.n0 a_14406_3692.t3 14.282
R5172 a_14406_3692.n0 a_14406_3692.t5 14.282
R5173 a_14406_3692.n3 a_14406_3692.t0 14.282
R5174 a_14406_3692.t2 a_14406_3692.n3 14.282
R5175 a_14406_3692.n2 a_14406_3692.n0 2.554
R5176 a_14406_3692.n3 a_14406_3692.n2 2.361
R5177 a_14406_3692.n2 a_14406_3692.n1 0.001
R5178 A[3].n8 A[3].n7 3150.3
R5179 A[3].t15 A[3].t8 575.234
R5180 A[3].t11 A[3].t6 437.233
R5181 A[3].n5 A[3].n4 412.11
R5182 A[3].n1 A[3].t2 394.151
R5183 A[3].n4 A[3].t0 294.653
R5184 A[3].n9 A[3].t19 284.688
R5185 A[3].n0 A[3].t9 269.523
R5186 A[3].t2 A[3].n0 269.523
R5187 A[3].n5 A[3].n3 224.13
R5188 A[3].n12 A[3].t11 221.268
R5189 A[3].n11 A[3].t1 214.686
R5190 A[3].t6 A[3].n11 214.686
R5191 A[3].n2 A[3].t12 198.043
R5192 A[3].n6 A[3].t5 185.301
R5193 A[3].n6 A[3].t16 185.301
R5194 A[3].n12 A[3].n10 182.757
R5195 A[3].n9 A[3].t7 160.666
R5196 A[3].n10 A[3].t15 160.666
R5197 A[3].n0 A[3].t4 160.666
R5198 A[3].n8 A[3].n5 141.789
R5199 A[3].n7 A[3].t17 140.583
R5200 A[3].n10 A[3].n9 115.593
R5201 A[3].n4 A[3].t3 111.663
R5202 A[3].n6 A[3].t18 107.646
R5203 A[3].n3 A[3].n1 97.816
R5204 A[3].n2 A[3].t13 93.989
R5205 A[3].n11 A[3].t10 80.333
R5206 A[3].n1 A[3].t14 80.333
R5207 A[3].n7 A[3].n6 61.856
R5208 A[3].n13 A[3].n12 30.336
R5209 A[3].n13 A[3].n8 13.792
R5210 A[3].n3 A[3].n2 6.615
R5211 A[3] A[3].n13 2.396
R5212 a_6961_n8094.t0 a_6961_n8094.t1 17.4
R5213 a_11156_n7386.n1 a_11156_n7386.t5 318.922
R5214 a_11156_n7386.n0 a_11156_n7386.t4 274.739
R5215 a_11156_n7386.n0 a_11156_n7386.t6 274.739
R5216 a_11156_n7386.n1 a_11156_n7386.t7 269.116
R5217 a_11156_n7386.t5 a_11156_n7386.n0 179.946
R5218 a_11156_n7386.n2 a_11156_n7386.n1 107.263
R5219 a_11156_n7386.n3 a_11156_n7386.t1 29.444
R5220 a_11156_n7386.t2 a_11156_n7386.n4 28.565
R5221 a_11156_n7386.n4 a_11156_n7386.t0 28.565
R5222 a_11156_n7386.n2 a_11156_n7386.t3 18.145
R5223 a_11156_n7386.n3 a_11156_n7386.n2 2.878
R5224 a_11156_n7386.n4 a_11156_n7386.n3 0.764
R5225 a_4657_n7364.n5 a_4657_n7364.n4 952.988
R5226 a_4657_n7364.n4 a_4657_n7364.t9 867.497
R5227 a_4657_n7364.n4 a_4657_n7364.t11 615.911
R5228 a_4657_n7364.n3 a_4657_n7364.t8 286.438
R5229 a_4657_n7364.n3 a_4657_n7364.t10 286.438
R5230 a_4657_n7364.t9 a_4657_n7364.n3 160.666
R5231 a_4657_n7364.n7 a_4657_n7364.n0 157.665
R5232 a_4657_n7364.n8 a_4657_n7364.n7 122.999
R5233 a_4657_n7364.n5 a_4657_n7364.n2 90.436
R5234 a_4657_n7364.n6 a_4657_n7364.n1 90.416
R5235 a_4657_n7364.n6 a_4657_n7364.n5 74.302
R5236 a_4657_n7364.n7 a_4657_n7364.n6 50.575
R5237 a_4657_n7364.n2 a_4657_n7364.t6 14.282
R5238 a_4657_n7364.n2 a_4657_n7364.t7 14.282
R5239 a_4657_n7364.n1 a_4657_n7364.t5 14.282
R5240 a_4657_n7364.n1 a_4657_n7364.t3 14.282
R5241 a_4657_n7364.n8 a_4657_n7364.t4 14.282
R5242 a_4657_n7364.t1 a_4657_n7364.n8 14.282
R5243 a_4657_n7364.n0 a_4657_n7364.t0 8.7
R5244 a_4657_n7364.n0 a_4657_n7364.t2 8.7
R5245 a_7073_n3722.n4 a_7073_n3722.n3 167.433
R5246 a_7073_n3722.n9 a_7073_n3722.n8 167.433
R5247 a_7073_n3722.n8 a_7073_n3722.t5 104.259
R5248 a_7073_n3722.n4 a_7073_n3722.t0 104.259
R5249 a_7073_n3722.n7 a_7073_n3722.n0 89.977
R5250 a_7073_n3722.n6 a_7073_n3722.n1 89.977
R5251 a_7073_n3722.n5 a_7073_n3722.n2 89.977
R5252 a_7073_n3722.n8 a_7073_n3722.n7 77.784
R5253 a_7073_n3722.n7 a_7073_n3722.n6 77.456
R5254 a_7073_n3722.n6 a_7073_n3722.n5 77.456
R5255 a_7073_n3722.n5 a_7073_n3722.n4 75.815
R5256 a_7073_n3722.n0 a_7073_n3722.t8 14.282
R5257 a_7073_n3722.n0 a_7073_n3722.t6 14.282
R5258 a_7073_n3722.n1 a_7073_n3722.t7 14.282
R5259 a_7073_n3722.n1 a_7073_n3722.t11 14.282
R5260 a_7073_n3722.n2 a_7073_n3722.t10 14.282
R5261 a_7073_n3722.n2 a_7073_n3722.t9 14.282
R5262 a_7073_n3722.n3 a_7073_n3722.t1 14.282
R5263 a_7073_n3722.n3 a_7073_n3722.t2 14.282
R5264 a_7073_n3722.t3 a_7073_n3722.n9 14.282
R5265 a_7073_n3722.n9 a_7073_n3722.t4 14.282
R5266 a_7422_n3722.n5 a_7422_n3722.t11 1527.4
R5267 a_7422_n3722.t11 a_7422_n3722.n4 657.379
R5268 a_7422_n3722.n7 a_7422_n3722.n0 258.161
R5269 a_7422_n3722.n2 a_7422_n3722.n1 258.161
R5270 a_7422_n3722.n3 a_7422_n3722.t10 206.421
R5271 a_7422_n3722.t9 a_7422_n3722.n3 206.421
R5272 a_7422_n3722.n5 a_7422_n3722.t9 200.029
R5273 a_7422_n3722.n6 a_7422_n3722.n5 97.614
R5274 a_7422_n3722.n3 a_7422_n3722.t8 80.333
R5275 a_7422_n3722.n2 a_7422_n3722.t0 14.283
R5276 a_7422_n3722.t4 a_7422_n3722.n7 14.283
R5277 a_7422_n3722.n0 a_7422_n3722.t7 14.282
R5278 a_7422_n3722.n0 a_7422_n3722.t5 14.282
R5279 a_7422_n3722.n1 a_7422_n3722.t1 14.282
R5280 a_7422_n3722.n1 a_7422_n3722.t2 14.282
R5281 a_7422_n3722.n4 a_7422_n3722.t6 8.7
R5282 a_7422_n3722.n4 a_7422_n3722.t3 8.7
R5283 a_7422_n3722.n7 a_7422_n3722.n6 4.366
R5284 a_7422_n3722.n6 a_7422_n3722.n2 0.852
R5285 a_19230_3112.t1 a_19230_3112.n0 28.565
R5286 a_19230_3112.n0 a_19230_3112.t3 28.565
R5287 a_19230_3112.n0 a_19230_3112.n2 100.24
R5288 a_19230_3112.n2 a_19230_3112.n3 566.188
R5289 a_19230_3112.n3 a_19230_3112.t4 408.211
R5290 a_19230_3112.n3 a_19230_3112.t7 990.34
R5291 a_19230_3112.t7 a_19230_3112.n4 160.666
R5292 a_19230_3112.n4 a_19230_3112.t6 286.438
R5293 a_19230_3112.n4 a_19230_3112.t5 286.438
R5294 a_19230_3112.n2 a_19230_3112.n1 100.603
R5295 a_19230_3112.n1 a_19230_3112.t2 28.568
R5296 a_19230_3112.n1 a_19230_3112.t0 17.64
R5297 a_20290_411.t0 a_20290_411.t1 17.4
R5298 a_3253_3699.n4 a_3253_3699.t7 214.335
R5299 a_3253_3699.t10 a_3253_3699.n4 214.335
R5300 a_3253_3699.n5 a_3253_3699.t10 143.851
R5301 a_3253_3699.n5 a_3253_3699.t8 135.658
R5302 a_3253_3699.n4 a_3253_3699.t9 80.333
R5303 a_3253_3699.n0 a_3253_3699.t3 28.565
R5304 a_3253_3699.n0 a_3253_3699.t4 28.565
R5305 a_3253_3699.n2 a_3253_3699.t0 28.565
R5306 a_3253_3699.n2 a_3253_3699.t5 28.565
R5307 a_3253_3699.t2 a_3253_3699.n7 28.565
R5308 a_3253_3699.n7 a_3253_3699.t1 28.565
R5309 a_3253_3699.n1 a_3253_3699.t6 9.714
R5310 a_3253_3699.n1 a_3253_3699.n0 1.003
R5311 a_3253_3699.n6 a_3253_3699.n3 0.833
R5312 a_3253_3699.n3 a_3253_3699.n2 0.653
R5313 a_3253_3699.n7 a_3253_3699.n6 0.653
R5314 a_3253_3699.n3 a_3253_3699.n1 0.341
R5315 a_3253_3699.n6 a_3253_3699.n5 0.032
R5316 a_3843_3262.t2 a_3843_3262.n0 28.568
R5317 a_3843_3262.n0 a_3843_3262.n4 192.754
R5318 a_3843_3262.n4 a_3843_3262.t0 28.565
R5319 a_3843_3262.n4 a_3843_3262.t1 28.565
R5320 a_3843_3262.n0 a_3843_3262.n1 1.123
R5321 a_3843_3262.n1 a_3843_3262.n2 22.54
R5322 a_3843_3262.n2 a_3843_3262.t5 615.911
R5323 a_3843_3262.n2 a_3843_3262.t4 867.497
R5324 a_3843_3262.t4 a_3843_3262.n3 160.666
R5325 a_3843_3262.n3 a_3843_3262.t7 286.438
R5326 a_3843_3262.n3 a_3843_3262.t6 286.438
R5327 a_3843_3262.n1 a_3843_3262.t3 18.726
R5328 a_238_n3726.n2 a_238_n3726.t6 448.382
R5329 a_238_n3726.n1 a_238_n3726.t5 286.438
R5330 a_238_n3726.n1 a_238_n3726.t7 286.438
R5331 a_238_n3726.n0 a_238_n3726.t4 247.69
R5332 a_238_n3726.n4 a_238_n3726.n3 182.117
R5333 a_238_n3726.t6 a_238_n3726.n1 160.666
R5334 a_238_n3726.n3 a_238_n3726.t0 28.568
R5335 a_238_n3726.n4 a_238_n3726.t1 28.565
R5336 a_238_n3726.t2 a_238_n3726.n4 28.565
R5337 a_238_n3726.n0 a_238_n3726.t3 18.127
R5338 a_238_n3726.n2 a_238_n3726.n0 4.039
R5339 a_238_n3726.n3 a_238_n3726.n2 0.937
R5340 a_13225_n7388.n1 a_13225_n7388.t6 318.922
R5341 a_13225_n7388.n0 a_13225_n7388.t5 274.739
R5342 a_13225_n7388.n0 a_13225_n7388.t7 274.739
R5343 a_13225_n7388.n1 a_13225_n7388.t4 269.116
R5344 a_13225_n7388.t6 a_13225_n7388.n0 179.946
R5345 a_13225_n7388.n2 a_13225_n7388.n1 107.263
R5346 a_13225_n7388.n3 a_13225_n7388.t0 29.444
R5347 a_13225_n7388.n4 a_13225_n7388.t1 28.565
R5348 a_13225_n7388.t2 a_13225_n7388.n4 28.565
R5349 a_13225_n7388.n2 a_13225_n7388.t3 18.145
R5350 a_13225_n7388.n3 a_13225_n7388.n2 2.878
R5351 a_13225_n7388.n4 a_13225_n7388.n3 0.764
R5352 a_12931_n8094.t0 a_12931_n8094.t1 380.209
R5353 a_12070_3694.n1 a_12070_3694.t1 14.282
R5354 a_12070_3694.n1 a_12070_3694.t3 14.282
R5355 a_12070_3694.n0 a_12070_3694.t2 14.282
R5356 a_12070_3694.n0 a_12070_3694.t4 14.282
R5357 a_12070_3694.t0 a_12070_3694.n3 14.282
R5358 a_12070_3694.n3 a_12070_3694.t5 14.282
R5359 a_12070_3694.n2 a_12070_3694.n0 2.538
R5360 a_12070_3694.n3 a_12070_3694.n2 2.375
R5361 a_12070_3694.n2 a_12070_3694.n1 0.001
R5362 a_13419_n3726.n4 a_13419_n3726.n3 167.433
R5363 a_13419_n3726.n9 a_13419_n3726.n8 167.433
R5364 a_13419_n3726.n4 a_13419_n3726.t9 104.259
R5365 a_13419_n3726.n8 a_13419_n3726.t1 104.259
R5366 a_13419_n3726.n5 a_13419_n3726.n2 89.977
R5367 a_13419_n3726.n6 a_13419_n3726.n1 89.977
R5368 a_13419_n3726.n7 a_13419_n3726.n0 89.977
R5369 a_13419_n3726.n5 a_13419_n3726.n4 77.784
R5370 a_13419_n3726.n6 a_13419_n3726.n5 77.456
R5371 a_13419_n3726.n7 a_13419_n3726.n6 77.456
R5372 a_13419_n3726.n8 a_13419_n3726.n7 75.815
R5373 a_13419_n3726.n3 a_13419_n3726.t3 14.282
R5374 a_13419_n3726.n3 a_13419_n3726.t8 14.282
R5375 a_13419_n3726.n2 a_13419_n3726.t5 14.282
R5376 a_13419_n3726.n2 a_13419_n3726.t6 14.282
R5377 a_13419_n3726.n1 a_13419_n3726.t4 14.282
R5378 a_13419_n3726.n1 a_13419_n3726.t10 14.282
R5379 a_13419_n3726.n0 a_13419_n3726.t7 14.282
R5380 a_13419_n3726.n0 a_13419_n3726.t11 14.282
R5381 a_13419_n3726.t0 a_13419_n3726.n9 14.282
R5382 a_13419_n3726.n9 a_13419_n3726.t2 14.282
R5383 a_307_3697.n2 a_307_3697.t9 214.335
R5384 a_307_3697.t7 a_307_3697.n2 214.335
R5385 a_307_3697.n3 a_307_3697.t7 143.851
R5386 a_307_3697.n3 a_307_3697.t8 135.658
R5387 a_307_3697.n2 a_307_3697.t10 80.333
R5388 a_307_3697.n4 a_307_3697.t6 28.565
R5389 a_307_3697.n4 a_307_3697.t5 28.565
R5390 a_307_3697.n0 a_307_3697.t3 28.565
R5391 a_307_3697.n0 a_307_3697.t2 28.565
R5392 a_307_3697.t0 a_307_3697.n7 28.565
R5393 a_307_3697.n7 a_307_3697.t1 28.565
R5394 a_307_3697.n1 a_307_3697.t4 9.714
R5395 a_307_3697.n1 a_307_3697.n0 1.003
R5396 a_307_3697.n6 a_307_3697.n5 0.833
R5397 a_307_3697.n5 a_307_3697.n4 0.653
R5398 a_307_3697.n7 a_307_3697.n6 0.653
R5399 a_307_3697.n6 a_307_3697.n1 0.341
R5400 a_307_3697.n5 a_307_3697.n3 0.032
R5401 a_20044_n3722.n4 a_20044_n3722.t9 1527.4
R5402 a_20044_n3722.t9 a_20044_n3722.n3 657.379
R5403 a_20044_n3722.n1 a_20044_n3722.n0 258.161
R5404 a_20044_n3722.n7 a_20044_n3722.n6 258.161
R5405 a_20044_n3722.n2 a_20044_n3722.t10 206.421
R5406 a_20044_n3722.t8 a_20044_n3722.n2 206.421
R5407 a_20044_n3722.n4 a_20044_n3722.t8 200.029
R5408 a_20044_n3722.n5 a_20044_n3722.n4 97.614
R5409 a_20044_n3722.n2 a_20044_n3722.t11 80.333
R5410 a_20044_n3722.n6 a_20044_n3722.t6 14.283
R5411 a_20044_n3722.n1 a_20044_n3722.t3 14.283
R5412 a_20044_n3722.n0 a_20044_n3722.t4 14.282
R5413 a_20044_n3722.n0 a_20044_n3722.t5 14.282
R5414 a_20044_n3722.t1 a_20044_n3722.n7 14.282
R5415 a_20044_n3722.n7 a_20044_n3722.t7 14.282
R5416 a_20044_n3722.n3 a_20044_n3722.t2 8.7
R5417 a_20044_n3722.n3 a_20044_n3722.t0 8.7
R5418 a_20044_n3722.n6 a_20044_n3722.n5 4.366
R5419 a_20044_n3722.n5 a_20044_n3722.n1 0.852
R5420 a_19645_n1016.t2 a_19645_n1016.n0 28.568
R5421 a_19645_n1016.n0 a_19645_n1016.n4 185.55
R5422 a_19645_n1016.n4 a_19645_n1016.t1 28.565
R5423 a_19645_n1016.n4 a_19645_n1016.t0 28.565
R5424 a_19645_n1016.n0 a_19645_n1016.n3 1.537
R5425 a_19645_n1016.n3 a_19645_n1016.t3 21.473
R5426 a_19645_n1016.n3 a_19645_n1016.n1 11.712
R5427 a_19645_n1016.n1 a_19645_n1016.t6 408.211
R5428 a_19645_n1016.n1 a_19645_n1016.t7 990.34
R5429 a_19645_n1016.t7 a_19645_n1016.n2 160.666
R5430 a_19645_n1016.n2 a_19645_n1016.t5 286.438
R5431 a_19645_n1016.n2 a_19645_n1016.t4 286.438
R5432 Y[0].n1 Y[0].n0 185.55
R5433 Y[0] Y[0].n2 33.128
R5434 Y[0].n1 Y[0].t2 28.568
R5435 Y[0].n0 Y[0].t1 28.565
R5436 Y[0].n0 Y[0].t0 28.565
R5437 Y[0].n2 Y[0].t3 21.373
R5438 Y[0].n2 Y[0].n1 1.637
R5439 a_19136_n3722.n2 a_19136_n3722.t5 448.382
R5440 a_19136_n3722.n1 a_19136_n3722.t4 286.438
R5441 a_19136_n3722.n1 a_19136_n3722.t6 286.438
R5442 a_19136_n3722.n0 a_19136_n3722.t7 247.69
R5443 a_19136_n3722.n4 a_19136_n3722.n3 182.117
R5444 a_19136_n3722.t5 a_19136_n3722.n1 160.666
R5445 a_19136_n3722.n3 a_19136_n3722.t0 28.568
R5446 a_19136_n3722.n4 a_19136_n3722.t1 28.565
R5447 a_19136_n3722.t2 a_19136_n3722.n4 28.565
R5448 a_19136_n3722.n0 a_19136_n3722.t3 18.127
R5449 a_19136_n3722.n2 a_19136_n3722.n0 4.039
R5450 a_19136_n3722.n3 a_19136_n3722.n2 0.937
R5451 a_19695_n3722.n2 a_19695_n3722.n1 167.433
R5452 a_19695_n3722.n6 a_19695_n3722.n5 167.433
R5453 a_19695_n3722.n2 a_19695_n3722.t3 104.259
R5454 a_19695_n3722.n6 a_19695_n3722.t9 104.259
R5455 a_19695_n3722.n3 a_19695_n3722.n0 89.977
R5456 a_19695_n3722.n7 a_19695_n3722.n4 89.977
R5457 a_19695_n3722.n9 a_19695_n3722.n8 89.977
R5458 a_19695_n3722.n3 a_19695_n3722.n2 77.784
R5459 a_19695_n3722.n8 a_19695_n3722.n3 77.456
R5460 a_19695_n3722.n8 a_19695_n3722.n7 77.456
R5461 a_19695_n3722.n7 a_19695_n3722.n6 75.815
R5462 a_19695_n3722.n1 a_19695_n3722.t4 14.282
R5463 a_19695_n3722.n1 a_19695_n3722.t5 14.282
R5464 a_19695_n3722.n0 a_19695_n3722.t0 14.282
R5465 a_19695_n3722.n0 a_19695_n3722.t1 14.282
R5466 a_19695_n3722.n4 a_19695_n3722.t7 14.282
R5467 a_19695_n3722.n4 a_19695_n3722.t8 14.282
R5468 a_19695_n3722.n5 a_19695_n3722.t10 14.282
R5469 a_19695_n3722.n5 a_19695_n3722.t11 14.282
R5470 a_19695_n3722.t2 a_19695_n3722.n9 14.282
R5471 a_19695_n3722.n9 a_19695_n3722.t6 14.282
R5472 a_6811_3260.t2 a_6811_3260.n0 28.565
R5473 a_6811_3260.n0 a_6811_3260.t0 28.565
R5474 a_6811_3260.n0 a_6811_3260.n1 192.754
R5475 a_6811_3260.n1 a_6811_3260.t1 28.568
R5476 a_6811_3260.n1 a_6811_3260.n2 1.123
R5477 a_6811_3260.n2 a_6811_3260.n3 27.985
R5478 a_6811_3260.n3 a_6811_3260.t6 615.911
R5479 a_6811_3260.n3 a_6811_3260.t7 867.497
R5480 a_6811_3260.t7 a_6811_3260.n4 160.666
R5481 a_6811_3260.n4 a_6811_3260.t5 286.438
R5482 a_6811_3260.n4 a_6811_3260.t4 286.438
R5483 a_6811_3260.n2 a_6811_3260.t3 18.726
R5484 a_23188_n3722.n4 a_23188_n3722.t8 1527.4
R5485 a_23188_n3722.t8 a_23188_n3722.n3 657.379
R5486 a_23188_n3722.n1 a_23188_n3722.n0 258.161
R5487 a_23188_n3722.n7 a_23188_n3722.n6 258.161
R5488 a_23188_n3722.n2 a_23188_n3722.t9 206.421
R5489 a_23188_n3722.t11 a_23188_n3722.n2 206.421
R5490 a_23188_n3722.n4 a_23188_n3722.t11 200.029
R5491 a_23188_n3722.n5 a_23188_n3722.n4 97.614
R5492 a_23188_n3722.n2 a_23188_n3722.t10 80.333
R5493 a_23188_n3722.n6 a_23188_n3722.t6 14.283
R5494 a_23188_n3722.n1 a_23188_n3722.t1 14.283
R5495 a_23188_n3722.n0 a_23188_n3722.t2 14.282
R5496 a_23188_n3722.n0 a_23188_n3722.t3 14.282
R5497 a_23188_n3722.n7 a_23188_n3722.t4 14.282
R5498 a_23188_n3722.t0 a_23188_n3722.n7 14.282
R5499 a_23188_n3722.n3 a_23188_n3722.t7 8.7
R5500 a_23188_n3722.n3 a_23188_n3722.t5 8.7
R5501 a_23188_n3722.n6 a_23188_n3722.n5 4.366
R5502 a_23188_n3722.n5 a_23188_n3722.n1 0.852
R5503 a_6607_n7362.n3 a_6607_n7362.n1 267.767
R5504 a_6607_n7362.n7 a_6607_n7362.t2 16.058
R5505 a_6607_n7362.t0 a_6607_n7362.n9 16.058
R5506 a_6607_n7362.n2 a_6607_n7362.t6 14.282
R5507 a_6607_n7362.n2 a_6607_n7362.t9 14.282
R5508 a_6607_n7362.n1 a_6607_n7362.t4 14.282
R5509 a_6607_n7362.n1 a_6607_n7362.t5 14.282
R5510 a_6607_n7362.n4 a_6607_n7362.t10 14.282
R5511 a_6607_n7362.n4 a_6607_n7362.t11 14.282
R5512 a_6607_n7362.n6 a_6607_n7362.t7 14.282
R5513 a_6607_n7362.n6 a_6607_n7362.t3 14.282
R5514 a_6607_n7362.n0 a_6607_n7362.t1 14.282
R5515 a_6607_n7362.n0 a_6607_n7362.t8 14.282
R5516 a_6607_n7362.n5 a_6607_n7362.n4 1.511
R5517 a_6607_n7362.n7 a_6607_n7362.n6 0.999
R5518 a_6607_n7362.n9 a_6607_n7362.n0 0.999
R5519 a_6607_n7362.n5 a_6607_n7362.n3 0.669
R5520 a_6607_n7362.n8 a_6607_n7362.n7 0.575
R5521 a_6607_n7362.n8 a_6607_n7362.n5 0.227
R5522 a_6607_n7362.n9 a_6607_n7362.n8 0.2
R5523 a_6607_n7362.n3 a_6607_n7362.n2 0.001
R5524 a_19705_n990.n3 a_19705_n990.n2 167.433
R5525 a_19705_n990.n7 a_19705_n990.n6 167.433
R5526 a_19705_n990.n3 a_19705_n990.t7 104.259
R5527 a_19705_n990.n7 a_19705_n990.t10 104.259
R5528 a_19705_n990.n4 a_19705_n990.n1 89.977
R5529 a_19705_n990.n5 a_19705_n990.n0 89.977
R5530 a_19705_n990.n9 a_19705_n990.n8 89.977
R5531 a_19705_n990.n4 a_19705_n990.n3 77.784
R5532 a_19705_n990.n5 a_19705_n990.n4 77.456
R5533 a_19705_n990.n8 a_19705_n990.n5 77.456
R5534 a_19705_n990.n8 a_19705_n990.n7 75.815
R5535 a_19705_n990.n2 a_19705_n990.t8 14.282
R5536 a_19705_n990.n2 a_19705_n990.t6 14.282
R5537 a_19705_n990.n1 a_19705_n990.t3 14.282
R5538 a_19705_n990.n1 a_19705_n990.t5 14.282
R5539 a_19705_n990.n0 a_19705_n990.t4 14.282
R5540 a_19705_n990.n0 a_19705_n990.t0 14.282
R5541 a_19705_n990.n6 a_19705_n990.t9 14.282
R5542 a_19705_n990.n6 a_19705_n990.t11 14.282
R5543 a_19705_n990.t2 a_19705_n990.n9 14.282
R5544 a_19705_n990.n9 a_19705_n990.t1 14.282
R5545 Y[3].n1 Y[3].n0 185.55
R5546 Y[3].n1 Y[3].t2 28.568
R5547 Y[3].n0 Y[3].t0 28.565
R5548 Y[3].n0 Y[3].t1 28.565
R5549 Y[3].n2 Y[3].t3 21.373
R5550 Y[3] Y[3].n2 20.004
R5551 Y[3].n2 Y[3].n1 1.637
R5552 a_19705_1744.n3 a_19705_1744.n2 167.433
R5553 a_19705_1744.n7 a_19705_1744.n6 167.433
R5554 a_19705_1744.n3 a_19705_1744.t10 104.259
R5555 a_19705_1744.n7 a_19705_1744.t4 104.259
R5556 a_19705_1744.n4 a_19705_1744.n1 89.977
R5557 a_19705_1744.n5 a_19705_1744.n0 89.977
R5558 a_19705_1744.n9 a_19705_1744.n8 89.977
R5559 a_19705_1744.n4 a_19705_1744.n3 77.784
R5560 a_19705_1744.n5 a_19705_1744.n4 77.456
R5561 a_19705_1744.n8 a_19705_1744.n5 77.456
R5562 a_19705_1744.n8 a_19705_1744.n7 75.815
R5563 a_19705_1744.n2 a_19705_1744.t11 14.282
R5564 a_19705_1744.n2 a_19705_1744.t9 14.282
R5565 a_19705_1744.n1 a_19705_1744.t0 14.282
R5566 a_19705_1744.n1 a_19705_1744.t2 14.282
R5567 a_19705_1744.n0 a_19705_1744.t1 14.282
R5568 a_19705_1744.n0 a_19705_1744.t7 14.282
R5569 a_19705_1744.n6 a_19705_1744.t3 14.282
R5570 a_19705_1744.n6 a_19705_1744.t5 14.282
R5571 a_19705_1744.n9 a_19705_1744.t8 14.282
R5572 a_19705_1744.t6 a_19705_1744.n9 14.282
R5573 a_10576_1744.n4 a_10576_1744.t8 1527.4
R5574 a_10576_1744.t8 a_10576_1744.n3 657.379
R5575 a_10576_1744.n1 a_10576_1744.n0 258.161
R5576 a_10576_1744.n7 a_10576_1744.n6 258.161
R5577 a_10576_1744.n2 a_10576_1744.t10 206.421
R5578 a_10576_1744.t9 a_10576_1744.n2 206.421
R5579 a_10576_1744.n4 a_10576_1744.t9 200.029
R5580 a_10576_1744.n5 a_10576_1744.n4 97.614
R5581 a_10576_1744.n2 a_10576_1744.t11 80.333
R5582 a_10576_1744.n6 a_10576_1744.t1 14.283
R5583 a_10576_1744.n1 a_10576_1744.t5 14.283
R5584 a_10576_1744.n0 a_10576_1744.t7 14.282
R5585 a_10576_1744.n0 a_10576_1744.t6 14.282
R5586 a_10576_1744.n7 a_10576_1744.t0 14.282
R5587 a_10576_1744.t2 a_10576_1744.n7 14.282
R5588 a_10576_1744.n3 a_10576_1744.t3 8.7
R5589 a_10576_1744.n3 a_10576_1744.t4 8.7
R5590 a_10576_1744.n6 a_10576_1744.n5 4.366
R5591 a_10576_1744.n5 a_10576_1744.n1 0.852
R5592 a_11101_n1475.t2 a_11101_n1475.n0 28.568
R5593 a_11101_n1475.n0 a_11101_n1475.n4 185.55
R5594 a_11101_n1475.n4 a_11101_n1475.t1 28.565
R5595 a_11101_n1475.n4 a_11101_n1475.t0 28.565
R5596 a_11101_n1475.n0 a_11101_n1475.n3 1.64
R5597 a_11101_n1475.n3 a_11101_n1475.t3 21.373
R5598 a_11101_n1475.n3 a_11101_n1475.n1 25.769
R5599 a_11101_n1475.n1 a_11101_n1475.t5 615.911
R5600 a_11101_n1475.n1 a_11101_n1475.t4 867.497
R5601 a_11101_n1475.t4 a_11101_n1475.n2 160.666
R5602 a_11101_n1475.n2 a_11101_n1475.t7 286.438
R5603 a_11101_n1475.n2 a_11101_n1475.t6 286.438
R5604 a_6180_n6669.n2 a_6180_n6669.t7 318.922
R5605 a_6180_n6669.n1 a_6180_n6669.t6 273.935
R5606 a_6180_n6669.n1 a_6180_n6669.t4 273.935
R5607 a_6180_n6669.n2 a_6180_n6669.t5 269.116
R5608 a_6180_n6669.n4 a_6180_n6669.n0 193.227
R5609 a_6180_n6669.t7 a_6180_n6669.n1 179.142
R5610 a_6180_n6669.n3 a_6180_n6669.n2 106.999
R5611 a_6180_n6669.t2 a_6180_n6669.n4 28.568
R5612 a_6180_n6669.n0 a_6180_n6669.t0 28.565
R5613 a_6180_n6669.n0 a_6180_n6669.t1 28.565
R5614 a_6180_n6669.n3 a_6180_n6669.t3 18.149
R5615 a_6180_n6669.n4 a_6180_n6669.n3 3.726
R5616 a_6524_n990.n2 a_6524_n990.t7 448.382
R5617 a_6524_n990.n1 a_6524_n990.t6 286.438
R5618 a_6524_n990.n1 a_6524_n990.t5 286.438
R5619 a_6524_n990.n0 a_6524_n990.t4 247.69
R5620 a_6524_n990.n4 a_6524_n990.n3 182.117
R5621 a_6524_n990.t7 a_6524_n990.n1 160.666
R5622 a_6524_n990.n3 a_6524_n990.t1 28.568
R5623 a_6524_n990.t2 a_6524_n990.n4 28.565
R5624 a_6524_n990.n4 a_6524_n990.t0 28.565
R5625 a_6524_n990.n0 a_6524_n990.t3 18.127
R5626 a_6524_n990.n2 a_6524_n990.n0 4.039
R5627 a_6524_n990.n3 a_6524_n990.n2 0.937
R5628 a_11205_3262.t2 a_11205_3262.n0 28.565
R5629 a_11205_3262.n0 a_11205_3262.t0 28.565
R5630 a_11205_3262.n0 a_11205_3262.n1 192.754
R5631 a_11205_3262.n1 a_11205_3262.t1 28.568
R5632 a_11205_3262.n1 a_11205_3262.n2 1.123
R5633 a_11205_3262.n2 a_11205_3262.n3 37.906
R5634 a_11205_3262.n3 a_11205_3262.t6 615.911
R5635 a_11205_3262.n3 a_11205_3262.t7 867.497
R5636 a_11205_3262.t7 a_11205_3262.n4 160.666
R5637 a_11205_3262.n4 a_11205_3262.t4 286.438
R5638 a_11205_3262.n4 a_11205_3262.t5 286.438
R5639 a_11205_3262.n2 a_11205_3262.t3 18.726
R5640 a_6524_1744.n2 a_6524_1744.t7 448.382
R5641 a_6524_1744.n1 a_6524_1744.t6 286.438
R5642 a_6524_1744.n1 a_6524_1744.t4 286.438
R5643 a_6524_1744.n0 a_6524_1744.t5 247.69
R5644 a_6524_1744.n4 a_6524_1744.n3 182.117
R5645 a_6524_1744.t7 a_6524_1744.n1 160.666
R5646 a_6524_1744.n3 a_6524_1744.t1 28.568
R5647 a_6524_1744.t2 a_6524_1744.n4 28.565
R5648 a_6524_1744.n4 a_6524_1744.t0 28.565
R5649 a_6524_1744.n0 a_6524_1744.t3 18.127
R5650 a_6524_1744.n2 a_6524_1744.n0 4.039
R5651 a_6524_1744.n3 a_6524_1744.n2 0.937
R5652 a_16573_1740.n2 a_16573_1740.n1 167.433
R5653 a_16573_1740.n6 a_16573_1740.n5 167.433
R5654 a_16573_1740.n2 a_16573_1740.t10 104.259
R5655 a_16573_1740.n6 a_16573_1740.t6 104.259
R5656 a_16573_1740.n3 a_16573_1740.n0 89.977
R5657 a_16573_1740.n7 a_16573_1740.n4 89.977
R5658 a_16573_1740.n9 a_16573_1740.n8 89.977
R5659 a_16573_1740.n3 a_16573_1740.n2 77.784
R5660 a_16573_1740.n8 a_16573_1740.n3 77.456
R5661 a_16573_1740.n8 a_16573_1740.n7 77.456
R5662 a_16573_1740.n7 a_16573_1740.n6 75.815
R5663 a_16573_1740.n1 a_16573_1740.t8 14.282
R5664 a_16573_1740.n1 a_16573_1740.t9 14.282
R5665 a_16573_1740.n0 a_16573_1740.t4 14.282
R5666 a_16573_1740.n0 a_16573_1740.t3 14.282
R5667 a_16573_1740.n4 a_16573_1740.t2 14.282
R5668 a_16573_1740.n4 a_16573_1740.t1 14.282
R5669 a_16573_1740.n5 a_16573_1740.t7 14.282
R5670 a_16573_1740.n5 a_16573_1740.t11 14.282
R5671 a_16573_1740.n9 a_16573_1740.t5 14.282
R5672 a_16573_1740.t0 a_16573_1740.n9 14.282
R5673 a_16922_1740.n4 a_16922_1740.t8 1527.4
R5674 a_16922_1740.t8 a_16922_1740.n3 657.379
R5675 a_16922_1740.n1 a_16922_1740.n0 258.161
R5676 a_16922_1740.n7 a_16922_1740.n6 258.161
R5677 a_16922_1740.n2 a_16922_1740.t11 206.421
R5678 a_16922_1740.t10 a_16922_1740.n2 206.421
R5679 a_16922_1740.n4 a_16922_1740.t10 200.029
R5680 a_16922_1740.n5 a_16922_1740.n4 97.614
R5681 a_16922_1740.n2 a_16922_1740.t9 80.333
R5682 a_16922_1740.n6 a_16922_1740.t2 14.283
R5683 a_16922_1740.n1 a_16922_1740.t5 14.283
R5684 a_16922_1740.n0 a_16922_1740.t6 14.282
R5685 a_16922_1740.n0 a_16922_1740.t7 14.282
R5686 a_16922_1740.n7 a_16922_1740.t1 14.282
R5687 a_16922_1740.t3 a_16922_1740.n7 14.282
R5688 a_16922_1740.n3 a_16922_1740.t0 8.7
R5689 a_16922_1740.n3 a_16922_1740.t4 8.7
R5690 a_16922_1740.n6 a_16922_1740.n5 4.366
R5691 a_16922_1740.n5 a_16922_1740.n1 0.852
R5692 a_10862_n7360.n7 a_10862_n7360.n1 1617.25
R5693 a_10862_n7360.n1 a_10862_n7360.t9 867.497
R5694 a_10862_n7360.n1 a_10862_n7360.t10 615.911
R5695 a_10862_n7360.n0 a_10862_n7360.t11 286.438
R5696 a_10862_n7360.n0 a_10862_n7360.t8 286.438
R5697 a_10862_n7360.t9 a_10862_n7360.n0 160.666
R5698 a_10862_n7360.n5 a_10862_n7360.n3 157.665
R5699 a_10862_n7360.n5 a_10862_n7360.n4 122.999
R5700 a_10862_n7360.n8 a_10862_n7360.n7 90.436
R5701 a_10862_n7360.n6 a_10862_n7360.n2 90.416
R5702 a_10862_n7360.n7 a_10862_n7360.n6 74.302
R5703 a_10862_n7360.n6 a_10862_n7360.n5 50.575
R5704 a_10862_n7360.n2 a_10862_n7360.t1 14.282
R5705 a_10862_n7360.n2 a_10862_n7360.t6 14.282
R5706 a_10862_n7360.n4 a_10862_n7360.t5 14.282
R5707 a_10862_n7360.n4 a_10862_n7360.t4 14.282
R5708 a_10862_n7360.t0 a_10862_n7360.n8 14.282
R5709 a_10862_n7360.n8 a_10862_n7360.t2 14.282
R5710 a_10862_n7360.n3 a_10862_n7360.t3 8.7
R5711 a_10862_n7360.n3 a_10862_n7360.t7 8.7
R5712 a_16563_n3726.n4 a_16563_n3726.n3 167.433
R5713 a_16563_n3726.n9 a_16563_n3726.n8 167.433
R5714 a_16563_n3726.n4 a_16563_n3726.t7 104.259
R5715 a_16563_n3726.t6 a_16563_n3726.n9 104.259
R5716 a_16563_n3726.n5 a_16563_n3726.n2 89.977
R5717 a_16563_n3726.n6 a_16563_n3726.n1 89.977
R5718 a_16563_n3726.n7 a_16563_n3726.n0 89.977
R5719 a_16563_n3726.n5 a_16563_n3726.n4 77.784
R5720 a_16563_n3726.n6 a_16563_n3726.n5 77.456
R5721 a_16563_n3726.n7 a_16563_n3726.n6 77.456
R5722 a_16563_n3726.n9 a_16563_n3726.n7 75.815
R5723 a_16563_n3726.n3 a_16563_n3726.t9 14.282
R5724 a_16563_n3726.n3 a_16563_n3726.t8 14.282
R5725 a_16563_n3726.n2 a_16563_n3726.t0 14.282
R5726 a_16563_n3726.n2 a_16563_n3726.t1 14.282
R5727 a_16563_n3726.n1 a_16563_n3726.t2 14.282
R5728 a_16563_n3726.n1 a_16563_n3726.t3 14.282
R5729 a_16563_n3726.n0 a_16563_n3726.t4 14.282
R5730 a_16563_n3726.n0 a_16563_n3726.t5 14.282
R5731 a_16563_n3726.n8 a_16563_n3726.t11 14.282
R5732 a_16563_n3726.n8 a_16563_n3726.t10 14.282
R5733 a_9088_n7388.n1 a_9088_n7388.t5 318.922
R5734 a_9088_n7388.n0 a_9088_n7388.t7 274.739
R5735 a_9088_n7388.n0 a_9088_n7388.t6 274.739
R5736 a_9088_n7388.n1 a_9088_n7388.t4 269.116
R5737 a_9088_n7388.t5 a_9088_n7388.n0 179.946
R5738 a_9088_n7388.n2 a_9088_n7388.n1 107.263
R5739 a_9088_n7388.n3 a_9088_n7388.t0 29.444
R5740 a_9088_n7388.n4 a_9088_n7388.t1 28.565
R5741 a_9088_n7388.t2 a_9088_n7388.n4 28.565
R5742 a_9088_n7388.n2 a_9088_n7388.t3 18.145
R5743 a_9088_n7388.n3 a_9088_n7388.n2 2.878
R5744 a_9088_n7388.n4 a_9088_n7388.n3 0.764
R5745 a_8794_n8094.t0 a_8794_n8094.t1 380.209
R5746 a_16573_n994.n3 a_16573_n994.n2 167.433
R5747 a_16573_n994.n7 a_16573_n994.n6 167.433
R5748 a_16573_n994.n3 a_16573_n994.t6 104.259
R5749 a_16573_n994.n7 a_16573_n994.t7 104.259
R5750 a_16573_n994.n4 a_16573_n994.n1 89.977
R5751 a_16573_n994.n5 a_16573_n994.n0 89.977
R5752 a_16573_n994.n9 a_16573_n994.n8 89.977
R5753 a_16573_n994.n4 a_16573_n994.n3 77.784
R5754 a_16573_n994.n5 a_16573_n994.n4 77.456
R5755 a_16573_n994.n8 a_16573_n994.n5 77.456
R5756 a_16573_n994.n8 a_16573_n994.n7 75.815
R5757 a_16573_n994.n2 a_16573_n994.t11 14.282
R5758 a_16573_n994.n2 a_16573_n994.t10 14.282
R5759 a_16573_n994.n1 a_16573_n994.t4 14.282
R5760 a_16573_n994.n1 a_16573_n994.t3 14.282
R5761 a_16573_n994.n0 a_16573_n994.t5 14.282
R5762 a_16573_n994.n0 a_16573_n994.t2 14.282
R5763 a_16573_n994.n6 a_16573_n994.t9 14.282
R5764 a_16573_n994.n6 a_16573_n994.t8 14.282
R5765 a_16573_n994.n9 a_16573_n994.t1 14.282
R5766 a_16573_n994.t0 a_16573_n994.n9 14.282
R5767 a_16922_n994.n2 a_16922_n994.t8 1527.4
R5768 a_16922_n994.t8 a_16922_n994.n1 657.379
R5769 a_16922_n994.n4 a_16922_n994.n3 258.161
R5770 a_16922_n994.n7 a_16922_n994.n6 258.161
R5771 a_16922_n994.n0 a_16922_n994.t11 206.421
R5772 a_16922_n994.t10 a_16922_n994.n0 206.421
R5773 a_16922_n994.n2 a_16922_n994.t10 200.029
R5774 a_16922_n994.n5 a_16922_n994.n2 97.614
R5775 a_16922_n994.n0 a_16922_n994.t9 80.333
R5776 a_16922_n994.n4 a_16922_n994.t2 14.283
R5777 a_16922_n994.n6 a_16922_n994.t7 14.283
R5778 a_16922_n994.n3 a_16922_n994.t1 14.282
R5779 a_16922_n994.n3 a_16922_n994.t3 14.282
R5780 a_16922_n994.n7 a_16922_n994.t6 14.282
R5781 a_16922_n994.t5 a_16922_n994.n7 14.282
R5782 a_16922_n994.n1 a_16922_n994.t0 8.7
R5783 a_16922_n994.n1 a_16922_n994.t4 8.7
R5784 a_16922_n994.n5 a_16922_n994.n4 4.366
R5785 a_16922_n994.n6 a_16922_n994.n5 0.852
R5786 a_10317_n6667.n1 a_10317_n6667.t5 318.922
R5787 a_10317_n6667.n0 a_10317_n6667.t4 273.935
R5788 a_10317_n6667.n0 a_10317_n6667.t7 273.935
R5789 a_10317_n6667.n1 a_10317_n6667.t6 269.116
R5790 a_10317_n6667.n4 a_10317_n6667.n3 193.227
R5791 a_10317_n6667.t5 a_10317_n6667.n0 179.142
R5792 a_10317_n6667.n2 a_10317_n6667.n1 106.999
R5793 a_10317_n6667.n3 a_10317_n6667.t1 28.568
R5794 a_10317_n6667.t2 a_10317_n6667.n4 28.565
R5795 a_10317_n6667.n4 a_10317_n6667.t0 28.565
R5796 a_10317_n6667.n2 a_10317_n6667.t3 18.149
R5797 a_10317_n6667.n3 a_10317_n6667.n2 3.726
R5798 a_10744_n7360.n2 a_10744_n7360.n0 267.767
R5799 a_10744_n7360.n6 a_10744_n7360.t11 16.058
R5800 a_10744_n7360.n8 a_10744_n7360.t0 16.058
R5801 a_10744_n7360.n1 a_10744_n7360.t4 14.282
R5802 a_10744_n7360.n1 a_10744_n7360.t8 14.282
R5803 a_10744_n7360.n0 a_10744_n7360.t5 14.282
R5804 a_10744_n7360.n0 a_10744_n7360.t3 14.282
R5805 a_10744_n7360.n3 a_10744_n7360.t6 14.282
R5806 a_10744_n7360.n3 a_10744_n7360.t7 14.282
R5807 a_10744_n7360.n5 a_10744_n7360.t9 14.282
R5808 a_10744_n7360.n5 a_10744_n7360.t10 14.282
R5809 a_10744_n7360.n9 a_10744_n7360.t1 14.282
R5810 a_10744_n7360.t2 a_10744_n7360.n9 14.282
R5811 a_10744_n7360.n4 a_10744_n7360.n3 1.511
R5812 a_10744_n7360.n6 a_10744_n7360.n5 0.999
R5813 a_10744_n7360.n9 a_10744_n7360.n8 0.999
R5814 a_10744_n7360.n4 a_10744_n7360.n2 0.669
R5815 a_10744_n7360.n7 a_10744_n7360.n6 0.575
R5816 a_10744_n7360.n7 a_10744_n7360.n4 0.227
R5817 a_10744_n7360.n8 a_10744_n7360.n7 0.2
R5818 a_10744_n7360.n2 a_10744_n7360.n1 0.001
R5819 a_17447_n1479.n0 a_17447_n1479.t0 28.565
R5820 a_17447_n1479.t2 a_17447_n1479.n0 28.565
R5821 a_17447_n1479.n0 a_17447_n1479.n1 185.55
R5822 a_17447_n1479.n1 a_17447_n1479.t1 28.568
R5823 a_17447_n1479.n1 a_17447_n1479.n4 1.628
R5824 a_17447_n1479.n4 a_17447_n1479.n2 25.436
R5825 a_17447_n1479.n2 a_17447_n1479.t5 615.911
R5826 a_17447_n1479.n2 a_17447_n1479.t6 867.497
R5827 a_17447_n1479.t6 a_17447_n1479.n3 160.666
R5828 a_17447_n1479.n3 a_17447_n1479.t7 286.438
R5829 a_17447_n1479.n3 a_17447_n1479.t4 286.438
R5830 a_17447_n1479.n4 a_17447_n1479.t3 22.074
R5831 a_18966_3696.t8 a_18966_3696.n2 406.978
R5832 a_18966_3696.n1 a_18966_3696.t6 207.38
R5833 a_18966_3696.n3 a_18966_3696.t8 136.943
R5834 a_18966_3696.n2 a_18966_3696.n1 112.003
R5835 a_18966_3696.n1 a_18966_3696.t7 80.333
R5836 a_18966_3696.n2 a_18966_3696.t5 80.333
R5837 a_18966_3696.n0 a_18966_3696.t0 17.4
R5838 a_18966_3696.n0 a_18966_3696.t2 17.4
R5839 a_18966_3696.n4 a_18966_3696.t3 15.036
R5840 a_18966_3696.n5 a_18966_3696.t4 14.282
R5841 a_18966_3696.t1 a_18966_3696.n5 14.282
R5842 a_18966_3696.n5 a_18966_3696.n4 1.654
R5843 a_18966_3696.n3 a_18966_3696.n0 0.672
R5844 a_18966_3696.n4 a_18966_3696.n3 0.665
R5845 a_19084_3696.n1 a_19084_3696.t1 14.282
R5846 a_19084_3696.n1 a_19084_3696.t5 14.282
R5847 a_19084_3696.n0 a_19084_3696.t4 14.282
R5848 a_19084_3696.n0 a_19084_3696.t3 14.282
R5849 a_19084_3696.n3 a_19084_3696.t0 14.282
R5850 a_19084_3696.t2 a_19084_3696.n3 14.282
R5851 a_19084_3696.n2 a_19084_3696.n0 2.538
R5852 a_19084_3696.n3 a_19084_3696.n2 2.375
R5853 a_19084_3696.n2 a_19084_3696.n1 0.001
R5854 a_6514_n3722.n2 a_6514_n3722.t6 448.382
R5855 a_6514_n3722.n1 a_6514_n3722.t4 286.438
R5856 a_6514_n3722.n1 a_6514_n3722.t7 286.438
R5857 a_6514_n3722.n0 a_6514_n3722.t5 247.69
R5858 a_6514_n3722.n4 a_6514_n3722.n3 182.117
R5859 a_6514_n3722.t6 a_6514_n3722.n1 160.666
R5860 a_6514_n3722.n3 a_6514_n3722.t1 28.568
R5861 a_6514_n3722.t2 a_6514_n3722.n4 28.565
R5862 a_6514_n3722.n4 a_6514_n3722.t0 28.565
R5863 a_6514_n3722.n0 a_6514_n3722.t3 18.127
R5864 a_6514_n3722.n2 a_6514_n3722.n0 4.039
R5865 a_6514_n3722.n3 a_6514_n3722.n2 0.937
R5866 a_1392_n2327.t0 a_1392_n2327.t1 17.4
R5867 a_2882_n7388.n1 a_2882_n7388.t6 318.922
R5868 a_2882_n7388.n0 a_2882_n7388.t4 274.739
R5869 a_2882_n7388.n0 a_2882_n7388.t7 274.739
R5870 a_2882_n7388.n1 a_2882_n7388.t5 269.116
R5871 a_2882_n7388.t6 a_2882_n7388.n0 179.946
R5872 a_2882_n7388.n2 a_2882_n7388.n1 107.263
R5873 a_2882_n7388.n3 a_2882_n7388.t0 29.444
R5874 a_2882_n7388.n4 a_2882_n7388.t1 28.565
R5875 a_2882_n7388.t2 a_2882_n7388.n4 28.565
R5876 a_2882_n7388.n2 a_2882_n7388.t3 18.145
R5877 a_2882_n7388.n3 a_2882_n7388.n2 2.878
R5878 a_2882_n7388.n4 a_2882_n7388.n3 0.764
R5879 a_7658_n5055.t0 a_7658_n5055.t1 17.4
R5880 a_16513_1714.t2 a_16513_1714.n0 28.568
R5881 a_16513_1714.n0 a_16513_1714.n2 97.311
R5882 a_16513_1714.n2 a_16513_1714.n3 903.039
R5883 a_16513_1714.n3 a_16513_1714.t4 408.211
R5884 a_16513_1714.n3 a_16513_1714.t5 990.34
R5885 a_16513_1714.t5 a_16513_1714.n4 160.666
R5886 a_16513_1714.n4 a_16513_1714.t7 286.438
R5887 a_16513_1714.n4 a_16513_1714.t6 286.438
R5888 a_16513_1714.n2 a_16513_1714.n1 94.754
R5889 a_16513_1714.n1 a_16513_1714.t0 28.565
R5890 a_16513_1714.n1 a_16513_1714.t1 28.565
R5891 a_16513_1714.n0 a_16513_1714.t3 17.64
R5892 a_797_n3726.n4 a_797_n3726.n3 167.433
R5893 a_797_n3726.n9 a_797_n3726.n8 167.433
R5894 a_797_n3726.n8 a_797_n3726.t0 104.259
R5895 a_797_n3726.n4 a_797_n3726.t9 104.259
R5896 a_797_n3726.n7 a_797_n3726.n0 89.977
R5897 a_797_n3726.n6 a_797_n3726.n1 89.977
R5898 a_797_n3726.n5 a_797_n3726.n2 89.977
R5899 a_797_n3726.n8 a_797_n3726.n7 77.784
R5900 a_797_n3726.n7 a_797_n3726.n6 77.456
R5901 a_797_n3726.n6 a_797_n3726.n5 77.456
R5902 a_797_n3726.n5 a_797_n3726.n4 75.815
R5903 a_797_n3726.n0 a_797_n3726.t3 14.282
R5904 a_797_n3726.n0 a_797_n3726.t4 14.282
R5905 a_797_n3726.n1 a_797_n3726.t5 14.282
R5906 a_797_n3726.n1 a_797_n3726.t6 14.282
R5907 a_797_n3726.n2 a_797_n3726.t7 14.282
R5908 a_797_n3726.n2 a_797_n3726.t8 14.282
R5909 a_797_n3726.n3 a_797_n3726.t10 14.282
R5910 a_797_n3726.n3 a_797_n3726.t11 14.282
R5911 a_797_n3726.n9 a_797_n3726.t1 14.282
R5912 a_797_n3726.t2 a_797_n3726.n9 14.282
R5913 a_10157_n3748.t2 a_10157_n3748.n0 28.568
R5914 a_10157_n3748.n0 a_10157_n3748.n4 197.272
R5915 a_10157_n3748.n4 a_10157_n3748.t1 28.565
R5916 a_10157_n3748.n4 a_10157_n3748.t0 28.565
R5917 a_10157_n3748.n0 a_10157_n3748.n1 0.459
R5918 a_10157_n3748.n1 a_10157_n3748.n2 32.171
R5919 a_10157_n3748.n2 a_10157_n3748.t7 408.211
R5920 a_10157_n3748.n2 a_10157_n3748.t5 990.34
R5921 a_10157_n3748.t5 a_10157_n3748.n3 160.666
R5922 a_10157_n3748.n3 a_10157_n3748.t6 286.438
R5923 a_10157_n3748.n3 a_10157_n3748.t4 286.438
R5924 a_10157_n3748.n1 a_10157_n3748.t3 18.103
R5925 B[0].t13 B[0].t5 802.481
R5926 B[0].n3 B[0].n1 653.738
R5927 B[0].n8 B[0].n7 592.056
R5928 B[0].t10 B[0].t6 415.315
R5929 B[0].t1 B[0].n5 313.873
R5930 B[0].n7 B[0].t14 294.986
R5931 B[0].n0 B[0].t15 284.688
R5932 B[0].n4 B[0].t4 272.288
R5933 B[0].n3 B[0].t10 218.406
R5934 B[0].n2 B[0].t7 214.335
R5935 B[0].t6 B[0].n2 214.335
R5936 B[0].n8 B[0].t2 204.68
R5937 B[0].n1 B[0].t13 192.799
R5938 B[0].n6 B[0].t1 190.152
R5939 B[0].n6 B[0].t3 190.152
R5940 B[0].n0 B[0].t8 160.666
R5941 B[0].n4 B[0].t9 160.666
R5942 B[0].n5 B[0].t11 160.666
R5943 B[0].n7 B[0].t0 110.859
R5944 B[0].n5 B[0].n4 96.129
R5945 B[0].n1 B[0].n0 91.889
R5946 B[0].n2 B[0].t12 80.333
R5947 B[0].t2 B[0].n6 80.333
R5948 B[0].n9 B[0].n8 49.449
R5949 B[0] B[0].n9 1.812
R5950 B[0].n9 B[0].n3 0.641
R5951 a_12870_1740.n2 a_12870_1740.t5 448.382
R5952 a_12870_1740.n1 a_12870_1740.t7 286.438
R5953 a_12870_1740.n1 a_12870_1740.t6 286.438
R5954 a_12870_1740.n0 a_12870_1740.t4 247.69
R5955 a_12870_1740.n4 a_12870_1740.n3 182.117
R5956 a_12870_1740.t5 a_12870_1740.n1 160.666
R5957 a_12870_1740.n3 a_12870_1740.t1 28.568
R5958 a_12870_1740.t2 a_12870_1740.n4 28.565
R5959 a_12870_1740.n4 a_12870_1740.t0 28.565
R5960 a_12870_1740.n0 a_12870_1740.t3 18.127
R5961 a_12870_1740.n2 a_12870_1740.n0 4.039
R5962 a_12870_1740.n3 a_12870_1740.n2 0.937
R5963 a_23424_n5055.t0 a_23424_n5055.t1 17.4
R5964 a_4938_3062.t0 a_4938_3062.t1 17.4
R5965 a_14004_n5059.t0 a_14004_n5059.t1 17.4
R5966 a_8676_n7362.n2 a_8676_n7362.n0 267.767
R5967 a_8676_n7362.n6 a_8676_n7362.t10 16.058
R5968 a_8676_n7362.n8 a_8676_n7362.t1 16.058
R5969 a_8676_n7362.n1 a_8676_n7362.t5 14.282
R5970 a_8676_n7362.n1 a_8676_n7362.t8 14.282
R5971 a_8676_n7362.n0 a_8676_n7362.t3 14.282
R5972 a_8676_n7362.n0 a_8676_n7362.t4 14.282
R5973 a_8676_n7362.n3 a_8676_n7362.t7 14.282
R5974 a_8676_n7362.n3 a_8676_n7362.t6 14.282
R5975 a_8676_n7362.n5 a_8676_n7362.t9 14.282
R5976 a_8676_n7362.n5 a_8676_n7362.t11 14.282
R5977 a_8676_n7362.n9 a_8676_n7362.t2 14.282
R5978 a_8676_n7362.t0 a_8676_n7362.n9 14.282
R5979 a_8676_n7362.n4 a_8676_n7362.n3 1.511
R5980 a_8676_n7362.n6 a_8676_n7362.n5 0.999
R5981 a_8676_n7362.n9 a_8676_n7362.n8 0.999
R5982 a_8676_n7362.n4 a_8676_n7362.n2 0.669
R5983 a_8676_n7362.n7 a_8676_n7362.n6 0.575
R5984 a_8676_n7362.n7 a_8676_n7362.n4 0.227
R5985 a_8676_n7362.n8 a_8676_n7362.n7 0.2
R5986 a_8676_n7362.n2 a_8676_n7362.n1 0.001
R5987 a_12870_n994.n2 a_12870_n994.t5 448.382
R5988 a_12870_n994.n1 a_12870_n994.t7 286.438
R5989 a_12870_n994.n1 a_12870_n994.t6 286.438
R5990 a_12870_n994.n0 a_12870_n994.t4 247.69
R5991 a_12870_n994.n4 a_12870_n994.n3 182.117
R5992 a_12870_n994.t5 a_12870_n994.n1 160.666
R5993 a_12870_n994.n3 a_12870_n994.t1 28.568
R5994 a_12870_n994.t2 a_12870_n994.n4 28.565
R5995 a_12870_n994.n4 a_12870_n994.t0 28.565
R5996 a_12870_n994.n0 a_12870_n994.t3 18.127
R5997 a_12870_n994.n2 a_12870_n994.n0 4.039
R5998 a_12870_n994.n3 a_12870_n994.n2 0.937
R5999 a_7894_n5055.t0 a_7894_n5055.t1 17.4
R6000 a_9404_3062.t0 a_9404_3062.t1 17.4
R6001 a_17148_n5059.t0 a_17148_n5059.t1 17.4
R6002 a_14999_n8092.t0 a_14999_n8092.t1 380.209
R6003 a_2345_3260.n0 a_2345_3260.t1 28.565
R6004 a_2345_3260.t2 a_2345_3260.n0 28.565
R6005 a_2345_3260.n0 a_2345_3260.n1 192.754
R6006 a_2345_3260.n1 a_2345_3260.t0 28.568
R6007 a_2345_3260.n1 a_2345_3260.n2 1.123
R6008 a_2345_3260.n2 a_2345_3260.n3 19.249
R6009 a_2345_3260.n3 a_2345_3260.t4 615.911
R6010 a_2345_3260.n3 a_2345_3260.t7 867.497
R6011 a_2345_3260.t7 a_2345_3260.n4 160.666
R6012 a_2345_3260.n4 a_2345_3260.t6 286.438
R6013 a_2345_3260.n4 a_2345_3260.t5 286.438
R6014 a_2345_3260.n2 a_2345_3260.t3 18.726
R6015 a_4772_407.t0 a_4772_407.t1 17.4
R6016 a_8794_n7362.n7 a_8794_n7362.n1 1401.24
R6017 a_8794_n7362.n1 a_8794_n7362.t9 867.497
R6018 a_8794_n7362.n1 a_8794_n7362.t10 615.911
R6019 a_8794_n7362.n0 a_8794_n7362.t8 286.438
R6020 a_8794_n7362.n0 a_8794_n7362.t11 286.438
R6021 a_8794_n7362.t9 a_8794_n7362.n0 160.666
R6022 a_8794_n7362.n5 a_8794_n7362.n3 157.665
R6023 a_8794_n7362.n5 a_8794_n7362.n4 122.999
R6024 a_8794_n7362.n8 a_8794_n7362.n7 90.436
R6025 a_8794_n7362.n6 a_8794_n7362.n2 90.416
R6026 a_8794_n7362.n7 a_8794_n7362.n6 74.302
R6027 a_8794_n7362.n6 a_8794_n7362.n5 50.575
R6028 a_8794_n7362.n2 a_8794_n7362.t0 14.282
R6029 a_8794_n7362.n2 a_8794_n7362.t5 14.282
R6030 a_8794_n7362.n4 a_8794_n7362.t6 14.282
R6031 a_8794_n7362.n4 a_8794_n7362.t7 14.282
R6032 a_8794_n7362.n8 a_8794_n7362.t1 14.282
R6033 a_8794_n7362.t2 a_8794_n7362.n8 14.282
R6034 a_8794_n7362.n3 a_8794_n7362.t3 8.7
R6035 a_8794_n7362.n3 a_8794_n7362.t4 8.7
R6036 a_13359_n3752.t2 a_13359_n3752.n0 28.565
R6037 a_13359_n3752.n0 a_13359_n3752.t1 28.565
R6038 a_13359_n3752.n0 a_13359_n3752.n1 197.272
R6039 a_13359_n3752.n1 a_13359_n3752.t0 28.568
R6040 a_13359_n3752.n1 a_13359_n3752.n2 0.459
R6041 a_13359_n3752.n2 a_13359_n3752.n3 25.659
R6042 a_13359_n3752.n3 a_13359_n3752.t4 408.211
R6043 a_13359_n3752.n3 a_13359_n3752.t6 990.34
R6044 a_13359_n3752.t6 a_13359_n3752.n4 160.666
R6045 a_13359_n3752.n4 a_13359_n3752.t7 286.438
R6046 a_13359_n3752.n4 a_13359_n3752.t5 286.438
R6047 a_13359_n3752.n2 a_13359_n3752.t3 18.103
R6048 a_12860_n3726.n2 a_12860_n3726.t7 448.382
R6049 a_12860_n3726.n1 a_12860_n3726.t6 286.438
R6050 a_12860_n3726.n1 a_12860_n3726.t5 286.438
R6051 a_12860_n3726.n0 a_12860_n3726.t4 247.69
R6052 a_12860_n3726.n4 a_12860_n3726.n3 182.117
R6053 a_12860_n3726.t7 a_12860_n3726.n1 160.666
R6054 a_12860_n3726.n3 a_12860_n3726.t0 28.568
R6055 a_12860_n3726.n4 a_12860_n3726.t1 28.565
R6056 a_12860_n3726.t2 a_12860_n3726.n4 28.565
R6057 a_12860_n3726.n0 a_12860_n3726.t3 18.127
R6058 a_12860_n3726.n2 a_12860_n3726.n0 4.039
R6059 a_12860_n3726.n3 a_12860_n3726.n2 0.937
R6060 a_14240_n5059.t0 a_14240_n5059.t1 17.4
R6061 a_4772_n2327.t0 a_4772_n2327.t1 17.4
R6062 a_19146_1744.n2 a_19146_1744.t4 448.382
R6063 a_19146_1744.n1 a_19146_1744.t6 286.438
R6064 a_19146_1744.n1 a_19146_1744.t7 286.438
R6065 a_19146_1744.n0 a_19146_1744.t5 247.69
R6066 a_19146_1744.n4 a_19146_1744.n3 182.117
R6067 a_19146_1744.t4 a_19146_1744.n1 160.666
R6068 a_19146_1744.n3 a_19146_1744.t1 28.568
R6069 a_19146_1744.n4 a_19146_1744.t0 28.565
R6070 a_19146_1744.t2 a_19146_1744.n4 28.565
R6071 a_19146_1744.n0 a_19146_1744.t3 18.127
R6072 a_19146_1744.n2 a_19146_1744.n0 4.039
R6073 a_19146_1744.n3 a_19146_1744.n2 0.937
R6074 a_17384_n5059.t0 a_17384_n5059.t1 17.4
R6075 a_15235_n8092.t0 a_15235_n8092.t1 17.4
R6076 a_20398_3112.t2 a_20398_3112.n0 28.568
R6077 a_20398_3112.n0 a_20398_3112.n4 149.031
R6078 a_20398_3112.n4 a_20398_3112.n3 67.391
R6079 a_20398_3112.n3 a_20398_3112.t0 28.565
R6080 a_20398_3112.n3 a_20398_3112.t1 28.565
R6081 a_20398_3112.n4 a_20398_3112.n1 1056.04
R6082 a_20398_3112.n1 a_20398_3112.t7 408.211
R6083 a_20398_3112.n1 a_20398_3112.t5 990.34
R6084 a_20398_3112.t5 a_20398_3112.n2 160.666
R6085 a_20398_3112.n2 a_20398_3112.t6 286.438
R6086 a_20398_3112.n2 a_20398_3112.t4 286.438
R6087 a_20398_3112.n0 a_20398_3112.t3 17.64
R6088 a_3490_3062.t0 a_3490_3062.t1 17.4
R6089 Y[7].n1 Y[7].n0 185.55
R6090 Y[7].n1 Y[7].t1 28.568
R6091 Y[7].n0 Y[7].t0 28.565
R6092 Y[7].n0 Y[7].t2 28.565
R6093 Y[7].n2 Y[7].t3 21.373
R6094 Y[7].n2 Y[7].n1 1.537
R6095 Y[7] Y[7].n2 0.312
R6096 a_11048_n2323.t0 a_11048_n2323.t1 17.4
R6097 a_7019_n7388.n1 a_7019_n7388.t6 318.922
R6098 a_7019_n7388.n0 a_7019_n7388.t5 274.739
R6099 a_7019_n7388.n0 a_7019_n7388.t7 274.739
R6100 a_7019_n7388.n1 a_7019_n7388.t4 269.116
R6101 a_7019_n7388.t6 a_7019_n7388.n0 179.946
R6102 a_7019_n7388.n2 a_7019_n7388.n1 107.263
R6103 a_7019_n7388.n3 a_7019_n7388.t0 29.444
R6104 a_7019_n7388.n4 a_7019_n7388.t1 28.565
R6105 a_7019_n7388.t2 a_7019_n7388.n4 28.565
R6106 a_7019_n7388.n2 a_7019_n7388.t3 18.145
R6107 a_7019_n7388.n3 a_7019_n7388.n2 2.878
R6108 a_7019_n7388.n4 a_7019_n7388.n3 0.764
R6109 a_6725_n8094.t0 a_6725_n8094.t1 380.209
R6110 a_544_3060.t0 a_544_3060.t1 17.4
R6111 a_6458_3060.t0 a_6458_3060.t1 17.4
R6112 a_22789_n1016.t2 a_22789_n1016.n0 28.565
R6113 a_22789_n1016.n0 a_22789_n1016.t1 28.565
R6114 a_22789_n1016.n1 a_22789_n1016.n2 0.002
R6115 a_22789_n1016.n0 a_22789_n1016.n1 185.55
R6116 a_22789_n1016.n1 a_22789_n1016.t0 28.568
R6117 a_22789_n1016.n2 a_22789_n1016.t3 23.414
R6118 a_22789_n1016.n2 a_22789_n1016.n3 12.317
R6119 a_22789_n1016.n3 a_22789_n1016.t5 408.211
R6120 a_22789_n1016.n3 a_22789_n1016.t6 990.34
R6121 a_22789_n1016.t6 a_22789_n1016.n4 160.666
R6122 a_22789_n1016.n4 a_22789_n1016.t7 286.438
R6123 a_22789_n1016.n4 a_22789_n1016.t4 286.438
R6124 a_1618_n5059.t0 a_1618_n5059.t1 17.4
R6125 a_4536_407.t0 a_4536_407.t1 17.4
R6126 a_22280_n3722.n3 a_22280_n3722.t6 448.382
R6127 a_22280_n3722.n2 a_22280_n3722.t5 286.438
R6128 a_22280_n3722.n2 a_22280_n3722.t7 286.438
R6129 a_22280_n3722.n1 a_22280_n3722.t4 247.69
R6130 a_22280_n3722.n4 a_22280_n3722.n0 182.117
R6131 a_22280_n3722.t6 a_22280_n3722.n2 160.666
R6132 a_22280_n3722.t2 a_22280_n3722.n4 28.568
R6133 a_22280_n3722.n0 a_22280_n3722.t0 28.565
R6134 a_22280_n3722.n0 a_22280_n3722.t1 28.565
R6135 a_22280_n3722.n1 a_22280_n3722.t3 18.127
R6136 a_22280_n3722.n3 a_22280_n3722.n1 4.039
R6137 a_22280_n3722.n4 a_22280_n3722.n3 0.937
R6138 a_17158_407.t0 a_17158_407.t1 17.4
R6139 a_14250_407.t0 a_14250_407.t1 17.4
R6140 Y[5].n1 Y[5].n0 185.55
R6141 Y[5].n1 Y[5].t1 28.568
R6142 Y[5].n0 Y[5].t2 28.565
R6143 Y[5].n0 Y[5].t0 28.565
R6144 Y[5].n2 Y[5].t3 21.373
R6145 Y[5] Y[5].n2 10.221
R6146 Y[5].n2 Y[5].n1 1.637
R6147 a_10862_n8092.t0 a_10862_n8092.t1 380.209
R6148 a_1628_407.t0 a_1628_407.t1 17.4
R6149 a_7668_n2323.t0 a_7668_n2323.t1 17.4
R6150 a_4539_n7364.n8 a_4539_n7364.n0 267.767
R6151 a_4539_n7364.n4 a_4539_n7364.t8 16.058
R6152 a_4539_n7364.n2 a_4539_n7364.t9 16.058
R6153 a_4539_n7364.n3 a_4539_n7364.t6 14.282
R6154 a_4539_n7364.n3 a_4539_n7364.t7 14.282
R6155 a_4539_n7364.n1 a_4539_n7364.t10 14.282
R6156 a_4539_n7364.n1 a_4539_n7364.t11 14.282
R6157 a_4539_n7364.n6 a_4539_n7364.t4 14.282
R6158 a_4539_n7364.n6 a_4539_n7364.t5 14.282
R6159 a_4539_n7364.n0 a_4539_n7364.t0 14.282
R6160 a_4539_n7364.n0 a_4539_n7364.t1 14.282
R6161 a_4539_n7364.t2 a_4539_n7364.n9 14.282
R6162 a_4539_n7364.n9 a_4539_n7364.t3 14.282
R6163 a_4539_n7364.n7 a_4539_n7364.n6 1.511
R6164 a_4539_n7364.n4 a_4539_n7364.n3 0.999
R6165 a_4539_n7364.n2 a_4539_n7364.n1 0.999
R6166 a_4539_n7364.n8 a_4539_n7364.n7 0.669
R6167 a_4539_n7364.n5 a_4539_n7364.n4 0.575
R6168 a_4539_n7364.n7 a_4539_n7364.n5 0.227
R6169 a_4539_n7364.n5 a_4539_n7364.n2 0.2
R6170 a_4539_n7364.n9 a_4539_n7364.n8 0.001
R6171 a_10812_411.t0 a_10812_411.t1 17.4
R6172 a_23434_n2323.t0 a_23434_n2323.t1 17.4
R6173 a_14014_n2327.t0 a_14014_n2327.t1 17.4
R6174 a_7904_n2323.t0 a_7904_n2323.t1 17.4
R6175 a_17394_n2327.t0 a_17394_n2327.t1 17.4
R6176 a_7904_411.t0 a_7904_411.t1 17.4
R6177 a_1628_n2327.t0 a_1628_n2327.t1 17.4
R6178 a_16503_n3752.t2 a_16503_n3752.n0 28.565
R6179 a_16503_n3752.n0 a_16503_n3752.t1 28.565
R6180 a_16503_n3752.n0 a_16503_n3752.n1 197.272
R6181 a_16503_n3752.n1 a_16503_n3752.t0 28.568
R6182 a_16503_n3752.n1 a_16503_n3752.n2 0.459
R6183 a_16503_n3752.n2 a_16503_n3752.n3 19.533
R6184 a_16503_n3752.n3 a_16503_n3752.t7 408.211
R6185 a_16503_n3752.n3 a_16503_n3752.t5 990.34
R6186 a_16503_n3752.t5 a_16503_n3752.n4 160.666
R6187 a_16503_n3752.n4 a_16503_n3752.t6 286.438
R6188 a_16503_n3752.n4 a_16503_n3752.t4 286.438
R6189 a_16503_n3752.n2 a_16503_n3752.t3 18.103
R6190 a_14014_407.t0 a_14014_407.t1 17.4
R6191 a_11098_n8092.t0 a_11098_n8092.t1 17.4
R6192 a_20280_n5055.t0 a_20280_n5055.t1 17.4
R6193 a_23670_411.t0 a_23670_411.t1 17.4
R6194 a_520_n8096.t0 a_520_n8096.t1 380.209
R6195 a_4657_n8096.t0 a_4657_n8096.t1 380.209
R6196 a_756_n8096.t0 a_756_n8096.t1 17.4
R6197 a_4893_n8096.t0 a_4893_n8096.t1 17.4
R6198 a_23660_n5055.t0 a_23660_n5055.t1 17.4
R6199 a_23434_411.t0 a_23434_411.t1 17.4
R6200 a_1992_3060.t0 a_1992_3060.t1 17.4
R6201 a_20526_411.t0 a_20526_411.t1 17.4
R6202 a_1392_407.t0 a_1392_407.t1 17.4
R6203 a_9030_n8094.t0 a_9030_n8094.t1 17.4
R6204 a_4526_n5059.t0 a_4526_n5059.t1 17.4
R6205 a_7668_411.t0 a_7668_411.t1 17.4
R6206 a_10802_n5055.t0 a_10802_n5055.t1 17.4
R6207 a_20516_n5055.t0 a_20516_n5055.t1 17.4
R6208 a_4536_n2327.t0 a_4536_n2327.t1 17.4
C0 VDD A[2] 2.75fF
C1 B[0] B[3] 0.08fF
C2 B[1] A[1] 17.11fF
C3 A[0] B[2] 0.11fF
C4 B[1] A[7] 0.07fF
C5 B[0] opcode[0] 0.27fF
C6 B[4] B[5] 3.11fF
C7 VDD opcode[1] 6.16fF
C8 A[1] A[5] 0.25fF
C9 A[0] A[6] 0.35fF
C10 B[2] B[7] 0.05fF
C11 B[3] B[6] 0.07fF
C12 A[2] A[4] 0.26fF
C13 Y[5] Y[7] 0.04fF
C14 B[5] Y[0] 0.10fF
C15 B[7] A[6] 0.21fF
C16 B[6] opcode[0] 0.30fF
C17 A[5] A[7] 0.20fF
C18 B[4] Y[2] 0.08fF
C19 A[4] opcode[1] 0.03fF
C20 opcode[1] Y[3] 0.19fF
C21 opcode[0] Y[4] 0.01fF
C22 Y[0] Y[2] 0.01fF
C23 B[1] B[3] 0.07fF
C24 A[0] A[1] 13.09fF
C25 VDD B[4] 4.36fF
C26 B[0] A[2] 0.23fF
C27 A[2] B[6] 0.11fF
C28 B[2] A[6] 0.10fF
C29 B[1] opcode[0] 0.33fF
C30 B[4] A[4] 22.46fF
C31 A[1] B[7] 0.13fF
C32 VDD Y[0] 4.45fF
C33 B[0] opcode[1] 0.08fF
C34 A[3] B[5] 0.18fF
C35 A[0] A[7] 0.38fF
C36 B[3] A[5] 0.07fF
C37 Y[6] Y[7] 0.10fF
C38 B[6] opcode[1] 0.15fF
C39 B[5] Y[1] 0.08fF
C40 A[5] opcode[0] 0.03fF
C41 B[7] A[7] 17.36fF
C42 opcode[1] Y[4] 0.21fF
C43 Y[1] Y[2] 11.31fF
C44 Y[0] Y[3] 0.00fF
C45 opcode[0] Y[5] 0.00fF
C46 VDD A[3] 2.77fF
C47 B[2] A[1] 0.19fF
C48 A[0] B[3] 0.11fF
C49 B[1] A[2] 14.94fF
C50 B[0] B[4] 0.09fF
C51 VDD Y[1] 2.18fF
C52 A[2] A[5] 0.29fF
C53 B[3] B[7] 0.04fF
C54 B[4] B[6] 0.06fF
C55 B[2] A[7] 0.10fF
C56 B[1] opcode[1] 0.16fF
C57 A[3] A[4] 27.66fF
C58 A[1] A[6] 0.28fF
C59 A[0] opcode[0] 0.25fF
C60 A[5] opcode[1] 0.02fF
C61 A[6] A[7] 28.57fF
C62 B[6] Y[0] 0.10fF
C63 B[5] Y[2] 0.10fF
C64 B[7] opcode[0] 0.35fF
C65 Y[1] Y[3] 0.01fF
C66 Y[0] Y[4] 0.00fF
C67 opcode[0] Y[6] 0.00fF
C68 opcode[1] Y[5] 0.23fF
C69 VDD B[5] 4.15fF
C70 A[0] A[2] 0.32fF
C71 B[0] A[3] 0.22fF
C72 B[2] B[3] 1.96fF
C73 B[1] B[4] 0.08fF
C74 A[1] A[7] 0.32fF
C75 A[2] B[7] 0.07fF
C76 A[0] opcode[1] 0.12fF
C77 B[4] A[5] 14.31fF
C78 B[2] opcode[0] 0.36fF
C79 B[3] A[6] 0.10fF
C80 VDD Y[2] 1.01fF
C81 B[5] A[4] 0.21fF
C82 B[1] Y[0] 0.10fF
C83 A[3] B[6] 0.18fF
C84 B[5] Y[3] 0.01fF
C85 A[6] opcode[0] 0.03fF
C86 B[7] opcode[1] 0.18fF
C87 B[6] Y[1] 0.08fF
C88 Y[1] Y[4] 0.01fF
C89 Y[2] Y[3] 1.97fF
C90 Y[0] Y[5] 0.00fF
C91 opcode[1] Y[6] 0.13fF
C92 B[2] A[2] 16.57fF
C93 VDD A[4] 2.16fF
C94 B[1] A[3] 0.10fF
C95 B[0] B[5] 0.08fF
C96 A[1] B[3] 0.13fF
C97 A[0] B[4] 0.11fF
C98 A[3] A[5] 0.19fF
C99 B[3] A[7] 0.10fF
C100 B[2] opcode[1] 0.19fF
C101 A[1] opcode[0] 1.76fF
C102 VDD Y[3] 1.09fF
C103 B[4] B[7] 0.03fF
C104 A[2] A[6] 0.35fF
C105 B[5] B[6] 3.75fF
C106 B[6] Y[2] 0.08fF
C107 B[7] Y[0] 0.10fF
C108 A[7] opcode[0] 0.04fF
C109 A[6] opcode[1] 0.03fF
C110 Y[2] Y[4] 0.01fF
C111 Y[1] Y[5] 0.01fF
C112 Y[0] Y[6] 0.00fF
C113 opcode[1] Y[7] 0.01fF
C114 VDD B[0] 2.68fF
C115 A[0] A[3] 0.34fF
C116 VDD B[6] 3.52fF
C117 B[2] B[4] 0.07fF
C118 B[1] B[5] 0.09fF
C119 B[0] A[4] 0.18fF
C120 A[1] A[2] 13.15fF
C121 A[4] B[6] 0.13fF
C122 B[5] A[5] 17.15fF
C123 B[4] A[6] 0.12fF
C124 B[3] opcode[0] 0.30fF
C125 A[2] A[7] 0.42fF
C126 A[3] B[7] 0.10fF
C127 B[2] Y[0] 0.12fF
C128 VDD Y[4] 0.88fF
C129 A[1] opcode[1] 0.03fF
C130 B[7] Y[1] 0.08fF
C131 A[7] opcode[1] 0.04fF
C132 B[6] Y[3] 0.11fF
C133 Y[3] Y[4] 3.83fF
C134 Y[0] Y[7] 0.00fF
C135 Y[1] Y[6] 0.01fF
C136 Y[2] Y[5] 0.01fF
C137 VDD B[1] 4.64fF
C138 A[1] B[4] 0.15fF
C139 A[0] B[5] 0.11fF
C140 VDD A[5] 1.98fF
C141 B[1] A[4] 0.08fF
C142 B[3] A[2] 0.18fF
C143 B[0] B[6] 0.08fF
C144 B[2] A[3] 19.89fF
C145 A[4] A[5] 22.87fF
C146 A[2] opcode[0] 0.04fF
C147 B[5] B[7] 0.04fF
C148 B[4] A[7] 0.12fF
C149 B[3] opcode[1] 0.14fF
C150 A[3] A[6] 0.23fF
C151 B[2] Y[1] 0.01fF
C152 B[7] Y[2] 0.08fF
C153 opcode[0] opcode[1] 0.43fF
C154 VDD Y[5] 0.83fF
C155 Y[2] Y[6] 0.01fF
C156 Y[3] Y[5] 0.01fF
C157 Y[1] Y[7] 0.00fF
C158 B[0] B[1] 0.33fF
C159 VDD A[0] 5.39fF
C160 B[2] B[5] 0.08fF
C161 A[0] A[4] 0.35fF
C162 VDD B[7] 3.94fF
C163 B[1] B[6] 0.08fF
C164 A[1] A[3] 0.22fF
C165 B[0] A[5] 0.13fF
C166 B[3] B[4] 2.60fF
C167 B[3] Y[0] 0.10fF
C168 A[3] A[7] 0.27fF
C169 B[6] A[5] 0.25fF
C170 A[4] B[7] 0.05fF
C171 B[4] opcode[0] 0.38fF
C172 B[5] A[6] 14.01fF
C173 A[2] opcode[1] 0.03fF
C174 opcode[0] Y[0] 1.61fF
C175 B[7] Y[3] 0.08fF
C176 VDD Y[6] 0.82fF
C177 Y[4] Y[5] 2.05fF
C178 Y[2] Y[7] 0.01fF
C179 Y[3] Y[6] 0.01fF
C180 B[0] A[0] 26.70fF
C181 VDD B[2] 4.32fF
C182 B[2] A[4] 0.08fF
C183 VDD A[6] 1.84fF
C184 B[0] B[7] 0.08fF
C185 A[2] B[4] 0.11fF
C186 B[3] A[3] 16.50fF
C187 A[0] B[6] 0.11fF
C188 A[1] B[5] 0.15fF
C189 B[1] A[5] 0.07fF
C190 B[4] opcode[1] 0.17fF
C191 B[5] A[7] 0.14fF
C192 A[3] opcode[0] 0.04fF
C193 B[3] Y[1] 0.13fF
C194 B[6] B[7] 3.78fF
C195 A[4] A[6] 0.19fF
C196 opcode[1] Y[0] 0.10fF
C197 opcode[0] Y[1] 0.08fF
C198 B[7] Y[4] 0.04fF
C199 VDD Y[7] 0.70fF
C200 Y[3] Y[7] 0.01fF
C201 Y[4] Y[6] 0.01fF
C202 B[1] A[0] 0.22fF
C203 VDD A[1] 3.21fF
C204 B[0] B[2] 0.08fF
C205 B[1] B[7] 0.09fF
C206 B[2] B[6] 0.08fF
C207 B[0] A[6] 0.10fF
C208 B[3] B[5] 0.06fF
C209 VDD A[7] 1.64fF
C210 A[0] A[5] 0.33fF
C211 A[2] A[3] 25.89fF
C212 A[1] A[4] 0.24fF
C213 B[6] A[6] 16.48fF
C214 B[5] opcode[0] 0.42fF
C215 A[4] A[7] 0.23fF
C216 B[4] Y[0] 0.10fF
C217 A[5] B[7] 0.06fF
C218 A[3] opcode[1] 0.03fF
C219 opcode[0] Y[2] 0.03fF
C220 opcode[1] Y[1] 0.15fF
C221 Y[4] Y[7] 0.01fF
C222 B[0] A[1] 15.95fF
C223 B[1] B[2] 0.20fF
C224 VDD B[3] 4.08fF
C225 B[0] A[7] 0.07fF
C226 A[1] B[6] 0.14fF
C227 B[4] A[3] 0.25fF
C228 B[2] A[5] 0.07fF
C229 B[1] A[6] 0.07fF
C230 VDD opcode[0] 12.62fF
C231 B[3] A[4] 14.53fF
C232 A[2] B[5] 0.11fF
C233 A[0] B[7] 0.15fF
C234 Y[5] Y[6] 1.45fF
C235 B[4] Y[1] 0.08fF
C236 A[5] A[6] 22.24fF
C237 A[4] opcode[0] 0.03fF
C238 B[6] A[7] 13.73fF
C239 B[5] opcode[1] 0.19fF
C240 Y[0] Y[1] 2.80fF
C241 opcode[1] Y[2] 0.17fF
C242 opcode[0] Y[3] 0.02fF
.ends

