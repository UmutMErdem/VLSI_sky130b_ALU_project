magic
tech sky130B
magscale 1 2
timestamp 1735469461
<< nwell >>
rect 1 6 1193 330
<< nmos >>
rect 332 -569 392 -169
rect 450 -569 510 -169
rect 685 -369 745 -169
<< pmos >>
rect 95 68 155 268
rect 213 68 273 268
rect 331 68 391 268
rect 449 68 509 268
rect 567 68 627 268
rect 685 68 745 268
rect 803 68 863 268
rect 921 68 981 268
rect 1039 68 1099 268
<< ndiff >>
rect 274 -181 332 -169
rect 274 -557 286 -181
rect 320 -557 332 -181
rect 274 -569 332 -557
rect 392 -181 450 -169
rect 392 -557 404 -181
rect 438 -557 450 -181
rect 392 -569 450 -557
rect 510 -181 568 -169
rect 510 -557 522 -181
rect 556 -557 568 -181
rect 627 -181 685 -169
rect 627 -357 639 -181
rect 673 -357 685 -181
rect 627 -369 685 -357
rect 745 -181 803 -169
rect 745 -357 757 -181
rect 791 -357 803 -181
rect 745 -369 803 -357
rect 510 -569 568 -557
<< pdiff >>
rect 37 256 95 268
rect 37 80 49 256
rect 83 80 95 256
rect 37 68 95 80
rect 155 256 213 268
rect 155 80 167 256
rect 201 80 213 256
rect 155 68 213 80
rect 273 256 331 268
rect 273 80 285 256
rect 319 80 331 256
rect 273 68 331 80
rect 391 256 449 268
rect 391 80 403 256
rect 437 80 449 256
rect 391 68 449 80
rect 509 256 567 268
rect 509 80 521 256
rect 555 80 567 256
rect 509 68 567 80
rect 627 256 685 268
rect 627 80 639 256
rect 673 80 685 256
rect 627 68 685 80
rect 745 256 803 268
rect 745 80 757 256
rect 791 80 803 256
rect 745 68 803 80
rect 863 256 921 268
rect 863 80 875 256
rect 909 80 921 256
rect 863 68 921 80
rect 981 256 1039 268
rect 981 80 993 256
rect 1027 80 1039 256
rect 981 68 1039 80
rect 1099 256 1157 268
rect 1099 80 1111 256
rect 1145 80 1157 256
rect 1099 68 1157 80
<< ndiffc >>
rect 286 -557 320 -181
rect 404 -557 438 -181
rect 522 -557 556 -181
rect 639 -357 673 -181
rect 757 -357 791 -181
<< pdiffc >>
rect 49 80 83 256
rect 167 80 201 256
rect 285 80 319 256
rect 403 80 437 256
rect 521 80 555 256
rect 639 80 673 256
rect 757 80 791 256
rect 875 80 909 256
rect 993 80 1027 256
rect 1111 80 1145 256
<< poly >>
rect 95 289 391 325
rect 95 268 155 289
rect 213 268 273 289
rect 331 268 391 289
rect 449 288 745 324
rect 449 268 509 288
rect 567 268 627 288
rect 685 268 745 288
rect 803 288 1099 324
rect 803 268 863 288
rect 921 268 981 288
rect 1039 268 1099 288
rect 95 42 155 68
rect 213 42 273 68
rect 331 42 391 68
rect 449 48 509 68
rect 449 42 510 48
rect 567 42 627 68
rect 685 42 745 68
rect 332 -143 390 42
rect 332 -169 392 -143
rect 450 -169 510 42
rect 803 36 863 68
rect 921 42 981 68
rect 1039 42 1099 68
rect 800 20 866 36
rect 800 -14 816 20
rect 850 -14 866 20
rect 800 -30 866 -14
rect 682 -97 748 -81
rect 682 -131 698 -97
rect 732 -131 748 -97
rect 682 -147 748 -131
rect 685 -169 745 -147
rect 685 -395 745 -369
rect 332 -591 392 -569
rect 450 -591 510 -569
rect 329 -607 395 -591
rect 329 -641 345 -607
rect 379 -641 395 -607
rect 329 -657 395 -641
rect 447 -607 513 -591
rect 447 -641 463 -607
rect 497 -641 513 -607
rect 447 -657 513 -641
<< polycont >>
rect 816 -14 850 20
rect 698 -131 732 -97
rect 345 -641 379 -607
rect 463 -641 497 -607
<< locali >>
rect 875 306 1145 340
rect 49 256 83 272
rect 49 64 83 80
rect 167 256 201 272
rect 167 64 201 80
rect 285 256 319 272
rect 285 64 319 80
rect 403 256 437 272
rect 403 64 437 80
rect 521 256 555 272
rect 521 64 555 80
rect 639 256 673 272
rect 639 64 673 80
rect 757 256 791 272
rect 757 64 791 80
rect 875 256 909 306
rect 875 64 909 80
rect 993 256 1027 272
rect 993 64 1027 80
rect 1111 256 1145 306
rect 1111 64 1145 80
rect 800 -14 816 20
rect 850 -14 866 20
rect 682 -131 698 -97
rect 732 -131 748 -97
rect 286 -181 320 -165
rect 286 -573 320 -557
rect 404 -181 438 -165
rect 404 -573 438 -557
rect 522 -181 556 -165
rect 639 -181 673 -165
rect 639 -373 673 -357
rect 757 -181 791 -165
rect 757 -373 791 -357
rect 522 -573 556 -557
rect 329 -641 345 -607
rect 379 -641 395 -607
rect 447 -641 463 -607
rect 497 -641 513 -607
<< viali >>
rect 49 80 83 256
rect 167 80 201 256
rect 285 80 319 256
rect 403 80 437 256
rect 521 80 555 256
rect 639 80 673 256
rect 757 80 791 256
rect 875 80 909 256
rect 993 80 1027 256
rect 1111 80 1145 256
rect 816 -14 850 20
rect 698 -131 732 -97
rect 286 -557 320 -181
rect 404 -557 438 -181
rect 522 -557 556 -181
rect 639 -357 673 -181
rect 757 -357 791 -181
rect 345 -641 379 -607
rect 463 -641 497 -607
<< metal1 >>
rect 322 536 522 552
rect 322 416 356 536
rect 492 416 522 536
rect 322 404 522 416
rect 50 374 1027 404
rect 50 268 82 374
rect 286 268 318 374
rect 522 268 554 374
rect 758 268 790 374
rect 993 268 1027 374
rect 43 256 89 268
rect 43 80 49 256
rect 83 80 89 256
rect 43 68 89 80
rect 161 256 207 268
rect 161 80 167 256
rect 201 80 207 256
rect 161 68 207 80
rect 279 256 325 268
rect 279 80 285 256
rect 319 80 325 256
rect 279 68 325 80
rect 397 256 443 268
rect 397 80 403 256
rect 437 80 443 256
rect 397 68 443 80
rect 515 256 561 268
rect 515 80 521 256
rect 555 80 561 256
rect 515 68 561 80
rect 633 256 679 268
rect 633 80 639 256
rect 673 80 679 256
rect 633 68 679 80
rect 751 256 797 268
rect 751 80 757 256
rect 791 80 797 256
rect 751 68 797 80
rect 869 256 915 268
rect 869 80 875 256
rect 909 80 915 256
rect 869 68 915 80
rect 987 256 1033 268
rect 987 80 993 256
rect 1027 80 1033 256
rect 987 68 1033 80
rect 1105 256 1151 268
rect 1105 80 1111 256
rect 1145 80 1151 256
rect 1105 68 1151 80
rect 166 -26 202 68
rect 402 -26 438 68
rect 638 -25 674 68
rect 800 20 866 27
rect 800 -14 816 20
rect 850 -14 866 20
rect 800 -25 866 -14
rect 638 -26 866 -25
rect 166 -55 866 -26
rect 166 -56 748 -55
rect 286 -169 320 -56
rect 682 -97 748 -56
rect 682 -131 698 -97
rect 732 -131 748 -97
rect 682 -138 748 -131
rect 1110 -165 1145 68
rect 756 -169 1145 -165
rect 280 -181 326 -169
rect 280 -557 286 -181
rect 320 -557 326 -181
rect 280 -569 326 -557
rect 398 -181 444 -169
rect 398 -557 404 -181
rect 438 -557 444 -181
rect 398 -569 444 -557
rect 516 -181 562 -169
rect 516 -557 522 -181
rect 556 -533 562 -181
rect 633 -181 679 -169
rect 633 -357 639 -181
rect 673 -357 679 -181
rect 633 -369 679 -357
rect 751 -181 1145 -169
rect 751 -357 757 -181
rect 791 -194 1145 -181
rect 791 -357 797 -194
rect 1041 -274 1145 -194
rect 751 -369 797 -357
rect 639 -533 674 -369
rect 718 -533 728 -525
rect 556 -557 728 -533
rect 516 -569 728 -557
rect 522 -573 728 -569
rect 58 -601 158 -573
rect 718 -585 728 -573
rect 788 -585 798 -525
rect 58 -607 395 -601
rect 58 -641 345 -607
rect 379 -641 395 -607
rect 58 -657 395 -641
rect 447 -607 513 -601
rect 447 -641 463 -607
rect 497 -641 513 -607
rect 58 -673 158 -657
rect 58 -737 158 -715
rect 447 -737 513 -641
rect 58 -785 513 -737
rect 58 -815 158 -785
<< via1 >>
rect 356 416 492 536
rect 728 -585 788 -525
<< metal2 >>
rect 356 536 492 546
rect 356 406 492 416
rect 718 -515 798 -505
rect 718 -605 798 -595
<< via2 >>
rect 356 416 492 536
rect 718 -525 798 -515
rect 718 -585 728 -525
rect 728 -585 788 -525
rect 788 -585 798 -525
rect 718 -595 798 -585
<< metal3 >>
rect 346 536 502 541
rect 346 416 356 536
rect 492 416 502 536
rect 346 411 502 416
rect 702 -533 708 -505
rect 698 -605 708 -533
rect 808 -605 818 -505
<< via3 >>
rect 356 416 492 536
rect 708 -515 808 -505
rect 708 -595 718 -515
rect 718 -595 798 -515
rect 798 -595 808 -515
rect 708 -605 808 -595
<< metal4 >>
rect 298 536 548 656
rect 298 436 356 536
rect 355 416 356 436
rect 492 436 548 536
rect 492 416 493 436
rect 355 415 493 416
rect 766 -504 934 -495
rect 707 -505 934 -504
rect 707 -605 708 -505
rect 808 -605 934 -505
rect 707 -606 934 -605
rect 766 -685 934 -606
<< labels >>
flabel metal4 322 498 522 640 1 FreeSans 480 0 0 0 VDD
port 4 n
flabel metal1 58 -815 158 -715 1 FreeSans 480 0 0 0 B
port 3 n
flabel metal1 58 -673 158 -573 1 FreeSans 480 0 0 0 A
port 2 n
flabel metal4 784 -645 904 -541 1 FreeSans 480 0 0 0 VSS
port 1 n
flabel metal1 1047 -264 1137 -179 1 FreeSans 240 0 0 0 Y
port 5 n
<< end >>
