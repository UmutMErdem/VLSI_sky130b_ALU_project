magic
tech sky130B
magscale 1 2
timestamp 1736796407
<< nwell >>
rect 8717 28151 9004 28152
rect 9864 28151 10099 28152
rect 6235 28097 6475 28098
rect 6232 27864 6475 28097
rect 6232 27682 6476 27864
rect 8714 27754 9004 28151
rect 9691 27758 10173 28151
rect 15230 28148 15517 28149
rect 16377 28148 16612 28149
rect 12748 28094 12988 28095
rect 5794 27358 6986 27682
rect 8119 27287 9004 27754
rect 8119 27234 9005 27287
rect 9261 27234 10173 27758
rect 12745 27861 12988 28094
rect 12745 27679 12989 27861
rect 15227 27751 15517 28148
rect 16204 27755 16686 28148
rect 28322 28147 28609 28148
rect 29469 28147 29704 28148
rect 21764 28143 22051 28144
rect 22911 28143 23146 28144
rect 19282 28089 19522 28090
rect 12307 27355 13499 27679
rect 8119 27230 9006 27234
rect 8548 26945 9006 27230
rect 9691 26975 10173 27234
rect 14632 27284 15517 27751
rect 14632 27231 15518 27284
rect 15774 27231 16686 27755
rect 19279 27856 19522 28089
rect 19279 27674 19523 27856
rect 21761 27746 22051 28143
rect 22738 27750 23220 28143
rect 25840 28093 26080 28094
rect 18841 27350 20033 27674
rect 14632 27227 15519 27231
rect 8548 26647 9032 26945
rect 9690 26651 10174 26975
rect 15061 26942 15519 27227
rect 16204 26972 16686 27231
rect 21166 27279 22051 27746
rect 21166 27226 22052 27279
rect 22308 27226 23220 27750
rect 25837 27860 26080 28093
rect 25837 27678 26081 27860
rect 28319 27750 28609 28147
rect 29296 27754 29778 28147
rect 25399 27354 26591 27678
rect 27724 27283 28609 27750
rect 27724 27230 28610 27283
rect 28866 27230 29778 27754
rect 27724 27226 28611 27230
rect 21166 27222 22053 27226
rect 15061 26644 15545 26942
rect 16203 26648 16687 26972
rect 21595 26937 22053 27222
rect 22738 26967 23220 27226
rect 21595 26639 22079 26937
rect 22737 26643 23221 26967
rect 28153 26941 28611 27226
rect 29296 26971 29778 27230
rect 28153 26643 28637 26941
rect 29295 26647 29779 26971
rect 6249 26447 6489 26448
rect 6246 26214 6489 26447
rect 12762 26444 13002 26445
rect 6246 26032 6490 26214
rect 12759 26211 13002 26444
rect 25854 26443 26094 26444
rect 19296 26439 19536 26440
rect 5808 25708 7000 26032
rect 9960 25615 10188 26105
rect 12759 26029 13003 26211
rect 19293 26206 19536 26439
rect 25851 26210 26094 26443
rect 12321 25705 13513 26029
rect 7271 25415 8594 25615
rect 9654 25415 10492 25615
rect 16473 25612 16701 26102
rect 19293 26024 19537 26206
rect 18855 25700 20047 26024
rect 7271 25091 10975 25415
rect 13784 25412 15107 25612
rect 16167 25412 17005 25612
rect 23007 25607 23235 26097
rect 25851 26028 26095 26210
rect 25413 25704 26605 26028
rect 29565 25611 29793 26101
rect 6244 24843 6484 24844
rect 6241 24610 6484 24843
rect 6241 24428 6485 24610
rect 5803 24104 6995 24428
rect 7699 24398 8537 25091
rect 9597 24398 10435 25091
rect 13784 25088 17488 25412
rect 20318 25407 21641 25607
rect 22701 25407 23539 25607
rect 26876 25411 28199 25611
rect 29259 25411 30097 25611
rect 12757 24840 12997 24841
rect 12754 24607 12997 24840
rect 12754 24425 12998 24607
rect 12316 24101 13508 24425
rect 14212 24395 15050 25088
rect 16110 24395 16948 25088
rect 20318 25083 24022 25407
rect 26876 25087 30580 25411
rect 19291 24835 19531 24836
rect 19288 24602 19531 24835
rect 19288 24420 19532 24602
rect 18850 24096 20042 24420
rect 20746 24390 21584 25083
rect 22644 24390 23482 25083
rect 25849 24839 26089 24840
rect 25846 24606 26089 24839
rect 25846 24424 26090 24606
rect 25408 24100 26600 24424
rect 27304 24394 28142 25087
rect 29202 24394 30040 25087
rect 36893 24755 37217 25196
rect 36403 22978 37217 24755
rect 36693 22977 37217 22978
rect 25410 22547 25645 22548
rect 26505 22547 26792 22548
rect 18897 22544 19132 22545
rect 19992 22544 20279 22545
rect 5805 22543 6040 22544
rect 6900 22543 7187 22544
rect 5731 22150 6213 22543
rect 5731 21626 6643 22150
rect 6900 22146 7190 22543
rect 12363 22539 12598 22540
rect 13458 22539 13745 22540
rect 9429 22489 9669 22490
rect 9429 22256 9672 22489
rect 6900 21679 7785 22146
rect 9428 22074 9672 22256
rect 12289 22146 12771 22539
rect 8918 21750 10110 22074
rect 6899 21626 7785 21679
rect 5731 21367 6213 21626
rect 6898 21622 7785 21626
rect 12289 21622 13201 22146
rect 13458 22142 13748 22539
rect 15987 22485 16227 22486
rect 15987 22252 16230 22485
rect 13458 21675 14343 22142
rect 15986 22070 16230 22252
rect 18823 22151 19305 22544
rect 15476 21746 16668 22070
rect 13457 21622 14343 21675
rect 5730 21043 6214 21367
rect 6898 21337 7356 21622
rect 12289 21363 12771 21622
rect 13456 21618 14343 21622
rect 18823 21627 19735 22151
rect 19992 22147 20282 22544
rect 22521 22490 22761 22491
rect 22521 22257 22764 22490
rect 19992 21680 20877 22147
rect 22520 22075 22764 22257
rect 25336 22154 25818 22547
rect 22010 21751 23202 22075
rect 19991 21627 20877 21680
rect 6872 21039 7356 21337
rect 12288 21039 12772 21363
rect 13456 21333 13914 21618
rect 18823 21368 19305 21627
rect 19990 21623 20877 21627
rect 25336 21630 26248 22154
rect 26505 22150 26795 22547
rect 36893 22504 37217 22977
rect 29034 22493 29274 22494
rect 29034 22260 29277 22493
rect 26505 21683 27390 22150
rect 29033 22078 29277 22260
rect 28523 21754 29715 22078
rect 26504 21630 27390 21683
rect 13430 21035 13914 21333
rect 18822 21044 19306 21368
rect 19990 21338 20448 21623
rect 25336 21371 25818 21630
rect 26503 21626 27390 21630
rect 19964 21040 20448 21338
rect 25335 21047 25819 21371
rect 26503 21341 26961 21626
rect 36893 21611 37217 22052
rect 26477 21043 26961 21341
rect 29020 20843 29260 20844
rect 22507 20840 22747 20841
rect 9415 20839 9655 20840
rect 9415 20606 9658 20839
rect 5716 20007 5944 20497
rect 9414 20424 9658 20606
rect 15973 20835 16213 20836
rect 15973 20602 16216 20835
rect 22507 20607 22750 20840
rect 29020 20610 29263 20843
rect 8904 20100 10096 20424
rect 5412 19807 6250 20007
rect 7310 19807 8633 20007
rect 12274 20003 12502 20493
rect 15972 20420 16216 20602
rect 15462 20096 16654 20420
rect 18808 20008 19036 20498
rect 22506 20425 22750 20607
rect 21996 20101 23188 20425
rect 25321 20011 25549 20501
rect 29019 20428 29263 20610
rect 28509 20104 29701 20428
rect 4929 19483 8633 19807
rect 11970 19803 12808 20003
rect 13868 19803 15191 20003
rect 18504 19808 19342 20008
rect 20402 19808 21725 20008
rect 25017 19811 25855 20011
rect 26915 19811 28238 20011
rect 36403 19834 37217 21611
rect 36693 19833 37217 19834
rect 5469 18790 6307 19483
rect 7367 18790 8205 19483
rect 11487 19479 15191 19803
rect 18021 19484 21725 19808
rect 24534 19487 28238 19811
rect 9420 19235 9660 19236
rect 9420 19002 9663 19235
rect 9419 18820 9663 19002
rect 8909 18496 10101 18820
rect 12027 18786 12865 19479
rect 13925 18786 14763 19479
rect 15978 19231 16218 19232
rect 15978 18998 16221 19231
rect 15977 18816 16221 18998
rect 15467 18492 16659 18816
rect 18561 18791 19399 19484
rect 20459 18791 21297 19484
rect 22512 19236 22752 19237
rect 22512 19003 22755 19236
rect 22511 18821 22755 19003
rect 22001 18497 23193 18821
rect 25074 18794 25912 19487
rect 26972 18794 27810 19487
rect 36893 19360 37217 19833
rect 29025 19239 29265 19240
rect 29025 19006 29268 19239
rect 29024 18824 29268 19006
rect 28514 18500 29706 18824
rect 36889 18479 37213 18920
rect 36399 16702 37213 18479
rect 36689 16701 37213 16702
rect -3666 15876 -3342 16303
rect 36889 16228 37213 16701
rect -3666 15822 -2649 15876
rect -3961 15632 -2649 15822
rect -4153 15156 -2649 15632
rect 7763 15298 8955 15544
rect 7763 15286 8956 15298
rect -3961 15038 -2649 15156
rect -3961 14978 -3342 15038
rect -3666 14498 -3342 14978
rect 7764 14974 8956 15286
rect 14312 15297 15504 15543
rect 20966 15318 22158 15564
rect 20966 15306 22159 15318
rect 14312 15285 15505 15297
rect 14313 14973 15505 15285
rect 20967 14994 22159 15306
rect 29619 15151 30811 15397
rect 29619 15139 30812 15151
rect 29620 14827 30812 15139
rect 32074 14989 32571 15446
rect 36889 15335 37213 15776
rect 31428 14743 34412 14989
rect 31428 14422 34413 14743
rect -3668 13808 -3344 14235
rect -3668 13754 -2651 13808
rect -3963 13564 -2651 13754
rect 31855 13729 32693 14422
rect 33221 14419 34413 14422
rect 13462 13688 13749 13689
rect 14609 13688 14844 13689
rect 26741 13688 27028 13689
rect 27888 13688 28123 13689
rect -4153 13088 -2651 13564
rect 1099 13398 2291 13644
rect 10980 13634 11220 13635
rect 6913 13600 7200 13601
rect 8060 13600 8295 13601
rect 4431 13546 4671 13547
rect 1099 13386 2292 13398
rect -3963 12970 -2651 13088
rect 1100 13074 2292 13386
rect 4428 13313 4671 13546
rect 4428 13131 4672 13313
rect 6910 13203 7200 13600
rect 7887 13207 8369 13600
rect 10977 13401 11220 13634
rect 10977 13219 11221 13401
rect 13459 13291 13749 13688
rect 14436 13295 14918 13688
rect 24259 13634 24499 13635
rect 20116 13620 20403 13621
rect 21263 13620 21498 13621
rect 17634 13566 17874 13567
rect -3963 12910 -3344 12970
rect -3668 12430 -3344 12910
rect 3990 12807 5182 13131
rect 6315 12736 7200 13203
rect 6315 12683 7201 12736
rect 7457 12683 8369 13207
rect 10539 12895 11731 13219
rect 12864 12824 13749 13291
rect 12864 12771 13750 12824
rect 14006 12771 14918 13295
rect 17631 13333 17874 13566
rect 17631 13151 17875 13333
rect 20113 13223 20403 13620
rect 21090 13227 21572 13620
rect 17193 12827 18385 13151
rect 12864 12767 13751 12771
rect 6315 12679 7202 12683
rect 6744 12394 7202 12679
rect 7887 12424 8369 12683
rect 13293 12482 13751 12767
rect 14436 12512 14918 12771
rect 19518 12756 20403 13223
rect 19518 12703 20404 12756
rect 20660 12703 21572 13227
rect 24256 13401 24499 13634
rect 24256 13219 24500 13401
rect 26738 13291 27028 13688
rect 27715 13295 28197 13688
rect 36399 13558 37213 15335
rect 36689 13557 37213 13558
rect 23818 12895 25010 13219
rect 26143 12824 27028 13291
rect 26143 12771 27029 12824
rect 27285 12771 28197 13295
rect 36889 13084 37213 13557
rect 26143 12767 27030 12771
rect 19518 12699 20405 12703
rect -3666 11739 -3342 12166
rect 6744 12096 7228 12394
rect 7886 12100 8370 12424
rect 13293 12184 13777 12482
rect 14435 12188 14919 12512
rect 19947 12414 20405 12699
rect 21090 12444 21572 12703
rect 26572 12482 27030 12767
rect 27715 12512 28197 12771
rect 29614 12580 30806 12826
rect 29614 12568 30807 12580
rect 19947 12116 20431 12414
rect 21089 12120 21573 12444
rect 26572 12184 27056 12482
rect 27714 12188 28198 12512
rect 29615 12256 30807 12568
rect 36893 12133 37217 12574
rect 10994 11984 11234 11985
rect 24273 11984 24513 11985
rect 4445 11896 4685 11897
rect -3666 11685 -2649 11739
rect -3961 11495 -2649 11685
rect -4153 11019 -2649 11495
rect 4442 11663 4685 11896
rect 10991 11751 11234 11984
rect 17648 11916 17888 11917
rect 4442 11481 4686 11663
rect 10991 11569 11235 11751
rect 17645 11683 17888 11916
rect 24270 11751 24513 11984
rect 4004 11157 5196 11481
rect 8156 11064 8384 11554
rect 10553 11245 11745 11569
rect 14705 11152 14933 11642
rect 17645 11501 17889 11683
rect 17207 11177 18399 11501
rect -3961 10901 -2649 11019
rect -3961 10841 -3342 10901
rect -3666 10361 -3342 10841
rect 1091 10813 2283 11059
rect 5467 10864 6790 11064
rect 7850 10864 8688 11064
rect 12016 10952 13339 11152
rect 14399 10952 15237 11152
rect 21359 11084 21587 11574
rect 24270 11569 24514 11751
rect 23832 11245 25024 11569
rect 27984 11152 28212 11642
rect 1091 10801 2284 10813
rect 1092 10489 2284 10801
rect 5467 10540 9171 10864
rect 12016 10628 15720 10952
rect 18670 10884 19993 11084
rect 21053 10884 21891 11084
rect 25295 10952 26618 11152
rect 27678 10952 28516 11152
rect 4440 10292 4680 10293
rect -3668 9671 -3344 10098
rect 4437 10059 4680 10292
rect 4437 9877 4681 10059
rect -3668 9617 -2651 9671
rect -3963 9427 -2651 9617
rect 3999 9553 5191 9877
rect 5895 9847 6733 10540
rect 7793 9847 8631 10540
rect 10989 10380 11229 10381
rect 10986 10147 11229 10380
rect 10986 9965 11230 10147
rect 10548 9641 11740 9965
rect 12444 9935 13282 10628
rect 14342 9935 15180 10628
rect 18670 10560 22374 10884
rect 25295 10628 28999 10952
rect 32076 10898 32573 11355
rect 31430 10652 34414 10898
rect 17643 10312 17883 10313
rect 17640 10079 17883 10312
rect 17640 9897 17884 10079
rect 17202 9573 18394 9897
rect 19098 9867 19936 10560
rect 20996 9867 21834 10560
rect 24268 10380 24508 10381
rect 24265 10147 24508 10380
rect 24265 9965 24509 10147
rect 23827 9641 25019 9965
rect 25723 9935 26561 10628
rect 27621 9935 28459 10628
rect 31430 10331 34415 10652
rect 36403 10356 37217 12133
rect 36693 10355 37217 10356
rect 29614 9547 30806 9793
rect 31857 9638 32695 10331
rect 33223 10328 34415 10331
rect 36893 9882 37217 10355
rect 29614 9535 30807 9547
rect -4153 8951 -2651 9427
rect 29615 9223 30807 9535
rect 36893 8989 37217 9430
rect -3963 8833 -2651 8951
rect -3963 8773 -3344 8833
rect -3668 8293 -3344 8773
rect -3668 7602 -3344 8029
rect 6905 7820 7192 7821
rect 8052 7820 8287 7821
rect 26733 7820 27020 7821
rect 27880 7820 28115 7821
rect -3668 7548 -2651 7602
rect -3963 7358 -2651 7548
rect 1072 7535 2264 7781
rect 4423 7766 4663 7767
rect 1072 7523 2265 7535
rect -4155 6882 -2651 7358
rect 1073 7211 2265 7523
rect 4420 7533 4663 7766
rect 4420 7351 4664 7533
rect 6902 7423 7192 7820
rect 7879 7427 8361 7820
rect 20111 7819 20398 7820
rect 21258 7819 21493 7820
rect 13456 7818 13743 7819
rect 14603 7818 14838 7819
rect 10974 7764 11214 7765
rect 3982 7027 5174 7351
rect 6307 6956 7192 7423
rect 6307 6903 7193 6956
rect 7449 6903 8361 7427
rect 10971 7531 11214 7764
rect 10971 7349 11215 7531
rect 13453 7421 13743 7818
rect 14430 7425 14912 7818
rect 17629 7765 17869 7766
rect 10533 7025 11725 7349
rect 6307 6899 7194 6903
rect -3963 6764 -2651 6882
rect -3963 6704 -3344 6764
rect -3668 6224 -3344 6704
rect 6736 6614 7194 6899
rect 7879 6644 8361 6903
rect 12858 6954 13743 7421
rect 12858 6901 13744 6954
rect 14000 6901 14912 7425
rect 17626 7532 17869 7765
rect 17626 7350 17870 7532
rect 20108 7422 20398 7819
rect 21085 7426 21567 7819
rect 24251 7766 24491 7767
rect 17188 7026 18380 7350
rect 12858 6897 13745 6901
rect 6736 6316 7220 6614
rect 7878 6320 8362 6644
rect 13287 6612 13745 6897
rect 14430 6642 14912 6901
rect 19513 6955 20398 7422
rect 19513 6902 20399 6955
rect 20655 6902 21567 7426
rect 24248 7533 24491 7766
rect 24248 7351 24492 7533
rect 26730 7423 27020 7820
rect 27707 7427 28189 7820
rect 29685 7627 30877 7873
rect 29685 7615 30878 7627
rect 23810 7027 25002 7351
rect 19513 6898 20400 6902
rect 13287 6314 13771 6612
rect 14429 6318 14913 6642
rect 19942 6613 20400 6898
rect 21085 6643 21567 6902
rect 26135 6956 27020 7423
rect 26135 6903 27021 6956
rect 27277 6903 28189 7427
rect 29686 7303 30878 7615
rect 32076 7403 32573 7860
rect 26135 6899 27022 6903
rect 19942 6315 20426 6613
rect 21084 6319 21568 6643
rect 26564 6614 27022 6899
rect 27707 6644 28189 6903
rect 31430 7157 34414 7403
rect 36403 7212 37217 8989
rect 36693 7211 37217 7212
rect 31430 6836 34415 7157
rect 26564 6316 27048 6614
rect 27706 6320 28190 6644
rect 31857 6143 32695 6836
rect 33223 6833 34415 6836
rect 36893 6738 37217 7211
rect 4437 6116 4677 6117
rect 24265 6116 24505 6117
rect -3670 5534 -3346 5961
rect 4434 5883 4677 6116
rect 17643 6115 17883 6116
rect 10988 6114 11228 6115
rect 4434 5701 4678 5883
rect 10985 5881 11228 6114
rect 17640 5882 17883 6115
rect 24262 5883 24505 6116
rect -3670 5480 -2653 5534
rect -3965 5290 -2653 5480
rect 3996 5377 5188 5701
rect -4155 4814 -2653 5290
rect 8148 5284 8376 5774
rect 10985 5699 11229 5881
rect 10547 5375 11739 5699
rect 5459 5084 6782 5284
rect 7842 5084 8680 5284
rect 14699 5282 14927 5772
rect 17640 5700 17884 5882
rect 17202 5376 18394 5700
rect 21354 5283 21582 5773
rect 24262 5701 24506 5883
rect 36889 5857 37213 6298
rect 23824 5377 25016 5701
rect 27976 5284 28204 5774
rect -3965 4696 -2653 4814
rect 1088 4775 2280 5021
rect 1088 4763 2281 4775
rect -3965 4636 -3346 4696
rect -3670 4156 -3346 4636
rect 1089 4451 2281 4763
rect 5459 4760 9163 5084
rect 12010 5082 13333 5282
rect 14393 5082 15231 5282
rect 18665 5083 19988 5283
rect 21048 5083 21886 5283
rect 25287 5084 26610 5284
rect 27670 5084 28508 5284
rect 4432 4512 4672 4513
rect 4429 4279 4672 4512
rect 4429 4097 4673 4279
rect -3668 3465 -3344 3892
rect 3991 3773 5183 4097
rect 5887 4067 6725 4760
rect 7785 4067 8623 4760
rect 12010 4758 15714 5082
rect 18665 4759 22369 5083
rect 25287 4760 28991 5084
rect 10983 4510 11223 4511
rect 10980 4277 11223 4510
rect 10980 4095 11224 4277
rect 10542 3771 11734 4095
rect 12438 4065 13276 4758
rect 14336 4065 15174 4758
rect 17638 4511 17878 4512
rect 17635 4278 17878 4511
rect 17635 4096 17879 4278
rect 17197 3772 18389 4096
rect 19093 4066 19931 4759
rect 20991 4066 21829 4759
rect 24260 4512 24500 4513
rect 24257 4279 24500 4512
rect 24257 4097 24501 4279
rect 23819 3773 25011 4097
rect 25715 4067 26553 4760
rect 27613 4067 28451 4760
rect 29682 4557 30874 4803
rect 29682 4545 30875 4557
rect 29683 4233 30875 4545
rect 36399 4080 37213 5857
rect 36689 4079 37213 4080
rect 36889 3606 37213 4079
rect -3668 3411 -2651 3465
rect -3963 3221 -2651 3411
rect -4155 2745 -2651 3221
rect 32076 3055 32573 3512
rect -3963 2627 -2651 2745
rect 31430 2809 34414 3055
rect -3963 2567 -3344 2627
rect -3668 2087 -3344 2567
rect 31430 2488 34415 2809
rect 36889 2713 37213 3154
rect -3670 1397 -3346 1824
rect 29689 1712 30881 1958
rect 31857 1795 32695 2488
rect 33223 2485 34415 2488
rect 29689 1700 30882 1712
rect -3670 1343 -2653 1397
rect -3965 1153 -2653 1343
rect 7799 1282 8991 1594
rect 14353 1287 15545 1599
rect -4155 677 -2653 1153
rect 7798 1270 8991 1282
rect 14352 1275 15545 1287
rect 21002 1275 22194 1587
rect 29690 1388 30882 1700
rect 7798 1024 8990 1270
rect 14352 1029 15544 1275
rect 21001 1263 22194 1275
rect 21001 1017 22193 1263
rect 36399 936 37213 2713
rect 36689 935 37213 936
rect -3965 559 -2653 677
rect -3965 499 -3346 559
rect -3670 19 -3346 499
rect 36889 462 37213 935
<< nmos >>
rect 6125 26783 6185 27183
rect 6243 26783 6303 27183
rect 6478 26983 6538 27183
rect 8123 26709 8183 26909
rect 8241 26709 8301 26909
rect 8359 26709 8419 26909
rect 9265 26713 9325 26913
rect 9383 26713 9443 26913
rect 9501 26713 9561 26913
rect 12638 26780 12698 27180
rect 12756 26780 12816 27180
rect 12991 26980 13051 27180
rect 14636 26706 14696 26906
rect 14754 26706 14814 26906
rect 14872 26706 14932 26906
rect 15778 26710 15838 26910
rect 15896 26710 15956 26910
rect 16014 26710 16074 26910
rect 19172 26775 19232 27175
rect 19290 26775 19350 27175
rect 19525 26975 19585 27175
rect 21170 26701 21230 26901
rect 21288 26701 21348 26901
rect 21406 26701 21466 26901
rect 22312 26705 22372 26905
rect 22430 26705 22490 26905
rect 22548 26705 22608 26905
rect 25730 26779 25790 27179
rect 25848 26779 25908 27179
rect 26083 26979 26143 27179
rect 27728 26705 27788 26905
rect 27846 26705 27906 26905
rect 27964 26705 28024 26905
rect 28870 26709 28930 26909
rect 28988 26709 29048 26909
rect 29106 26709 29166 26909
rect 6139 25133 6199 25533
rect 6257 25133 6317 25533
rect 6492 25333 6552 25533
rect 12652 25130 12712 25530
rect 12770 25130 12830 25530
rect 13005 25330 13065 25530
rect 6134 23529 6194 23929
rect 6252 23529 6312 23929
rect 6487 23729 6547 23929
rect 7491 23928 7551 24128
rect 7911 23728 7971 24128
rect 8029 23728 8089 24128
rect 8147 23728 8207 24128
rect 8265 23728 8325 24128
rect 8789 23928 8849 24128
rect 9389 23928 9449 24128
rect 9809 23728 9869 24128
rect 9927 23728 9987 24128
rect 10045 23728 10105 24128
rect 10163 23728 10223 24128
rect 10687 23928 10747 24128
rect 19186 25125 19246 25525
rect 19304 25125 19364 25525
rect 19539 25325 19599 25525
rect 12647 23526 12707 23926
rect 12765 23526 12825 23926
rect 13000 23726 13060 23926
rect 14004 23925 14064 24125
rect 14424 23725 14484 24125
rect 14542 23725 14602 24125
rect 14660 23725 14720 24125
rect 14778 23725 14838 24125
rect 15302 23925 15362 24125
rect 15902 23925 15962 24125
rect 16322 23725 16382 24125
rect 16440 23725 16500 24125
rect 16558 23725 16618 24125
rect 16676 23725 16736 24125
rect 17200 23925 17260 24125
rect 25744 25129 25804 25529
rect 25862 25129 25922 25529
rect 26097 25329 26157 25529
rect 19181 23521 19241 23921
rect 19299 23521 19359 23921
rect 19534 23721 19594 23921
rect 20538 23920 20598 24120
rect 20958 23720 21018 24120
rect 21076 23720 21136 24120
rect 21194 23720 21254 24120
rect 21312 23720 21372 24120
rect 21836 23920 21896 24120
rect 22436 23920 22496 24120
rect 22856 23720 22916 24120
rect 22974 23720 23034 24120
rect 23092 23720 23152 24120
rect 23210 23720 23270 24120
rect 23734 23920 23794 24120
rect 25739 23525 25799 23925
rect 25857 23525 25917 23925
rect 26092 23725 26152 23925
rect 27096 23924 27156 24124
rect 27516 23724 27576 24124
rect 27634 23724 27694 24124
rect 27752 23724 27812 24124
rect 27870 23724 27930 24124
rect 28394 23924 28454 24124
rect 28994 23924 29054 24124
rect 29414 23724 29474 24124
rect 29532 23724 29592 24124
rect 29650 23724 29710 24124
rect 29768 23724 29828 24124
rect 30292 23924 30352 24124
rect 38088 24208 38288 24268
rect 38088 24016 38488 24076
rect 38088 23898 38488 23958
rect 38088 23780 38488 23840
rect 38088 23662 38488 23722
rect 38088 23466 38288 23526
rect 6343 21105 6403 21305
rect 6461 21105 6521 21305
rect 6579 21105 6639 21305
rect 9366 21375 9426 21575
rect 7485 21101 7545 21301
rect 7603 21101 7663 21301
rect 7721 21101 7781 21301
rect 9601 21175 9661 21575
rect 9719 21175 9779 21575
rect 12901 21101 12961 21301
rect 13019 21101 13079 21301
rect 13137 21101 13197 21301
rect 15924 21371 15984 21571
rect 14043 21097 14103 21297
rect 14161 21097 14221 21297
rect 14279 21097 14339 21297
rect 16159 21171 16219 21571
rect 16277 21171 16337 21571
rect 19435 21106 19495 21306
rect 19553 21106 19613 21306
rect 19671 21106 19731 21306
rect 22458 21376 22518 21576
rect 20577 21102 20637 21302
rect 20695 21102 20755 21302
rect 20813 21102 20873 21302
rect 22693 21176 22753 21576
rect 22811 21176 22871 21576
rect 25948 21109 26008 21309
rect 26066 21109 26126 21309
rect 26184 21109 26244 21309
rect 28971 21379 29031 21579
rect 27090 21105 27150 21305
rect 27208 21105 27268 21305
rect 27326 21105 27386 21305
rect 29206 21179 29266 21579
rect 29324 21179 29384 21579
rect 38088 21064 38288 21124
rect 38088 20872 38488 20932
rect 38088 20754 38488 20814
rect 38088 20636 38488 20696
rect 38088 20518 38488 20578
rect 9352 19725 9412 19925
rect 9587 19525 9647 19925
rect 9705 19525 9765 19925
rect 15910 19721 15970 19921
rect 5157 18320 5217 18520
rect 5681 18120 5741 18520
rect 5799 18120 5859 18520
rect 5917 18120 5977 18520
rect 6035 18120 6095 18520
rect 6455 18320 6515 18520
rect 7055 18320 7115 18520
rect 7579 18120 7639 18520
rect 7697 18120 7757 18520
rect 7815 18120 7875 18520
rect 7933 18120 7993 18520
rect 8353 18320 8413 18520
rect 16145 19521 16205 19921
rect 16263 19521 16323 19921
rect 22444 19726 22504 19926
rect 9357 18121 9417 18321
rect 9592 17921 9652 18321
rect 9710 17921 9770 18321
rect 11715 18316 11775 18516
rect 12239 18116 12299 18516
rect 12357 18116 12417 18516
rect 12475 18116 12535 18516
rect 12593 18116 12653 18516
rect 13013 18316 13073 18516
rect 13613 18316 13673 18516
rect 14137 18116 14197 18516
rect 14255 18116 14315 18516
rect 14373 18116 14433 18516
rect 14491 18116 14551 18516
rect 14911 18316 14971 18516
rect 22679 19526 22739 19926
rect 22797 19526 22857 19926
rect 38088 20322 38288 20382
rect 28957 19729 29017 19929
rect 18249 18321 18309 18521
rect 15915 18117 15975 18317
rect 16150 17917 16210 18317
rect 16268 17917 16328 18317
rect 18773 18121 18833 18521
rect 18891 18121 18951 18521
rect 19009 18121 19069 18521
rect 19127 18121 19187 18521
rect 19547 18321 19607 18521
rect 20147 18321 20207 18521
rect 20671 18121 20731 18521
rect 20789 18121 20849 18521
rect 20907 18121 20967 18521
rect 21025 18121 21085 18521
rect 21445 18321 21505 18521
rect 29192 19529 29252 19929
rect 29310 19529 29370 19929
rect 24762 18324 24822 18524
rect 22449 18122 22509 18322
rect 22684 17922 22744 18322
rect 22802 17922 22862 18322
rect 25286 18124 25346 18524
rect 25404 18124 25464 18524
rect 25522 18124 25582 18524
rect 25640 18124 25700 18524
rect 26060 18324 26120 18524
rect 26660 18324 26720 18524
rect 27184 18124 27244 18524
rect 27302 18124 27362 18524
rect 27420 18124 27480 18524
rect 27538 18124 27598 18524
rect 27958 18324 28018 18524
rect 28962 18125 29022 18325
rect 29197 17925 29257 18325
rect 29315 17925 29375 18325
rect 38084 17932 38284 17992
rect 38084 17740 38484 17800
rect 38084 17622 38484 17682
rect 38084 17504 38484 17564
rect 38084 17386 38484 17446
rect 38084 17190 38284 17250
rect -2379 16024 -2179 16084
rect -2379 15604 -1979 15664
rect -2379 15486 -1979 15546
rect -2379 15368 -1979 15428
rect -2379 15250 -1979 15310
rect -2379 14726 -2179 14786
rect 8095 14399 8155 14799
rect 8213 14399 8273 14799
rect 8448 14599 8508 14799
rect 14644 14398 14704 14798
rect 14762 14398 14822 14798
rect 14997 14598 15057 14798
rect 21298 14419 21358 14819
rect 21416 14419 21476 14819
rect 21651 14619 21711 14819
rect 29951 14252 30011 14652
rect 30069 14252 30129 14652
rect 30304 14452 30364 14652
rect 38084 14788 38284 14848
rect 38084 14596 38484 14656
rect -2381 13956 -2181 14016
rect -2381 13536 -1981 13596
rect -2381 13418 -1981 13478
rect -2381 13300 -1981 13360
rect -2381 13182 -1981 13242
rect 38084 14478 38484 14538
rect 38084 14360 38484 14420
rect 33552 13844 33612 14244
rect 33670 13844 33730 14244
rect 33905 14044 33965 14244
rect 38084 14242 38484 14302
rect 38084 14046 38284 14106
rect -2381 12658 -2181 12718
rect 1431 12499 1491 12899
rect 1549 12499 1609 12899
rect 1784 12699 1844 12899
rect 4321 12232 4381 12632
rect 4439 12232 4499 12632
rect 4674 12432 4734 12632
rect 31647 13259 31707 13459
rect 6319 12158 6379 12358
rect 6437 12158 6497 12358
rect 6555 12158 6615 12358
rect 7461 12162 7521 12362
rect 7579 12162 7639 12362
rect 7697 12162 7757 12362
rect 10870 12320 10930 12720
rect 10988 12320 11048 12720
rect 11223 12520 11283 12720
rect 12868 12246 12928 12446
rect 12986 12246 13046 12446
rect 13104 12246 13164 12446
rect 14010 12250 14070 12450
rect 14128 12250 14188 12450
rect 14246 12250 14306 12450
rect 17524 12252 17584 12652
rect 17642 12252 17702 12652
rect 17877 12452 17937 12652
rect 32067 13059 32127 13459
rect 32185 13059 32245 13459
rect 32303 13059 32363 13459
rect 32421 13059 32481 13459
rect 32945 13259 33005 13459
rect 19522 12178 19582 12378
rect 19640 12178 19700 12378
rect 19758 12178 19818 12378
rect 20664 12182 20724 12382
rect 20782 12182 20842 12382
rect 20900 12182 20960 12382
rect 24149 12320 24209 12720
rect 24267 12320 24327 12720
rect 24502 12520 24562 12720
rect 26147 12246 26207 12446
rect 26265 12246 26325 12446
rect 26383 12246 26443 12446
rect 27289 12250 27349 12450
rect 27407 12250 27467 12450
rect 27525 12250 27585 12450
rect -2379 11887 -2179 11947
rect 29946 11681 30006 12081
rect 30064 11681 30124 12081
rect 30299 11881 30359 12081
rect -2379 11467 -1979 11527
rect -2379 11349 -1979 11409
rect -2379 11231 -1979 11291
rect -2379 11113 -1979 11173
rect 38088 11586 38288 11646
rect 38088 11394 38488 11454
rect -2379 10589 -2179 10649
rect 4335 10582 4395 10982
rect 4453 10582 4513 10982
rect 4688 10782 4748 10982
rect 10884 10670 10944 11070
rect 11002 10670 11062 11070
rect 11237 10870 11297 11070
rect 1423 9914 1483 10314
rect 1541 9914 1601 10314
rect 1776 10114 1836 10314
rect -2381 9819 -2181 9879
rect -2381 9399 -1981 9459
rect 38088 11276 38488 11336
rect 38088 11158 38488 11218
rect -2381 9281 -1981 9341
rect -2381 9163 -1981 9223
rect -2381 9045 -1981 9105
rect 4330 8978 4390 9378
rect 4448 8978 4508 9378
rect 4683 9178 4743 9378
rect 5687 9377 5747 9577
rect 6107 9177 6167 9577
rect 6225 9177 6285 9577
rect 6343 9177 6403 9577
rect 6461 9177 6521 9577
rect 6985 9377 7045 9577
rect 7585 9377 7645 9577
rect 8005 9177 8065 9577
rect 8123 9177 8183 9577
rect 8241 9177 8301 9577
rect 8359 9177 8419 9577
rect 8883 9377 8943 9577
rect 17538 10602 17598 11002
rect 17656 10602 17716 11002
rect 17891 10802 17951 11002
rect 24163 10670 24223 11070
rect 24281 10670 24341 11070
rect 24516 10870 24576 11070
rect 10879 9066 10939 9466
rect 10997 9066 11057 9466
rect 11232 9266 11292 9466
rect 12236 9465 12296 9665
rect 12656 9265 12716 9665
rect 12774 9265 12834 9665
rect 12892 9265 12952 9665
rect 13010 9265 13070 9665
rect 13534 9465 13594 9665
rect 14134 9465 14194 9665
rect 14554 9265 14614 9665
rect 14672 9265 14732 9665
rect 14790 9265 14850 9665
rect 14908 9265 14968 9665
rect 15432 9465 15492 9665
rect 38088 11040 38488 11100
rect 17533 8998 17593 9398
rect 17651 8998 17711 9398
rect 17886 9198 17946 9398
rect 18890 9397 18950 9597
rect 19310 9197 19370 9597
rect 19428 9197 19488 9597
rect 19546 9197 19606 9597
rect 19664 9197 19724 9597
rect 20188 9397 20248 9597
rect 20788 9397 20848 9597
rect 21208 9197 21268 9597
rect 21326 9197 21386 9597
rect 21444 9197 21504 9597
rect 21562 9197 21622 9597
rect 22086 9397 22146 9597
rect 38088 10844 38288 10904
rect 24158 9066 24218 9466
rect 24276 9066 24336 9466
rect 24511 9266 24571 9466
rect 25515 9465 25575 9665
rect 25935 9265 25995 9665
rect 26053 9265 26113 9665
rect 26171 9265 26231 9665
rect 26289 9265 26349 9665
rect 26813 9465 26873 9665
rect 27413 9465 27473 9665
rect 27833 9265 27893 9665
rect 27951 9265 28011 9665
rect 28069 9265 28129 9665
rect 28187 9265 28247 9665
rect 28711 9465 28771 9665
rect 33554 9753 33614 10153
rect 33672 9753 33732 10153
rect 33907 9953 33967 10153
rect 31649 9168 31709 9368
rect 29946 8648 30006 9048
rect 30064 8648 30124 9048
rect 30299 8848 30359 9048
rect 32069 8968 32129 9368
rect 32187 8968 32247 9368
rect 32305 8968 32365 9368
rect 32423 8968 32483 9368
rect 32947 9168 33007 9368
rect -2381 8521 -2181 8581
rect 38088 8442 38288 8502
rect 38088 8250 38488 8310
rect 38088 8132 38488 8192
rect 38088 8014 38488 8074
rect 38088 7896 38488 7956
rect -2381 7750 -2181 7810
rect -2381 7330 -1981 7390
rect -2381 7212 -1981 7272
rect -2381 7094 -1981 7154
rect -2381 6976 -1981 7036
rect 1404 6636 1464 7036
rect 1522 6636 1582 7036
rect 1757 6836 1817 7036
rect -2381 6452 -2181 6512
rect 4313 6452 4373 6852
rect 4431 6452 4491 6852
rect 4666 6652 4726 6852
rect 6311 6378 6371 6578
rect 6429 6378 6489 6578
rect 6547 6378 6607 6578
rect 7453 6382 7513 6582
rect 7571 6382 7631 6582
rect 7689 6382 7749 6582
rect 10864 6450 10924 6850
rect 10982 6450 11042 6850
rect 11217 6650 11277 6850
rect 38088 7700 38288 7760
rect 12862 6376 12922 6576
rect 12980 6376 13040 6576
rect 13098 6376 13158 6576
rect 14004 6380 14064 6580
rect 14122 6380 14182 6580
rect 14240 6380 14300 6580
rect 17519 6451 17579 6851
rect 17637 6451 17697 6851
rect 17872 6651 17932 6851
rect 19517 6377 19577 6577
rect 19635 6377 19695 6577
rect 19753 6377 19813 6577
rect 20659 6381 20719 6581
rect 20777 6381 20837 6581
rect 20895 6381 20955 6581
rect 24141 6452 24201 6852
rect 24259 6452 24319 6852
rect 24494 6652 24554 6852
rect 30017 6728 30077 7128
rect 30135 6728 30195 7128
rect 30370 6928 30430 7128
rect 26139 6378 26199 6578
rect 26257 6378 26317 6578
rect 26375 6378 26435 6578
rect 27281 6382 27341 6582
rect 27399 6382 27459 6582
rect 27517 6382 27577 6582
rect 33554 6258 33614 6658
rect 33672 6258 33732 6658
rect 33907 6458 33967 6658
rect -2383 5682 -2183 5742
rect -2383 5262 -1983 5322
rect -2383 5144 -1983 5204
rect 31649 5673 31709 5873
rect 32069 5473 32129 5873
rect 32187 5473 32247 5873
rect 32305 5473 32365 5873
rect 32423 5473 32483 5873
rect 32947 5673 33007 5873
rect -2383 5026 -1983 5086
rect -2383 4908 -1983 4968
rect 4327 4802 4387 5202
rect 4445 4802 4505 5202
rect 4680 5002 4740 5202
rect -2383 4384 -2183 4444
rect 1420 3876 1480 4276
rect 1538 3876 1598 4276
rect 1773 4076 1833 4276
rect -2381 3613 -2181 3673
rect 10878 4800 10938 5200
rect 10996 4800 11056 5200
rect 11231 5000 11291 5200
rect -2381 3193 -1981 3253
rect 4322 3198 4382 3598
rect 4440 3198 4500 3598
rect 4675 3398 4735 3598
rect 5679 3597 5739 3797
rect 6099 3397 6159 3797
rect 6217 3397 6277 3797
rect 6335 3397 6395 3797
rect 6453 3397 6513 3797
rect 6977 3597 7037 3797
rect 7577 3597 7637 3797
rect 7997 3397 8057 3797
rect 8115 3397 8175 3797
rect 8233 3397 8293 3797
rect 8351 3397 8411 3797
rect 8875 3597 8935 3797
rect 17533 4801 17593 5201
rect 17651 4801 17711 5201
rect 17886 5001 17946 5201
rect -2381 3075 -1981 3135
rect 10873 3196 10933 3596
rect 10991 3196 11051 3596
rect 11226 3396 11286 3596
rect 12230 3595 12290 3795
rect 12650 3395 12710 3795
rect 12768 3395 12828 3795
rect 12886 3395 12946 3795
rect 13004 3395 13064 3795
rect 13528 3595 13588 3795
rect 14128 3595 14188 3795
rect 14548 3395 14608 3795
rect 14666 3395 14726 3795
rect 14784 3395 14844 3795
rect 14902 3395 14962 3795
rect 15426 3595 15486 3795
rect 24155 4802 24215 5202
rect 24273 4802 24333 5202
rect 24508 5002 24568 5202
rect 38084 5310 38284 5370
rect 38084 5118 38484 5178
rect 38084 5000 38484 5060
rect -2381 2957 -1981 3017
rect 17528 3197 17588 3597
rect 17646 3197 17706 3597
rect 17881 3397 17941 3597
rect 18885 3596 18945 3796
rect 19305 3396 19365 3796
rect 19423 3396 19483 3796
rect 19541 3396 19601 3796
rect 19659 3396 19719 3796
rect 20183 3596 20243 3796
rect 20783 3596 20843 3796
rect 21203 3396 21263 3796
rect 21321 3396 21381 3796
rect 21439 3396 21499 3796
rect 21557 3396 21617 3796
rect 22081 3596 22141 3796
rect 38084 4882 38484 4942
rect 38084 4764 38484 4824
rect 38084 4568 38284 4628
rect 24150 3198 24210 3598
rect 24268 3198 24328 3598
rect 24503 3398 24563 3598
rect 25507 3597 25567 3797
rect 25927 3397 25987 3797
rect 26045 3397 26105 3797
rect 26163 3397 26223 3797
rect 26281 3397 26341 3797
rect 26805 3597 26865 3797
rect 27405 3597 27465 3797
rect 27825 3397 27885 3797
rect 27943 3397 28003 3797
rect 28061 3397 28121 3797
rect 28179 3397 28239 3797
rect 28703 3597 28763 3797
rect 30014 3658 30074 4058
rect 30132 3658 30192 4058
rect 30367 3858 30427 4058
rect -2381 2839 -1981 2899
rect -2381 2315 -2181 2375
rect 8130 1769 8190 2169
rect 8248 1769 8308 2169
rect 8483 1769 8543 1969
rect 14684 1774 14744 2174
rect 14802 1774 14862 2174
rect 15037 1774 15097 1974
rect -2383 1545 -2183 1605
rect 21333 1762 21393 2162
rect 21451 1762 21511 2162
rect 21686 1762 21746 1962
rect 33554 1910 33614 2310
rect 33672 1910 33732 2310
rect 33907 2110 33967 2310
rect 38084 2166 38284 2226
rect 38084 1974 38484 2034
rect 38084 1856 38484 1916
rect 38084 1738 38484 1798
rect 38084 1620 38484 1680
rect 31649 1325 31709 1525
rect -2383 1125 -1983 1185
rect -2383 1007 -1983 1067
rect -2383 889 -1983 949
rect -2383 771 -1983 831
rect 30021 813 30081 1213
rect 30139 813 30199 1213
rect 30374 1013 30434 1213
rect 32069 1125 32129 1525
rect 32187 1125 32247 1525
rect 32305 1125 32365 1525
rect 32423 1125 32483 1525
rect 32947 1325 33007 1525
rect 38084 1424 38284 1484
rect -2383 247 -2183 307
<< pmos >>
rect 5888 27420 5948 27620
rect 6006 27420 6066 27620
rect 6124 27420 6184 27620
rect 6242 27420 6302 27620
rect 6360 27420 6420 27620
rect 6478 27420 6538 27620
rect 6596 27420 6656 27620
rect 6714 27420 6774 27620
rect 6832 27420 6892 27620
rect 8213 27292 8273 27692
rect 8331 27292 8391 27692
rect 8449 27292 8509 27692
rect 8567 27292 8627 27692
rect 8685 27292 8745 27692
rect 8803 27292 8863 27692
rect 9355 27296 9415 27696
rect 9473 27296 9533 27696
rect 9591 27296 9651 27696
rect 9709 27296 9769 27696
rect 9827 27296 9887 27696
rect 9945 27296 10005 27696
rect 12401 27417 12461 27617
rect 12519 27417 12579 27617
rect 12637 27417 12697 27617
rect 12755 27417 12815 27617
rect 12873 27417 12933 27617
rect 12991 27417 13051 27617
rect 13109 27417 13169 27617
rect 13227 27417 13287 27617
rect 13345 27417 13405 27617
rect 14726 27289 14786 27689
rect 14844 27289 14904 27689
rect 14962 27289 15022 27689
rect 15080 27289 15140 27689
rect 15198 27289 15258 27689
rect 15316 27289 15376 27689
rect 15868 27293 15928 27693
rect 15986 27293 16046 27693
rect 16104 27293 16164 27693
rect 16222 27293 16282 27693
rect 16340 27293 16400 27693
rect 16458 27293 16518 27693
rect 18935 27412 18995 27612
rect 19053 27412 19113 27612
rect 19171 27412 19231 27612
rect 19289 27412 19349 27612
rect 19407 27412 19467 27612
rect 19525 27412 19585 27612
rect 19643 27412 19703 27612
rect 19761 27412 19821 27612
rect 19879 27412 19939 27612
rect 8642 26709 8702 26909
rect 8760 26709 8820 26909
rect 8878 26709 8938 26909
rect 9784 26713 9844 26913
rect 9902 26713 9962 26913
rect 10020 26713 10080 26913
rect 21260 27284 21320 27684
rect 21378 27284 21438 27684
rect 21496 27284 21556 27684
rect 21614 27284 21674 27684
rect 21732 27284 21792 27684
rect 21850 27284 21910 27684
rect 22402 27288 22462 27688
rect 22520 27288 22580 27688
rect 22638 27288 22698 27688
rect 22756 27288 22816 27688
rect 22874 27288 22934 27688
rect 22992 27288 23052 27688
rect 25493 27416 25553 27616
rect 25611 27416 25671 27616
rect 25729 27416 25789 27616
rect 25847 27416 25907 27616
rect 25965 27416 26025 27616
rect 26083 27416 26143 27616
rect 26201 27416 26261 27616
rect 26319 27416 26379 27616
rect 26437 27416 26497 27616
rect 15155 26706 15215 26906
rect 15273 26706 15333 26906
rect 15391 26706 15451 26906
rect 16297 26710 16357 26910
rect 16415 26710 16475 26910
rect 16533 26710 16593 26910
rect 27818 27288 27878 27688
rect 27936 27288 27996 27688
rect 28054 27288 28114 27688
rect 28172 27288 28232 27688
rect 28290 27288 28350 27688
rect 28408 27288 28468 27688
rect 28960 27292 29020 27692
rect 29078 27292 29138 27692
rect 29196 27292 29256 27692
rect 29314 27292 29374 27692
rect 29432 27292 29492 27692
rect 29550 27292 29610 27692
rect 21689 26701 21749 26901
rect 21807 26701 21867 26901
rect 21925 26701 21985 26901
rect 22831 26705 22891 26905
rect 22949 26705 23009 26905
rect 23067 26705 23127 26905
rect 28247 26705 28307 26905
rect 28365 26705 28425 26905
rect 28483 26705 28543 26905
rect 29389 26709 29449 26909
rect 29507 26709 29567 26909
rect 29625 26709 29685 26909
rect 5902 25770 5962 25970
rect 6020 25770 6080 25970
rect 6138 25770 6198 25970
rect 6256 25770 6316 25970
rect 6374 25770 6434 25970
rect 6492 25770 6552 25970
rect 6610 25770 6670 25970
rect 6728 25770 6788 25970
rect 6846 25770 6906 25970
rect 12415 25767 12475 25967
rect 12533 25767 12593 25967
rect 12651 25767 12711 25967
rect 12769 25767 12829 25967
rect 12887 25767 12947 25967
rect 13005 25767 13065 25967
rect 13123 25767 13183 25967
rect 13241 25767 13301 25967
rect 13359 25767 13419 25967
rect 7366 25153 7426 25353
rect 7484 25153 7544 25353
rect 7602 25153 7662 25353
rect 7850 25153 7910 25553
rect 7968 25153 8028 25553
rect 8086 25153 8146 25553
rect 8204 25153 8264 25553
rect 8322 25153 8382 25553
rect 8440 25153 8500 25553
rect 8687 25153 8747 25353
rect 8805 25153 8865 25353
rect 8923 25153 8983 25353
rect 9264 25153 9324 25353
rect 9382 25153 9442 25353
rect 9500 25153 9560 25353
rect 9748 25153 9808 25553
rect 9866 25153 9926 25553
rect 9984 25153 10044 25553
rect 10102 25153 10162 25553
rect 10220 25153 10280 25553
rect 10338 25153 10398 25553
rect 18949 25762 19009 25962
rect 19067 25762 19127 25962
rect 19185 25762 19245 25962
rect 19303 25762 19363 25962
rect 19421 25762 19481 25962
rect 19539 25762 19599 25962
rect 19657 25762 19717 25962
rect 19775 25762 19835 25962
rect 19893 25762 19953 25962
rect 25507 25766 25567 25966
rect 25625 25766 25685 25966
rect 25743 25766 25803 25966
rect 25861 25766 25921 25966
rect 25979 25766 26039 25966
rect 26097 25766 26157 25966
rect 26215 25766 26275 25966
rect 26333 25766 26393 25966
rect 26451 25766 26511 25966
rect 10585 25153 10645 25353
rect 10703 25153 10763 25353
rect 10821 25153 10881 25353
rect 5897 24166 5957 24366
rect 6015 24166 6075 24366
rect 6133 24166 6193 24366
rect 6251 24166 6311 24366
rect 6369 24166 6429 24366
rect 6487 24166 6547 24366
rect 6605 24166 6665 24366
rect 6723 24166 6783 24366
rect 6841 24166 6901 24366
rect 7793 24460 7853 24860
rect 7911 24460 7971 24860
rect 8029 24460 8089 24860
rect 8147 24460 8207 24860
rect 8265 24460 8325 24860
rect 8383 24460 8443 24860
rect 13879 25150 13939 25350
rect 13997 25150 14057 25350
rect 14115 25150 14175 25350
rect 14363 25150 14423 25550
rect 14481 25150 14541 25550
rect 14599 25150 14659 25550
rect 14717 25150 14777 25550
rect 14835 25150 14895 25550
rect 14953 25150 15013 25550
rect 15200 25150 15260 25350
rect 15318 25150 15378 25350
rect 15436 25150 15496 25350
rect 15777 25150 15837 25350
rect 15895 25150 15955 25350
rect 16013 25150 16073 25350
rect 16261 25150 16321 25550
rect 16379 25150 16439 25550
rect 16497 25150 16557 25550
rect 16615 25150 16675 25550
rect 16733 25150 16793 25550
rect 16851 25150 16911 25550
rect 17098 25150 17158 25350
rect 17216 25150 17276 25350
rect 17334 25150 17394 25350
rect 9691 24460 9751 24860
rect 9809 24460 9869 24860
rect 9927 24460 9987 24860
rect 10045 24460 10105 24860
rect 10163 24460 10223 24860
rect 10281 24460 10341 24860
rect 12410 24163 12470 24363
rect 12528 24163 12588 24363
rect 12646 24163 12706 24363
rect 12764 24163 12824 24363
rect 12882 24163 12942 24363
rect 13000 24163 13060 24363
rect 13118 24163 13178 24363
rect 13236 24163 13296 24363
rect 13354 24163 13414 24363
rect 14306 24457 14366 24857
rect 14424 24457 14484 24857
rect 14542 24457 14602 24857
rect 14660 24457 14720 24857
rect 14778 24457 14838 24857
rect 14896 24457 14956 24857
rect 20413 25145 20473 25345
rect 20531 25145 20591 25345
rect 20649 25145 20709 25345
rect 20897 25145 20957 25545
rect 21015 25145 21075 25545
rect 21133 25145 21193 25545
rect 21251 25145 21311 25545
rect 21369 25145 21429 25545
rect 21487 25145 21547 25545
rect 21734 25145 21794 25345
rect 21852 25145 21912 25345
rect 21970 25145 22030 25345
rect 22311 25145 22371 25345
rect 22429 25145 22489 25345
rect 22547 25145 22607 25345
rect 22795 25145 22855 25545
rect 22913 25145 22973 25545
rect 23031 25145 23091 25545
rect 23149 25145 23209 25545
rect 23267 25145 23327 25545
rect 23385 25145 23445 25545
rect 23632 25145 23692 25345
rect 23750 25145 23810 25345
rect 23868 25145 23928 25345
rect 16204 24457 16264 24857
rect 16322 24457 16382 24857
rect 16440 24457 16500 24857
rect 16558 24457 16618 24857
rect 16676 24457 16736 24857
rect 16794 24457 16854 24857
rect 18944 24158 19004 24358
rect 19062 24158 19122 24358
rect 19180 24158 19240 24358
rect 19298 24158 19358 24358
rect 19416 24158 19476 24358
rect 19534 24158 19594 24358
rect 19652 24158 19712 24358
rect 19770 24158 19830 24358
rect 19888 24158 19948 24358
rect 20840 24452 20900 24852
rect 20958 24452 21018 24852
rect 21076 24452 21136 24852
rect 21194 24452 21254 24852
rect 21312 24452 21372 24852
rect 21430 24452 21490 24852
rect 26971 25149 27031 25349
rect 27089 25149 27149 25349
rect 27207 25149 27267 25349
rect 27455 25149 27515 25549
rect 27573 25149 27633 25549
rect 27691 25149 27751 25549
rect 27809 25149 27869 25549
rect 27927 25149 27987 25549
rect 28045 25149 28105 25549
rect 28292 25149 28352 25349
rect 28410 25149 28470 25349
rect 28528 25149 28588 25349
rect 28869 25149 28929 25349
rect 28987 25149 29047 25349
rect 29105 25149 29165 25349
rect 29353 25149 29413 25549
rect 29471 25149 29531 25549
rect 29589 25149 29649 25549
rect 29707 25149 29767 25549
rect 29825 25149 29885 25549
rect 29943 25149 30003 25549
rect 30190 25149 30250 25349
rect 30308 25149 30368 25349
rect 30426 25149 30486 25349
rect 22738 24452 22798 24852
rect 22856 24452 22916 24852
rect 22974 24452 23034 24852
rect 23092 24452 23152 24852
rect 23210 24452 23270 24852
rect 23328 24452 23388 24852
rect 25502 24162 25562 24362
rect 25620 24162 25680 24362
rect 25738 24162 25798 24362
rect 25856 24162 25916 24362
rect 25974 24162 26034 24362
rect 26092 24162 26152 24362
rect 26210 24162 26270 24362
rect 26328 24162 26388 24362
rect 26446 24162 26506 24362
rect 27398 24456 27458 24856
rect 27516 24456 27576 24856
rect 27634 24456 27694 24856
rect 27752 24456 27812 24856
rect 27870 24456 27930 24856
rect 27988 24456 28048 24856
rect 36955 25042 37155 25102
rect 29296 24456 29356 24856
rect 29414 24456 29474 24856
rect 29532 24456 29592 24856
rect 29650 24456 29710 24856
rect 29768 24456 29828 24856
rect 29886 24456 29946 24856
rect 36955 24924 37155 24984
rect 36955 24806 37155 24866
rect 36755 24601 37155 24661
rect 36755 24483 37155 24543
rect 36755 24365 37155 24425
rect 36755 24134 37155 24194
rect 36755 24016 37155 24076
rect 36755 23898 37155 23958
rect 36755 23780 37155 23840
rect 36755 23662 37155 23722
rect 36755 23544 37155 23604
rect 36755 23307 37155 23367
rect 36755 23189 37155 23249
rect 36755 23071 37155 23131
rect 36955 22834 37155 22894
rect 36955 22716 37155 22776
rect 36955 22598 37155 22658
rect 5899 21688 5959 22088
rect 6017 21688 6077 22088
rect 6135 21688 6195 22088
rect 6253 21688 6313 22088
rect 6371 21688 6431 22088
rect 6489 21688 6549 22088
rect 7041 21684 7101 22084
rect 7159 21684 7219 22084
rect 7277 21684 7337 22084
rect 7395 21684 7455 22084
rect 7513 21684 7573 22084
rect 7631 21684 7691 22084
rect 9012 21812 9072 22012
rect 9130 21812 9190 22012
rect 9248 21812 9308 22012
rect 9366 21812 9426 22012
rect 9484 21812 9544 22012
rect 9602 21812 9662 22012
rect 9720 21812 9780 22012
rect 9838 21812 9898 22012
rect 9956 21812 10016 22012
rect 12457 21684 12517 22084
rect 12575 21684 12635 22084
rect 12693 21684 12753 22084
rect 12811 21684 12871 22084
rect 12929 21684 12989 22084
rect 13047 21684 13107 22084
rect 5824 21105 5884 21305
rect 5942 21105 6002 21305
rect 6060 21105 6120 21305
rect 6966 21101 7026 21301
rect 7084 21101 7144 21301
rect 7202 21101 7262 21301
rect 13599 21680 13659 22080
rect 13717 21680 13777 22080
rect 13835 21680 13895 22080
rect 13953 21680 14013 22080
rect 14071 21680 14131 22080
rect 14189 21680 14249 22080
rect 15570 21808 15630 22008
rect 15688 21808 15748 22008
rect 15806 21808 15866 22008
rect 15924 21808 15984 22008
rect 16042 21808 16102 22008
rect 16160 21808 16220 22008
rect 16278 21808 16338 22008
rect 16396 21808 16456 22008
rect 16514 21808 16574 22008
rect 18991 21689 19051 22089
rect 19109 21689 19169 22089
rect 19227 21689 19287 22089
rect 19345 21689 19405 22089
rect 19463 21689 19523 22089
rect 19581 21689 19641 22089
rect 12382 21101 12442 21301
rect 12500 21101 12560 21301
rect 12618 21101 12678 21301
rect 13524 21097 13584 21297
rect 13642 21097 13702 21297
rect 13760 21097 13820 21297
rect 20133 21685 20193 22085
rect 20251 21685 20311 22085
rect 20369 21685 20429 22085
rect 20487 21685 20547 22085
rect 20605 21685 20665 22085
rect 20723 21685 20783 22085
rect 22104 21813 22164 22013
rect 22222 21813 22282 22013
rect 22340 21813 22400 22013
rect 22458 21813 22518 22013
rect 22576 21813 22636 22013
rect 22694 21813 22754 22013
rect 22812 21813 22872 22013
rect 22930 21813 22990 22013
rect 23048 21813 23108 22013
rect 25504 21692 25564 22092
rect 25622 21692 25682 22092
rect 25740 21692 25800 22092
rect 25858 21692 25918 22092
rect 25976 21692 26036 22092
rect 26094 21692 26154 22092
rect 18916 21106 18976 21306
rect 19034 21106 19094 21306
rect 19152 21106 19212 21306
rect 20058 21102 20118 21302
rect 20176 21102 20236 21302
rect 20294 21102 20354 21302
rect 26646 21688 26706 22088
rect 26764 21688 26824 22088
rect 26882 21688 26942 22088
rect 27000 21688 27060 22088
rect 27118 21688 27178 22088
rect 27236 21688 27296 22088
rect 28617 21816 28677 22016
rect 28735 21816 28795 22016
rect 28853 21816 28913 22016
rect 28971 21816 29031 22016
rect 29089 21816 29149 22016
rect 29207 21816 29267 22016
rect 29325 21816 29385 22016
rect 29443 21816 29503 22016
rect 29561 21816 29621 22016
rect 36955 21898 37155 21958
rect 36955 21780 37155 21840
rect 36955 21662 37155 21722
rect 25429 21109 25489 21309
rect 25547 21109 25607 21309
rect 25665 21109 25725 21309
rect 26571 21105 26631 21305
rect 26689 21105 26749 21305
rect 26807 21105 26867 21305
rect 36755 21457 37155 21517
rect 36755 21339 37155 21399
rect 36755 21221 37155 21281
rect 36755 20990 37155 21050
rect 36755 20872 37155 20932
rect 36755 20754 37155 20814
rect 36755 20636 37155 20696
rect 36755 20518 37155 20578
rect 8998 20162 9058 20362
rect 9116 20162 9176 20362
rect 9234 20162 9294 20362
rect 9352 20162 9412 20362
rect 9470 20162 9530 20362
rect 9588 20162 9648 20362
rect 9706 20162 9766 20362
rect 9824 20162 9884 20362
rect 9942 20162 10002 20362
rect 15556 20158 15616 20358
rect 15674 20158 15734 20358
rect 15792 20158 15852 20358
rect 15910 20158 15970 20358
rect 16028 20158 16088 20358
rect 16146 20158 16206 20358
rect 16264 20158 16324 20358
rect 16382 20158 16442 20358
rect 16500 20158 16560 20358
rect 22090 20163 22150 20363
rect 22208 20163 22268 20363
rect 22326 20163 22386 20363
rect 22444 20163 22504 20363
rect 22562 20163 22622 20363
rect 22680 20163 22740 20363
rect 22798 20163 22858 20363
rect 22916 20163 22976 20363
rect 23034 20163 23094 20363
rect 36755 20400 37155 20460
rect 28603 20166 28663 20366
rect 28721 20166 28781 20366
rect 28839 20166 28899 20366
rect 28957 20166 29017 20366
rect 29075 20166 29135 20366
rect 29193 20166 29253 20366
rect 29311 20166 29371 20366
rect 29429 20166 29489 20366
rect 29547 20166 29607 20366
rect 5023 19545 5083 19745
rect 5141 19545 5201 19745
rect 5259 19545 5319 19745
rect 5506 19545 5566 19945
rect 5624 19545 5684 19945
rect 5742 19545 5802 19945
rect 5860 19545 5920 19945
rect 5978 19545 6038 19945
rect 6096 19545 6156 19945
rect 6344 19545 6404 19745
rect 6462 19545 6522 19745
rect 6580 19545 6640 19745
rect 6921 19545 6981 19745
rect 7039 19545 7099 19745
rect 7157 19545 7217 19745
rect 7404 19545 7464 19945
rect 7522 19545 7582 19945
rect 7640 19545 7700 19945
rect 7758 19545 7818 19945
rect 7876 19545 7936 19945
rect 7994 19545 8054 19945
rect 8242 19545 8302 19745
rect 8360 19545 8420 19745
rect 8478 19545 8538 19745
rect 5563 18852 5623 19252
rect 5681 18852 5741 19252
rect 5799 18852 5859 19252
rect 5917 18852 5977 19252
rect 6035 18852 6095 19252
rect 6153 18852 6213 19252
rect 11581 19541 11641 19741
rect 11699 19541 11759 19741
rect 11817 19541 11877 19741
rect 12064 19541 12124 19941
rect 12182 19541 12242 19941
rect 12300 19541 12360 19941
rect 12418 19541 12478 19941
rect 12536 19541 12596 19941
rect 12654 19541 12714 19941
rect 12902 19541 12962 19741
rect 13020 19541 13080 19741
rect 13138 19541 13198 19741
rect 13479 19541 13539 19741
rect 13597 19541 13657 19741
rect 13715 19541 13775 19741
rect 13962 19541 14022 19941
rect 14080 19541 14140 19941
rect 14198 19541 14258 19941
rect 14316 19541 14376 19941
rect 14434 19541 14494 19941
rect 14552 19541 14612 19941
rect 14800 19541 14860 19741
rect 14918 19541 14978 19741
rect 15036 19541 15096 19741
rect 7461 18852 7521 19252
rect 7579 18852 7639 19252
rect 7697 18852 7757 19252
rect 7815 18852 7875 19252
rect 7933 18852 7993 19252
rect 8051 18852 8111 19252
rect 9003 18558 9063 18758
rect 9121 18558 9181 18758
rect 9239 18558 9299 18758
rect 9357 18558 9417 18758
rect 9475 18558 9535 18758
rect 9593 18558 9653 18758
rect 9711 18558 9771 18758
rect 9829 18558 9889 18758
rect 9947 18558 10007 18758
rect 12121 18848 12181 19248
rect 12239 18848 12299 19248
rect 12357 18848 12417 19248
rect 12475 18848 12535 19248
rect 12593 18848 12653 19248
rect 12711 18848 12771 19248
rect 18115 19546 18175 19746
rect 18233 19546 18293 19746
rect 18351 19546 18411 19746
rect 18598 19546 18658 19946
rect 18716 19546 18776 19946
rect 18834 19546 18894 19946
rect 18952 19546 19012 19946
rect 19070 19546 19130 19946
rect 19188 19546 19248 19946
rect 19436 19546 19496 19746
rect 19554 19546 19614 19746
rect 19672 19546 19732 19746
rect 20013 19546 20073 19746
rect 20131 19546 20191 19746
rect 20249 19546 20309 19746
rect 20496 19546 20556 19946
rect 20614 19546 20674 19946
rect 20732 19546 20792 19946
rect 20850 19546 20910 19946
rect 20968 19546 21028 19946
rect 21086 19546 21146 19946
rect 36755 20163 37155 20223
rect 21334 19546 21394 19746
rect 21452 19546 21512 19746
rect 21570 19546 21630 19746
rect 14019 18848 14079 19248
rect 14137 18848 14197 19248
rect 14255 18848 14315 19248
rect 14373 18848 14433 19248
rect 14491 18848 14551 19248
rect 14609 18848 14669 19248
rect 15561 18554 15621 18754
rect 15679 18554 15739 18754
rect 15797 18554 15857 18754
rect 15915 18554 15975 18754
rect 16033 18554 16093 18754
rect 16151 18554 16211 18754
rect 16269 18554 16329 18754
rect 16387 18554 16447 18754
rect 16505 18554 16565 18754
rect 18655 18853 18715 19253
rect 18773 18853 18833 19253
rect 18891 18853 18951 19253
rect 19009 18853 19069 19253
rect 19127 18853 19187 19253
rect 19245 18853 19305 19253
rect 24628 19549 24688 19749
rect 24746 19549 24806 19749
rect 24864 19549 24924 19749
rect 25111 19549 25171 19949
rect 25229 19549 25289 19949
rect 25347 19549 25407 19949
rect 25465 19549 25525 19949
rect 25583 19549 25643 19949
rect 25701 19549 25761 19949
rect 25949 19549 26009 19749
rect 26067 19549 26127 19749
rect 26185 19549 26245 19749
rect 26526 19549 26586 19749
rect 26644 19549 26704 19749
rect 26762 19549 26822 19749
rect 27009 19549 27069 19949
rect 27127 19549 27187 19949
rect 27245 19549 27305 19949
rect 27363 19549 27423 19949
rect 27481 19549 27541 19949
rect 27599 19549 27659 19949
rect 36755 20045 37155 20105
rect 27847 19549 27907 19749
rect 27965 19549 28025 19749
rect 28083 19549 28143 19749
rect 20553 18853 20613 19253
rect 20671 18853 20731 19253
rect 20789 18853 20849 19253
rect 20907 18853 20967 19253
rect 21025 18853 21085 19253
rect 21143 18853 21203 19253
rect 22095 18559 22155 18759
rect 22213 18559 22273 18759
rect 22331 18559 22391 18759
rect 22449 18559 22509 18759
rect 22567 18559 22627 18759
rect 22685 18559 22745 18759
rect 22803 18559 22863 18759
rect 22921 18559 22981 18759
rect 23039 18559 23099 18759
rect 25168 18856 25228 19256
rect 25286 18856 25346 19256
rect 25404 18856 25464 19256
rect 25522 18856 25582 19256
rect 25640 18856 25700 19256
rect 25758 18856 25818 19256
rect 36755 19927 37155 19987
rect 36955 19690 37155 19750
rect 36955 19572 37155 19632
rect 36955 19454 37155 19514
rect 27066 18856 27126 19256
rect 27184 18856 27244 19256
rect 27302 18856 27362 19256
rect 27420 18856 27480 19256
rect 27538 18856 27598 19256
rect 27656 18856 27716 19256
rect 36951 18766 37151 18826
rect 28608 18562 28668 18762
rect 28726 18562 28786 18762
rect 28844 18562 28904 18762
rect 28962 18562 29022 18762
rect 29080 18562 29140 18762
rect 29198 18562 29258 18762
rect 29316 18562 29376 18762
rect 29434 18562 29494 18762
rect 29552 18562 29612 18762
rect 36951 18648 37151 18708
rect 36951 18530 37151 18590
rect 36751 18325 37151 18385
rect 36751 18207 37151 18267
rect 36751 18089 37151 18149
rect 36751 17858 37151 17918
rect 36751 17740 37151 17800
rect 36751 17622 37151 17682
rect 36751 17504 37151 17564
rect 36751 17386 37151 17446
rect 36751 17268 37151 17328
rect 36751 17031 37151 17091
rect 36751 16913 37151 16973
rect 36751 16795 37151 16855
rect 36951 16558 37151 16618
rect 36951 16440 37151 16500
rect 36951 16322 37151 16382
rect -3604 16149 -3404 16209
rect -3604 16031 -3404 16091
rect -3604 15913 -3404 15973
rect -3804 15665 -3404 15725
rect -3111 15722 -2711 15782
rect -3804 15547 -3404 15607
rect -3111 15604 -2711 15664
rect 36951 15622 37151 15682
rect -3804 15429 -3404 15489
rect -3111 15486 -2711 15546
rect -3804 15311 -3404 15371
rect -3804 15193 -3404 15253
rect -3804 15075 -3404 15135
rect -3111 15368 -2711 15428
rect 36951 15504 37151 15564
rect 36951 15386 37151 15446
rect -3111 15250 -2711 15310
rect -3111 15132 -2711 15192
rect 7858 15036 7918 15236
rect 7976 15036 8036 15236
rect 8094 15036 8154 15236
rect 8212 15036 8272 15236
rect 8330 15036 8390 15236
rect 8448 15036 8508 15236
rect 8566 15036 8626 15236
rect 8684 15036 8744 15236
rect 8802 15036 8862 15236
rect -3604 14828 -3404 14888
rect 14407 15035 14467 15235
rect 14525 15035 14585 15235
rect 14643 15035 14703 15235
rect 14761 15035 14821 15235
rect 14879 15035 14939 15235
rect 14997 15035 15057 15235
rect 15115 15035 15175 15235
rect 15233 15035 15293 15235
rect 15351 15035 15411 15235
rect 21061 15056 21121 15256
rect 21179 15056 21239 15256
rect 21297 15056 21357 15256
rect 21415 15056 21475 15256
rect 21533 15056 21593 15256
rect 21651 15056 21711 15256
rect 21769 15056 21829 15256
rect 21887 15056 21947 15256
rect 22005 15056 22065 15256
rect 36751 15181 37151 15241
rect -3604 14710 -3404 14770
rect -3604 14592 -3404 14652
rect 29714 14889 29774 15089
rect 29832 14889 29892 15089
rect 29950 14889 30010 15089
rect 30068 14889 30128 15089
rect 30186 14889 30246 15089
rect 30304 14889 30364 15089
rect 30422 14889 30482 15089
rect 30540 14889 30600 15089
rect 30658 14889 30718 15089
rect 36751 15063 37151 15123
rect 36751 14945 37151 15005
rect 31522 14484 31582 14684
rect 31640 14484 31700 14684
rect 31758 14484 31818 14684
rect 32006 14484 32066 14884
rect 32124 14484 32184 14884
rect 32242 14484 32302 14884
rect 32360 14484 32420 14884
rect 32478 14484 32538 14884
rect 32596 14484 32656 14884
rect 32843 14484 32903 14684
rect 32961 14484 33021 14684
rect 33079 14484 33139 14684
rect 36751 14714 37151 14774
rect 33315 14481 33375 14681
rect 33433 14481 33493 14681
rect 33551 14481 33611 14681
rect 33669 14481 33729 14681
rect 33787 14481 33847 14681
rect 33905 14481 33965 14681
rect 34023 14481 34083 14681
rect 34141 14481 34201 14681
rect 34259 14481 34319 14681
rect 36751 14596 37151 14656
rect -3606 14081 -3406 14141
rect -3606 13963 -3406 14023
rect -3606 13845 -3406 13905
rect -3806 13597 -3406 13657
rect -3113 13654 -2713 13714
rect -3806 13479 -3406 13539
rect -3113 13536 -2713 13596
rect -3806 13361 -3406 13421
rect -3113 13418 -2713 13478
rect -3806 13243 -3406 13303
rect -3806 13125 -3406 13185
rect -3806 13007 -3406 13067
rect -3113 13300 -2713 13360
rect -3113 13182 -2713 13242
rect -3113 13064 -2713 13124
rect 1194 13136 1254 13336
rect 1312 13136 1372 13336
rect 1430 13136 1490 13336
rect 1548 13136 1608 13336
rect 1666 13136 1726 13336
rect 1784 13136 1844 13336
rect 1902 13136 1962 13336
rect 2020 13136 2080 13336
rect 2138 13136 2198 13336
rect 31949 13791 32009 14191
rect 32067 13791 32127 14191
rect 32185 13791 32245 14191
rect 32303 13791 32363 14191
rect 32421 13791 32481 14191
rect 32539 13791 32599 14191
rect 36751 14478 37151 14538
rect 36751 14360 37151 14420
rect 36751 14242 37151 14302
rect 36751 14124 37151 14184
rect 36751 13887 37151 13947
rect 36751 13769 37151 13829
rect 36751 13651 37151 13711
rect -3606 12760 -3406 12820
rect -3606 12642 -3406 12702
rect -3606 12524 -3406 12584
rect 4084 12869 4144 13069
rect 4202 12869 4262 13069
rect 4320 12869 4380 13069
rect 4438 12869 4498 13069
rect 4556 12869 4616 13069
rect 4674 12869 4734 13069
rect 4792 12869 4852 13069
rect 4910 12869 4970 13069
rect 5028 12869 5088 13069
rect 6409 12741 6469 13141
rect 6527 12741 6587 13141
rect 6645 12741 6705 13141
rect 6763 12741 6823 13141
rect 6881 12741 6941 13141
rect 6999 12741 7059 13141
rect 7551 12745 7611 13145
rect 7669 12745 7729 13145
rect 7787 12745 7847 13145
rect 7905 12745 7965 13145
rect 8023 12745 8083 13145
rect 8141 12745 8201 13145
rect 10633 12957 10693 13157
rect 10751 12957 10811 13157
rect 10869 12957 10929 13157
rect 10987 12957 11047 13157
rect 11105 12957 11165 13157
rect 11223 12957 11283 13157
rect 11341 12957 11401 13157
rect 11459 12957 11519 13157
rect 11577 12957 11637 13157
rect 12958 12829 13018 13229
rect 13076 12829 13136 13229
rect 13194 12829 13254 13229
rect 13312 12829 13372 13229
rect 13430 12829 13490 13229
rect 13548 12829 13608 13229
rect 14100 12833 14160 13233
rect 14218 12833 14278 13233
rect 14336 12833 14396 13233
rect 14454 12833 14514 13233
rect 14572 12833 14632 13233
rect 14690 12833 14750 13233
rect 17287 12889 17347 13089
rect 17405 12889 17465 13089
rect 17523 12889 17583 13089
rect 17641 12889 17701 13089
rect 17759 12889 17819 13089
rect 17877 12889 17937 13089
rect 17995 12889 18055 13089
rect 18113 12889 18173 13089
rect 18231 12889 18291 13089
rect 6838 12158 6898 12358
rect 6956 12158 7016 12358
rect 7074 12158 7134 12358
rect 7980 12162 8040 12362
rect 8098 12162 8158 12362
rect 8216 12162 8276 12362
rect 19612 12761 19672 13161
rect 19730 12761 19790 13161
rect 19848 12761 19908 13161
rect 19966 12761 20026 13161
rect 20084 12761 20144 13161
rect 20202 12761 20262 13161
rect 20754 12765 20814 13165
rect 20872 12765 20932 13165
rect 20990 12765 21050 13165
rect 21108 12765 21168 13165
rect 21226 12765 21286 13165
rect 21344 12765 21404 13165
rect 23912 12957 23972 13157
rect 24030 12957 24090 13157
rect 24148 12957 24208 13157
rect 24266 12957 24326 13157
rect 24384 12957 24444 13157
rect 24502 12957 24562 13157
rect 24620 12957 24680 13157
rect 24738 12957 24798 13157
rect 24856 12957 24916 13157
rect 13387 12246 13447 12446
rect 13505 12246 13565 12446
rect 13623 12246 13683 12446
rect 14529 12250 14589 12450
rect 14647 12250 14707 12450
rect 14765 12250 14825 12450
rect 26237 12829 26297 13229
rect 26355 12829 26415 13229
rect 26473 12829 26533 13229
rect 26591 12829 26651 13229
rect 26709 12829 26769 13229
rect 26827 12829 26887 13229
rect 27379 12833 27439 13233
rect 27497 12833 27557 13233
rect 27615 12833 27675 13233
rect 27733 12833 27793 13233
rect 27851 12833 27911 13233
rect 27969 12833 28029 13233
rect 36951 13414 37151 13474
rect 36951 13296 37151 13356
rect 36951 13178 37151 13238
rect 20041 12178 20101 12378
rect 20159 12178 20219 12378
rect 20277 12178 20337 12378
rect 21183 12182 21243 12382
rect 21301 12182 21361 12382
rect 21419 12182 21479 12382
rect 26666 12246 26726 12446
rect 26784 12246 26844 12446
rect 26902 12246 26962 12446
rect 27808 12250 27868 12450
rect 27926 12250 27986 12450
rect 28044 12250 28104 12450
rect 29709 12318 29769 12518
rect 29827 12318 29887 12518
rect 29945 12318 30005 12518
rect 30063 12318 30123 12518
rect 30181 12318 30241 12518
rect 30299 12318 30359 12518
rect 30417 12318 30477 12518
rect 30535 12318 30595 12518
rect 30653 12318 30713 12518
rect 36955 12420 37155 12480
rect -3604 12012 -3404 12072
rect -3604 11894 -3404 11954
rect 36955 12302 37155 12362
rect 36955 12184 37155 12244
rect -3604 11776 -3404 11836
rect -3804 11528 -3404 11588
rect -3111 11585 -2711 11645
rect 36755 11979 37155 12039
rect 36755 11861 37155 11921
rect 36755 11743 37155 11803
rect -3804 11410 -3404 11470
rect -3111 11467 -2711 11527
rect -3804 11292 -3404 11352
rect -3111 11349 -2711 11409
rect -3804 11174 -3404 11234
rect -3804 11056 -3404 11116
rect -3804 10938 -3404 10998
rect -3111 11231 -2711 11291
rect 4098 11219 4158 11419
rect 4216 11219 4276 11419
rect 4334 11219 4394 11419
rect 4452 11219 4512 11419
rect 4570 11219 4630 11419
rect 4688 11219 4748 11419
rect 4806 11219 4866 11419
rect 4924 11219 4984 11419
rect 5042 11219 5102 11419
rect 10647 11307 10707 11507
rect 10765 11307 10825 11507
rect 10883 11307 10943 11507
rect 11001 11307 11061 11507
rect 11119 11307 11179 11507
rect 11237 11307 11297 11507
rect 11355 11307 11415 11507
rect 11473 11307 11533 11507
rect 11591 11307 11651 11507
rect -3111 11113 -2711 11173
rect -3111 10995 -2711 11055
rect 17301 11239 17361 11439
rect 17419 11239 17479 11439
rect 17537 11239 17597 11439
rect 17655 11239 17715 11439
rect 17773 11239 17833 11439
rect 17891 11239 17951 11439
rect 18009 11239 18069 11439
rect 18127 11239 18187 11439
rect 18245 11239 18305 11439
rect 23926 11307 23986 11507
rect 24044 11307 24104 11507
rect 24162 11307 24222 11507
rect 24280 11307 24340 11507
rect 24398 11307 24458 11507
rect 24516 11307 24576 11507
rect 24634 11307 24694 11507
rect 24752 11307 24812 11507
rect 24870 11307 24930 11507
rect 36755 11512 37155 11572
rect 36755 11394 37155 11454
rect -3604 10691 -3404 10751
rect -3604 10573 -3404 10633
rect 1186 10551 1246 10751
rect 1304 10551 1364 10751
rect 1422 10551 1482 10751
rect 1540 10551 1600 10751
rect 1658 10551 1718 10751
rect 1776 10551 1836 10751
rect 1894 10551 1954 10751
rect 2012 10551 2072 10751
rect 2130 10551 2190 10751
rect -3604 10455 -3404 10515
rect 5562 10602 5622 10802
rect 5680 10602 5740 10802
rect 5798 10602 5858 10802
rect 6046 10602 6106 11002
rect 6164 10602 6224 11002
rect 6282 10602 6342 11002
rect 6400 10602 6460 11002
rect 6518 10602 6578 11002
rect 6636 10602 6696 11002
rect 6883 10602 6943 10802
rect 7001 10602 7061 10802
rect 7119 10602 7179 10802
rect 7460 10602 7520 10802
rect 7578 10602 7638 10802
rect 7696 10602 7756 10802
rect 7944 10602 8004 11002
rect 8062 10602 8122 11002
rect 8180 10602 8240 11002
rect 8298 10602 8358 11002
rect 8416 10602 8476 11002
rect 8534 10602 8594 11002
rect 8781 10602 8841 10802
rect 8899 10602 8959 10802
rect 9017 10602 9077 10802
rect -3606 9944 -3406 10004
rect -3606 9826 -3406 9886
rect -3606 9708 -3406 9768
rect 4093 9615 4153 9815
rect 4211 9615 4271 9815
rect 4329 9615 4389 9815
rect 4447 9615 4507 9815
rect 4565 9615 4625 9815
rect 4683 9615 4743 9815
rect 4801 9615 4861 9815
rect 4919 9615 4979 9815
rect 5037 9615 5097 9815
rect 5989 9909 6049 10309
rect 6107 9909 6167 10309
rect 6225 9909 6285 10309
rect 6343 9909 6403 10309
rect 6461 9909 6521 10309
rect 6579 9909 6639 10309
rect -3806 9460 -3406 9520
rect -3113 9517 -2713 9577
rect -3806 9342 -3406 9402
rect -3113 9399 -2713 9459
rect 12111 10690 12171 10890
rect 12229 10690 12289 10890
rect 12347 10690 12407 10890
rect 12595 10690 12655 11090
rect 12713 10690 12773 11090
rect 12831 10690 12891 11090
rect 12949 10690 13009 11090
rect 13067 10690 13127 11090
rect 13185 10690 13245 11090
rect 13432 10690 13492 10890
rect 13550 10690 13610 10890
rect 13668 10690 13728 10890
rect 14009 10690 14069 10890
rect 14127 10690 14187 10890
rect 14245 10690 14305 10890
rect 14493 10690 14553 11090
rect 14611 10690 14671 11090
rect 14729 10690 14789 11090
rect 14847 10690 14907 11090
rect 14965 10690 15025 11090
rect 15083 10690 15143 11090
rect 36755 11276 37155 11336
rect 36755 11158 37155 11218
rect 15330 10690 15390 10890
rect 15448 10690 15508 10890
rect 15566 10690 15626 10890
rect 7887 9909 7947 10309
rect 8005 9909 8065 10309
rect 8123 9909 8183 10309
rect 8241 9909 8301 10309
rect 8359 9909 8419 10309
rect 8477 9909 8537 10309
rect 10642 9703 10702 9903
rect 10760 9703 10820 9903
rect 10878 9703 10938 9903
rect 10996 9703 11056 9903
rect 11114 9703 11174 9903
rect 11232 9703 11292 9903
rect 11350 9703 11410 9903
rect 11468 9703 11528 9903
rect 11586 9703 11646 9903
rect 12538 9997 12598 10397
rect 12656 9997 12716 10397
rect 12774 9997 12834 10397
rect 12892 9997 12952 10397
rect 13010 9997 13070 10397
rect 13128 9997 13188 10397
rect -3806 9224 -3406 9284
rect -3113 9281 -2713 9341
rect -3806 9106 -3406 9166
rect -3806 8988 -3406 9048
rect -3806 8870 -3406 8930
rect -3113 9163 -2713 9223
rect -3113 9045 -2713 9105
rect -3113 8927 -2713 8987
rect 18765 10622 18825 10822
rect 18883 10622 18943 10822
rect 19001 10622 19061 10822
rect 19249 10622 19309 11022
rect 19367 10622 19427 11022
rect 19485 10622 19545 11022
rect 19603 10622 19663 11022
rect 19721 10622 19781 11022
rect 19839 10622 19899 11022
rect 20086 10622 20146 10822
rect 20204 10622 20264 10822
rect 20322 10622 20382 10822
rect 20663 10622 20723 10822
rect 20781 10622 20841 10822
rect 20899 10622 20959 10822
rect 21147 10622 21207 11022
rect 21265 10622 21325 11022
rect 21383 10622 21443 11022
rect 21501 10622 21561 11022
rect 21619 10622 21679 11022
rect 21737 10622 21797 11022
rect 21984 10622 22044 10822
rect 22102 10622 22162 10822
rect 22220 10622 22280 10822
rect 14436 9997 14496 10397
rect 14554 9997 14614 10397
rect 14672 9997 14732 10397
rect 14790 9997 14850 10397
rect 14908 9997 14968 10397
rect 15026 9997 15086 10397
rect 17296 9635 17356 9835
rect 17414 9635 17474 9835
rect 17532 9635 17592 9835
rect 17650 9635 17710 9835
rect 17768 9635 17828 9835
rect 17886 9635 17946 9835
rect 18004 9635 18064 9835
rect 18122 9635 18182 9835
rect 18240 9635 18300 9835
rect 19192 9929 19252 10329
rect 19310 9929 19370 10329
rect 19428 9929 19488 10329
rect 19546 9929 19606 10329
rect 19664 9929 19724 10329
rect 19782 9929 19842 10329
rect 25390 10690 25450 10890
rect 25508 10690 25568 10890
rect 25626 10690 25686 10890
rect 25874 10690 25934 11090
rect 25992 10690 26052 11090
rect 26110 10690 26170 11090
rect 26228 10690 26288 11090
rect 26346 10690 26406 11090
rect 26464 10690 26524 11090
rect 26711 10690 26771 10890
rect 26829 10690 26889 10890
rect 26947 10690 27007 10890
rect 27288 10690 27348 10890
rect 27406 10690 27466 10890
rect 27524 10690 27584 10890
rect 27772 10690 27832 11090
rect 27890 10690 27950 11090
rect 28008 10690 28068 11090
rect 28126 10690 28186 11090
rect 28244 10690 28304 11090
rect 28362 10690 28422 11090
rect 36755 11040 37155 11100
rect 36755 10922 37155 10982
rect 28609 10690 28669 10890
rect 28727 10690 28787 10890
rect 28845 10690 28905 10890
rect 21090 9929 21150 10329
rect 21208 9929 21268 10329
rect 21326 9929 21386 10329
rect 21444 9929 21504 10329
rect 21562 9929 21622 10329
rect 21680 9929 21740 10329
rect 23921 9703 23981 9903
rect 24039 9703 24099 9903
rect 24157 9703 24217 9903
rect 24275 9703 24335 9903
rect 24393 9703 24453 9903
rect 24511 9703 24571 9903
rect 24629 9703 24689 9903
rect 24747 9703 24807 9903
rect 24865 9703 24925 9903
rect 25817 9997 25877 10397
rect 25935 9997 25995 10397
rect 26053 9997 26113 10397
rect 26171 9997 26231 10397
rect 26289 9997 26349 10397
rect 26407 9997 26467 10397
rect 27715 9997 27775 10397
rect 27833 9997 27893 10397
rect 27951 9997 28011 10397
rect 28069 9997 28129 10397
rect 28187 9997 28247 10397
rect 28305 9997 28365 10397
rect 31524 10393 31584 10593
rect 31642 10393 31702 10593
rect 31760 10393 31820 10593
rect 32008 10393 32068 10793
rect 32126 10393 32186 10793
rect 32244 10393 32304 10793
rect 32362 10393 32422 10793
rect 32480 10393 32540 10793
rect 32598 10393 32658 10793
rect 36755 10685 37155 10745
rect 32845 10393 32905 10593
rect 32963 10393 33023 10593
rect 33081 10393 33141 10593
rect 33317 10390 33377 10590
rect 33435 10390 33495 10590
rect 33553 10390 33613 10590
rect 33671 10390 33731 10590
rect 33789 10390 33849 10590
rect 33907 10390 33967 10590
rect 34025 10390 34085 10590
rect 34143 10390 34203 10590
rect 34261 10390 34321 10590
rect 36755 10567 37155 10627
rect 36755 10449 37155 10509
rect 29709 9285 29769 9485
rect 29827 9285 29887 9485
rect 29945 9285 30005 9485
rect 30063 9285 30123 9485
rect 30181 9285 30241 9485
rect 30299 9285 30359 9485
rect 30417 9285 30477 9485
rect 30535 9285 30595 9485
rect 30653 9285 30713 9485
rect 31951 9700 32011 10100
rect 32069 9700 32129 10100
rect 32187 9700 32247 10100
rect 32305 9700 32365 10100
rect 32423 9700 32483 10100
rect 32541 9700 32601 10100
rect 36955 10212 37155 10272
rect 36955 10094 37155 10154
rect 36955 9976 37155 10036
rect -3606 8623 -3406 8683
rect 36955 9276 37155 9336
rect 36955 9158 37155 9218
rect 36955 9040 37155 9100
rect 36755 8835 37155 8895
rect 36755 8717 37155 8777
rect -3606 8505 -3406 8565
rect 36755 8599 37155 8659
rect -3606 8387 -3406 8447
rect 36755 8368 37155 8428
rect 36755 8250 37155 8310
rect 36755 8132 37155 8192
rect -3606 7875 -3406 7935
rect -3606 7757 -3406 7817
rect 36755 8014 37155 8074
rect 36755 7896 37155 7956
rect -3606 7639 -3406 7699
rect -3806 7391 -3406 7451
rect -3113 7448 -2713 7508
rect -3806 7273 -3406 7333
rect -3113 7330 -2713 7390
rect -3806 7155 -3406 7215
rect -3113 7212 -2713 7272
rect 1167 7273 1227 7473
rect 1285 7273 1345 7473
rect 1403 7273 1463 7473
rect 1521 7273 1581 7473
rect 1639 7273 1699 7473
rect 1757 7273 1817 7473
rect 1875 7273 1935 7473
rect 1993 7273 2053 7473
rect 2111 7273 2171 7473
rect -3806 7037 -3406 7097
rect -3806 6919 -3406 6979
rect -3806 6801 -3406 6861
rect -3113 7094 -2713 7154
rect 4076 7089 4136 7289
rect 4194 7089 4254 7289
rect 4312 7089 4372 7289
rect 4430 7089 4490 7289
rect 4548 7089 4608 7289
rect 4666 7089 4726 7289
rect 4784 7089 4844 7289
rect 4902 7089 4962 7289
rect 5020 7089 5080 7289
rect -3113 6976 -2713 7036
rect -3113 6858 -2713 6918
rect 6401 6961 6461 7361
rect 6519 6961 6579 7361
rect 6637 6961 6697 7361
rect 6755 6961 6815 7361
rect 6873 6961 6933 7361
rect 6991 6961 7051 7361
rect 7543 6965 7603 7365
rect 7661 6965 7721 7365
rect 7779 6965 7839 7365
rect 7897 6965 7957 7365
rect 8015 6965 8075 7365
rect 8133 6965 8193 7365
rect 36755 7778 37155 7838
rect 10627 7087 10687 7287
rect 10745 7087 10805 7287
rect 10863 7087 10923 7287
rect 10981 7087 11041 7287
rect 11099 7087 11159 7287
rect 11217 7087 11277 7287
rect 11335 7087 11395 7287
rect 11453 7087 11513 7287
rect 11571 7087 11631 7287
rect -3606 6554 -3406 6614
rect -3606 6436 -3406 6496
rect 12952 6959 13012 7359
rect 13070 6959 13130 7359
rect 13188 6959 13248 7359
rect 13306 6959 13366 7359
rect 13424 6959 13484 7359
rect 13542 6959 13602 7359
rect 14094 6963 14154 7363
rect 14212 6963 14272 7363
rect 14330 6963 14390 7363
rect 14448 6963 14508 7363
rect 14566 6963 14626 7363
rect 14684 6963 14744 7363
rect 17282 7088 17342 7288
rect 17400 7088 17460 7288
rect 17518 7088 17578 7288
rect 17636 7088 17696 7288
rect 17754 7088 17814 7288
rect 17872 7088 17932 7288
rect 17990 7088 18050 7288
rect 18108 7088 18168 7288
rect 18226 7088 18286 7288
rect -3606 6318 -3406 6378
rect 6830 6378 6890 6578
rect 6948 6378 7008 6578
rect 7066 6378 7126 6578
rect 7972 6382 8032 6582
rect 8090 6382 8150 6582
rect 8208 6382 8268 6582
rect 19607 6960 19667 7360
rect 19725 6960 19785 7360
rect 19843 6960 19903 7360
rect 19961 6960 20021 7360
rect 20079 6960 20139 7360
rect 20197 6960 20257 7360
rect 20749 6964 20809 7364
rect 20867 6964 20927 7364
rect 20985 6964 21045 7364
rect 21103 6964 21163 7364
rect 21221 6964 21281 7364
rect 21339 6964 21399 7364
rect 29780 7365 29840 7565
rect 29898 7365 29958 7565
rect 30016 7365 30076 7565
rect 30134 7365 30194 7565
rect 30252 7365 30312 7565
rect 30370 7365 30430 7565
rect 30488 7365 30548 7565
rect 30606 7365 30666 7565
rect 30724 7365 30784 7565
rect 36755 7541 37155 7601
rect 36755 7423 37155 7483
rect 23904 7089 23964 7289
rect 24022 7089 24082 7289
rect 24140 7089 24200 7289
rect 24258 7089 24318 7289
rect 24376 7089 24436 7289
rect 24494 7089 24554 7289
rect 24612 7089 24672 7289
rect 24730 7089 24790 7289
rect 24848 7089 24908 7289
rect 13381 6376 13441 6576
rect 13499 6376 13559 6576
rect 13617 6376 13677 6576
rect 14523 6380 14583 6580
rect 14641 6380 14701 6580
rect 14759 6380 14819 6580
rect 26229 6961 26289 7361
rect 26347 6961 26407 7361
rect 26465 6961 26525 7361
rect 26583 6961 26643 7361
rect 26701 6961 26761 7361
rect 26819 6961 26879 7361
rect 27371 6965 27431 7365
rect 27489 6965 27549 7365
rect 27607 6965 27667 7365
rect 27725 6965 27785 7365
rect 27843 6965 27903 7365
rect 27961 6965 28021 7365
rect 20036 6377 20096 6577
rect 20154 6377 20214 6577
rect 20272 6377 20332 6577
rect 21178 6381 21238 6581
rect 21296 6381 21356 6581
rect 21414 6381 21474 6581
rect 31524 6898 31584 7098
rect 31642 6898 31702 7098
rect 31760 6898 31820 7098
rect 32008 6898 32068 7298
rect 32126 6898 32186 7298
rect 32244 6898 32304 7298
rect 32362 6898 32422 7298
rect 32480 6898 32540 7298
rect 32598 6898 32658 7298
rect 36755 7305 37155 7365
rect 32845 6898 32905 7098
rect 32963 6898 33023 7098
rect 33081 6898 33141 7098
rect 33317 6895 33377 7095
rect 33435 6895 33495 7095
rect 33553 6895 33613 7095
rect 33671 6895 33731 7095
rect 33789 6895 33849 7095
rect 33907 6895 33967 7095
rect 34025 6895 34085 7095
rect 34143 6895 34203 7095
rect 34261 6895 34321 7095
rect 36955 7068 37155 7128
rect 36955 6950 37155 7010
rect 26658 6378 26718 6578
rect 26776 6378 26836 6578
rect 26894 6378 26954 6578
rect 27800 6382 27860 6582
rect 27918 6382 27978 6582
rect 28036 6382 28096 6582
rect -3608 5807 -3408 5867
rect -3608 5689 -3408 5749
rect 31951 6205 32011 6605
rect 32069 6205 32129 6605
rect 32187 6205 32247 6605
rect 32305 6205 32365 6605
rect 32423 6205 32483 6605
rect 32541 6205 32601 6605
rect 36955 6832 37155 6892
rect 36951 6144 37151 6204
rect 36951 6026 37151 6086
rect 36951 5908 37151 5968
rect -3608 5571 -3408 5631
rect -3808 5323 -3408 5383
rect -3115 5380 -2715 5440
rect 4090 5439 4150 5639
rect 4208 5439 4268 5639
rect 4326 5439 4386 5639
rect 4444 5439 4504 5639
rect 4562 5439 4622 5639
rect 4680 5439 4740 5639
rect 4798 5439 4858 5639
rect 4916 5439 4976 5639
rect 5034 5439 5094 5639
rect -3808 5205 -3408 5265
rect -3115 5262 -2715 5322
rect -3808 5087 -3408 5147
rect -3115 5144 -2715 5204
rect 10641 5437 10701 5637
rect 10759 5437 10819 5637
rect 10877 5437 10937 5637
rect 10995 5437 11055 5637
rect 11113 5437 11173 5637
rect 11231 5437 11291 5637
rect 11349 5437 11409 5637
rect 11467 5437 11527 5637
rect 11585 5437 11645 5637
rect 17296 5438 17356 5638
rect 17414 5438 17474 5638
rect 17532 5438 17592 5638
rect 17650 5438 17710 5638
rect 17768 5438 17828 5638
rect 17886 5438 17946 5638
rect 18004 5438 18064 5638
rect 18122 5438 18182 5638
rect 18240 5438 18300 5638
rect 23918 5439 23978 5639
rect 24036 5439 24096 5639
rect 24154 5439 24214 5639
rect 24272 5439 24332 5639
rect 24390 5439 24450 5639
rect 24508 5439 24568 5639
rect 24626 5439 24686 5639
rect 24744 5439 24804 5639
rect 24862 5439 24922 5639
rect 36751 5703 37151 5763
rect 36751 5585 37151 5645
rect 36751 5467 37151 5527
rect -3808 4969 -3408 5029
rect -3808 4851 -3408 4911
rect -3808 4733 -3408 4793
rect -3115 5026 -2715 5086
rect -3115 4908 -2715 4968
rect -3115 4790 -2715 4850
rect 5554 4822 5614 5022
rect 5672 4822 5732 5022
rect 5790 4822 5850 5022
rect 6038 4822 6098 5222
rect 6156 4822 6216 5222
rect 6274 4822 6334 5222
rect 6392 4822 6452 5222
rect 6510 4822 6570 5222
rect 6628 4822 6688 5222
rect 6875 4822 6935 5022
rect 6993 4822 7053 5022
rect 7111 4822 7171 5022
rect 7452 4822 7512 5022
rect 7570 4822 7630 5022
rect 7688 4822 7748 5022
rect 7936 4822 7996 5222
rect 8054 4822 8114 5222
rect 8172 4822 8232 5222
rect 8290 4822 8350 5222
rect 8408 4822 8468 5222
rect 8526 4822 8586 5222
rect 8773 4822 8833 5022
rect 8891 4822 8951 5022
rect 9009 4822 9069 5022
rect -3608 4486 -3408 4546
rect 1183 4513 1243 4713
rect 1301 4513 1361 4713
rect 1419 4513 1479 4713
rect 1537 4513 1597 4713
rect 1655 4513 1715 4713
rect 1773 4513 1833 4713
rect 1891 4513 1951 4713
rect 2009 4513 2069 4713
rect 2127 4513 2187 4713
rect -3608 4368 -3408 4428
rect -3608 4250 -3408 4310
rect -3606 3738 -3406 3798
rect -3606 3620 -3406 3680
rect 4085 3835 4145 4035
rect 4203 3835 4263 4035
rect 4321 3835 4381 4035
rect 4439 3835 4499 4035
rect 4557 3835 4617 4035
rect 4675 3835 4735 4035
rect 4793 3835 4853 4035
rect 4911 3835 4971 4035
rect 5029 3835 5089 4035
rect 5981 4129 6041 4529
rect 6099 4129 6159 4529
rect 6217 4129 6277 4529
rect 6335 4129 6395 4529
rect 6453 4129 6513 4529
rect 6571 4129 6631 4529
rect -3606 3502 -3406 3562
rect 12105 4820 12165 5020
rect 12223 4820 12283 5020
rect 12341 4820 12401 5020
rect 12589 4820 12649 5220
rect 12707 4820 12767 5220
rect 12825 4820 12885 5220
rect 12943 4820 13003 5220
rect 13061 4820 13121 5220
rect 13179 4820 13239 5220
rect 13426 4820 13486 5020
rect 13544 4820 13604 5020
rect 13662 4820 13722 5020
rect 14003 4820 14063 5020
rect 14121 4820 14181 5020
rect 14239 4820 14299 5020
rect 14487 4820 14547 5220
rect 14605 4820 14665 5220
rect 14723 4820 14783 5220
rect 14841 4820 14901 5220
rect 14959 4820 15019 5220
rect 15077 4820 15137 5220
rect 15324 4820 15384 5020
rect 15442 4820 15502 5020
rect 15560 4820 15620 5020
rect 7879 4129 7939 4529
rect 7997 4129 8057 4529
rect 8115 4129 8175 4529
rect 8233 4129 8293 4529
rect 8351 4129 8411 4529
rect 8469 4129 8529 4529
rect 10636 3833 10696 4033
rect 10754 3833 10814 4033
rect 10872 3833 10932 4033
rect 10990 3833 11050 4033
rect 11108 3833 11168 4033
rect 11226 3833 11286 4033
rect 11344 3833 11404 4033
rect 11462 3833 11522 4033
rect 11580 3833 11640 4033
rect 12532 4127 12592 4527
rect 12650 4127 12710 4527
rect 12768 4127 12828 4527
rect 12886 4127 12946 4527
rect 13004 4127 13064 4527
rect 13122 4127 13182 4527
rect -3806 3254 -3406 3314
rect -3113 3311 -2713 3371
rect -3806 3136 -3406 3196
rect -3113 3193 -2713 3253
rect 18760 4821 18820 5021
rect 18878 4821 18938 5021
rect 18996 4821 19056 5021
rect 19244 4821 19304 5221
rect 19362 4821 19422 5221
rect 19480 4821 19540 5221
rect 19598 4821 19658 5221
rect 19716 4821 19776 5221
rect 19834 4821 19894 5221
rect 20081 4821 20141 5021
rect 20199 4821 20259 5021
rect 20317 4821 20377 5021
rect 20658 4821 20718 5021
rect 20776 4821 20836 5021
rect 20894 4821 20954 5021
rect 21142 4821 21202 5221
rect 21260 4821 21320 5221
rect 21378 4821 21438 5221
rect 21496 4821 21556 5221
rect 21614 4821 21674 5221
rect 21732 4821 21792 5221
rect 21979 4821 22039 5021
rect 22097 4821 22157 5021
rect 22215 4821 22275 5021
rect 14430 4127 14490 4527
rect 14548 4127 14608 4527
rect 14666 4127 14726 4527
rect 14784 4127 14844 4527
rect 14902 4127 14962 4527
rect 15020 4127 15080 4527
rect 17291 3834 17351 4034
rect 17409 3834 17469 4034
rect 17527 3834 17587 4034
rect 17645 3834 17705 4034
rect 17763 3834 17823 4034
rect 17881 3834 17941 4034
rect 17999 3834 18059 4034
rect 18117 3834 18177 4034
rect 18235 3834 18295 4034
rect 19187 4128 19247 4528
rect 19305 4128 19365 4528
rect 19423 4128 19483 4528
rect 19541 4128 19601 4528
rect 19659 4128 19719 4528
rect 19777 4128 19837 4528
rect -3806 3018 -3406 3078
rect -3113 3075 -2713 3135
rect 25382 4822 25442 5022
rect 25500 4822 25560 5022
rect 25618 4822 25678 5022
rect 25866 4822 25926 5222
rect 25984 4822 26044 5222
rect 26102 4822 26162 5222
rect 26220 4822 26280 5222
rect 26338 4822 26398 5222
rect 26456 4822 26516 5222
rect 26703 4822 26763 5022
rect 26821 4822 26881 5022
rect 26939 4822 26999 5022
rect 27280 4822 27340 5022
rect 27398 4822 27458 5022
rect 27516 4822 27576 5022
rect 27764 4822 27824 5222
rect 27882 4822 27942 5222
rect 28000 4822 28060 5222
rect 28118 4822 28178 5222
rect 28236 4822 28296 5222
rect 28354 4822 28414 5222
rect 36751 5236 37151 5296
rect 36751 5118 37151 5178
rect 28601 4822 28661 5022
rect 28719 4822 28779 5022
rect 28837 4822 28897 5022
rect 36751 5000 37151 5060
rect 21085 4128 21145 4528
rect 21203 4128 21263 4528
rect 21321 4128 21381 4528
rect 21439 4128 21499 4528
rect 21557 4128 21617 4528
rect 21675 4128 21735 4528
rect 23913 3835 23973 4035
rect 24031 3835 24091 4035
rect 24149 3835 24209 4035
rect 24267 3835 24327 4035
rect 24385 3835 24445 4035
rect 24503 3835 24563 4035
rect 24621 3835 24681 4035
rect 24739 3835 24799 4035
rect 24857 3835 24917 4035
rect 25809 4129 25869 4529
rect 25927 4129 25987 4529
rect 26045 4129 26105 4529
rect 26163 4129 26223 4529
rect 26281 4129 26341 4529
rect 26399 4129 26459 4529
rect -3806 2900 -3406 2960
rect -3806 2782 -3406 2842
rect -3806 2664 -3406 2724
rect -3113 2957 -2713 3017
rect 36751 4882 37151 4942
rect 36751 4764 37151 4824
rect 36751 4646 37151 4706
rect 27707 4129 27767 4529
rect 27825 4129 27885 4529
rect 27943 4129 28003 4529
rect 28061 4129 28121 4529
rect 28179 4129 28239 4529
rect 28297 4129 28357 4529
rect 29777 4295 29837 4495
rect 29895 4295 29955 4495
rect 30013 4295 30073 4495
rect 30131 4295 30191 4495
rect 30249 4295 30309 4495
rect 30367 4295 30427 4495
rect 30485 4295 30545 4495
rect 30603 4295 30663 4495
rect 30721 4295 30781 4495
rect 36751 4409 37151 4469
rect 36751 4291 37151 4351
rect 36751 4173 37151 4233
rect 36951 3936 37151 3996
rect 36951 3818 37151 3878
rect 36951 3700 37151 3760
rect -3113 2839 -2713 2899
rect -3113 2721 -2713 2781
rect 31524 2550 31584 2750
rect 31642 2550 31702 2750
rect 31760 2550 31820 2750
rect 32008 2550 32068 2950
rect 32126 2550 32186 2950
rect 32244 2550 32304 2950
rect 32362 2550 32422 2950
rect 32480 2550 32540 2950
rect 32598 2550 32658 2950
rect 36951 3000 37151 3060
rect 36951 2882 37151 2942
rect 32845 2550 32905 2750
rect 32963 2550 33023 2750
rect 33081 2550 33141 2750
rect 36951 2764 37151 2824
rect -3606 2417 -3406 2477
rect -3606 2299 -3406 2359
rect 33317 2547 33377 2747
rect 33435 2547 33495 2747
rect 33553 2547 33613 2747
rect 33671 2547 33731 2747
rect 33789 2547 33849 2747
rect 33907 2547 33967 2747
rect 34025 2547 34085 2747
rect 34143 2547 34203 2747
rect 34261 2547 34321 2747
rect 36751 2559 37151 2619
rect -3606 2181 -3406 2241
rect -3608 1670 -3408 1730
rect -3608 1552 -3408 1612
rect -3608 1434 -3408 1494
rect 7893 1332 7953 1532
rect 8011 1332 8071 1532
rect 8129 1332 8189 1532
rect 8247 1332 8307 1532
rect 8365 1332 8425 1532
rect 8483 1332 8543 1532
rect 8601 1332 8661 1532
rect 8719 1332 8779 1532
rect 8837 1332 8897 1532
rect 14447 1337 14507 1537
rect 14565 1337 14625 1537
rect 14683 1337 14743 1537
rect 14801 1337 14861 1537
rect 14919 1337 14979 1537
rect 15037 1337 15097 1537
rect 15155 1337 15215 1537
rect 15273 1337 15333 1537
rect 15391 1337 15451 1537
rect -3808 1186 -3408 1246
rect -3115 1243 -2715 1303
rect 21096 1325 21156 1525
rect 21214 1325 21274 1525
rect 21332 1325 21392 1525
rect 21450 1325 21510 1525
rect 21568 1325 21628 1525
rect 21686 1325 21746 1525
rect 21804 1325 21864 1525
rect 21922 1325 21982 1525
rect 22040 1325 22100 1525
rect 29784 1450 29844 1650
rect 29902 1450 29962 1650
rect 30020 1450 30080 1650
rect 30138 1450 30198 1650
rect 30256 1450 30316 1650
rect 30374 1450 30434 1650
rect 30492 1450 30552 1650
rect 30610 1450 30670 1650
rect 30728 1450 30788 1650
rect 31951 1857 32011 2257
rect 32069 1857 32129 2257
rect 32187 1857 32247 2257
rect 32305 1857 32365 2257
rect 32423 1857 32483 2257
rect 32541 1857 32601 2257
rect 36751 2441 37151 2501
rect 36751 2323 37151 2383
rect 36751 2092 37151 2152
rect 36751 1974 37151 2034
rect 36751 1856 37151 1916
rect 36751 1738 37151 1798
rect 36751 1620 37151 1680
rect -3808 1068 -3408 1128
rect -3115 1125 -2715 1185
rect -3808 950 -3408 1010
rect -3115 1007 -2715 1067
rect -3808 832 -3408 892
rect -3808 714 -3408 774
rect -3808 596 -3408 656
rect -3115 889 -2715 949
rect -3115 771 -2715 831
rect 36751 1502 37151 1562
rect 36751 1265 37151 1325
rect 36751 1147 37151 1207
rect 36751 1029 37151 1089
rect 36951 792 37151 852
rect -3115 653 -2715 713
rect 36951 674 37151 734
rect 36951 556 37151 616
rect -3608 349 -3408 409
rect -3608 231 -3408 291
rect -3608 113 -3408 173
<< ndiff >>
rect 6067 27171 6125 27183
rect 6067 26795 6079 27171
rect 6113 26795 6125 27171
rect 6067 26783 6125 26795
rect 6185 27171 6243 27183
rect 6185 26795 6197 27171
rect 6231 26795 6243 27171
rect 6185 26783 6243 26795
rect 6303 27171 6361 27183
rect 6303 26795 6315 27171
rect 6349 26795 6361 27171
rect 6420 27171 6478 27183
rect 6420 26995 6432 27171
rect 6466 26995 6478 27171
rect 6420 26983 6478 26995
rect 6538 27171 6596 27183
rect 6538 26995 6550 27171
rect 6584 26995 6596 27171
rect 6538 26983 6596 26995
rect 12580 27168 12638 27180
rect 8065 26897 8123 26909
rect 6303 26783 6361 26795
rect 8065 26721 8077 26897
rect 8111 26721 8123 26897
rect 8065 26709 8123 26721
rect 8183 26897 8241 26909
rect 8183 26721 8195 26897
rect 8229 26721 8241 26897
rect 8183 26709 8241 26721
rect 8301 26897 8359 26909
rect 8301 26721 8313 26897
rect 8347 26721 8359 26897
rect 8301 26709 8359 26721
rect 8419 26897 8477 26909
rect 8419 26721 8431 26897
rect 8465 26721 8477 26897
rect 8419 26709 8477 26721
rect 9207 26901 9265 26913
rect 9207 26725 9219 26901
rect 9253 26725 9265 26901
rect 9207 26713 9265 26725
rect 9325 26901 9383 26913
rect 9325 26725 9337 26901
rect 9371 26725 9383 26901
rect 9325 26713 9383 26725
rect 9443 26901 9501 26913
rect 9443 26725 9455 26901
rect 9489 26725 9501 26901
rect 9443 26713 9501 26725
rect 9561 26901 9619 26913
rect 9561 26725 9573 26901
rect 9607 26725 9619 26901
rect 9561 26713 9619 26725
rect 12580 26792 12592 27168
rect 12626 26792 12638 27168
rect 12580 26780 12638 26792
rect 12698 27168 12756 27180
rect 12698 26792 12710 27168
rect 12744 26792 12756 27168
rect 12698 26780 12756 26792
rect 12816 27168 12874 27180
rect 12816 26792 12828 27168
rect 12862 26792 12874 27168
rect 12933 27168 12991 27180
rect 12933 26992 12945 27168
rect 12979 26992 12991 27168
rect 12933 26980 12991 26992
rect 13051 27168 13109 27180
rect 13051 26992 13063 27168
rect 13097 26992 13109 27168
rect 13051 26980 13109 26992
rect 19114 27163 19172 27175
rect 14578 26894 14636 26906
rect 12816 26780 12874 26792
rect 14578 26718 14590 26894
rect 14624 26718 14636 26894
rect 14578 26706 14636 26718
rect 14696 26894 14754 26906
rect 14696 26718 14708 26894
rect 14742 26718 14754 26894
rect 14696 26706 14754 26718
rect 14814 26894 14872 26906
rect 14814 26718 14826 26894
rect 14860 26718 14872 26894
rect 14814 26706 14872 26718
rect 14932 26894 14990 26906
rect 14932 26718 14944 26894
rect 14978 26718 14990 26894
rect 14932 26706 14990 26718
rect 15720 26898 15778 26910
rect 15720 26722 15732 26898
rect 15766 26722 15778 26898
rect 15720 26710 15778 26722
rect 15838 26898 15896 26910
rect 15838 26722 15850 26898
rect 15884 26722 15896 26898
rect 15838 26710 15896 26722
rect 15956 26898 16014 26910
rect 15956 26722 15968 26898
rect 16002 26722 16014 26898
rect 15956 26710 16014 26722
rect 16074 26898 16132 26910
rect 16074 26722 16086 26898
rect 16120 26722 16132 26898
rect 16074 26710 16132 26722
rect 19114 26787 19126 27163
rect 19160 26787 19172 27163
rect 19114 26775 19172 26787
rect 19232 27163 19290 27175
rect 19232 26787 19244 27163
rect 19278 26787 19290 27163
rect 19232 26775 19290 26787
rect 19350 27163 19408 27175
rect 19350 26787 19362 27163
rect 19396 26787 19408 27163
rect 19467 27163 19525 27175
rect 19467 26987 19479 27163
rect 19513 26987 19525 27163
rect 19467 26975 19525 26987
rect 19585 27163 19643 27175
rect 19585 26987 19597 27163
rect 19631 26987 19643 27163
rect 19585 26975 19643 26987
rect 25672 27167 25730 27179
rect 21112 26889 21170 26901
rect 19350 26775 19408 26787
rect 21112 26713 21124 26889
rect 21158 26713 21170 26889
rect 21112 26701 21170 26713
rect 21230 26889 21288 26901
rect 21230 26713 21242 26889
rect 21276 26713 21288 26889
rect 21230 26701 21288 26713
rect 21348 26889 21406 26901
rect 21348 26713 21360 26889
rect 21394 26713 21406 26889
rect 21348 26701 21406 26713
rect 21466 26889 21524 26901
rect 21466 26713 21478 26889
rect 21512 26713 21524 26889
rect 21466 26701 21524 26713
rect 22254 26893 22312 26905
rect 22254 26717 22266 26893
rect 22300 26717 22312 26893
rect 22254 26705 22312 26717
rect 22372 26893 22430 26905
rect 22372 26717 22384 26893
rect 22418 26717 22430 26893
rect 22372 26705 22430 26717
rect 22490 26893 22548 26905
rect 22490 26717 22502 26893
rect 22536 26717 22548 26893
rect 22490 26705 22548 26717
rect 22608 26893 22666 26905
rect 22608 26717 22620 26893
rect 22654 26717 22666 26893
rect 22608 26705 22666 26717
rect 25672 26791 25684 27167
rect 25718 26791 25730 27167
rect 25672 26779 25730 26791
rect 25790 27167 25848 27179
rect 25790 26791 25802 27167
rect 25836 26791 25848 27167
rect 25790 26779 25848 26791
rect 25908 27167 25966 27179
rect 25908 26791 25920 27167
rect 25954 26791 25966 27167
rect 26025 27167 26083 27179
rect 26025 26991 26037 27167
rect 26071 26991 26083 27167
rect 26025 26979 26083 26991
rect 26143 27167 26201 27179
rect 26143 26991 26155 27167
rect 26189 26991 26201 27167
rect 26143 26979 26201 26991
rect 27670 26893 27728 26905
rect 25908 26779 25966 26791
rect 27670 26717 27682 26893
rect 27716 26717 27728 26893
rect 27670 26705 27728 26717
rect 27788 26893 27846 26905
rect 27788 26717 27800 26893
rect 27834 26717 27846 26893
rect 27788 26705 27846 26717
rect 27906 26893 27964 26905
rect 27906 26717 27918 26893
rect 27952 26717 27964 26893
rect 27906 26705 27964 26717
rect 28024 26893 28082 26905
rect 28024 26717 28036 26893
rect 28070 26717 28082 26893
rect 28024 26705 28082 26717
rect 28812 26897 28870 26909
rect 28812 26721 28824 26897
rect 28858 26721 28870 26897
rect 28812 26709 28870 26721
rect 28930 26897 28988 26909
rect 28930 26721 28942 26897
rect 28976 26721 28988 26897
rect 28930 26709 28988 26721
rect 29048 26897 29106 26909
rect 29048 26721 29060 26897
rect 29094 26721 29106 26897
rect 29048 26709 29106 26721
rect 29166 26897 29224 26909
rect 29166 26721 29178 26897
rect 29212 26721 29224 26897
rect 29166 26709 29224 26721
rect 6081 25521 6139 25533
rect 6081 25145 6093 25521
rect 6127 25145 6139 25521
rect 6081 25133 6139 25145
rect 6199 25521 6257 25533
rect 6199 25145 6211 25521
rect 6245 25145 6257 25521
rect 6199 25133 6257 25145
rect 6317 25521 6375 25533
rect 6317 25145 6329 25521
rect 6363 25145 6375 25521
rect 6434 25521 6492 25533
rect 6434 25345 6446 25521
rect 6480 25345 6492 25521
rect 6434 25333 6492 25345
rect 6552 25521 6610 25533
rect 6552 25345 6564 25521
rect 6598 25345 6610 25521
rect 6552 25333 6610 25345
rect 6317 25133 6375 25145
rect 12594 25518 12652 25530
rect 12594 25142 12606 25518
rect 12640 25142 12652 25518
rect 12594 25130 12652 25142
rect 12712 25518 12770 25530
rect 12712 25142 12724 25518
rect 12758 25142 12770 25518
rect 12712 25130 12770 25142
rect 12830 25518 12888 25530
rect 12830 25142 12842 25518
rect 12876 25142 12888 25518
rect 12947 25518 13005 25530
rect 12947 25342 12959 25518
rect 12993 25342 13005 25518
rect 12947 25330 13005 25342
rect 13065 25518 13123 25530
rect 13065 25342 13077 25518
rect 13111 25342 13123 25518
rect 13065 25330 13123 25342
rect 12830 25130 12888 25142
rect 19128 25513 19186 25525
rect 7433 24116 7491 24128
rect 7433 23940 7445 24116
rect 7479 23940 7491 24116
rect 6076 23917 6134 23929
rect 6076 23541 6088 23917
rect 6122 23541 6134 23917
rect 6076 23529 6134 23541
rect 6194 23917 6252 23929
rect 6194 23541 6206 23917
rect 6240 23541 6252 23917
rect 6194 23529 6252 23541
rect 6312 23917 6370 23929
rect 6312 23541 6324 23917
rect 6358 23541 6370 23917
rect 6429 23917 6487 23929
rect 6429 23741 6441 23917
rect 6475 23741 6487 23917
rect 6429 23729 6487 23741
rect 6547 23917 6605 23929
rect 7433 23928 7491 23940
rect 7551 24116 7609 24128
rect 7551 23940 7563 24116
rect 7597 23940 7609 24116
rect 7551 23928 7609 23940
rect 7853 24116 7911 24128
rect 6547 23741 6559 23917
rect 6593 23741 6605 23917
rect 6547 23729 6605 23741
rect 7853 23740 7865 24116
rect 7899 23740 7911 24116
rect 7853 23728 7911 23740
rect 7971 24116 8029 24128
rect 7971 23740 7983 24116
rect 8017 23740 8029 24116
rect 7971 23728 8029 23740
rect 8089 24116 8147 24128
rect 8089 23740 8101 24116
rect 8135 23740 8147 24116
rect 8089 23728 8147 23740
rect 8207 24116 8265 24128
rect 8207 23740 8219 24116
rect 8253 23740 8265 24116
rect 8207 23728 8265 23740
rect 8325 24116 8383 24128
rect 8325 23740 8337 24116
rect 8371 23740 8383 24116
rect 8731 24116 8789 24128
rect 8731 23940 8743 24116
rect 8777 23940 8789 24116
rect 8731 23928 8789 23940
rect 8849 24116 8907 24128
rect 8849 23940 8861 24116
rect 8895 23940 8907 24116
rect 8849 23928 8907 23940
rect 9331 24116 9389 24128
rect 9331 23940 9343 24116
rect 9377 23940 9389 24116
rect 9331 23928 9389 23940
rect 9449 24116 9507 24128
rect 9449 23940 9461 24116
rect 9495 23940 9507 24116
rect 9449 23928 9507 23940
rect 9751 24116 9809 24128
rect 8325 23728 8383 23740
rect 9751 23740 9763 24116
rect 9797 23740 9809 24116
rect 9751 23728 9809 23740
rect 9869 24116 9927 24128
rect 9869 23740 9881 24116
rect 9915 23740 9927 24116
rect 9869 23728 9927 23740
rect 9987 24116 10045 24128
rect 9987 23740 9999 24116
rect 10033 23740 10045 24116
rect 9987 23728 10045 23740
rect 10105 24116 10163 24128
rect 10105 23740 10117 24116
rect 10151 23740 10163 24116
rect 10105 23728 10163 23740
rect 10223 24116 10281 24128
rect 10223 23740 10235 24116
rect 10269 23740 10281 24116
rect 10629 24116 10687 24128
rect 10629 23940 10641 24116
rect 10675 23940 10687 24116
rect 10629 23928 10687 23940
rect 10747 24116 10805 24128
rect 10747 23940 10759 24116
rect 10793 23940 10805 24116
rect 10747 23928 10805 23940
rect 19128 25137 19140 25513
rect 19174 25137 19186 25513
rect 19128 25125 19186 25137
rect 19246 25513 19304 25525
rect 19246 25137 19258 25513
rect 19292 25137 19304 25513
rect 19246 25125 19304 25137
rect 19364 25513 19422 25525
rect 19364 25137 19376 25513
rect 19410 25137 19422 25513
rect 19481 25513 19539 25525
rect 19481 25337 19493 25513
rect 19527 25337 19539 25513
rect 19481 25325 19539 25337
rect 19599 25513 19657 25525
rect 19599 25337 19611 25513
rect 19645 25337 19657 25513
rect 19599 25325 19657 25337
rect 19364 25125 19422 25137
rect 25686 25517 25744 25529
rect 13946 24113 14004 24125
rect 13946 23937 13958 24113
rect 13992 23937 14004 24113
rect 12589 23914 12647 23926
rect 10223 23728 10281 23740
rect 6312 23529 6370 23541
rect 12589 23538 12601 23914
rect 12635 23538 12647 23914
rect 12589 23526 12647 23538
rect 12707 23914 12765 23926
rect 12707 23538 12719 23914
rect 12753 23538 12765 23914
rect 12707 23526 12765 23538
rect 12825 23914 12883 23926
rect 12825 23538 12837 23914
rect 12871 23538 12883 23914
rect 12942 23914 13000 23926
rect 12942 23738 12954 23914
rect 12988 23738 13000 23914
rect 12942 23726 13000 23738
rect 13060 23914 13118 23926
rect 13946 23925 14004 23937
rect 14064 24113 14122 24125
rect 14064 23937 14076 24113
rect 14110 23937 14122 24113
rect 14064 23925 14122 23937
rect 14366 24113 14424 24125
rect 13060 23738 13072 23914
rect 13106 23738 13118 23914
rect 13060 23726 13118 23738
rect 14366 23737 14378 24113
rect 14412 23737 14424 24113
rect 14366 23725 14424 23737
rect 14484 24113 14542 24125
rect 14484 23737 14496 24113
rect 14530 23737 14542 24113
rect 14484 23725 14542 23737
rect 14602 24113 14660 24125
rect 14602 23737 14614 24113
rect 14648 23737 14660 24113
rect 14602 23725 14660 23737
rect 14720 24113 14778 24125
rect 14720 23737 14732 24113
rect 14766 23737 14778 24113
rect 14720 23725 14778 23737
rect 14838 24113 14896 24125
rect 14838 23737 14850 24113
rect 14884 23737 14896 24113
rect 15244 24113 15302 24125
rect 15244 23937 15256 24113
rect 15290 23937 15302 24113
rect 15244 23925 15302 23937
rect 15362 24113 15420 24125
rect 15362 23937 15374 24113
rect 15408 23937 15420 24113
rect 15362 23925 15420 23937
rect 15844 24113 15902 24125
rect 15844 23937 15856 24113
rect 15890 23937 15902 24113
rect 15844 23925 15902 23937
rect 15962 24113 16020 24125
rect 15962 23937 15974 24113
rect 16008 23937 16020 24113
rect 15962 23925 16020 23937
rect 16264 24113 16322 24125
rect 14838 23725 14896 23737
rect 16264 23737 16276 24113
rect 16310 23737 16322 24113
rect 16264 23725 16322 23737
rect 16382 24113 16440 24125
rect 16382 23737 16394 24113
rect 16428 23737 16440 24113
rect 16382 23725 16440 23737
rect 16500 24113 16558 24125
rect 16500 23737 16512 24113
rect 16546 23737 16558 24113
rect 16500 23725 16558 23737
rect 16618 24113 16676 24125
rect 16618 23737 16630 24113
rect 16664 23737 16676 24113
rect 16618 23725 16676 23737
rect 16736 24113 16794 24125
rect 16736 23737 16748 24113
rect 16782 23737 16794 24113
rect 17142 24113 17200 24125
rect 17142 23937 17154 24113
rect 17188 23937 17200 24113
rect 17142 23925 17200 23937
rect 17260 24113 17318 24125
rect 17260 23937 17272 24113
rect 17306 23937 17318 24113
rect 17260 23925 17318 23937
rect 25686 25141 25698 25517
rect 25732 25141 25744 25517
rect 25686 25129 25744 25141
rect 25804 25517 25862 25529
rect 25804 25141 25816 25517
rect 25850 25141 25862 25517
rect 25804 25129 25862 25141
rect 25922 25517 25980 25529
rect 25922 25141 25934 25517
rect 25968 25141 25980 25517
rect 26039 25517 26097 25529
rect 26039 25341 26051 25517
rect 26085 25341 26097 25517
rect 26039 25329 26097 25341
rect 26157 25517 26215 25529
rect 26157 25341 26169 25517
rect 26203 25341 26215 25517
rect 26157 25329 26215 25341
rect 25922 25129 25980 25141
rect 20480 24108 20538 24120
rect 20480 23932 20492 24108
rect 20526 23932 20538 24108
rect 19123 23909 19181 23921
rect 16736 23725 16794 23737
rect 12825 23526 12883 23538
rect 19123 23533 19135 23909
rect 19169 23533 19181 23909
rect 19123 23521 19181 23533
rect 19241 23909 19299 23921
rect 19241 23533 19253 23909
rect 19287 23533 19299 23909
rect 19241 23521 19299 23533
rect 19359 23909 19417 23921
rect 19359 23533 19371 23909
rect 19405 23533 19417 23909
rect 19476 23909 19534 23921
rect 19476 23733 19488 23909
rect 19522 23733 19534 23909
rect 19476 23721 19534 23733
rect 19594 23909 19652 23921
rect 20480 23920 20538 23932
rect 20598 24108 20656 24120
rect 20598 23932 20610 24108
rect 20644 23932 20656 24108
rect 20598 23920 20656 23932
rect 20900 24108 20958 24120
rect 19594 23733 19606 23909
rect 19640 23733 19652 23909
rect 19594 23721 19652 23733
rect 20900 23732 20912 24108
rect 20946 23732 20958 24108
rect 20900 23720 20958 23732
rect 21018 24108 21076 24120
rect 21018 23732 21030 24108
rect 21064 23732 21076 24108
rect 21018 23720 21076 23732
rect 21136 24108 21194 24120
rect 21136 23732 21148 24108
rect 21182 23732 21194 24108
rect 21136 23720 21194 23732
rect 21254 24108 21312 24120
rect 21254 23732 21266 24108
rect 21300 23732 21312 24108
rect 21254 23720 21312 23732
rect 21372 24108 21430 24120
rect 21372 23732 21384 24108
rect 21418 23732 21430 24108
rect 21778 24108 21836 24120
rect 21778 23932 21790 24108
rect 21824 23932 21836 24108
rect 21778 23920 21836 23932
rect 21896 24108 21954 24120
rect 21896 23932 21908 24108
rect 21942 23932 21954 24108
rect 21896 23920 21954 23932
rect 22378 24108 22436 24120
rect 22378 23932 22390 24108
rect 22424 23932 22436 24108
rect 22378 23920 22436 23932
rect 22496 24108 22554 24120
rect 22496 23932 22508 24108
rect 22542 23932 22554 24108
rect 22496 23920 22554 23932
rect 22798 24108 22856 24120
rect 21372 23720 21430 23732
rect 22798 23732 22810 24108
rect 22844 23732 22856 24108
rect 22798 23720 22856 23732
rect 22916 24108 22974 24120
rect 22916 23732 22928 24108
rect 22962 23732 22974 24108
rect 22916 23720 22974 23732
rect 23034 24108 23092 24120
rect 23034 23732 23046 24108
rect 23080 23732 23092 24108
rect 23034 23720 23092 23732
rect 23152 24108 23210 24120
rect 23152 23732 23164 24108
rect 23198 23732 23210 24108
rect 23152 23720 23210 23732
rect 23270 24108 23328 24120
rect 23270 23732 23282 24108
rect 23316 23732 23328 24108
rect 23676 24108 23734 24120
rect 23676 23932 23688 24108
rect 23722 23932 23734 24108
rect 23676 23920 23734 23932
rect 23794 24108 23852 24120
rect 23794 23932 23806 24108
rect 23840 23932 23852 24108
rect 23794 23920 23852 23932
rect 27038 24112 27096 24124
rect 27038 23936 27050 24112
rect 27084 23936 27096 24112
rect 25681 23913 25739 23925
rect 23270 23720 23328 23732
rect 19359 23521 19417 23533
rect 25681 23537 25693 23913
rect 25727 23537 25739 23913
rect 25681 23525 25739 23537
rect 25799 23913 25857 23925
rect 25799 23537 25811 23913
rect 25845 23537 25857 23913
rect 25799 23525 25857 23537
rect 25917 23913 25975 23925
rect 25917 23537 25929 23913
rect 25963 23537 25975 23913
rect 26034 23913 26092 23925
rect 26034 23737 26046 23913
rect 26080 23737 26092 23913
rect 26034 23725 26092 23737
rect 26152 23913 26210 23925
rect 27038 23924 27096 23936
rect 27156 24112 27214 24124
rect 27156 23936 27168 24112
rect 27202 23936 27214 24112
rect 27156 23924 27214 23936
rect 27458 24112 27516 24124
rect 26152 23737 26164 23913
rect 26198 23737 26210 23913
rect 26152 23725 26210 23737
rect 27458 23736 27470 24112
rect 27504 23736 27516 24112
rect 27458 23724 27516 23736
rect 27576 24112 27634 24124
rect 27576 23736 27588 24112
rect 27622 23736 27634 24112
rect 27576 23724 27634 23736
rect 27694 24112 27752 24124
rect 27694 23736 27706 24112
rect 27740 23736 27752 24112
rect 27694 23724 27752 23736
rect 27812 24112 27870 24124
rect 27812 23736 27824 24112
rect 27858 23736 27870 24112
rect 27812 23724 27870 23736
rect 27930 24112 27988 24124
rect 27930 23736 27942 24112
rect 27976 23736 27988 24112
rect 28336 24112 28394 24124
rect 28336 23936 28348 24112
rect 28382 23936 28394 24112
rect 28336 23924 28394 23936
rect 28454 24112 28512 24124
rect 28454 23936 28466 24112
rect 28500 23936 28512 24112
rect 28454 23924 28512 23936
rect 28936 24112 28994 24124
rect 28936 23936 28948 24112
rect 28982 23936 28994 24112
rect 28936 23924 28994 23936
rect 29054 24112 29112 24124
rect 29054 23936 29066 24112
rect 29100 23936 29112 24112
rect 29054 23924 29112 23936
rect 29356 24112 29414 24124
rect 27930 23724 27988 23736
rect 29356 23736 29368 24112
rect 29402 23736 29414 24112
rect 29356 23724 29414 23736
rect 29474 24112 29532 24124
rect 29474 23736 29486 24112
rect 29520 23736 29532 24112
rect 29474 23724 29532 23736
rect 29592 24112 29650 24124
rect 29592 23736 29604 24112
rect 29638 23736 29650 24112
rect 29592 23724 29650 23736
rect 29710 24112 29768 24124
rect 29710 23736 29722 24112
rect 29756 23736 29768 24112
rect 29710 23724 29768 23736
rect 29828 24112 29886 24124
rect 29828 23736 29840 24112
rect 29874 23736 29886 24112
rect 30234 24112 30292 24124
rect 30234 23936 30246 24112
rect 30280 23936 30292 24112
rect 30234 23924 30292 23936
rect 30352 24112 30410 24124
rect 30352 23936 30364 24112
rect 30398 23936 30410 24112
rect 38088 24314 38288 24326
rect 38088 24280 38100 24314
rect 38276 24280 38288 24314
rect 38088 24268 38288 24280
rect 38088 24196 38288 24208
rect 38088 24162 38100 24196
rect 38276 24162 38288 24196
rect 38088 24134 38288 24162
rect 38088 24122 38488 24134
rect 38088 24088 38100 24122
rect 38476 24088 38488 24122
rect 38088 24076 38488 24088
rect 30352 23924 30410 23936
rect 29828 23724 29886 23736
rect 38088 24004 38488 24016
rect 38088 23970 38100 24004
rect 38476 23970 38488 24004
rect 38088 23958 38488 23970
rect 38088 23886 38488 23898
rect 38088 23852 38100 23886
rect 38476 23852 38488 23886
rect 38088 23840 38488 23852
rect 38088 23768 38488 23780
rect 38088 23734 38100 23768
rect 38476 23734 38488 23768
rect 38088 23722 38488 23734
rect 25917 23525 25975 23537
rect 38088 23650 38488 23662
rect 38088 23616 38100 23650
rect 38476 23616 38488 23650
rect 38088 23604 38488 23616
rect 38088 23572 38288 23604
rect 38088 23538 38100 23572
rect 38276 23538 38288 23572
rect 38088 23526 38288 23538
rect 38088 23454 38288 23466
rect 38088 23420 38100 23454
rect 38276 23420 38288 23454
rect 38088 23408 38288 23420
rect 6285 21293 6343 21305
rect 6285 21117 6297 21293
rect 6331 21117 6343 21293
rect 6285 21105 6343 21117
rect 6403 21293 6461 21305
rect 6403 21117 6415 21293
rect 6449 21117 6461 21293
rect 6403 21105 6461 21117
rect 6521 21293 6579 21305
rect 6521 21117 6533 21293
rect 6567 21117 6579 21293
rect 6521 21105 6579 21117
rect 6639 21293 6697 21305
rect 9308 21563 9366 21575
rect 9308 21387 9320 21563
rect 9354 21387 9366 21563
rect 9308 21375 9366 21387
rect 9426 21563 9484 21575
rect 9426 21387 9438 21563
rect 9472 21387 9484 21563
rect 9426 21375 9484 21387
rect 9543 21563 9601 21575
rect 6639 21117 6651 21293
rect 6685 21117 6697 21293
rect 6639 21105 6697 21117
rect 7427 21289 7485 21301
rect 7427 21113 7439 21289
rect 7473 21113 7485 21289
rect 7427 21101 7485 21113
rect 7545 21289 7603 21301
rect 7545 21113 7557 21289
rect 7591 21113 7603 21289
rect 7545 21101 7603 21113
rect 7663 21289 7721 21301
rect 7663 21113 7675 21289
rect 7709 21113 7721 21289
rect 7663 21101 7721 21113
rect 7781 21289 7839 21301
rect 7781 21113 7793 21289
rect 7827 21113 7839 21289
rect 9543 21187 9555 21563
rect 9589 21187 9601 21563
rect 9543 21175 9601 21187
rect 9661 21563 9719 21575
rect 9661 21187 9673 21563
rect 9707 21187 9719 21563
rect 9661 21175 9719 21187
rect 9779 21563 9837 21575
rect 9779 21187 9791 21563
rect 9825 21187 9837 21563
rect 9779 21175 9837 21187
rect 7781 21101 7839 21113
rect 12843 21289 12901 21301
rect 12843 21113 12855 21289
rect 12889 21113 12901 21289
rect 12843 21101 12901 21113
rect 12961 21289 13019 21301
rect 12961 21113 12973 21289
rect 13007 21113 13019 21289
rect 12961 21101 13019 21113
rect 13079 21289 13137 21301
rect 13079 21113 13091 21289
rect 13125 21113 13137 21289
rect 13079 21101 13137 21113
rect 13197 21289 13255 21301
rect 15866 21559 15924 21571
rect 15866 21383 15878 21559
rect 15912 21383 15924 21559
rect 15866 21371 15924 21383
rect 15984 21559 16042 21571
rect 15984 21383 15996 21559
rect 16030 21383 16042 21559
rect 15984 21371 16042 21383
rect 16101 21559 16159 21571
rect 13197 21113 13209 21289
rect 13243 21113 13255 21289
rect 13197 21101 13255 21113
rect 13985 21285 14043 21297
rect 13985 21109 13997 21285
rect 14031 21109 14043 21285
rect 13985 21097 14043 21109
rect 14103 21285 14161 21297
rect 14103 21109 14115 21285
rect 14149 21109 14161 21285
rect 14103 21097 14161 21109
rect 14221 21285 14279 21297
rect 14221 21109 14233 21285
rect 14267 21109 14279 21285
rect 14221 21097 14279 21109
rect 14339 21285 14397 21297
rect 14339 21109 14351 21285
rect 14385 21109 14397 21285
rect 16101 21183 16113 21559
rect 16147 21183 16159 21559
rect 16101 21171 16159 21183
rect 16219 21559 16277 21571
rect 16219 21183 16231 21559
rect 16265 21183 16277 21559
rect 16219 21171 16277 21183
rect 16337 21559 16395 21571
rect 16337 21183 16349 21559
rect 16383 21183 16395 21559
rect 16337 21171 16395 21183
rect 14339 21097 14397 21109
rect 19377 21294 19435 21306
rect 19377 21118 19389 21294
rect 19423 21118 19435 21294
rect 19377 21106 19435 21118
rect 19495 21294 19553 21306
rect 19495 21118 19507 21294
rect 19541 21118 19553 21294
rect 19495 21106 19553 21118
rect 19613 21294 19671 21306
rect 19613 21118 19625 21294
rect 19659 21118 19671 21294
rect 19613 21106 19671 21118
rect 19731 21294 19789 21306
rect 22400 21564 22458 21576
rect 22400 21388 22412 21564
rect 22446 21388 22458 21564
rect 22400 21376 22458 21388
rect 22518 21564 22576 21576
rect 22518 21388 22530 21564
rect 22564 21388 22576 21564
rect 22518 21376 22576 21388
rect 22635 21564 22693 21576
rect 19731 21118 19743 21294
rect 19777 21118 19789 21294
rect 19731 21106 19789 21118
rect 20519 21290 20577 21302
rect 20519 21114 20531 21290
rect 20565 21114 20577 21290
rect 20519 21102 20577 21114
rect 20637 21290 20695 21302
rect 20637 21114 20649 21290
rect 20683 21114 20695 21290
rect 20637 21102 20695 21114
rect 20755 21290 20813 21302
rect 20755 21114 20767 21290
rect 20801 21114 20813 21290
rect 20755 21102 20813 21114
rect 20873 21290 20931 21302
rect 20873 21114 20885 21290
rect 20919 21114 20931 21290
rect 22635 21188 22647 21564
rect 22681 21188 22693 21564
rect 22635 21176 22693 21188
rect 22753 21564 22811 21576
rect 22753 21188 22765 21564
rect 22799 21188 22811 21564
rect 22753 21176 22811 21188
rect 22871 21564 22929 21576
rect 22871 21188 22883 21564
rect 22917 21188 22929 21564
rect 22871 21176 22929 21188
rect 20873 21102 20931 21114
rect 25890 21297 25948 21309
rect 25890 21121 25902 21297
rect 25936 21121 25948 21297
rect 25890 21109 25948 21121
rect 26008 21297 26066 21309
rect 26008 21121 26020 21297
rect 26054 21121 26066 21297
rect 26008 21109 26066 21121
rect 26126 21297 26184 21309
rect 26126 21121 26138 21297
rect 26172 21121 26184 21297
rect 26126 21109 26184 21121
rect 26244 21297 26302 21309
rect 28913 21567 28971 21579
rect 28913 21391 28925 21567
rect 28959 21391 28971 21567
rect 28913 21379 28971 21391
rect 29031 21567 29089 21579
rect 29031 21391 29043 21567
rect 29077 21391 29089 21567
rect 29031 21379 29089 21391
rect 29148 21567 29206 21579
rect 26244 21121 26256 21297
rect 26290 21121 26302 21297
rect 26244 21109 26302 21121
rect 27032 21293 27090 21305
rect 27032 21117 27044 21293
rect 27078 21117 27090 21293
rect 27032 21105 27090 21117
rect 27150 21293 27208 21305
rect 27150 21117 27162 21293
rect 27196 21117 27208 21293
rect 27150 21105 27208 21117
rect 27268 21293 27326 21305
rect 27268 21117 27280 21293
rect 27314 21117 27326 21293
rect 27268 21105 27326 21117
rect 27386 21293 27444 21305
rect 27386 21117 27398 21293
rect 27432 21117 27444 21293
rect 29148 21191 29160 21567
rect 29194 21191 29206 21567
rect 29148 21179 29206 21191
rect 29266 21567 29324 21579
rect 29266 21191 29278 21567
rect 29312 21191 29324 21567
rect 29266 21179 29324 21191
rect 29384 21567 29442 21579
rect 29384 21191 29396 21567
rect 29430 21191 29442 21567
rect 29384 21179 29442 21191
rect 27386 21105 27444 21117
rect 38088 21170 38288 21182
rect 38088 21136 38100 21170
rect 38276 21136 38288 21170
rect 38088 21124 38288 21136
rect 38088 21052 38288 21064
rect 38088 21018 38100 21052
rect 38276 21018 38288 21052
rect 38088 20990 38288 21018
rect 38088 20978 38488 20990
rect 38088 20944 38100 20978
rect 38476 20944 38488 20978
rect 38088 20932 38488 20944
rect 38088 20860 38488 20872
rect 38088 20826 38100 20860
rect 38476 20826 38488 20860
rect 38088 20814 38488 20826
rect 38088 20742 38488 20754
rect 38088 20708 38100 20742
rect 38476 20708 38488 20742
rect 38088 20696 38488 20708
rect 38088 20624 38488 20636
rect 38088 20590 38100 20624
rect 38476 20590 38488 20624
rect 38088 20578 38488 20590
rect 9294 19913 9352 19925
rect 9294 19737 9306 19913
rect 9340 19737 9352 19913
rect 9294 19725 9352 19737
rect 9412 19913 9470 19925
rect 9412 19737 9424 19913
rect 9458 19737 9470 19913
rect 9412 19725 9470 19737
rect 9529 19913 9587 19925
rect 9529 19537 9541 19913
rect 9575 19537 9587 19913
rect 9529 19525 9587 19537
rect 9647 19913 9705 19925
rect 9647 19537 9659 19913
rect 9693 19537 9705 19913
rect 9647 19525 9705 19537
rect 9765 19913 9823 19925
rect 9765 19537 9777 19913
rect 9811 19537 9823 19913
rect 15852 19909 15910 19921
rect 15852 19733 15864 19909
rect 15898 19733 15910 19909
rect 15852 19721 15910 19733
rect 15970 19909 16028 19921
rect 15970 19733 15982 19909
rect 16016 19733 16028 19909
rect 15970 19721 16028 19733
rect 16087 19909 16145 19921
rect 9765 19525 9823 19537
rect 5099 18508 5157 18520
rect 5099 18332 5111 18508
rect 5145 18332 5157 18508
rect 5099 18320 5157 18332
rect 5217 18508 5275 18520
rect 5217 18332 5229 18508
rect 5263 18332 5275 18508
rect 5217 18320 5275 18332
rect 5623 18508 5681 18520
rect 5623 18132 5635 18508
rect 5669 18132 5681 18508
rect 5623 18120 5681 18132
rect 5741 18508 5799 18520
rect 5741 18132 5753 18508
rect 5787 18132 5799 18508
rect 5741 18120 5799 18132
rect 5859 18508 5917 18520
rect 5859 18132 5871 18508
rect 5905 18132 5917 18508
rect 5859 18120 5917 18132
rect 5977 18508 6035 18520
rect 5977 18132 5989 18508
rect 6023 18132 6035 18508
rect 5977 18120 6035 18132
rect 6095 18508 6153 18520
rect 6095 18132 6107 18508
rect 6141 18132 6153 18508
rect 6397 18508 6455 18520
rect 6397 18332 6409 18508
rect 6443 18332 6455 18508
rect 6397 18320 6455 18332
rect 6515 18508 6573 18520
rect 6515 18332 6527 18508
rect 6561 18332 6573 18508
rect 6515 18320 6573 18332
rect 6997 18508 7055 18520
rect 6997 18332 7009 18508
rect 7043 18332 7055 18508
rect 6997 18320 7055 18332
rect 7115 18508 7173 18520
rect 7115 18332 7127 18508
rect 7161 18332 7173 18508
rect 7115 18320 7173 18332
rect 7521 18508 7579 18520
rect 6095 18120 6153 18132
rect 7521 18132 7533 18508
rect 7567 18132 7579 18508
rect 7521 18120 7579 18132
rect 7639 18508 7697 18520
rect 7639 18132 7651 18508
rect 7685 18132 7697 18508
rect 7639 18120 7697 18132
rect 7757 18508 7815 18520
rect 7757 18132 7769 18508
rect 7803 18132 7815 18508
rect 7757 18120 7815 18132
rect 7875 18508 7933 18520
rect 7875 18132 7887 18508
rect 7921 18132 7933 18508
rect 7875 18120 7933 18132
rect 7993 18508 8051 18520
rect 7993 18132 8005 18508
rect 8039 18132 8051 18508
rect 8295 18508 8353 18520
rect 8295 18332 8307 18508
rect 8341 18332 8353 18508
rect 8295 18320 8353 18332
rect 8413 18508 8471 18520
rect 8413 18332 8425 18508
rect 8459 18332 8471 18508
rect 8413 18320 8471 18332
rect 16087 19533 16099 19909
rect 16133 19533 16145 19909
rect 16087 19521 16145 19533
rect 16205 19909 16263 19921
rect 16205 19533 16217 19909
rect 16251 19533 16263 19909
rect 16205 19521 16263 19533
rect 16323 19909 16381 19921
rect 16323 19533 16335 19909
rect 16369 19533 16381 19909
rect 22386 19914 22444 19926
rect 22386 19738 22398 19914
rect 22432 19738 22444 19914
rect 22386 19726 22444 19738
rect 22504 19914 22562 19926
rect 22504 19738 22516 19914
rect 22550 19738 22562 19914
rect 22504 19726 22562 19738
rect 22621 19914 22679 19926
rect 16323 19521 16381 19533
rect 11657 18504 11715 18516
rect 11657 18328 11669 18504
rect 11703 18328 11715 18504
rect 9299 18309 9357 18321
rect 7993 18120 8051 18132
rect 9299 18133 9311 18309
rect 9345 18133 9357 18309
rect 9299 18121 9357 18133
rect 9417 18309 9475 18321
rect 9417 18133 9429 18309
rect 9463 18133 9475 18309
rect 9417 18121 9475 18133
rect 9534 18309 9592 18321
rect 9534 17933 9546 18309
rect 9580 17933 9592 18309
rect 9534 17921 9592 17933
rect 9652 18309 9710 18321
rect 9652 17933 9664 18309
rect 9698 17933 9710 18309
rect 9652 17921 9710 17933
rect 9770 18309 9828 18321
rect 11657 18316 11715 18328
rect 11775 18504 11833 18516
rect 11775 18328 11787 18504
rect 11821 18328 11833 18504
rect 11775 18316 11833 18328
rect 12181 18504 12239 18516
rect 9770 17933 9782 18309
rect 9816 17933 9828 18309
rect 12181 18128 12193 18504
rect 12227 18128 12239 18504
rect 12181 18116 12239 18128
rect 12299 18504 12357 18516
rect 12299 18128 12311 18504
rect 12345 18128 12357 18504
rect 12299 18116 12357 18128
rect 12417 18504 12475 18516
rect 12417 18128 12429 18504
rect 12463 18128 12475 18504
rect 12417 18116 12475 18128
rect 12535 18504 12593 18516
rect 12535 18128 12547 18504
rect 12581 18128 12593 18504
rect 12535 18116 12593 18128
rect 12653 18504 12711 18516
rect 12653 18128 12665 18504
rect 12699 18128 12711 18504
rect 12955 18504 13013 18516
rect 12955 18328 12967 18504
rect 13001 18328 13013 18504
rect 12955 18316 13013 18328
rect 13073 18504 13131 18516
rect 13073 18328 13085 18504
rect 13119 18328 13131 18504
rect 13073 18316 13131 18328
rect 13555 18504 13613 18516
rect 13555 18328 13567 18504
rect 13601 18328 13613 18504
rect 13555 18316 13613 18328
rect 13673 18504 13731 18516
rect 13673 18328 13685 18504
rect 13719 18328 13731 18504
rect 13673 18316 13731 18328
rect 14079 18504 14137 18516
rect 12653 18116 12711 18128
rect 14079 18128 14091 18504
rect 14125 18128 14137 18504
rect 14079 18116 14137 18128
rect 14197 18504 14255 18516
rect 14197 18128 14209 18504
rect 14243 18128 14255 18504
rect 14197 18116 14255 18128
rect 14315 18504 14373 18516
rect 14315 18128 14327 18504
rect 14361 18128 14373 18504
rect 14315 18116 14373 18128
rect 14433 18504 14491 18516
rect 14433 18128 14445 18504
rect 14479 18128 14491 18504
rect 14433 18116 14491 18128
rect 14551 18504 14609 18516
rect 14551 18128 14563 18504
rect 14597 18128 14609 18504
rect 14853 18504 14911 18516
rect 14853 18328 14865 18504
rect 14899 18328 14911 18504
rect 14853 18316 14911 18328
rect 14971 18504 15029 18516
rect 14971 18328 14983 18504
rect 15017 18328 15029 18504
rect 14971 18316 15029 18328
rect 22621 19538 22633 19914
rect 22667 19538 22679 19914
rect 22621 19526 22679 19538
rect 22739 19914 22797 19926
rect 22739 19538 22751 19914
rect 22785 19538 22797 19914
rect 22739 19526 22797 19538
rect 22857 19914 22915 19926
rect 22857 19538 22869 19914
rect 22903 19538 22915 19914
rect 38088 20506 38488 20518
rect 38088 20472 38100 20506
rect 38476 20472 38488 20506
rect 38088 20460 38488 20472
rect 38088 20428 38288 20460
rect 38088 20394 38100 20428
rect 38276 20394 38288 20428
rect 38088 20382 38288 20394
rect 28899 19917 28957 19929
rect 28899 19741 28911 19917
rect 28945 19741 28957 19917
rect 28899 19729 28957 19741
rect 29017 19917 29075 19929
rect 29017 19741 29029 19917
rect 29063 19741 29075 19917
rect 29017 19729 29075 19741
rect 29134 19917 29192 19929
rect 22857 19526 22915 19538
rect 18191 18509 18249 18521
rect 18191 18333 18203 18509
rect 18237 18333 18249 18509
rect 18191 18321 18249 18333
rect 18309 18509 18367 18521
rect 18309 18333 18321 18509
rect 18355 18333 18367 18509
rect 18309 18321 18367 18333
rect 18715 18509 18773 18521
rect 15857 18305 15915 18317
rect 14551 18116 14609 18128
rect 15857 18129 15869 18305
rect 15903 18129 15915 18305
rect 15857 18117 15915 18129
rect 15975 18305 16033 18317
rect 15975 18129 15987 18305
rect 16021 18129 16033 18305
rect 15975 18117 16033 18129
rect 16092 18305 16150 18317
rect 9770 17921 9828 17933
rect 16092 17929 16104 18305
rect 16138 17929 16150 18305
rect 16092 17917 16150 17929
rect 16210 18305 16268 18317
rect 16210 17929 16222 18305
rect 16256 17929 16268 18305
rect 16210 17917 16268 17929
rect 16328 18305 16386 18317
rect 16328 17929 16340 18305
rect 16374 17929 16386 18305
rect 18715 18133 18727 18509
rect 18761 18133 18773 18509
rect 18715 18121 18773 18133
rect 18833 18509 18891 18521
rect 18833 18133 18845 18509
rect 18879 18133 18891 18509
rect 18833 18121 18891 18133
rect 18951 18509 19009 18521
rect 18951 18133 18963 18509
rect 18997 18133 19009 18509
rect 18951 18121 19009 18133
rect 19069 18509 19127 18521
rect 19069 18133 19081 18509
rect 19115 18133 19127 18509
rect 19069 18121 19127 18133
rect 19187 18509 19245 18521
rect 19187 18133 19199 18509
rect 19233 18133 19245 18509
rect 19489 18509 19547 18521
rect 19489 18333 19501 18509
rect 19535 18333 19547 18509
rect 19489 18321 19547 18333
rect 19607 18509 19665 18521
rect 19607 18333 19619 18509
rect 19653 18333 19665 18509
rect 19607 18321 19665 18333
rect 20089 18509 20147 18521
rect 20089 18333 20101 18509
rect 20135 18333 20147 18509
rect 20089 18321 20147 18333
rect 20207 18509 20265 18521
rect 20207 18333 20219 18509
rect 20253 18333 20265 18509
rect 20207 18321 20265 18333
rect 20613 18509 20671 18521
rect 19187 18121 19245 18133
rect 20613 18133 20625 18509
rect 20659 18133 20671 18509
rect 20613 18121 20671 18133
rect 20731 18509 20789 18521
rect 20731 18133 20743 18509
rect 20777 18133 20789 18509
rect 20731 18121 20789 18133
rect 20849 18509 20907 18521
rect 20849 18133 20861 18509
rect 20895 18133 20907 18509
rect 20849 18121 20907 18133
rect 20967 18509 21025 18521
rect 20967 18133 20979 18509
rect 21013 18133 21025 18509
rect 20967 18121 21025 18133
rect 21085 18509 21143 18521
rect 21085 18133 21097 18509
rect 21131 18133 21143 18509
rect 21387 18509 21445 18521
rect 21387 18333 21399 18509
rect 21433 18333 21445 18509
rect 21387 18321 21445 18333
rect 21505 18509 21563 18521
rect 21505 18333 21517 18509
rect 21551 18333 21563 18509
rect 21505 18321 21563 18333
rect 29134 19541 29146 19917
rect 29180 19541 29192 19917
rect 29134 19529 29192 19541
rect 29252 19917 29310 19929
rect 29252 19541 29264 19917
rect 29298 19541 29310 19917
rect 29252 19529 29310 19541
rect 29370 19917 29428 19929
rect 29370 19541 29382 19917
rect 29416 19541 29428 19917
rect 29370 19529 29428 19541
rect 38088 20310 38288 20322
rect 38088 20276 38100 20310
rect 38276 20276 38288 20310
rect 38088 20264 38288 20276
rect 24704 18512 24762 18524
rect 24704 18336 24716 18512
rect 24750 18336 24762 18512
rect 24704 18324 24762 18336
rect 24822 18512 24880 18524
rect 24822 18336 24834 18512
rect 24868 18336 24880 18512
rect 24822 18324 24880 18336
rect 25228 18512 25286 18524
rect 22391 18310 22449 18322
rect 21085 18121 21143 18133
rect 22391 18134 22403 18310
rect 22437 18134 22449 18310
rect 22391 18122 22449 18134
rect 22509 18310 22567 18322
rect 22509 18134 22521 18310
rect 22555 18134 22567 18310
rect 22509 18122 22567 18134
rect 22626 18310 22684 18322
rect 16328 17917 16386 17929
rect 22626 17934 22638 18310
rect 22672 17934 22684 18310
rect 22626 17922 22684 17934
rect 22744 18310 22802 18322
rect 22744 17934 22756 18310
rect 22790 17934 22802 18310
rect 22744 17922 22802 17934
rect 22862 18310 22920 18322
rect 22862 17934 22874 18310
rect 22908 17934 22920 18310
rect 25228 18136 25240 18512
rect 25274 18136 25286 18512
rect 25228 18124 25286 18136
rect 25346 18512 25404 18524
rect 25346 18136 25358 18512
rect 25392 18136 25404 18512
rect 25346 18124 25404 18136
rect 25464 18512 25522 18524
rect 25464 18136 25476 18512
rect 25510 18136 25522 18512
rect 25464 18124 25522 18136
rect 25582 18512 25640 18524
rect 25582 18136 25594 18512
rect 25628 18136 25640 18512
rect 25582 18124 25640 18136
rect 25700 18512 25758 18524
rect 25700 18136 25712 18512
rect 25746 18136 25758 18512
rect 26002 18512 26060 18524
rect 26002 18336 26014 18512
rect 26048 18336 26060 18512
rect 26002 18324 26060 18336
rect 26120 18512 26178 18524
rect 26120 18336 26132 18512
rect 26166 18336 26178 18512
rect 26120 18324 26178 18336
rect 26602 18512 26660 18524
rect 26602 18336 26614 18512
rect 26648 18336 26660 18512
rect 26602 18324 26660 18336
rect 26720 18512 26778 18524
rect 26720 18336 26732 18512
rect 26766 18336 26778 18512
rect 26720 18324 26778 18336
rect 27126 18512 27184 18524
rect 25700 18124 25758 18136
rect 27126 18136 27138 18512
rect 27172 18136 27184 18512
rect 27126 18124 27184 18136
rect 27244 18512 27302 18524
rect 27244 18136 27256 18512
rect 27290 18136 27302 18512
rect 27244 18124 27302 18136
rect 27362 18512 27420 18524
rect 27362 18136 27374 18512
rect 27408 18136 27420 18512
rect 27362 18124 27420 18136
rect 27480 18512 27538 18524
rect 27480 18136 27492 18512
rect 27526 18136 27538 18512
rect 27480 18124 27538 18136
rect 27598 18512 27656 18524
rect 27598 18136 27610 18512
rect 27644 18136 27656 18512
rect 27900 18512 27958 18524
rect 27900 18336 27912 18512
rect 27946 18336 27958 18512
rect 27900 18324 27958 18336
rect 28018 18512 28076 18524
rect 28018 18336 28030 18512
rect 28064 18336 28076 18512
rect 28018 18324 28076 18336
rect 28904 18313 28962 18325
rect 27598 18124 27656 18136
rect 28904 18137 28916 18313
rect 28950 18137 28962 18313
rect 28904 18125 28962 18137
rect 29022 18313 29080 18325
rect 29022 18137 29034 18313
rect 29068 18137 29080 18313
rect 29022 18125 29080 18137
rect 29139 18313 29197 18325
rect 22862 17922 22920 17934
rect 29139 17937 29151 18313
rect 29185 17937 29197 18313
rect 29139 17925 29197 17937
rect 29257 18313 29315 18325
rect 29257 17937 29269 18313
rect 29303 17937 29315 18313
rect 29257 17925 29315 17937
rect 29375 18313 29433 18325
rect 29375 17937 29387 18313
rect 29421 17937 29433 18313
rect 29375 17925 29433 17937
rect 38084 18038 38284 18050
rect 38084 18004 38096 18038
rect 38272 18004 38284 18038
rect 38084 17992 38284 18004
rect 38084 17920 38284 17932
rect 38084 17886 38096 17920
rect 38272 17886 38284 17920
rect 38084 17858 38284 17886
rect 38084 17846 38484 17858
rect 38084 17812 38096 17846
rect 38472 17812 38484 17846
rect 38084 17800 38484 17812
rect 38084 17728 38484 17740
rect 38084 17694 38096 17728
rect 38472 17694 38484 17728
rect 38084 17682 38484 17694
rect 38084 17610 38484 17622
rect 38084 17576 38096 17610
rect 38472 17576 38484 17610
rect 38084 17564 38484 17576
rect 38084 17492 38484 17504
rect 38084 17458 38096 17492
rect 38472 17458 38484 17492
rect 38084 17446 38484 17458
rect 38084 17374 38484 17386
rect 38084 17340 38096 17374
rect 38472 17340 38484 17374
rect 38084 17328 38484 17340
rect 38084 17296 38284 17328
rect 38084 17262 38096 17296
rect 38272 17262 38284 17296
rect 38084 17250 38284 17262
rect 38084 17178 38284 17190
rect 38084 17144 38096 17178
rect 38272 17144 38284 17178
rect 38084 17132 38284 17144
rect -2379 16130 -2179 16142
rect -2379 16096 -2367 16130
rect -2191 16096 -2179 16130
rect -2379 16084 -2179 16096
rect -2379 16012 -2179 16024
rect -2379 15978 -2367 16012
rect -2191 15978 -2179 16012
rect -2379 15966 -2179 15978
rect -2379 15710 -1979 15722
rect -2379 15676 -2367 15710
rect -1991 15676 -1979 15710
rect -2379 15664 -1979 15676
rect -2379 15592 -1979 15604
rect -2379 15558 -2367 15592
rect -1991 15558 -1979 15592
rect -2379 15546 -1979 15558
rect -2379 15474 -1979 15486
rect -2379 15440 -2367 15474
rect -1991 15440 -1979 15474
rect -2379 15428 -1979 15440
rect -2379 15356 -1979 15368
rect -2379 15322 -2367 15356
rect -1991 15322 -1979 15356
rect -2379 15310 -1979 15322
rect -2379 15238 -1979 15250
rect -2379 15204 -2367 15238
rect -1991 15204 -1979 15238
rect -2379 15192 -1979 15204
rect -2379 14832 -2179 14844
rect -2379 14798 -2367 14832
rect -2191 14798 -2179 14832
rect -2379 14786 -2179 14798
rect 8037 14787 8095 14799
rect -2379 14714 -2179 14726
rect -2379 14680 -2367 14714
rect -2191 14680 -2179 14714
rect -2379 14668 -2179 14680
rect 8037 14411 8049 14787
rect 8083 14411 8095 14787
rect 8037 14399 8095 14411
rect 8155 14787 8213 14799
rect 8155 14411 8167 14787
rect 8201 14411 8213 14787
rect 8155 14399 8213 14411
rect 8273 14787 8331 14799
rect 8273 14411 8285 14787
rect 8319 14411 8331 14787
rect 8390 14787 8448 14799
rect 8390 14611 8402 14787
rect 8436 14611 8448 14787
rect 8390 14599 8448 14611
rect 8508 14787 8566 14799
rect 21240 14807 21298 14819
rect 8508 14611 8520 14787
rect 8554 14611 8566 14787
rect 8508 14599 8566 14611
rect 14586 14786 14644 14798
rect 8273 14399 8331 14411
rect 14586 14410 14598 14786
rect 14632 14410 14644 14786
rect 14586 14398 14644 14410
rect 14704 14786 14762 14798
rect 14704 14410 14716 14786
rect 14750 14410 14762 14786
rect 14704 14398 14762 14410
rect 14822 14786 14880 14798
rect 14822 14410 14834 14786
rect 14868 14410 14880 14786
rect 14939 14786 14997 14798
rect 14939 14610 14951 14786
rect 14985 14610 14997 14786
rect 14939 14598 14997 14610
rect 15057 14786 15115 14798
rect 15057 14610 15069 14786
rect 15103 14610 15115 14786
rect 15057 14598 15115 14610
rect 21240 14431 21252 14807
rect 21286 14431 21298 14807
rect 21240 14419 21298 14431
rect 21358 14807 21416 14819
rect 21358 14431 21370 14807
rect 21404 14431 21416 14807
rect 21358 14419 21416 14431
rect 21476 14807 21534 14819
rect 21476 14431 21488 14807
rect 21522 14431 21534 14807
rect 21593 14807 21651 14819
rect 21593 14631 21605 14807
rect 21639 14631 21651 14807
rect 21593 14619 21651 14631
rect 21711 14807 21769 14819
rect 21711 14631 21723 14807
rect 21757 14631 21769 14807
rect 21711 14619 21769 14631
rect 29893 14640 29951 14652
rect 21476 14419 21534 14431
rect 14822 14398 14880 14410
rect 29893 14264 29905 14640
rect 29939 14264 29951 14640
rect 29893 14252 29951 14264
rect 30011 14640 30069 14652
rect 30011 14264 30023 14640
rect 30057 14264 30069 14640
rect 30011 14252 30069 14264
rect 30129 14640 30187 14652
rect 30129 14264 30141 14640
rect 30175 14264 30187 14640
rect 30246 14640 30304 14652
rect 30246 14464 30258 14640
rect 30292 14464 30304 14640
rect 30246 14452 30304 14464
rect 30364 14640 30422 14652
rect 30364 14464 30376 14640
rect 30410 14464 30422 14640
rect 30364 14452 30422 14464
rect 30129 14252 30187 14264
rect 38084 14894 38284 14906
rect 38084 14860 38096 14894
rect 38272 14860 38284 14894
rect 38084 14848 38284 14860
rect 38084 14776 38284 14788
rect 38084 14742 38096 14776
rect 38272 14742 38284 14776
rect 38084 14714 38284 14742
rect 38084 14702 38484 14714
rect 38084 14668 38096 14702
rect 38472 14668 38484 14702
rect 38084 14656 38484 14668
rect -2381 14062 -2181 14074
rect -2381 14028 -2369 14062
rect -2193 14028 -2181 14062
rect -2381 14016 -2181 14028
rect -2381 13944 -2181 13956
rect -2381 13910 -2369 13944
rect -2193 13910 -2181 13944
rect -2381 13898 -2181 13910
rect -2381 13642 -1981 13654
rect -2381 13608 -2369 13642
rect -1993 13608 -1981 13642
rect -2381 13596 -1981 13608
rect -2381 13524 -1981 13536
rect -2381 13490 -2369 13524
rect -1993 13490 -1981 13524
rect -2381 13478 -1981 13490
rect -2381 13406 -1981 13418
rect -2381 13372 -2369 13406
rect -1993 13372 -1981 13406
rect -2381 13360 -1981 13372
rect -2381 13288 -1981 13300
rect -2381 13254 -2369 13288
rect -1993 13254 -1981 13288
rect -2381 13242 -1981 13254
rect -2381 13170 -1981 13182
rect -2381 13136 -2369 13170
rect -1993 13136 -1981 13170
rect 38084 14584 38484 14596
rect 38084 14550 38096 14584
rect 38472 14550 38484 14584
rect 38084 14538 38484 14550
rect 38084 14466 38484 14478
rect 38084 14432 38096 14466
rect 38472 14432 38484 14466
rect 38084 14420 38484 14432
rect 38084 14348 38484 14360
rect 38084 14314 38096 14348
rect 38472 14314 38484 14348
rect 33494 14232 33552 14244
rect 33494 13856 33506 14232
rect 33540 13856 33552 14232
rect 33494 13844 33552 13856
rect 33612 14232 33670 14244
rect 33612 13856 33624 14232
rect 33658 13856 33670 14232
rect 33612 13844 33670 13856
rect 33730 14232 33788 14244
rect 33730 13856 33742 14232
rect 33776 13856 33788 14232
rect 33847 14232 33905 14244
rect 33847 14056 33859 14232
rect 33893 14056 33905 14232
rect 33847 14044 33905 14056
rect 33965 14232 34023 14244
rect 33965 14056 33977 14232
rect 34011 14056 34023 14232
rect 38084 14302 38484 14314
rect 33965 14044 34023 14056
rect 33730 13844 33788 13856
rect 38084 14230 38484 14242
rect 38084 14196 38096 14230
rect 38472 14196 38484 14230
rect 38084 14184 38484 14196
rect 38084 14152 38284 14184
rect 38084 14118 38096 14152
rect 38272 14118 38284 14152
rect 38084 14106 38284 14118
rect 31589 13447 31647 13459
rect -2381 13124 -1981 13136
rect 1373 12887 1431 12899
rect -2381 12764 -2181 12776
rect -2381 12730 -2369 12764
rect -2193 12730 -2181 12764
rect -2381 12718 -2181 12730
rect -2381 12646 -2181 12658
rect -2381 12612 -2369 12646
rect -2193 12612 -2181 12646
rect -2381 12600 -2181 12612
rect 1373 12511 1385 12887
rect 1419 12511 1431 12887
rect 1373 12499 1431 12511
rect 1491 12887 1549 12899
rect 1491 12511 1503 12887
rect 1537 12511 1549 12887
rect 1491 12499 1549 12511
rect 1609 12887 1667 12899
rect 1609 12511 1621 12887
rect 1655 12511 1667 12887
rect 1726 12887 1784 12899
rect 1726 12711 1738 12887
rect 1772 12711 1784 12887
rect 1726 12699 1784 12711
rect 1844 12887 1902 12899
rect 1844 12711 1856 12887
rect 1890 12711 1902 12887
rect 1844 12699 1902 12711
rect 1609 12499 1667 12511
rect 4263 12620 4321 12632
rect 4263 12244 4275 12620
rect 4309 12244 4321 12620
rect 4263 12232 4321 12244
rect 4381 12620 4439 12632
rect 4381 12244 4393 12620
rect 4427 12244 4439 12620
rect 4381 12232 4439 12244
rect 4499 12620 4557 12632
rect 4499 12244 4511 12620
rect 4545 12244 4557 12620
rect 4616 12620 4674 12632
rect 4616 12444 4628 12620
rect 4662 12444 4674 12620
rect 4616 12432 4674 12444
rect 4734 12620 4792 12632
rect 4734 12444 4746 12620
rect 4780 12444 4792 12620
rect 4734 12432 4792 12444
rect 31589 13271 31601 13447
rect 31635 13271 31647 13447
rect 31589 13259 31647 13271
rect 31707 13447 31765 13459
rect 31707 13271 31719 13447
rect 31753 13271 31765 13447
rect 31707 13259 31765 13271
rect 32009 13447 32067 13459
rect 10812 12708 10870 12720
rect 6261 12346 6319 12358
rect 4499 12232 4557 12244
rect 6261 12170 6273 12346
rect 6307 12170 6319 12346
rect 6261 12158 6319 12170
rect 6379 12346 6437 12358
rect 6379 12170 6391 12346
rect 6425 12170 6437 12346
rect 6379 12158 6437 12170
rect 6497 12346 6555 12358
rect 6497 12170 6509 12346
rect 6543 12170 6555 12346
rect 6497 12158 6555 12170
rect 6615 12346 6673 12358
rect 6615 12170 6627 12346
rect 6661 12170 6673 12346
rect 6615 12158 6673 12170
rect 7403 12350 7461 12362
rect 7403 12174 7415 12350
rect 7449 12174 7461 12350
rect 7403 12162 7461 12174
rect 7521 12350 7579 12362
rect 7521 12174 7533 12350
rect 7567 12174 7579 12350
rect 7521 12162 7579 12174
rect 7639 12350 7697 12362
rect 7639 12174 7651 12350
rect 7685 12174 7697 12350
rect 7639 12162 7697 12174
rect 7757 12350 7815 12362
rect 7757 12174 7769 12350
rect 7803 12174 7815 12350
rect 7757 12162 7815 12174
rect 10812 12332 10824 12708
rect 10858 12332 10870 12708
rect 10812 12320 10870 12332
rect 10930 12708 10988 12720
rect 10930 12332 10942 12708
rect 10976 12332 10988 12708
rect 10930 12320 10988 12332
rect 11048 12708 11106 12720
rect 11048 12332 11060 12708
rect 11094 12332 11106 12708
rect 11165 12708 11223 12720
rect 11165 12532 11177 12708
rect 11211 12532 11223 12708
rect 11165 12520 11223 12532
rect 11283 12708 11341 12720
rect 11283 12532 11295 12708
rect 11329 12532 11341 12708
rect 11283 12520 11341 12532
rect 17466 12640 17524 12652
rect 12810 12434 12868 12446
rect 11048 12320 11106 12332
rect 12810 12258 12822 12434
rect 12856 12258 12868 12434
rect 12810 12246 12868 12258
rect 12928 12434 12986 12446
rect 12928 12258 12940 12434
rect 12974 12258 12986 12434
rect 12928 12246 12986 12258
rect 13046 12434 13104 12446
rect 13046 12258 13058 12434
rect 13092 12258 13104 12434
rect 13046 12246 13104 12258
rect 13164 12434 13222 12446
rect 13164 12258 13176 12434
rect 13210 12258 13222 12434
rect 13164 12246 13222 12258
rect 13952 12438 14010 12450
rect 13952 12262 13964 12438
rect 13998 12262 14010 12438
rect 13952 12250 14010 12262
rect 14070 12438 14128 12450
rect 14070 12262 14082 12438
rect 14116 12262 14128 12438
rect 14070 12250 14128 12262
rect 14188 12438 14246 12450
rect 14188 12262 14200 12438
rect 14234 12262 14246 12438
rect 14188 12250 14246 12262
rect 14306 12438 14364 12450
rect 14306 12262 14318 12438
rect 14352 12262 14364 12438
rect 14306 12250 14364 12262
rect 17466 12264 17478 12640
rect 17512 12264 17524 12640
rect 17466 12252 17524 12264
rect 17584 12640 17642 12652
rect 17584 12264 17596 12640
rect 17630 12264 17642 12640
rect 17584 12252 17642 12264
rect 17702 12640 17760 12652
rect 17702 12264 17714 12640
rect 17748 12264 17760 12640
rect 17819 12640 17877 12652
rect 17819 12464 17831 12640
rect 17865 12464 17877 12640
rect 17819 12452 17877 12464
rect 17937 12640 17995 12652
rect 17937 12464 17949 12640
rect 17983 12464 17995 12640
rect 17937 12452 17995 12464
rect 32009 13071 32021 13447
rect 32055 13071 32067 13447
rect 32009 13059 32067 13071
rect 32127 13447 32185 13459
rect 32127 13071 32139 13447
rect 32173 13071 32185 13447
rect 32127 13059 32185 13071
rect 32245 13447 32303 13459
rect 32245 13071 32257 13447
rect 32291 13071 32303 13447
rect 32245 13059 32303 13071
rect 32363 13447 32421 13459
rect 32363 13071 32375 13447
rect 32409 13071 32421 13447
rect 32363 13059 32421 13071
rect 32481 13447 32539 13459
rect 32481 13071 32493 13447
rect 32527 13071 32539 13447
rect 32887 13447 32945 13459
rect 32887 13271 32899 13447
rect 32933 13271 32945 13447
rect 32887 13259 32945 13271
rect 33005 13447 33063 13459
rect 33005 13271 33017 13447
rect 33051 13271 33063 13447
rect 33005 13259 33063 13271
rect 38084 14034 38284 14046
rect 38084 14000 38096 14034
rect 38272 14000 38284 14034
rect 38084 13988 38284 14000
rect 32481 13059 32539 13071
rect 24091 12708 24149 12720
rect 19464 12366 19522 12378
rect 17702 12252 17760 12264
rect 19464 12190 19476 12366
rect 19510 12190 19522 12366
rect 19464 12178 19522 12190
rect 19582 12366 19640 12378
rect 19582 12190 19594 12366
rect 19628 12190 19640 12366
rect 19582 12178 19640 12190
rect 19700 12366 19758 12378
rect 19700 12190 19712 12366
rect 19746 12190 19758 12366
rect 19700 12178 19758 12190
rect 19818 12366 19876 12378
rect 19818 12190 19830 12366
rect 19864 12190 19876 12366
rect 19818 12178 19876 12190
rect 20606 12370 20664 12382
rect 20606 12194 20618 12370
rect 20652 12194 20664 12370
rect 20606 12182 20664 12194
rect 20724 12370 20782 12382
rect 20724 12194 20736 12370
rect 20770 12194 20782 12370
rect 20724 12182 20782 12194
rect 20842 12370 20900 12382
rect 20842 12194 20854 12370
rect 20888 12194 20900 12370
rect 20842 12182 20900 12194
rect 20960 12370 21018 12382
rect 20960 12194 20972 12370
rect 21006 12194 21018 12370
rect 20960 12182 21018 12194
rect 24091 12332 24103 12708
rect 24137 12332 24149 12708
rect 24091 12320 24149 12332
rect 24209 12708 24267 12720
rect 24209 12332 24221 12708
rect 24255 12332 24267 12708
rect 24209 12320 24267 12332
rect 24327 12708 24385 12720
rect 24327 12332 24339 12708
rect 24373 12332 24385 12708
rect 24444 12708 24502 12720
rect 24444 12532 24456 12708
rect 24490 12532 24502 12708
rect 24444 12520 24502 12532
rect 24562 12708 24620 12720
rect 24562 12532 24574 12708
rect 24608 12532 24620 12708
rect 24562 12520 24620 12532
rect 26089 12434 26147 12446
rect 24327 12320 24385 12332
rect 26089 12258 26101 12434
rect 26135 12258 26147 12434
rect 26089 12246 26147 12258
rect 26207 12434 26265 12446
rect 26207 12258 26219 12434
rect 26253 12258 26265 12434
rect 26207 12246 26265 12258
rect 26325 12434 26383 12446
rect 26325 12258 26337 12434
rect 26371 12258 26383 12434
rect 26325 12246 26383 12258
rect 26443 12434 26501 12446
rect 26443 12258 26455 12434
rect 26489 12258 26501 12434
rect 26443 12246 26501 12258
rect 27231 12438 27289 12450
rect 27231 12262 27243 12438
rect 27277 12262 27289 12438
rect 27231 12250 27289 12262
rect 27349 12438 27407 12450
rect 27349 12262 27361 12438
rect 27395 12262 27407 12438
rect 27349 12250 27407 12262
rect 27467 12438 27525 12450
rect 27467 12262 27479 12438
rect 27513 12262 27525 12438
rect 27467 12250 27525 12262
rect 27585 12438 27643 12450
rect 27585 12262 27597 12438
rect 27631 12262 27643 12438
rect 27585 12250 27643 12262
rect 29888 12069 29946 12081
rect -2379 11993 -2179 12005
rect -2379 11959 -2367 11993
rect -2191 11959 -2179 11993
rect -2379 11947 -2179 11959
rect -2379 11875 -2179 11887
rect -2379 11841 -2367 11875
rect -2191 11841 -2179 11875
rect -2379 11829 -2179 11841
rect 29888 11693 29900 12069
rect 29934 11693 29946 12069
rect 29888 11681 29946 11693
rect 30006 12069 30064 12081
rect 30006 11693 30018 12069
rect 30052 11693 30064 12069
rect 30006 11681 30064 11693
rect 30124 12069 30182 12081
rect 30124 11693 30136 12069
rect 30170 11693 30182 12069
rect 30241 12069 30299 12081
rect 30241 11893 30253 12069
rect 30287 11893 30299 12069
rect 30241 11881 30299 11893
rect 30359 12069 30417 12081
rect 30359 11893 30371 12069
rect 30405 11893 30417 12069
rect 30359 11881 30417 11893
rect 30124 11681 30182 11693
rect -2379 11573 -1979 11585
rect -2379 11539 -2367 11573
rect -1991 11539 -1979 11573
rect -2379 11527 -1979 11539
rect -2379 11455 -1979 11467
rect -2379 11421 -2367 11455
rect -1991 11421 -1979 11455
rect -2379 11409 -1979 11421
rect -2379 11337 -1979 11349
rect -2379 11303 -2367 11337
rect -1991 11303 -1979 11337
rect -2379 11291 -1979 11303
rect -2379 11219 -1979 11231
rect -2379 11185 -2367 11219
rect -1991 11185 -1979 11219
rect -2379 11173 -1979 11185
rect -2379 11101 -1979 11113
rect -2379 11067 -2367 11101
rect -1991 11067 -1979 11101
rect -2379 11055 -1979 11067
rect 38088 11692 38288 11704
rect 38088 11658 38100 11692
rect 38276 11658 38288 11692
rect 38088 11646 38288 11658
rect 38088 11574 38288 11586
rect 38088 11540 38100 11574
rect 38276 11540 38288 11574
rect 38088 11512 38288 11540
rect 38088 11500 38488 11512
rect 38088 11466 38100 11500
rect 38476 11466 38488 11500
rect 38088 11454 38488 11466
rect 10826 11058 10884 11070
rect 4277 10970 4335 10982
rect -2379 10695 -2179 10707
rect -2379 10661 -2367 10695
rect -2191 10661 -2179 10695
rect -2379 10649 -2179 10661
rect -2379 10577 -2179 10589
rect -2379 10543 -2367 10577
rect -2191 10543 -2179 10577
rect 4277 10594 4289 10970
rect 4323 10594 4335 10970
rect 4277 10582 4335 10594
rect 4395 10970 4453 10982
rect 4395 10594 4407 10970
rect 4441 10594 4453 10970
rect 4395 10582 4453 10594
rect 4513 10970 4571 10982
rect 4513 10594 4525 10970
rect 4559 10594 4571 10970
rect 4630 10970 4688 10982
rect 4630 10794 4642 10970
rect 4676 10794 4688 10970
rect 4630 10782 4688 10794
rect 4748 10970 4806 10982
rect 4748 10794 4760 10970
rect 4794 10794 4806 10970
rect 4748 10782 4806 10794
rect 4513 10582 4571 10594
rect -2379 10531 -2179 10543
rect 10826 10682 10838 11058
rect 10872 10682 10884 11058
rect 10826 10670 10884 10682
rect 10944 11058 11002 11070
rect 10944 10682 10956 11058
rect 10990 10682 11002 11058
rect 10944 10670 11002 10682
rect 11062 11058 11120 11070
rect 11062 10682 11074 11058
rect 11108 10682 11120 11058
rect 11179 11058 11237 11070
rect 11179 10882 11191 11058
rect 11225 10882 11237 11058
rect 11179 10870 11237 10882
rect 11297 11058 11355 11070
rect 11297 10882 11309 11058
rect 11343 10882 11355 11058
rect 11297 10870 11355 10882
rect 11062 10670 11120 10682
rect 1365 10302 1423 10314
rect -2381 9925 -2181 9937
rect -2381 9891 -2369 9925
rect -2193 9891 -2181 9925
rect 1365 9926 1377 10302
rect 1411 9926 1423 10302
rect 1365 9914 1423 9926
rect 1483 10302 1541 10314
rect 1483 9926 1495 10302
rect 1529 9926 1541 10302
rect 1483 9914 1541 9926
rect 1601 10302 1659 10314
rect 1601 9926 1613 10302
rect 1647 9926 1659 10302
rect 1718 10302 1776 10314
rect 1718 10126 1730 10302
rect 1764 10126 1776 10302
rect 1718 10114 1776 10126
rect 1836 10302 1894 10314
rect 1836 10126 1848 10302
rect 1882 10126 1894 10302
rect 1836 10114 1894 10126
rect 1601 9914 1659 9926
rect -2381 9879 -2181 9891
rect -2381 9807 -2181 9819
rect -2381 9773 -2369 9807
rect -2193 9773 -2181 9807
rect -2381 9761 -2181 9773
rect -2381 9505 -1981 9517
rect -2381 9471 -2369 9505
rect -1993 9471 -1981 9505
rect -2381 9459 -1981 9471
rect -2381 9387 -1981 9399
rect -2381 9353 -2369 9387
rect -1993 9353 -1981 9387
rect 38088 11382 38488 11394
rect 38088 11348 38100 11382
rect 38476 11348 38488 11382
rect 38088 11336 38488 11348
rect 38088 11264 38488 11276
rect 38088 11230 38100 11264
rect 38476 11230 38488 11264
rect 38088 11218 38488 11230
rect 38088 11146 38488 11158
rect 38088 11112 38100 11146
rect 38476 11112 38488 11146
rect 24105 11058 24163 11070
rect 17480 10990 17538 11002
rect 5629 9565 5687 9577
rect 5629 9389 5641 9565
rect 5675 9389 5687 9565
rect -2381 9341 -1981 9353
rect -2381 9269 -1981 9281
rect -2381 9235 -2369 9269
rect -1993 9235 -1981 9269
rect -2381 9223 -1981 9235
rect -2381 9151 -1981 9163
rect -2381 9117 -2369 9151
rect -1993 9117 -1981 9151
rect 4272 9366 4330 9378
rect -2381 9105 -1981 9117
rect -2381 9033 -1981 9045
rect -2381 8999 -2369 9033
rect -1993 8999 -1981 9033
rect -2381 8987 -1981 8999
rect 4272 8990 4284 9366
rect 4318 8990 4330 9366
rect 4272 8978 4330 8990
rect 4390 9366 4448 9378
rect 4390 8990 4402 9366
rect 4436 8990 4448 9366
rect 4390 8978 4448 8990
rect 4508 9366 4566 9378
rect 4508 8990 4520 9366
rect 4554 8990 4566 9366
rect 4625 9366 4683 9378
rect 4625 9190 4637 9366
rect 4671 9190 4683 9366
rect 4625 9178 4683 9190
rect 4743 9366 4801 9378
rect 5629 9377 5687 9389
rect 5747 9565 5805 9577
rect 5747 9389 5759 9565
rect 5793 9389 5805 9565
rect 5747 9377 5805 9389
rect 6049 9565 6107 9577
rect 4743 9190 4755 9366
rect 4789 9190 4801 9366
rect 4743 9178 4801 9190
rect 6049 9189 6061 9565
rect 6095 9189 6107 9565
rect 6049 9177 6107 9189
rect 6167 9565 6225 9577
rect 6167 9189 6179 9565
rect 6213 9189 6225 9565
rect 6167 9177 6225 9189
rect 6285 9565 6343 9577
rect 6285 9189 6297 9565
rect 6331 9189 6343 9565
rect 6285 9177 6343 9189
rect 6403 9565 6461 9577
rect 6403 9189 6415 9565
rect 6449 9189 6461 9565
rect 6403 9177 6461 9189
rect 6521 9565 6579 9577
rect 6521 9189 6533 9565
rect 6567 9189 6579 9565
rect 6927 9565 6985 9577
rect 6927 9389 6939 9565
rect 6973 9389 6985 9565
rect 6927 9377 6985 9389
rect 7045 9565 7103 9577
rect 7045 9389 7057 9565
rect 7091 9389 7103 9565
rect 7045 9377 7103 9389
rect 7527 9565 7585 9577
rect 7527 9389 7539 9565
rect 7573 9389 7585 9565
rect 7527 9377 7585 9389
rect 7645 9565 7703 9577
rect 7645 9389 7657 9565
rect 7691 9389 7703 9565
rect 7645 9377 7703 9389
rect 7947 9565 8005 9577
rect 6521 9177 6579 9189
rect 7947 9189 7959 9565
rect 7993 9189 8005 9565
rect 7947 9177 8005 9189
rect 8065 9565 8123 9577
rect 8065 9189 8077 9565
rect 8111 9189 8123 9565
rect 8065 9177 8123 9189
rect 8183 9565 8241 9577
rect 8183 9189 8195 9565
rect 8229 9189 8241 9565
rect 8183 9177 8241 9189
rect 8301 9565 8359 9577
rect 8301 9189 8313 9565
rect 8347 9189 8359 9565
rect 8301 9177 8359 9189
rect 8419 9565 8477 9577
rect 8419 9189 8431 9565
rect 8465 9189 8477 9565
rect 8825 9565 8883 9577
rect 8825 9389 8837 9565
rect 8871 9389 8883 9565
rect 8825 9377 8883 9389
rect 8943 9565 9001 9577
rect 8943 9389 8955 9565
rect 8989 9389 9001 9565
rect 17480 10614 17492 10990
rect 17526 10614 17538 10990
rect 17480 10602 17538 10614
rect 17598 10990 17656 11002
rect 17598 10614 17610 10990
rect 17644 10614 17656 10990
rect 17598 10602 17656 10614
rect 17716 10990 17774 11002
rect 17716 10614 17728 10990
rect 17762 10614 17774 10990
rect 17833 10990 17891 11002
rect 17833 10814 17845 10990
rect 17879 10814 17891 10990
rect 17833 10802 17891 10814
rect 17951 10990 18009 11002
rect 17951 10814 17963 10990
rect 17997 10814 18009 10990
rect 17951 10802 18009 10814
rect 17716 10602 17774 10614
rect 24105 10682 24117 11058
rect 24151 10682 24163 11058
rect 24105 10670 24163 10682
rect 24223 11058 24281 11070
rect 24223 10682 24235 11058
rect 24269 10682 24281 11058
rect 24223 10670 24281 10682
rect 24341 11058 24399 11070
rect 24341 10682 24353 11058
rect 24387 10682 24399 11058
rect 24458 11058 24516 11070
rect 24458 10882 24470 11058
rect 24504 10882 24516 11058
rect 24458 10870 24516 10882
rect 24576 11058 24634 11070
rect 24576 10882 24588 11058
rect 24622 10882 24634 11058
rect 24576 10870 24634 10882
rect 24341 10670 24399 10682
rect 12178 9653 12236 9665
rect 12178 9477 12190 9653
rect 12224 9477 12236 9653
rect 8943 9377 9001 9389
rect 10821 9454 10879 9466
rect 8419 9177 8477 9189
rect 10821 9078 10833 9454
rect 10867 9078 10879 9454
rect 4508 8978 4566 8990
rect 10821 9066 10879 9078
rect 10939 9454 10997 9466
rect 10939 9078 10951 9454
rect 10985 9078 10997 9454
rect 10939 9066 10997 9078
rect 11057 9454 11115 9466
rect 11057 9078 11069 9454
rect 11103 9078 11115 9454
rect 11174 9454 11232 9466
rect 11174 9278 11186 9454
rect 11220 9278 11232 9454
rect 11174 9266 11232 9278
rect 11292 9454 11350 9466
rect 12178 9465 12236 9477
rect 12296 9653 12354 9665
rect 12296 9477 12308 9653
rect 12342 9477 12354 9653
rect 12296 9465 12354 9477
rect 12598 9653 12656 9665
rect 11292 9278 11304 9454
rect 11338 9278 11350 9454
rect 11292 9266 11350 9278
rect 12598 9277 12610 9653
rect 12644 9277 12656 9653
rect 12598 9265 12656 9277
rect 12716 9653 12774 9665
rect 12716 9277 12728 9653
rect 12762 9277 12774 9653
rect 12716 9265 12774 9277
rect 12834 9653 12892 9665
rect 12834 9277 12846 9653
rect 12880 9277 12892 9653
rect 12834 9265 12892 9277
rect 12952 9653 13010 9665
rect 12952 9277 12964 9653
rect 12998 9277 13010 9653
rect 12952 9265 13010 9277
rect 13070 9653 13128 9665
rect 13070 9277 13082 9653
rect 13116 9277 13128 9653
rect 13476 9653 13534 9665
rect 13476 9477 13488 9653
rect 13522 9477 13534 9653
rect 13476 9465 13534 9477
rect 13594 9653 13652 9665
rect 13594 9477 13606 9653
rect 13640 9477 13652 9653
rect 13594 9465 13652 9477
rect 14076 9653 14134 9665
rect 14076 9477 14088 9653
rect 14122 9477 14134 9653
rect 14076 9465 14134 9477
rect 14194 9653 14252 9665
rect 14194 9477 14206 9653
rect 14240 9477 14252 9653
rect 14194 9465 14252 9477
rect 14496 9653 14554 9665
rect 13070 9265 13128 9277
rect 14496 9277 14508 9653
rect 14542 9277 14554 9653
rect 14496 9265 14554 9277
rect 14614 9653 14672 9665
rect 14614 9277 14626 9653
rect 14660 9277 14672 9653
rect 14614 9265 14672 9277
rect 14732 9653 14790 9665
rect 14732 9277 14744 9653
rect 14778 9277 14790 9653
rect 14732 9265 14790 9277
rect 14850 9653 14908 9665
rect 14850 9277 14862 9653
rect 14896 9277 14908 9653
rect 14850 9265 14908 9277
rect 14968 9653 15026 9665
rect 14968 9277 14980 9653
rect 15014 9277 15026 9653
rect 15374 9653 15432 9665
rect 15374 9477 15386 9653
rect 15420 9477 15432 9653
rect 15374 9465 15432 9477
rect 15492 9653 15550 9665
rect 15492 9477 15504 9653
rect 15538 9477 15550 9653
rect 15492 9465 15550 9477
rect 38088 11100 38488 11112
rect 18832 9585 18890 9597
rect 18832 9409 18844 9585
rect 18878 9409 18890 9585
rect 14968 9265 15026 9277
rect 17475 9386 17533 9398
rect 11057 9066 11115 9078
rect 17475 9010 17487 9386
rect 17521 9010 17533 9386
rect 17475 8998 17533 9010
rect 17593 9386 17651 9398
rect 17593 9010 17605 9386
rect 17639 9010 17651 9386
rect 17593 8998 17651 9010
rect 17711 9386 17769 9398
rect 17711 9010 17723 9386
rect 17757 9010 17769 9386
rect 17828 9386 17886 9398
rect 17828 9210 17840 9386
rect 17874 9210 17886 9386
rect 17828 9198 17886 9210
rect 17946 9386 18004 9398
rect 18832 9397 18890 9409
rect 18950 9585 19008 9597
rect 18950 9409 18962 9585
rect 18996 9409 19008 9585
rect 18950 9397 19008 9409
rect 19252 9585 19310 9597
rect 17946 9210 17958 9386
rect 17992 9210 18004 9386
rect 17946 9198 18004 9210
rect 19252 9209 19264 9585
rect 19298 9209 19310 9585
rect 19252 9197 19310 9209
rect 19370 9585 19428 9597
rect 19370 9209 19382 9585
rect 19416 9209 19428 9585
rect 19370 9197 19428 9209
rect 19488 9585 19546 9597
rect 19488 9209 19500 9585
rect 19534 9209 19546 9585
rect 19488 9197 19546 9209
rect 19606 9585 19664 9597
rect 19606 9209 19618 9585
rect 19652 9209 19664 9585
rect 19606 9197 19664 9209
rect 19724 9585 19782 9597
rect 19724 9209 19736 9585
rect 19770 9209 19782 9585
rect 20130 9585 20188 9597
rect 20130 9409 20142 9585
rect 20176 9409 20188 9585
rect 20130 9397 20188 9409
rect 20248 9585 20306 9597
rect 20248 9409 20260 9585
rect 20294 9409 20306 9585
rect 20248 9397 20306 9409
rect 20730 9585 20788 9597
rect 20730 9409 20742 9585
rect 20776 9409 20788 9585
rect 20730 9397 20788 9409
rect 20848 9585 20906 9597
rect 20848 9409 20860 9585
rect 20894 9409 20906 9585
rect 20848 9397 20906 9409
rect 21150 9585 21208 9597
rect 19724 9197 19782 9209
rect 21150 9209 21162 9585
rect 21196 9209 21208 9585
rect 21150 9197 21208 9209
rect 21268 9585 21326 9597
rect 21268 9209 21280 9585
rect 21314 9209 21326 9585
rect 21268 9197 21326 9209
rect 21386 9585 21444 9597
rect 21386 9209 21398 9585
rect 21432 9209 21444 9585
rect 21386 9197 21444 9209
rect 21504 9585 21562 9597
rect 21504 9209 21516 9585
rect 21550 9209 21562 9585
rect 21504 9197 21562 9209
rect 21622 9585 21680 9597
rect 21622 9209 21634 9585
rect 21668 9209 21680 9585
rect 22028 9585 22086 9597
rect 22028 9409 22040 9585
rect 22074 9409 22086 9585
rect 22028 9397 22086 9409
rect 22146 9585 22204 9597
rect 22146 9409 22158 9585
rect 22192 9409 22204 9585
rect 38088 11028 38488 11040
rect 38088 10994 38100 11028
rect 38476 10994 38488 11028
rect 38088 10982 38488 10994
rect 38088 10950 38288 10982
rect 38088 10916 38100 10950
rect 38276 10916 38288 10950
rect 38088 10904 38288 10916
rect 25457 9653 25515 9665
rect 25457 9477 25469 9653
rect 25503 9477 25515 9653
rect 22146 9397 22204 9409
rect 24100 9454 24158 9466
rect 21622 9197 21680 9209
rect 17711 8998 17769 9010
rect 24100 9078 24112 9454
rect 24146 9078 24158 9454
rect 24100 9066 24158 9078
rect 24218 9454 24276 9466
rect 24218 9078 24230 9454
rect 24264 9078 24276 9454
rect 24218 9066 24276 9078
rect 24336 9454 24394 9466
rect 24336 9078 24348 9454
rect 24382 9078 24394 9454
rect 24453 9454 24511 9466
rect 24453 9278 24465 9454
rect 24499 9278 24511 9454
rect 24453 9266 24511 9278
rect 24571 9454 24629 9466
rect 25457 9465 25515 9477
rect 25575 9653 25633 9665
rect 25575 9477 25587 9653
rect 25621 9477 25633 9653
rect 25575 9465 25633 9477
rect 25877 9653 25935 9665
rect 24571 9278 24583 9454
rect 24617 9278 24629 9454
rect 24571 9266 24629 9278
rect 25877 9277 25889 9653
rect 25923 9277 25935 9653
rect 25877 9265 25935 9277
rect 25995 9653 26053 9665
rect 25995 9277 26007 9653
rect 26041 9277 26053 9653
rect 25995 9265 26053 9277
rect 26113 9653 26171 9665
rect 26113 9277 26125 9653
rect 26159 9277 26171 9653
rect 26113 9265 26171 9277
rect 26231 9653 26289 9665
rect 26231 9277 26243 9653
rect 26277 9277 26289 9653
rect 26231 9265 26289 9277
rect 26349 9653 26407 9665
rect 26349 9277 26361 9653
rect 26395 9277 26407 9653
rect 26755 9653 26813 9665
rect 26755 9477 26767 9653
rect 26801 9477 26813 9653
rect 26755 9465 26813 9477
rect 26873 9653 26931 9665
rect 26873 9477 26885 9653
rect 26919 9477 26931 9653
rect 26873 9465 26931 9477
rect 27355 9653 27413 9665
rect 27355 9477 27367 9653
rect 27401 9477 27413 9653
rect 27355 9465 27413 9477
rect 27473 9653 27531 9665
rect 27473 9477 27485 9653
rect 27519 9477 27531 9653
rect 27473 9465 27531 9477
rect 27775 9653 27833 9665
rect 26349 9265 26407 9277
rect 27775 9277 27787 9653
rect 27821 9277 27833 9653
rect 27775 9265 27833 9277
rect 27893 9653 27951 9665
rect 27893 9277 27905 9653
rect 27939 9277 27951 9653
rect 27893 9265 27951 9277
rect 28011 9653 28069 9665
rect 28011 9277 28023 9653
rect 28057 9277 28069 9653
rect 28011 9265 28069 9277
rect 28129 9653 28187 9665
rect 28129 9277 28141 9653
rect 28175 9277 28187 9653
rect 28129 9265 28187 9277
rect 28247 9653 28305 9665
rect 28247 9277 28259 9653
rect 28293 9277 28305 9653
rect 28653 9653 28711 9665
rect 28653 9477 28665 9653
rect 28699 9477 28711 9653
rect 28653 9465 28711 9477
rect 28771 9653 28829 9665
rect 28771 9477 28783 9653
rect 28817 9477 28829 9653
rect 28771 9465 28829 9477
rect 33496 10141 33554 10153
rect 33496 9765 33508 10141
rect 33542 9765 33554 10141
rect 33496 9753 33554 9765
rect 33614 10141 33672 10153
rect 33614 9765 33626 10141
rect 33660 9765 33672 10141
rect 33614 9753 33672 9765
rect 33732 10141 33790 10153
rect 33732 9765 33744 10141
rect 33778 9765 33790 10141
rect 33849 10141 33907 10153
rect 33849 9965 33861 10141
rect 33895 9965 33907 10141
rect 33849 9953 33907 9965
rect 33967 10141 34025 10153
rect 33967 9965 33979 10141
rect 34013 9965 34025 10141
rect 38088 10832 38288 10844
rect 38088 10798 38100 10832
rect 38276 10798 38288 10832
rect 38088 10786 38288 10798
rect 33967 9953 34025 9965
rect 33732 9753 33790 9765
rect 31591 9356 31649 9368
rect 28247 9265 28305 9277
rect 24336 9066 24394 9078
rect 31591 9180 31603 9356
rect 31637 9180 31649 9356
rect 31591 9168 31649 9180
rect 31709 9356 31767 9368
rect 31709 9180 31721 9356
rect 31755 9180 31767 9356
rect 31709 9168 31767 9180
rect 32011 9356 32069 9368
rect 29888 9036 29946 9048
rect 29888 8660 29900 9036
rect 29934 8660 29946 9036
rect 29888 8648 29946 8660
rect 30006 9036 30064 9048
rect 30006 8660 30018 9036
rect 30052 8660 30064 9036
rect 30006 8648 30064 8660
rect 30124 9036 30182 9048
rect 30124 8660 30136 9036
rect 30170 8660 30182 9036
rect 30241 9036 30299 9048
rect 30241 8860 30253 9036
rect 30287 8860 30299 9036
rect 30241 8848 30299 8860
rect 30359 9036 30417 9048
rect 30359 8860 30371 9036
rect 30405 8860 30417 9036
rect 32011 8980 32023 9356
rect 32057 8980 32069 9356
rect 32011 8968 32069 8980
rect 32129 9356 32187 9368
rect 32129 8980 32141 9356
rect 32175 8980 32187 9356
rect 32129 8968 32187 8980
rect 32247 9356 32305 9368
rect 32247 8980 32259 9356
rect 32293 8980 32305 9356
rect 32247 8968 32305 8980
rect 32365 9356 32423 9368
rect 32365 8980 32377 9356
rect 32411 8980 32423 9356
rect 32365 8968 32423 8980
rect 32483 9356 32541 9368
rect 32483 8980 32495 9356
rect 32529 8980 32541 9356
rect 32889 9356 32947 9368
rect 32889 9180 32901 9356
rect 32935 9180 32947 9356
rect 32889 9168 32947 9180
rect 33007 9356 33065 9368
rect 33007 9180 33019 9356
rect 33053 9180 33065 9356
rect 33007 9168 33065 9180
rect 32483 8968 32541 8980
rect 30359 8848 30417 8860
rect 30124 8648 30182 8660
rect -2381 8627 -2181 8639
rect -2381 8593 -2369 8627
rect -2193 8593 -2181 8627
rect -2381 8581 -2181 8593
rect -2381 8509 -2181 8521
rect -2381 8475 -2369 8509
rect -2193 8475 -2181 8509
rect -2381 8463 -2181 8475
rect 38088 8548 38288 8560
rect 38088 8514 38100 8548
rect 38276 8514 38288 8548
rect 38088 8502 38288 8514
rect 38088 8430 38288 8442
rect 38088 8396 38100 8430
rect 38276 8396 38288 8430
rect 38088 8368 38288 8396
rect 38088 8356 38488 8368
rect 38088 8322 38100 8356
rect 38476 8322 38488 8356
rect 38088 8310 38488 8322
rect 38088 8238 38488 8250
rect 38088 8204 38100 8238
rect 38476 8204 38488 8238
rect 38088 8192 38488 8204
rect 38088 8120 38488 8132
rect 38088 8086 38100 8120
rect 38476 8086 38488 8120
rect 38088 8074 38488 8086
rect 38088 8002 38488 8014
rect 38088 7968 38100 8002
rect 38476 7968 38488 8002
rect 38088 7956 38488 7968
rect -2381 7856 -2181 7868
rect -2381 7822 -2369 7856
rect -2193 7822 -2181 7856
rect -2381 7810 -2181 7822
rect -2381 7738 -2181 7750
rect -2381 7704 -2369 7738
rect -2193 7704 -2181 7738
rect -2381 7692 -2181 7704
rect -2381 7436 -1981 7448
rect -2381 7402 -2369 7436
rect -1993 7402 -1981 7436
rect -2381 7390 -1981 7402
rect -2381 7318 -1981 7330
rect -2381 7284 -2369 7318
rect -1993 7284 -1981 7318
rect -2381 7272 -1981 7284
rect -2381 7200 -1981 7212
rect -2381 7166 -2369 7200
rect -1993 7166 -1981 7200
rect -2381 7154 -1981 7166
rect -2381 7082 -1981 7094
rect -2381 7048 -2369 7082
rect -1993 7048 -1981 7082
rect -2381 7036 -1981 7048
rect 1346 7024 1404 7036
rect -2381 6964 -1981 6976
rect -2381 6930 -2369 6964
rect -1993 6930 -1981 6964
rect -2381 6918 -1981 6930
rect 1346 6648 1358 7024
rect 1392 6648 1404 7024
rect 1346 6636 1404 6648
rect 1464 7024 1522 7036
rect 1464 6648 1476 7024
rect 1510 6648 1522 7024
rect 1464 6636 1522 6648
rect 1582 7024 1640 7036
rect 1582 6648 1594 7024
rect 1628 6648 1640 7024
rect 1699 7024 1757 7036
rect 1699 6848 1711 7024
rect 1745 6848 1757 7024
rect 1699 6836 1757 6848
rect 1817 7024 1875 7036
rect 1817 6848 1829 7024
rect 1863 6848 1875 7024
rect 1817 6836 1875 6848
rect 4255 6840 4313 6852
rect 1582 6636 1640 6648
rect -2381 6558 -2181 6570
rect -2381 6524 -2369 6558
rect -2193 6524 -2181 6558
rect -2381 6512 -2181 6524
rect -2381 6440 -2181 6452
rect -2381 6406 -2369 6440
rect -2193 6406 -2181 6440
rect 4255 6464 4267 6840
rect 4301 6464 4313 6840
rect 4255 6452 4313 6464
rect 4373 6840 4431 6852
rect 4373 6464 4385 6840
rect 4419 6464 4431 6840
rect 4373 6452 4431 6464
rect 4491 6840 4549 6852
rect 4491 6464 4503 6840
rect 4537 6464 4549 6840
rect 4608 6840 4666 6852
rect 4608 6664 4620 6840
rect 4654 6664 4666 6840
rect 4608 6652 4666 6664
rect 4726 6840 4784 6852
rect 4726 6664 4738 6840
rect 4772 6664 4784 6840
rect 4726 6652 4784 6664
rect 10806 6838 10864 6850
rect 6253 6566 6311 6578
rect 4491 6452 4549 6464
rect -2381 6394 -2181 6406
rect 6253 6390 6265 6566
rect 6299 6390 6311 6566
rect 6253 6378 6311 6390
rect 6371 6566 6429 6578
rect 6371 6390 6383 6566
rect 6417 6390 6429 6566
rect 6371 6378 6429 6390
rect 6489 6566 6547 6578
rect 6489 6390 6501 6566
rect 6535 6390 6547 6566
rect 6489 6378 6547 6390
rect 6607 6566 6665 6578
rect 6607 6390 6619 6566
rect 6653 6390 6665 6566
rect 6607 6378 6665 6390
rect 7395 6570 7453 6582
rect 7395 6394 7407 6570
rect 7441 6394 7453 6570
rect 7395 6382 7453 6394
rect 7513 6570 7571 6582
rect 7513 6394 7525 6570
rect 7559 6394 7571 6570
rect 7513 6382 7571 6394
rect 7631 6570 7689 6582
rect 7631 6394 7643 6570
rect 7677 6394 7689 6570
rect 7631 6382 7689 6394
rect 7749 6570 7807 6582
rect 7749 6394 7761 6570
rect 7795 6394 7807 6570
rect 7749 6382 7807 6394
rect 10806 6462 10818 6838
rect 10852 6462 10864 6838
rect 10806 6450 10864 6462
rect 10924 6838 10982 6850
rect 10924 6462 10936 6838
rect 10970 6462 10982 6838
rect 10924 6450 10982 6462
rect 11042 6838 11100 6850
rect 11042 6462 11054 6838
rect 11088 6462 11100 6838
rect 11159 6838 11217 6850
rect 11159 6662 11171 6838
rect 11205 6662 11217 6838
rect 11159 6650 11217 6662
rect 11277 6838 11335 6850
rect 11277 6662 11289 6838
rect 11323 6662 11335 6838
rect 11277 6650 11335 6662
rect 38088 7884 38488 7896
rect 38088 7850 38100 7884
rect 38476 7850 38488 7884
rect 38088 7838 38488 7850
rect 38088 7806 38288 7838
rect 38088 7772 38100 7806
rect 38276 7772 38288 7806
rect 38088 7760 38288 7772
rect 17461 6839 17519 6851
rect 12804 6564 12862 6576
rect 11042 6450 11100 6462
rect 12804 6388 12816 6564
rect 12850 6388 12862 6564
rect 12804 6376 12862 6388
rect 12922 6564 12980 6576
rect 12922 6388 12934 6564
rect 12968 6388 12980 6564
rect 12922 6376 12980 6388
rect 13040 6564 13098 6576
rect 13040 6388 13052 6564
rect 13086 6388 13098 6564
rect 13040 6376 13098 6388
rect 13158 6564 13216 6576
rect 13158 6388 13170 6564
rect 13204 6388 13216 6564
rect 13158 6376 13216 6388
rect 13946 6568 14004 6580
rect 13946 6392 13958 6568
rect 13992 6392 14004 6568
rect 13946 6380 14004 6392
rect 14064 6568 14122 6580
rect 14064 6392 14076 6568
rect 14110 6392 14122 6568
rect 14064 6380 14122 6392
rect 14182 6568 14240 6580
rect 14182 6392 14194 6568
rect 14228 6392 14240 6568
rect 14182 6380 14240 6392
rect 14300 6568 14358 6580
rect 14300 6392 14312 6568
rect 14346 6392 14358 6568
rect 14300 6380 14358 6392
rect 17461 6463 17473 6839
rect 17507 6463 17519 6839
rect 17461 6451 17519 6463
rect 17579 6839 17637 6851
rect 17579 6463 17591 6839
rect 17625 6463 17637 6839
rect 17579 6451 17637 6463
rect 17697 6839 17755 6851
rect 17697 6463 17709 6839
rect 17743 6463 17755 6839
rect 17814 6839 17872 6851
rect 17814 6663 17826 6839
rect 17860 6663 17872 6839
rect 17814 6651 17872 6663
rect 17932 6839 17990 6851
rect 17932 6663 17944 6839
rect 17978 6663 17990 6839
rect 17932 6651 17990 6663
rect 29959 7116 30017 7128
rect 24083 6840 24141 6852
rect 19459 6565 19517 6577
rect 17697 6451 17755 6463
rect 19459 6389 19471 6565
rect 19505 6389 19517 6565
rect 19459 6377 19517 6389
rect 19577 6565 19635 6577
rect 19577 6389 19589 6565
rect 19623 6389 19635 6565
rect 19577 6377 19635 6389
rect 19695 6565 19753 6577
rect 19695 6389 19707 6565
rect 19741 6389 19753 6565
rect 19695 6377 19753 6389
rect 19813 6565 19871 6577
rect 19813 6389 19825 6565
rect 19859 6389 19871 6565
rect 19813 6377 19871 6389
rect 20601 6569 20659 6581
rect 20601 6393 20613 6569
rect 20647 6393 20659 6569
rect 20601 6381 20659 6393
rect 20719 6569 20777 6581
rect 20719 6393 20731 6569
rect 20765 6393 20777 6569
rect 20719 6381 20777 6393
rect 20837 6569 20895 6581
rect 20837 6393 20849 6569
rect 20883 6393 20895 6569
rect 20837 6381 20895 6393
rect 20955 6569 21013 6581
rect 20955 6393 20967 6569
rect 21001 6393 21013 6569
rect 20955 6381 21013 6393
rect 24083 6464 24095 6840
rect 24129 6464 24141 6840
rect 24083 6452 24141 6464
rect 24201 6840 24259 6852
rect 24201 6464 24213 6840
rect 24247 6464 24259 6840
rect 24201 6452 24259 6464
rect 24319 6840 24377 6852
rect 24319 6464 24331 6840
rect 24365 6464 24377 6840
rect 24436 6840 24494 6852
rect 24436 6664 24448 6840
rect 24482 6664 24494 6840
rect 24436 6652 24494 6664
rect 24554 6840 24612 6852
rect 24554 6664 24566 6840
rect 24600 6664 24612 6840
rect 24554 6652 24612 6664
rect 29959 6740 29971 7116
rect 30005 6740 30017 7116
rect 29959 6728 30017 6740
rect 30077 7116 30135 7128
rect 30077 6740 30089 7116
rect 30123 6740 30135 7116
rect 30077 6728 30135 6740
rect 30195 7116 30253 7128
rect 30195 6740 30207 7116
rect 30241 6740 30253 7116
rect 30312 7116 30370 7128
rect 30312 6940 30324 7116
rect 30358 6940 30370 7116
rect 30312 6928 30370 6940
rect 30430 7116 30488 7128
rect 30430 6940 30442 7116
rect 30476 6940 30488 7116
rect 30430 6928 30488 6940
rect 30195 6728 30253 6740
rect 26081 6566 26139 6578
rect 24319 6452 24377 6464
rect 26081 6390 26093 6566
rect 26127 6390 26139 6566
rect 26081 6378 26139 6390
rect 26199 6566 26257 6578
rect 26199 6390 26211 6566
rect 26245 6390 26257 6566
rect 26199 6378 26257 6390
rect 26317 6566 26375 6578
rect 26317 6390 26329 6566
rect 26363 6390 26375 6566
rect 26317 6378 26375 6390
rect 26435 6566 26493 6578
rect 26435 6390 26447 6566
rect 26481 6390 26493 6566
rect 26435 6378 26493 6390
rect 27223 6570 27281 6582
rect 27223 6394 27235 6570
rect 27269 6394 27281 6570
rect 27223 6382 27281 6394
rect 27341 6570 27399 6582
rect 27341 6394 27353 6570
rect 27387 6394 27399 6570
rect 27341 6382 27399 6394
rect 27459 6570 27517 6582
rect 27459 6394 27471 6570
rect 27505 6394 27517 6570
rect 27459 6382 27517 6394
rect 27577 6570 27635 6582
rect 27577 6394 27589 6570
rect 27623 6394 27635 6570
rect 27577 6382 27635 6394
rect 38088 7688 38288 7700
rect 38088 7654 38100 7688
rect 38276 7654 38288 7688
rect 38088 7642 38288 7654
rect 33496 6646 33554 6658
rect 33496 6270 33508 6646
rect 33542 6270 33554 6646
rect 33496 6258 33554 6270
rect 33614 6646 33672 6658
rect 33614 6270 33626 6646
rect 33660 6270 33672 6646
rect 33614 6258 33672 6270
rect 33732 6646 33790 6658
rect 33732 6270 33744 6646
rect 33778 6270 33790 6646
rect 33849 6646 33907 6658
rect 33849 6470 33861 6646
rect 33895 6470 33907 6646
rect 33849 6458 33907 6470
rect 33967 6646 34025 6658
rect 33967 6470 33979 6646
rect 34013 6470 34025 6646
rect 33967 6458 34025 6470
rect 33732 6258 33790 6270
rect 31591 5861 31649 5873
rect -2383 5788 -2183 5800
rect -2383 5754 -2371 5788
rect -2195 5754 -2183 5788
rect -2383 5742 -2183 5754
rect -2383 5670 -2183 5682
rect -2383 5636 -2371 5670
rect -2195 5636 -2183 5670
rect -2383 5624 -2183 5636
rect -2383 5368 -1983 5380
rect -2383 5334 -2371 5368
rect -1995 5334 -1983 5368
rect -2383 5322 -1983 5334
rect -2383 5250 -1983 5262
rect -2383 5216 -2371 5250
rect -1995 5216 -1983 5250
rect -2383 5204 -1983 5216
rect 31591 5685 31603 5861
rect 31637 5685 31649 5861
rect 31591 5673 31649 5685
rect 31709 5861 31767 5873
rect 31709 5685 31721 5861
rect 31755 5685 31767 5861
rect 31709 5673 31767 5685
rect 32011 5861 32069 5873
rect 32011 5485 32023 5861
rect 32057 5485 32069 5861
rect 32011 5473 32069 5485
rect 32129 5861 32187 5873
rect 32129 5485 32141 5861
rect 32175 5485 32187 5861
rect 32129 5473 32187 5485
rect 32247 5861 32305 5873
rect 32247 5485 32259 5861
rect 32293 5485 32305 5861
rect 32247 5473 32305 5485
rect 32365 5861 32423 5873
rect 32365 5485 32377 5861
rect 32411 5485 32423 5861
rect 32365 5473 32423 5485
rect 32483 5861 32541 5873
rect 32483 5485 32495 5861
rect 32529 5485 32541 5861
rect 32889 5861 32947 5873
rect 32889 5685 32901 5861
rect 32935 5685 32947 5861
rect 32889 5673 32947 5685
rect 33007 5861 33065 5873
rect 33007 5685 33019 5861
rect 33053 5685 33065 5861
rect 33007 5673 33065 5685
rect 32483 5473 32541 5485
rect -2383 5132 -1983 5144
rect -2383 5098 -2371 5132
rect -1995 5098 -1983 5132
rect -2383 5086 -1983 5098
rect -2383 5014 -1983 5026
rect -2383 4980 -2371 5014
rect -1995 4980 -1983 5014
rect 4269 5190 4327 5202
rect -2383 4968 -1983 4980
rect -2383 4896 -1983 4908
rect -2383 4862 -2371 4896
rect -1995 4862 -1983 4896
rect -2383 4850 -1983 4862
rect 4269 4814 4281 5190
rect 4315 4814 4327 5190
rect 4269 4802 4327 4814
rect 4387 5190 4445 5202
rect 4387 4814 4399 5190
rect 4433 4814 4445 5190
rect 4387 4802 4445 4814
rect 4505 5190 4563 5202
rect 4505 4814 4517 5190
rect 4551 4814 4563 5190
rect 4622 5190 4680 5202
rect 4622 5014 4634 5190
rect 4668 5014 4680 5190
rect 4622 5002 4680 5014
rect 4740 5190 4798 5202
rect 4740 5014 4752 5190
rect 4786 5014 4798 5190
rect 4740 5002 4798 5014
rect 4505 4802 4563 4814
rect 10820 5188 10878 5200
rect -2383 4490 -2183 4502
rect -2383 4456 -2371 4490
rect -2195 4456 -2183 4490
rect -2383 4444 -2183 4456
rect -2383 4372 -2183 4384
rect -2383 4338 -2371 4372
rect -2195 4338 -2183 4372
rect -2383 4326 -2183 4338
rect 1362 4264 1420 4276
rect 1362 3888 1374 4264
rect 1408 3888 1420 4264
rect 1362 3876 1420 3888
rect 1480 4264 1538 4276
rect 1480 3888 1492 4264
rect 1526 3888 1538 4264
rect 1480 3876 1538 3888
rect 1598 4264 1656 4276
rect 1598 3888 1610 4264
rect 1644 3888 1656 4264
rect 1715 4264 1773 4276
rect 1715 4088 1727 4264
rect 1761 4088 1773 4264
rect 1715 4076 1773 4088
rect 1833 4264 1891 4276
rect 1833 4088 1845 4264
rect 1879 4088 1891 4264
rect 1833 4076 1891 4088
rect 1598 3876 1656 3888
rect -2381 3719 -2181 3731
rect -2381 3685 -2369 3719
rect -2193 3685 -2181 3719
rect -2381 3673 -2181 3685
rect -2381 3601 -2181 3613
rect -2381 3567 -2369 3601
rect -2193 3567 -2181 3601
rect 10820 4812 10832 5188
rect 10866 4812 10878 5188
rect 10820 4800 10878 4812
rect 10938 5188 10996 5200
rect 10938 4812 10950 5188
rect 10984 4812 10996 5188
rect 10938 4800 10996 4812
rect 11056 5188 11114 5200
rect 11056 4812 11068 5188
rect 11102 4812 11114 5188
rect 11173 5188 11231 5200
rect 11173 5012 11185 5188
rect 11219 5012 11231 5188
rect 11173 5000 11231 5012
rect 11291 5188 11349 5200
rect 11291 5012 11303 5188
rect 11337 5012 11349 5188
rect 11291 5000 11349 5012
rect 11056 4800 11114 4812
rect 17475 5189 17533 5201
rect 5621 3785 5679 3797
rect 5621 3609 5633 3785
rect 5667 3609 5679 3785
rect -2381 3555 -2181 3567
rect 4264 3586 4322 3598
rect -2381 3299 -1981 3311
rect -2381 3265 -2369 3299
rect -1993 3265 -1981 3299
rect -2381 3253 -1981 3265
rect 4264 3210 4276 3586
rect 4310 3210 4322 3586
rect 4264 3198 4322 3210
rect 4382 3586 4440 3598
rect 4382 3210 4394 3586
rect 4428 3210 4440 3586
rect 4382 3198 4440 3210
rect 4500 3586 4558 3598
rect 4500 3210 4512 3586
rect 4546 3210 4558 3586
rect 4617 3586 4675 3598
rect 4617 3410 4629 3586
rect 4663 3410 4675 3586
rect 4617 3398 4675 3410
rect 4735 3586 4793 3598
rect 5621 3597 5679 3609
rect 5739 3785 5797 3797
rect 5739 3609 5751 3785
rect 5785 3609 5797 3785
rect 5739 3597 5797 3609
rect 6041 3785 6099 3797
rect 4735 3410 4747 3586
rect 4781 3410 4793 3586
rect 4735 3398 4793 3410
rect 6041 3409 6053 3785
rect 6087 3409 6099 3785
rect 6041 3397 6099 3409
rect 6159 3785 6217 3797
rect 6159 3409 6171 3785
rect 6205 3409 6217 3785
rect 6159 3397 6217 3409
rect 6277 3785 6335 3797
rect 6277 3409 6289 3785
rect 6323 3409 6335 3785
rect 6277 3397 6335 3409
rect 6395 3785 6453 3797
rect 6395 3409 6407 3785
rect 6441 3409 6453 3785
rect 6395 3397 6453 3409
rect 6513 3785 6571 3797
rect 6513 3409 6525 3785
rect 6559 3409 6571 3785
rect 6919 3785 6977 3797
rect 6919 3609 6931 3785
rect 6965 3609 6977 3785
rect 6919 3597 6977 3609
rect 7037 3785 7095 3797
rect 7037 3609 7049 3785
rect 7083 3609 7095 3785
rect 7037 3597 7095 3609
rect 7519 3785 7577 3797
rect 7519 3609 7531 3785
rect 7565 3609 7577 3785
rect 7519 3597 7577 3609
rect 7637 3785 7695 3797
rect 7637 3609 7649 3785
rect 7683 3609 7695 3785
rect 7637 3597 7695 3609
rect 7939 3785 7997 3797
rect 6513 3397 6571 3409
rect 7939 3409 7951 3785
rect 7985 3409 7997 3785
rect 7939 3397 7997 3409
rect 8057 3785 8115 3797
rect 8057 3409 8069 3785
rect 8103 3409 8115 3785
rect 8057 3397 8115 3409
rect 8175 3785 8233 3797
rect 8175 3409 8187 3785
rect 8221 3409 8233 3785
rect 8175 3397 8233 3409
rect 8293 3785 8351 3797
rect 8293 3409 8305 3785
rect 8339 3409 8351 3785
rect 8293 3397 8351 3409
rect 8411 3785 8469 3797
rect 8411 3409 8423 3785
rect 8457 3409 8469 3785
rect 8817 3785 8875 3797
rect 8817 3609 8829 3785
rect 8863 3609 8875 3785
rect 8817 3597 8875 3609
rect 8935 3785 8993 3797
rect 8935 3609 8947 3785
rect 8981 3609 8993 3785
rect 8935 3597 8993 3609
rect 17475 4813 17487 5189
rect 17521 4813 17533 5189
rect 17475 4801 17533 4813
rect 17593 5189 17651 5201
rect 17593 4813 17605 5189
rect 17639 4813 17651 5189
rect 17593 4801 17651 4813
rect 17711 5189 17769 5201
rect 17711 4813 17723 5189
rect 17757 4813 17769 5189
rect 17828 5189 17886 5201
rect 17828 5013 17840 5189
rect 17874 5013 17886 5189
rect 17828 5001 17886 5013
rect 17946 5189 18004 5201
rect 17946 5013 17958 5189
rect 17992 5013 18004 5189
rect 17946 5001 18004 5013
rect 17711 4801 17769 4813
rect 24097 5190 24155 5202
rect 12172 3783 12230 3795
rect 12172 3607 12184 3783
rect 12218 3607 12230 3783
rect 10815 3584 10873 3596
rect 8411 3397 8469 3409
rect 4500 3198 4558 3210
rect -2381 3181 -1981 3193
rect -2381 3147 -2369 3181
rect -1993 3147 -1981 3181
rect -2381 3135 -1981 3147
rect 10815 3208 10827 3584
rect 10861 3208 10873 3584
rect 10815 3196 10873 3208
rect 10933 3584 10991 3596
rect 10933 3208 10945 3584
rect 10979 3208 10991 3584
rect 10933 3196 10991 3208
rect 11051 3584 11109 3596
rect 11051 3208 11063 3584
rect 11097 3208 11109 3584
rect 11168 3584 11226 3596
rect 11168 3408 11180 3584
rect 11214 3408 11226 3584
rect 11168 3396 11226 3408
rect 11286 3584 11344 3596
rect 12172 3595 12230 3607
rect 12290 3783 12348 3795
rect 12290 3607 12302 3783
rect 12336 3607 12348 3783
rect 12290 3595 12348 3607
rect 12592 3783 12650 3795
rect 11286 3408 11298 3584
rect 11332 3408 11344 3584
rect 11286 3396 11344 3408
rect 12592 3407 12604 3783
rect 12638 3407 12650 3783
rect 12592 3395 12650 3407
rect 12710 3783 12768 3795
rect 12710 3407 12722 3783
rect 12756 3407 12768 3783
rect 12710 3395 12768 3407
rect 12828 3783 12886 3795
rect 12828 3407 12840 3783
rect 12874 3407 12886 3783
rect 12828 3395 12886 3407
rect 12946 3783 13004 3795
rect 12946 3407 12958 3783
rect 12992 3407 13004 3783
rect 12946 3395 13004 3407
rect 13064 3783 13122 3795
rect 13064 3407 13076 3783
rect 13110 3407 13122 3783
rect 13470 3783 13528 3795
rect 13470 3607 13482 3783
rect 13516 3607 13528 3783
rect 13470 3595 13528 3607
rect 13588 3783 13646 3795
rect 13588 3607 13600 3783
rect 13634 3607 13646 3783
rect 13588 3595 13646 3607
rect 14070 3783 14128 3795
rect 14070 3607 14082 3783
rect 14116 3607 14128 3783
rect 14070 3595 14128 3607
rect 14188 3783 14246 3795
rect 14188 3607 14200 3783
rect 14234 3607 14246 3783
rect 14188 3595 14246 3607
rect 14490 3783 14548 3795
rect 13064 3395 13122 3407
rect 14490 3407 14502 3783
rect 14536 3407 14548 3783
rect 14490 3395 14548 3407
rect 14608 3783 14666 3795
rect 14608 3407 14620 3783
rect 14654 3407 14666 3783
rect 14608 3395 14666 3407
rect 14726 3783 14784 3795
rect 14726 3407 14738 3783
rect 14772 3407 14784 3783
rect 14726 3395 14784 3407
rect 14844 3783 14902 3795
rect 14844 3407 14856 3783
rect 14890 3407 14902 3783
rect 14844 3395 14902 3407
rect 14962 3783 15020 3795
rect 14962 3407 14974 3783
rect 15008 3407 15020 3783
rect 15368 3783 15426 3795
rect 15368 3607 15380 3783
rect 15414 3607 15426 3783
rect 15368 3595 15426 3607
rect 15486 3783 15544 3795
rect 15486 3607 15498 3783
rect 15532 3607 15544 3783
rect 15486 3595 15544 3607
rect 24097 4814 24109 5190
rect 24143 4814 24155 5190
rect 24097 4802 24155 4814
rect 24215 5190 24273 5202
rect 24215 4814 24227 5190
rect 24261 4814 24273 5190
rect 24215 4802 24273 4814
rect 24333 5190 24391 5202
rect 24333 4814 24345 5190
rect 24379 4814 24391 5190
rect 24450 5190 24508 5202
rect 24450 5014 24462 5190
rect 24496 5014 24508 5190
rect 24450 5002 24508 5014
rect 24568 5190 24626 5202
rect 24568 5014 24580 5190
rect 24614 5014 24626 5190
rect 24568 5002 24626 5014
rect 24333 4802 24391 4814
rect 38084 5416 38284 5428
rect 38084 5382 38096 5416
rect 38272 5382 38284 5416
rect 38084 5370 38284 5382
rect 38084 5298 38284 5310
rect 38084 5264 38096 5298
rect 38272 5264 38284 5298
rect 38084 5236 38284 5264
rect 38084 5224 38484 5236
rect 38084 5190 38096 5224
rect 38472 5190 38484 5224
rect 38084 5178 38484 5190
rect 38084 5106 38484 5118
rect 38084 5072 38096 5106
rect 38472 5072 38484 5106
rect 38084 5060 38484 5072
rect 18827 3784 18885 3796
rect 18827 3608 18839 3784
rect 18873 3608 18885 3784
rect 17470 3585 17528 3597
rect 14962 3395 15020 3407
rect 11051 3196 11109 3208
rect -2381 3063 -1981 3075
rect -2381 3029 -2369 3063
rect -1993 3029 -1981 3063
rect -2381 3017 -1981 3029
rect -2381 2945 -1981 2957
rect -2381 2911 -2369 2945
rect -1993 2911 -1981 2945
rect 17470 3209 17482 3585
rect 17516 3209 17528 3585
rect 17470 3197 17528 3209
rect 17588 3585 17646 3597
rect 17588 3209 17600 3585
rect 17634 3209 17646 3585
rect 17588 3197 17646 3209
rect 17706 3585 17764 3597
rect 17706 3209 17718 3585
rect 17752 3209 17764 3585
rect 17823 3585 17881 3597
rect 17823 3409 17835 3585
rect 17869 3409 17881 3585
rect 17823 3397 17881 3409
rect 17941 3585 17999 3597
rect 18827 3596 18885 3608
rect 18945 3784 19003 3796
rect 18945 3608 18957 3784
rect 18991 3608 19003 3784
rect 18945 3596 19003 3608
rect 19247 3784 19305 3796
rect 17941 3409 17953 3585
rect 17987 3409 17999 3585
rect 17941 3397 17999 3409
rect 19247 3408 19259 3784
rect 19293 3408 19305 3784
rect 19247 3396 19305 3408
rect 19365 3784 19423 3796
rect 19365 3408 19377 3784
rect 19411 3408 19423 3784
rect 19365 3396 19423 3408
rect 19483 3784 19541 3796
rect 19483 3408 19495 3784
rect 19529 3408 19541 3784
rect 19483 3396 19541 3408
rect 19601 3784 19659 3796
rect 19601 3408 19613 3784
rect 19647 3408 19659 3784
rect 19601 3396 19659 3408
rect 19719 3784 19777 3796
rect 19719 3408 19731 3784
rect 19765 3408 19777 3784
rect 20125 3784 20183 3796
rect 20125 3608 20137 3784
rect 20171 3608 20183 3784
rect 20125 3596 20183 3608
rect 20243 3784 20301 3796
rect 20243 3608 20255 3784
rect 20289 3608 20301 3784
rect 20243 3596 20301 3608
rect 20725 3784 20783 3796
rect 20725 3608 20737 3784
rect 20771 3608 20783 3784
rect 20725 3596 20783 3608
rect 20843 3784 20901 3796
rect 20843 3608 20855 3784
rect 20889 3608 20901 3784
rect 20843 3596 20901 3608
rect 21145 3784 21203 3796
rect 19719 3396 19777 3408
rect 21145 3408 21157 3784
rect 21191 3408 21203 3784
rect 21145 3396 21203 3408
rect 21263 3784 21321 3796
rect 21263 3408 21275 3784
rect 21309 3408 21321 3784
rect 21263 3396 21321 3408
rect 21381 3784 21439 3796
rect 21381 3408 21393 3784
rect 21427 3408 21439 3784
rect 21381 3396 21439 3408
rect 21499 3784 21557 3796
rect 21499 3408 21511 3784
rect 21545 3408 21557 3784
rect 21499 3396 21557 3408
rect 21617 3784 21675 3796
rect 21617 3408 21629 3784
rect 21663 3408 21675 3784
rect 22023 3784 22081 3796
rect 22023 3608 22035 3784
rect 22069 3608 22081 3784
rect 22023 3596 22081 3608
rect 22141 3784 22199 3796
rect 22141 3608 22153 3784
rect 22187 3608 22199 3784
rect 22141 3596 22199 3608
rect 38084 4988 38484 5000
rect 38084 4954 38096 4988
rect 38472 4954 38484 4988
rect 38084 4942 38484 4954
rect 38084 4870 38484 4882
rect 38084 4836 38096 4870
rect 38472 4836 38484 4870
rect 38084 4824 38484 4836
rect 38084 4752 38484 4764
rect 38084 4718 38096 4752
rect 38472 4718 38484 4752
rect 38084 4706 38484 4718
rect 38084 4674 38284 4706
rect 38084 4640 38096 4674
rect 38272 4640 38284 4674
rect 38084 4628 38284 4640
rect 29956 4046 30014 4058
rect 25449 3785 25507 3797
rect 25449 3609 25461 3785
rect 25495 3609 25507 3785
rect 24092 3586 24150 3598
rect 21617 3396 21675 3408
rect 17706 3197 17764 3209
rect 24092 3210 24104 3586
rect 24138 3210 24150 3586
rect 24092 3198 24150 3210
rect 24210 3586 24268 3598
rect 24210 3210 24222 3586
rect 24256 3210 24268 3586
rect 24210 3198 24268 3210
rect 24328 3586 24386 3598
rect 24328 3210 24340 3586
rect 24374 3210 24386 3586
rect 24445 3586 24503 3598
rect 24445 3410 24457 3586
rect 24491 3410 24503 3586
rect 24445 3398 24503 3410
rect 24563 3586 24621 3598
rect 25449 3597 25507 3609
rect 25567 3785 25625 3797
rect 25567 3609 25579 3785
rect 25613 3609 25625 3785
rect 25567 3597 25625 3609
rect 25869 3785 25927 3797
rect 24563 3410 24575 3586
rect 24609 3410 24621 3586
rect 24563 3398 24621 3410
rect 25869 3409 25881 3785
rect 25915 3409 25927 3785
rect 25869 3397 25927 3409
rect 25987 3785 26045 3797
rect 25987 3409 25999 3785
rect 26033 3409 26045 3785
rect 25987 3397 26045 3409
rect 26105 3785 26163 3797
rect 26105 3409 26117 3785
rect 26151 3409 26163 3785
rect 26105 3397 26163 3409
rect 26223 3785 26281 3797
rect 26223 3409 26235 3785
rect 26269 3409 26281 3785
rect 26223 3397 26281 3409
rect 26341 3785 26399 3797
rect 26341 3409 26353 3785
rect 26387 3409 26399 3785
rect 26747 3785 26805 3797
rect 26747 3609 26759 3785
rect 26793 3609 26805 3785
rect 26747 3597 26805 3609
rect 26865 3785 26923 3797
rect 26865 3609 26877 3785
rect 26911 3609 26923 3785
rect 26865 3597 26923 3609
rect 27347 3785 27405 3797
rect 27347 3609 27359 3785
rect 27393 3609 27405 3785
rect 27347 3597 27405 3609
rect 27465 3785 27523 3797
rect 27465 3609 27477 3785
rect 27511 3609 27523 3785
rect 27465 3597 27523 3609
rect 27767 3785 27825 3797
rect 26341 3397 26399 3409
rect 27767 3409 27779 3785
rect 27813 3409 27825 3785
rect 27767 3397 27825 3409
rect 27885 3785 27943 3797
rect 27885 3409 27897 3785
rect 27931 3409 27943 3785
rect 27885 3397 27943 3409
rect 28003 3785 28061 3797
rect 28003 3409 28015 3785
rect 28049 3409 28061 3785
rect 28003 3397 28061 3409
rect 28121 3785 28179 3797
rect 28121 3409 28133 3785
rect 28167 3409 28179 3785
rect 28121 3397 28179 3409
rect 28239 3785 28297 3797
rect 28239 3409 28251 3785
rect 28285 3409 28297 3785
rect 28645 3785 28703 3797
rect 28645 3609 28657 3785
rect 28691 3609 28703 3785
rect 28645 3597 28703 3609
rect 28763 3785 28821 3797
rect 28763 3609 28775 3785
rect 28809 3609 28821 3785
rect 29956 3670 29968 4046
rect 30002 3670 30014 4046
rect 29956 3658 30014 3670
rect 30074 4046 30132 4058
rect 30074 3670 30086 4046
rect 30120 3670 30132 4046
rect 30074 3658 30132 3670
rect 30192 4046 30250 4058
rect 30192 3670 30204 4046
rect 30238 3670 30250 4046
rect 30309 4046 30367 4058
rect 30309 3870 30321 4046
rect 30355 3870 30367 4046
rect 30309 3858 30367 3870
rect 30427 4046 30485 4058
rect 30427 3870 30439 4046
rect 30473 3870 30485 4046
rect 30427 3858 30485 3870
rect 38084 4556 38284 4568
rect 38084 4522 38096 4556
rect 38272 4522 38284 4556
rect 38084 4510 38284 4522
rect 30192 3658 30250 3670
rect 28763 3597 28821 3609
rect 28239 3397 28297 3409
rect 24328 3198 24386 3210
rect -2381 2899 -1981 2911
rect -2381 2827 -1981 2839
rect -2381 2793 -2369 2827
rect -1993 2793 -1981 2827
rect -2381 2781 -1981 2793
rect -2381 2421 -2181 2433
rect -2381 2387 -2369 2421
rect -2193 2387 -2181 2421
rect -2381 2375 -2181 2387
rect -2381 2303 -2181 2315
rect -2381 2269 -2369 2303
rect -2193 2269 -2181 2303
rect -2381 2257 -2181 2269
rect 8072 2157 8130 2169
rect 8072 1781 8084 2157
rect 8118 1781 8130 2157
rect 8072 1769 8130 1781
rect 8190 2157 8248 2169
rect 8190 1781 8202 2157
rect 8236 1781 8248 2157
rect 8190 1769 8248 1781
rect 8308 2157 8366 2169
rect 8308 1781 8320 2157
rect 8354 1781 8366 2157
rect 14626 2162 14684 2174
rect 8308 1769 8366 1781
rect 8425 1957 8483 1969
rect 8425 1781 8437 1957
rect 8471 1781 8483 1957
rect 8425 1769 8483 1781
rect 8543 1957 8601 1969
rect 8543 1781 8555 1957
rect 8589 1781 8601 1957
rect 8543 1769 8601 1781
rect 14626 1786 14638 2162
rect 14672 1786 14684 2162
rect 14626 1774 14684 1786
rect 14744 2162 14802 2174
rect 14744 1786 14756 2162
rect 14790 1786 14802 2162
rect 14744 1774 14802 1786
rect 14862 2162 14920 2174
rect 14862 1786 14874 2162
rect 14908 1786 14920 2162
rect 21275 2150 21333 2162
rect 14862 1774 14920 1786
rect 14979 1962 15037 1974
rect 14979 1786 14991 1962
rect 15025 1786 15037 1962
rect 14979 1774 15037 1786
rect 15097 1962 15155 1974
rect 15097 1786 15109 1962
rect 15143 1786 15155 1962
rect 15097 1774 15155 1786
rect 21275 1774 21287 2150
rect 21321 1774 21333 2150
rect -2383 1651 -2183 1663
rect -2383 1617 -2371 1651
rect -2195 1617 -2183 1651
rect -2383 1605 -2183 1617
rect -2383 1533 -2183 1545
rect -2383 1499 -2371 1533
rect -2195 1499 -2183 1533
rect 21275 1762 21333 1774
rect 21393 2150 21451 2162
rect 21393 1774 21405 2150
rect 21439 1774 21451 2150
rect 21393 1762 21451 1774
rect 21511 2150 21569 2162
rect 21511 1774 21523 2150
rect 21557 1774 21569 2150
rect 21511 1762 21569 1774
rect 21628 1950 21686 1962
rect 21628 1774 21640 1950
rect 21674 1774 21686 1950
rect 21628 1762 21686 1774
rect 21746 1950 21804 1962
rect 21746 1774 21758 1950
rect 21792 1774 21804 1950
rect 21746 1762 21804 1774
rect -2383 1487 -2183 1499
rect 33496 2298 33554 2310
rect 33496 1922 33508 2298
rect 33542 1922 33554 2298
rect 33496 1910 33554 1922
rect 33614 2298 33672 2310
rect 33614 1922 33626 2298
rect 33660 1922 33672 2298
rect 33614 1910 33672 1922
rect 33732 2298 33790 2310
rect 33732 1922 33744 2298
rect 33778 1922 33790 2298
rect 33849 2298 33907 2310
rect 33849 2122 33861 2298
rect 33895 2122 33907 2298
rect 33849 2110 33907 2122
rect 33967 2298 34025 2310
rect 33967 2122 33979 2298
rect 34013 2122 34025 2298
rect 33967 2110 34025 2122
rect 38084 2272 38284 2284
rect 38084 2238 38096 2272
rect 38272 2238 38284 2272
rect 38084 2226 38284 2238
rect 38084 2154 38284 2166
rect 38084 2120 38096 2154
rect 38272 2120 38284 2154
rect 38084 2092 38284 2120
rect 38084 2080 38484 2092
rect 38084 2046 38096 2080
rect 38472 2046 38484 2080
rect 38084 2034 38484 2046
rect 33732 1910 33790 1922
rect 38084 1962 38484 1974
rect 38084 1928 38096 1962
rect 38472 1928 38484 1962
rect 38084 1916 38484 1928
rect 38084 1844 38484 1856
rect 38084 1810 38096 1844
rect 38472 1810 38484 1844
rect 38084 1798 38484 1810
rect 38084 1726 38484 1738
rect 38084 1692 38096 1726
rect 38472 1692 38484 1726
rect 38084 1680 38484 1692
rect 31591 1513 31649 1525
rect -2383 1231 -1983 1243
rect -2383 1197 -2371 1231
rect -1995 1197 -1983 1231
rect 31591 1337 31603 1513
rect 31637 1337 31649 1513
rect 31591 1325 31649 1337
rect 31709 1513 31767 1525
rect 31709 1337 31721 1513
rect 31755 1337 31767 1513
rect 31709 1325 31767 1337
rect 32011 1513 32069 1525
rect 29963 1201 30021 1213
rect -2383 1185 -1983 1197
rect -2383 1113 -1983 1125
rect -2383 1079 -2371 1113
rect -1995 1079 -1983 1113
rect -2383 1067 -1983 1079
rect -2383 995 -1983 1007
rect -2383 961 -2371 995
rect -1995 961 -1983 995
rect -2383 949 -1983 961
rect -2383 877 -1983 889
rect -2383 843 -2371 877
rect -1995 843 -1983 877
rect -2383 831 -1983 843
rect 29963 825 29975 1201
rect 30009 825 30021 1201
rect 29963 813 30021 825
rect 30081 1201 30139 1213
rect 30081 825 30093 1201
rect 30127 825 30139 1201
rect 30081 813 30139 825
rect 30199 1201 30257 1213
rect 30199 825 30211 1201
rect 30245 825 30257 1201
rect 30316 1201 30374 1213
rect 30316 1025 30328 1201
rect 30362 1025 30374 1201
rect 30316 1013 30374 1025
rect 30434 1201 30492 1213
rect 30434 1025 30446 1201
rect 30480 1025 30492 1201
rect 32011 1137 32023 1513
rect 32057 1137 32069 1513
rect 32011 1125 32069 1137
rect 32129 1513 32187 1525
rect 32129 1137 32141 1513
rect 32175 1137 32187 1513
rect 32129 1125 32187 1137
rect 32247 1513 32305 1525
rect 32247 1137 32259 1513
rect 32293 1137 32305 1513
rect 32247 1125 32305 1137
rect 32365 1513 32423 1525
rect 32365 1137 32377 1513
rect 32411 1137 32423 1513
rect 32365 1125 32423 1137
rect 32483 1513 32541 1525
rect 32483 1137 32495 1513
rect 32529 1137 32541 1513
rect 32889 1513 32947 1525
rect 32889 1337 32901 1513
rect 32935 1337 32947 1513
rect 32889 1325 32947 1337
rect 33007 1513 33065 1525
rect 33007 1337 33019 1513
rect 33053 1337 33065 1513
rect 33007 1325 33065 1337
rect 32483 1125 32541 1137
rect 38084 1608 38484 1620
rect 38084 1574 38096 1608
rect 38472 1574 38484 1608
rect 38084 1562 38484 1574
rect 38084 1530 38284 1562
rect 38084 1496 38096 1530
rect 38272 1496 38284 1530
rect 38084 1484 38284 1496
rect 30434 1013 30492 1025
rect 30199 813 30257 825
rect -2383 759 -1983 771
rect -2383 725 -2371 759
rect -1995 725 -1983 759
rect -2383 713 -1983 725
rect 38084 1412 38284 1424
rect 38084 1378 38096 1412
rect 38272 1378 38284 1412
rect 38084 1366 38284 1378
rect -2383 353 -2183 365
rect -2383 319 -2371 353
rect -2195 319 -2183 353
rect -2383 307 -2183 319
rect -2383 235 -2183 247
rect -2383 201 -2371 235
rect -2195 201 -2183 235
rect -2383 189 -2183 201
<< pdiff >>
rect 8155 27680 8213 27692
rect 5830 27608 5888 27620
rect 5830 27432 5842 27608
rect 5876 27432 5888 27608
rect 5830 27420 5888 27432
rect 5948 27608 6006 27620
rect 5948 27432 5960 27608
rect 5994 27432 6006 27608
rect 5948 27420 6006 27432
rect 6066 27608 6124 27620
rect 6066 27432 6078 27608
rect 6112 27432 6124 27608
rect 6066 27420 6124 27432
rect 6184 27608 6242 27620
rect 6184 27432 6196 27608
rect 6230 27432 6242 27608
rect 6184 27420 6242 27432
rect 6302 27608 6360 27620
rect 6302 27432 6314 27608
rect 6348 27432 6360 27608
rect 6302 27420 6360 27432
rect 6420 27608 6478 27620
rect 6420 27432 6432 27608
rect 6466 27432 6478 27608
rect 6420 27420 6478 27432
rect 6538 27608 6596 27620
rect 6538 27432 6550 27608
rect 6584 27432 6596 27608
rect 6538 27420 6596 27432
rect 6656 27608 6714 27620
rect 6656 27432 6668 27608
rect 6702 27432 6714 27608
rect 6656 27420 6714 27432
rect 6774 27608 6832 27620
rect 6774 27432 6786 27608
rect 6820 27432 6832 27608
rect 6774 27420 6832 27432
rect 6892 27608 6950 27620
rect 6892 27432 6904 27608
rect 6938 27432 6950 27608
rect 6892 27420 6950 27432
rect 8155 27304 8167 27680
rect 8201 27304 8213 27680
rect 8155 27292 8213 27304
rect 8273 27680 8331 27692
rect 8273 27304 8285 27680
rect 8319 27304 8331 27680
rect 8273 27292 8331 27304
rect 8391 27680 8449 27692
rect 8391 27304 8403 27680
rect 8437 27304 8449 27680
rect 8391 27292 8449 27304
rect 8509 27680 8567 27692
rect 8509 27304 8521 27680
rect 8555 27304 8567 27680
rect 8509 27292 8567 27304
rect 8627 27680 8685 27692
rect 8627 27304 8639 27680
rect 8673 27304 8685 27680
rect 8627 27292 8685 27304
rect 8745 27680 8803 27692
rect 8745 27304 8757 27680
rect 8791 27304 8803 27680
rect 8745 27292 8803 27304
rect 8863 27680 8921 27692
rect 8863 27304 8875 27680
rect 8909 27304 8921 27680
rect 8863 27292 8921 27304
rect 9297 27684 9355 27696
rect 9297 27308 9309 27684
rect 9343 27308 9355 27684
rect 9297 27296 9355 27308
rect 9415 27684 9473 27696
rect 9415 27308 9427 27684
rect 9461 27308 9473 27684
rect 9415 27296 9473 27308
rect 9533 27684 9591 27696
rect 9533 27308 9545 27684
rect 9579 27308 9591 27684
rect 9533 27296 9591 27308
rect 9651 27684 9709 27696
rect 9651 27308 9663 27684
rect 9697 27308 9709 27684
rect 9651 27296 9709 27308
rect 9769 27684 9827 27696
rect 9769 27308 9781 27684
rect 9815 27308 9827 27684
rect 9769 27296 9827 27308
rect 9887 27684 9945 27696
rect 9887 27308 9899 27684
rect 9933 27308 9945 27684
rect 9887 27296 9945 27308
rect 10005 27684 10063 27696
rect 10005 27308 10017 27684
rect 10051 27308 10063 27684
rect 14668 27677 14726 27689
rect 12343 27605 12401 27617
rect 12343 27429 12355 27605
rect 12389 27429 12401 27605
rect 12343 27417 12401 27429
rect 12461 27605 12519 27617
rect 12461 27429 12473 27605
rect 12507 27429 12519 27605
rect 12461 27417 12519 27429
rect 12579 27605 12637 27617
rect 12579 27429 12591 27605
rect 12625 27429 12637 27605
rect 12579 27417 12637 27429
rect 12697 27605 12755 27617
rect 12697 27429 12709 27605
rect 12743 27429 12755 27605
rect 12697 27417 12755 27429
rect 12815 27605 12873 27617
rect 12815 27429 12827 27605
rect 12861 27429 12873 27605
rect 12815 27417 12873 27429
rect 12933 27605 12991 27617
rect 12933 27429 12945 27605
rect 12979 27429 12991 27605
rect 12933 27417 12991 27429
rect 13051 27605 13109 27617
rect 13051 27429 13063 27605
rect 13097 27429 13109 27605
rect 13051 27417 13109 27429
rect 13169 27605 13227 27617
rect 13169 27429 13181 27605
rect 13215 27429 13227 27605
rect 13169 27417 13227 27429
rect 13287 27605 13345 27617
rect 13287 27429 13299 27605
rect 13333 27429 13345 27605
rect 13287 27417 13345 27429
rect 13405 27605 13463 27617
rect 13405 27429 13417 27605
rect 13451 27429 13463 27605
rect 13405 27417 13463 27429
rect 10005 27296 10063 27308
rect 14668 27301 14680 27677
rect 14714 27301 14726 27677
rect 14668 27289 14726 27301
rect 14786 27677 14844 27689
rect 14786 27301 14798 27677
rect 14832 27301 14844 27677
rect 14786 27289 14844 27301
rect 14904 27677 14962 27689
rect 14904 27301 14916 27677
rect 14950 27301 14962 27677
rect 14904 27289 14962 27301
rect 15022 27677 15080 27689
rect 15022 27301 15034 27677
rect 15068 27301 15080 27677
rect 15022 27289 15080 27301
rect 15140 27677 15198 27689
rect 15140 27301 15152 27677
rect 15186 27301 15198 27677
rect 15140 27289 15198 27301
rect 15258 27677 15316 27689
rect 15258 27301 15270 27677
rect 15304 27301 15316 27677
rect 15258 27289 15316 27301
rect 15376 27677 15434 27689
rect 15376 27301 15388 27677
rect 15422 27301 15434 27677
rect 15376 27289 15434 27301
rect 15810 27681 15868 27693
rect 15810 27305 15822 27681
rect 15856 27305 15868 27681
rect 15810 27293 15868 27305
rect 15928 27681 15986 27693
rect 15928 27305 15940 27681
rect 15974 27305 15986 27681
rect 15928 27293 15986 27305
rect 16046 27681 16104 27693
rect 16046 27305 16058 27681
rect 16092 27305 16104 27681
rect 16046 27293 16104 27305
rect 16164 27681 16222 27693
rect 16164 27305 16176 27681
rect 16210 27305 16222 27681
rect 16164 27293 16222 27305
rect 16282 27681 16340 27693
rect 16282 27305 16294 27681
rect 16328 27305 16340 27681
rect 16282 27293 16340 27305
rect 16400 27681 16458 27693
rect 16400 27305 16412 27681
rect 16446 27305 16458 27681
rect 16400 27293 16458 27305
rect 16518 27681 16576 27693
rect 16518 27305 16530 27681
rect 16564 27305 16576 27681
rect 21202 27672 21260 27684
rect 18877 27600 18935 27612
rect 18877 27424 18889 27600
rect 18923 27424 18935 27600
rect 18877 27412 18935 27424
rect 18995 27600 19053 27612
rect 18995 27424 19007 27600
rect 19041 27424 19053 27600
rect 18995 27412 19053 27424
rect 19113 27600 19171 27612
rect 19113 27424 19125 27600
rect 19159 27424 19171 27600
rect 19113 27412 19171 27424
rect 19231 27600 19289 27612
rect 19231 27424 19243 27600
rect 19277 27424 19289 27600
rect 19231 27412 19289 27424
rect 19349 27600 19407 27612
rect 19349 27424 19361 27600
rect 19395 27424 19407 27600
rect 19349 27412 19407 27424
rect 19467 27600 19525 27612
rect 19467 27424 19479 27600
rect 19513 27424 19525 27600
rect 19467 27412 19525 27424
rect 19585 27600 19643 27612
rect 19585 27424 19597 27600
rect 19631 27424 19643 27600
rect 19585 27412 19643 27424
rect 19703 27600 19761 27612
rect 19703 27424 19715 27600
rect 19749 27424 19761 27600
rect 19703 27412 19761 27424
rect 19821 27600 19879 27612
rect 19821 27424 19833 27600
rect 19867 27424 19879 27600
rect 19821 27412 19879 27424
rect 19939 27600 19997 27612
rect 19939 27424 19951 27600
rect 19985 27424 19997 27600
rect 19939 27412 19997 27424
rect 16518 27293 16576 27305
rect 8584 26897 8642 26909
rect 8584 26721 8596 26897
rect 8630 26721 8642 26897
rect 8584 26709 8642 26721
rect 8702 26897 8760 26909
rect 8702 26721 8714 26897
rect 8748 26721 8760 26897
rect 8702 26709 8760 26721
rect 8820 26897 8878 26909
rect 8820 26721 8832 26897
rect 8866 26721 8878 26897
rect 8820 26709 8878 26721
rect 8938 26897 8996 26909
rect 8938 26721 8950 26897
rect 8984 26721 8996 26897
rect 8938 26709 8996 26721
rect 9726 26901 9784 26913
rect 9726 26725 9738 26901
rect 9772 26725 9784 26901
rect 9726 26713 9784 26725
rect 9844 26901 9902 26913
rect 9844 26725 9856 26901
rect 9890 26725 9902 26901
rect 9844 26713 9902 26725
rect 9962 26901 10020 26913
rect 9962 26725 9974 26901
rect 10008 26725 10020 26901
rect 9962 26713 10020 26725
rect 10080 26901 10138 26913
rect 10080 26725 10092 26901
rect 10126 26725 10138 26901
rect 21202 27296 21214 27672
rect 21248 27296 21260 27672
rect 21202 27284 21260 27296
rect 21320 27672 21378 27684
rect 21320 27296 21332 27672
rect 21366 27296 21378 27672
rect 21320 27284 21378 27296
rect 21438 27672 21496 27684
rect 21438 27296 21450 27672
rect 21484 27296 21496 27672
rect 21438 27284 21496 27296
rect 21556 27672 21614 27684
rect 21556 27296 21568 27672
rect 21602 27296 21614 27672
rect 21556 27284 21614 27296
rect 21674 27672 21732 27684
rect 21674 27296 21686 27672
rect 21720 27296 21732 27672
rect 21674 27284 21732 27296
rect 21792 27672 21850 27684
rect 21792 27296 21804 27672
rect 21838 27296 21850 27672
rect 21792 27284 21850 27296
rect 21910 27672 21968 27684
rect 21910 27296 21922 27672
rect 21956 27296 21968 27672
rect 21910 27284 21968 27296
rect 22344 27676 22402 27688
rect 22344 27300 22356 27676
rect 22390 27300 22402 27676
rect 22344 27288 22402 27300
rect 22462 27676 22520 27688
rect 22462 27300 22474 27676
rect 22508 27300 22520 27676
rect 22462 27288 22520 27300
rect 22580 27676 22638 27688
rect 22580 27300 22592 27676
rect 22626 27300 22638 27676
rect 22580 27288 22638 27300
rect 22698 27676 22756 27688
rect 22698 27300 22710 27676
rect 22744 27300 22756 27676
rect 22698 27288 22756 27300
rect 22816 27676 22874 27688
rect 22816 27300 22828 27676
rect 22862 27300 22874 27676
rect 22816 27288 22874 27300
rect 22934 27676 22992 27688
rect 22934 27300 22946 27676
rect 22980 27300 22992 27676
rect 22934 27288 22992 27300
rect 23052 27676 23110 27688
rect 23052 27300 23064 27676
rect 23098 27300 23110 27676
rect 27760 27676 27818 27688
rect 25435 27604 25493 27616
rect 25435 27428 25447 27604
rect 25481 27428 25493 27604
rect 25435 27416 25493 27428
rect 25553 27604 25611 27616
rect 25553 27428 25565 27604
rect 25599 27428 25611 27604
rect 25553 27416 25611 27428
rect 25671 27604 25729 27616
rect 25671 27428 25683 27604
rect 25717 27428 25729 27604
rect 25671 27416 25729 27428
rect 25789 27604 25847 27616
rect 25789 27428 25801 27604
rect 25835 27428 25847 27604
rect 25789 27416 25847 27428
rect 25907 27604 25965 27616
rect 25907 27428 25919 27604
rect 25953 27428 25965 27604
rect 25907 27416 25965 27428
rect 26025 27604 26083 27616
rect 26025 27428 26037 27604
rect 26071 27428 26083 27604
rect 26025 27416 26083 27428
rect 26143 27604 26201 27616
rect 26143 27428 26155 27604
rect 26189 27428 26201 27604
rect 26143 27416 26201 27428
rect 26261 27604 26319 27616
rect 26261 27428 26273 27604
rect 26307 27428 26319 27604
rect 26261 27416 26319 27428
rect 26379 27604 26437 27616
rect 26379 27428 26391 27604
rect 26425 27428 26437 27604
rect 26379 27416 26437 27428
rect 26497 27604 26555 27616
rect 26497 27428 26509 27604
rect 26543 27428 26555 27604
rect 26497 27416 26555 27428
rect 23052 27288 23110 27300
rect 10080 26713 10138 26725
rect 15097 26894 15155 26906
rect 15097 26718 15109 26894
rect 15143 26718 15155 26894
rect 15097 26706 15155 26718
rect 15215 26894 15273 26906
rect 15215 26718 15227 26894
rect 15261 26718 15273 26894
rect 15215 26706 15273 26718
rect 15333 26894 15391 26906
rect 15333 26718 15345 26894
rect 15379 26718 15391 26894
rect 15333 26706 15391 26718
rect 15451 26894 15509 26906
rect 15451 26718 15463 26894
rect 15497 26718 15509 26894
rect 15451 26706 15509 26718
rect 16239 26898 16297 26910
rect 16239 26722 16251 26898
rect 16285 26722 16297 26898
rect 16239 26710 16297 26722
rect 16357 26898 16415 26910
rect 16357 26722 16369 26898
rect 16403 26722 16415 26898
rect 16357 26710 16415 26722
rect 16475 26898 16533 26910
rect 16475 26722 16487 26898
rect 16521 26722 16533 26898
rect 16475 26710 16533 26722
rect 16593 26898 16651 26910
rect 16593 26722 16605 26898
rect 16639 26722 16651 26898
rect 27760 27300 27772 27676
rect 27806 27300 27818 27676
rect 27760 27288 27818 27300
rect 27878 27676 27936 27688
rect 27878 27300 27890 27676
rect 27924 27300 27936 27676
rect 27878 27288 27936 27300
rect 27996 27676 28054 27688
rect 27996 27300 28008 27676
rect 28042 27300 28054 27676
rect 27996 27288 28054 27300
rect 28114 27676 28172 27688
rect 28114 27300 28126 27676
rect 28160 27300 28172 27676
rect 28114 27288 28172 27300
rect 28232 27676 28290 27688
rect 28232 27300 28244 27676
rect 28278 27300 28290 27676
rect 28232 27288 28290 27300
rect 28350 27676 28408 27688
rect 28350 27300 28362 27676
rect 28396 27300 28408 27676
rect 28350 27288 28408 27300
rect 28468 27676 28526 27688
rect 28468 27300 28480 27676
rect 28514 27300 28526 27676
rect 28468 27288 28526 27300
rect 28902 27680 28960 27692
rect 28902 27304 28914 27680
rect 28948 27304 28960 27680
rect 28902 27292 28960 27304
rect 29020 27680 29078 27692
rect 29020 27304 29032 27680
rect 29066 27304 29078 27680
rect 29020 27292 29078 27304
rect 29138 27680 29196 27692
rect 29138 27304 29150 27680
rect 29184 27304 29196 27680
rect 29138 27292 29196 27304
rect 29256 27680 29314 27692
rect 29256 27304 29268 27680
rect 29302 27304 29314 27680
rect 29256 27292 29314 27304
rect 29374 27680 29432 27692
rect 29374 27304 29386 27680
rect 29420 27304 29432 27680
rect 29374 27292 29432 27304
rect 29492 27680 29550 27692
rect 29492 27304 29504 27680
rect 29538 27304 29550 27680
rect 29492 27292 29550 27304
rect 29610 27680 29668 27692
rect 29610 27304 29622 27680
rect 29656 27304 29668 27680
rect 29610 27292 29668 27304
rect 16593 26710 16651 26722
rect 21631 26889 21689 26901
rect 21631 26713 21643 26889
rect 21677 26713 21689 26889
rect 21631 26701 21689 26713
rect 21749 26889 21807 26901
rect 21749 26713 21761 26889
rect 21795 26713 21807 26889
rect 21749 26701 21807 26713
rect 21867 26889 21925 26901
rect 21867 26713 21879 26889
rect 21913 26713 21925 26889
rect 21867 26701 21925 26713
rect 21985 26889 22043 26901
rect 21985 26713 21997 26889
rect 22031 26713 22043 26889
rect 21985 26701 22043 26713
rect 22773 26893 22831 26905
rect 22773 26717 22785 26893
rect 22819 26717 22831 26893
rect 22773 26705 22831 26717
rect 22891 26893 22949 26905
rect 22891 26717 22903 26893
rect 22937 26717 22949 26893
rect 22891 26705 22949 26717
rect 23009 26893 23067 26905
rect 23009 26717 23021 26893
rect 23055 26717 23067 26893
rect 23009 26705 23067 26717
rect 23127 26893 23185 26905
rect 23127 26717 23139 26893
rect 23173 26717 23185 26893
rect 23127 26705 23185 26717
rect 28189 26893 28247 26905
rect 28189 26717 28201 26893
rect 28235 26717 28247 26893
rect 28189 26705 28247 26717
rect 28307 26893 28365 26905
rect 28307 26717 28319 26893
rect 28353 26717 28365 26893
rect 28307 26705 28365 26717
rect 28425 26893 28483 26905
rect 28425 26717 28437 26893
rect 28471 26717 28483 26893
rect 28425 26705 28483 26717
rect 28543 26893 28601 26905
rect 28543 26717 28555 26893
rect 28589 26717 28601 26893
rect 28543 26705 28601 26717
rect 29331 26897 29389 26909
rect 29331 26721 29343 26897
rect 29377 26721 29389 26897
rect 29331 26709 29389 26721
rect 29449 26897 29507 26909
rect 29449 26721 29461 26897
rect 29495 26721 29507 26897
rect 29449 26709 29507 26721
rect 29567 26897 29625 26909
rect 29567 26721 29579 26897
rect 29613 26721 29625 26897
rect 29567 26709 29625 26721
rect 29685 26897 29743 26909
rect 29685 26721 29697 26897
rect 29731 26721 29743 26897
rect 29685 26709 29743 26721
rect 5844 25958 5902 25970
rect 5844 25782 5856 25958
rect 5890 25782 5902 25958
rect 5844 25770 5902 25782
rect 5962 25958 6020 25970
rect 5962 25782 5974 25958
rect 6008 25782 6020 25958
rect 5962 25770 6020 25782
rect 6080 25958 6138 25970
rect 6080 25782 6092 25958
rect 6126 25782 6138 25958
rect 6080 25770 6138 25782
rect 6198 25958 6256 25970
rect 6198 25782 6210 25958
rect 6244 25782 6256 25958
rect 6198 25770 6256 25782
rect 6316 25958 6374 25970
rect 6316 25782 6328 25958
rect 6362 25782 6374 25958
rect 6316 25770 6374 25782
rect 6434 25958 6492 25970
rect 6434 25782 6446 25958
rect 6480 25782 6492 25958
rect 6434 25770 6492 25782
rect 6552 25958 6610 25970
rect 6552 25782 6564 25958
rect 6598 25782 6610 25958
rect 6552 25770 6610 25782
rect 6670 25958 6728 25970
rect 6670 25782 6682 25958
rect 6716 25782 6728 25958
rect 6670 25770 6728 25782
rect 6788 25958 6846 25970
rect 6788 25782 6800 25958
rect 6834 25782 6846 25958
rect 6788 25770 6846 25782
rect 6906 25958 6964 25970
rect 6906 25782 6918 25958
rect 6952 25782 6964 25958
rect 12357 25955 12415 25967
rect 6906 25770 6964 25782
rect 12357 25779 12369 25955
rect 12403 25779 12415 25955
rect 12357 25767 12415 25779
rect 12475 25955 12533 25967
rect 12475 25779 12487 25955
rect 12521 25779 12533 25955
rect 12475 25767 12533 25779
rect 12593 25955 12651 25967
rect 12593 25779 12605 25955
rect 12639 25779 12651 25955
rect 12593 25767 12651 25779
rect 12711 25955 12769 25967
rect 12711 25779 12723 25955
rect 12757 25779 12769 25955
rect 12711 25767 12769 25779
rect 12829 25955 12887 25967
rect 12829 25779 12841 25955
rect 12875 25779 12887 25955
rect 12829 25767 12887 25779
rect 12947 25955 13005 25967
rect 12947 25779 12959 25955
rect 12993 25779 13005 25955
rect 12947 25767 13005 25779
rect 13065 25955 13123 25967
rect 13065 25779 13077 25955
rect 13111 25779 13123 25955
rect 13065 25767 13123 25779
rect 13183 25955 13241 25967
rect 13183 25779 13195 25955
rect 13229 25779 13241 25955
rect 13183 25767 13241 25779
rect 13301 25955 13359 25967
rect 13301 25779 13313 25955
rect 13347 25779 13359 25955
rect 13301 25767 13359 25779
rect 13419 25955 13477 25967
rect 13419 25779 13431 25955
rect 13465 25779 13477 25955
rect 18891 25950 18949 25962
rect 13419 25767 13477 25779
rect 18891 25774 18903 25950
rect 18937 25774 18949 25950
rect 7792 25541 7850 25553
rect 7308 25341 7366 25353
rect 7308 25165 7320 25341
rect 7354 25165 7366 25341
rect 7308 25153 7366 25165
rect 7426 25341 7484 25353
rect 7426 25165 7438 25341
rect 7472 25165 7484 25341
rect 7426 25153 7484 25165
rect 7544 25341 7602 25353
rect 7544 25165 7556 25341
rect 7590 25165 7602 25341
rect 7544 25153 7602 25165
rect 7662 25341 7720 25353
rect 7662 25165 7674 25341
rect 7708 25165 7720 25341
rect 7662 25153 7720 25165
rect 7792 25165 7804 25541
rect 7838 25165 7850 25541
rect 7792 25153 7850 25165
rect 7910 25541 7968 25553
rect 7910 25165 7922 25541
rect 7956 25165 7968 25541
rect 7910 25153 7968 25165
rect 8028 25541 8086 25553
rect 8028 25165 8040 25541
rect 8074 25165 8086 25541
rect 8028 25153 8086 25165
rect 8146 25541 8204 25553
rect 8146 25165 8158 25541
rect 8192 25165 8204 25541
rect 8146 25153 8204 25165
rect 8264 25541 8322 25553
rect 8264 25165 8276 25541
rect 8310 25165 8322 25541
rect 8264 25153 8322 25165
rect 8382 25541 8440 25553
rect 8382 25165 8394 25541
rect 8428 25165 8440 25541
rect 8382 25153 8440 25165
rect 8500 25541 8558 25553
rect 8500 25165 8512 25541
rect 8546 25165 8558 25541
rect 9690 25541 9748 25553
rect 8500 25153 8558 25165
rect 8629 25341 8687 25353
rect 8629 25165 8641 25341
rect 8675 25165 8687 25341
rect 8629 25153 8687 25165
rect 8747 25341 8805 25353
rect 8747 25165 8759 25341
rect 8793 25165 8805 25341
rect 8747 25153 8805 25165
rect 8865 25341 8923 25353
rect 8865 25165 8877 25341
rect 8911 25165 8923 25341
rect 8865 25153 8923 25165
rect 8983 25341 9041 25353
rect 8983 25165 8995 25341
rect 9029 25165 9041 25341
rect 8983 25153 9041 25165
rect 9206 25341 9264 25353
rect 9206 25165 9218 25341
rect 9252 25165 9264 25341
rect 9206 25153 9264 25165
rect 9324 25341 9382 25353
rect 9324 25165 9336 25341
rect 9370 25165 9382 25341
rect 9324 25153 9382 25165
rect 9442 25341 9500 25353
rect 9442 25165 9454 25341
rect 9488 25165 9500 25341
rect 9442 25153 9500 25165
rect 9560 25341 9618 25353
rect 9560 25165 9572 25341
rect 9606 25165 9618 25341
rect 9560 25153 9618 25165
rect 9690 25165 9702 25541
rect 9736 25165 9748 25541
rect 9690 25153 9748 25165
rect 9808 25541 9866 25553
rect 9808 25165 9820 25541
rect 9854 25165 9866 25541
rect 9808 25153 9866 25165
rect 9926 25541 9984 25553
rect 9926 25165 9938 25541
rect 9972 25165 9984 25541
rect 9926 25153 9984 25165
rect 10044 25541 10102 25553
rect 10044 25165 10056 25541
rect 10090 25165 10102 25541
rect 10044 25153 10102 25165
rect 10162 25541 10220 25553
rect 10162 25165 10174 25541
rect 10208 25165 10220 25541
rect 10162 25153 10220 25165
rect 10280 25541 10338 25553
rect 10280 25165 10292 25541
rect 10326 25165 10338 25541
rect 10280 25153 10338 25165
rect 10398 25541 10456 25553
rect 10398 25165 10410 25541
rect 10444 25165 10456 25541
rect 18891 25762 18949 25774
rect 19009 25950 19067 25962
rect 19009 25774 19021 25950
rect 19055 25774 19067 25950
rect 19009 25762 19067 25774
rect 19127 25950 19185 25962
rect 19127 25774 19139 25950
rect 19173 25774 19185 25950
rect 19127 25762 19185 25774
rect 19245 25950 19303 25962
rect 19245 25774 19257 25950
rect 19291 25774 19303 25950
rect 19245 25762 19303 25774
rect 19363 25950 19421 25962
rect 19363 25774 19375 25950
rect 19409 25774 19421 25950
rect 19363 25762 19421 25774
rect 19481 25950 19539 25962
rect 19481 25774 19493 25950
rect 19527 25774 19539 25950
rect 19481 25762 19539 25774
rect 19599 25950 19657 25962
rect 19599 25774 19611 25950
rect 19645 25774 19657 25950
rect 19599 25762 19657 25774
rect 19717 25950 19775 25962
rect 19717 25774 19729 25950
rect 19763 25774 19775 25950
rect 19717 25762 19775 25774
rect 19835 25950 19893 25962
rect 19835 25774 19847 25950
rect 19881 25774 19893 25950
rect 19835 25762 19893 25774
rect 19953 25950 20011 25962
rect 19953 25774 19965 25950
rect 19999 25774 20011 25950
rect 25449 25954 25507 25966
rect 19953 25762 20011 25774
rect 25449 25778 25461 25954
rect 25495 25778 25507 25954
rect 25449 25766 25507 25778
rect 25567 25954 25625 25966
rect 25567 25778 25579 25954
rect 25613 25778 25625 25954
rect 25567 25766 25625 25778
rect 25685 25954 25743 25966
rect 25685 25778 25697 25954
rect 25731 25778 25743 25954
rect 25685 25766 25743 25778
rect 25803 25954 25861 25966
rect 25803 25778 25815 25954
rect 25849 25778 25861 25954
rect 25803 25766 25861 25778
rect 25921 25954 25979 25966
rect 25921 25778 25933 25954
rect 25967 25778 25979 25954
rect 25921 25766 25979 25778
rect 26039 25954 26097 25966
rect 26039 25778 26051 25954
rect 26085 25778 26097 25954
rect 26039 25766 26097 25778
rect 26157 25954 26215 25966
rect 26157 25778 26169 25954
rect 26203 25778 26215 25954
rect 26157 25766 26215 25778
rect 26275 25954 26333 25966
rect 26275 25778 26287 25954
rect 26321 25778 26333 25954
rect 26275 25766 26333 25778
rect 26393 25954 26451 25966
rect 26393 25778 26405 25954
rect 26439 25778 26451 25954
rect 26393 25766 26451 25778
rect 26511 25954 26569 25966
rect 26511 25778 26523 25954
rect 26557 25778 26569 25954
rect 26511 25766 26569 25778
rect 14305 25538 14363 25550
rect 10398 25153 10456 25165
rect 10527 25341 10585 25353
rect 10527 25165 10539 25341
rect 10573 25165 10585 25341
rect 10527 25153 10585 25165
rect 10645 25341 10703 25353
rect 10645 25165 10657 25341
rect 10691 25165 10703 25341
rect 10645 25153 10703 25165
rect 10763 25341 10821 25353
rect 10763 25165 10775 25341
rect 10809 25165 10821 25341
rect 10763 25153 10821 25165
rect 10881 25341 10939 25353
rect 10881 25165 10893 25341
rect 10927 25165 10939 25341
rect 10881 25153 10939 25165
rect 5839 24354 5897 24366
rect 5839 24178 5851 24354
rect 5885 24178 5897 24354
rect 5839 24166 5897 24178
rect 5957 24354 6015 24366
rect 5957 24178 5969 24354
rect 6003 24178 6015 24354
rect 5957 24166 6015 24178
rect 6075 24354 6133 24366
rect 6075 24178 6087 24354
rect 6121 24178 6133 24354
rect 6075 24166 6133 24178
rect 6193 24354 6251 24366
rect 6193 24178 6205 24354
rect 6239 24178 6251 24354
rect 6193 24166 6251 24178
rect 6311 24354 6369 24366
rect 6311 24178 6323 24354
rect 6357 24178 6369 24354
rect 6311 24166 6369 24178
rect 6429 24354 6487 24366
rect 6429 24178 6441 24354
rect 6475 24178 6487 24354
rect 6429 24166 6487 24178
rect 6547 24354 6605 24366
rect 6547 24178 6559 24354
rect 6593 24178 6605 24354
rect 6547 24166 6605 24178
rect 6665 24354 6723 24366
rect 6665 24178 6677 24354
rect 6711 24178 6723 24354
rect 6665 24166 6723 24178
rect 6783 24354 6841 24366
rect 6783 24178 6795 24354
rect 6829 24178 6841 24354
rect 6783 24166 6841 24178
rect 6901 24354 6959 24366
rect 6901 24178 6913 24354
rect 6947 24178 6959 24354
rect 6901 24166 6959 24178
rect 7735 24848 7793 24860
rect 7735 24472 7747 24848
rect 7781 24472 7793 24848
rect 7735 24460 7793 24472
rect 7853 24848 7911 24860
rect 7853 24472 7865 24848
rect 7899 24472 7911 24848
rect 7853 24460 7911 24472
rect 7971 24848 8029 24860
rect 7971 24472 7983 24848
rect 8017 24472 8029 24848
rect 7971 24460 8029 24472
rect 8089 24848 8147 24860
rect 8089 24472 8101 24848
rect 8135 24472 8147 24848
rect 8089 24460 8147 24472
rect 8207 24848 8265 24860
rect 8207 24472 8219 24848
rect 8253 24472 8265 24848
rect 8207 24460 8265 24472
rect 8325 24848 8383 24860
rect 8325 24472 8337 24848
rect 8371 24472 8383 24848
rect 8325 24460 8383 24472
rect 8443 24848 8501 24860
rect 8443 24472 8455 24848
rect 8489 24472 8501 24848
rect 8443 24460 8501 24472
rect 13821 25338 13879 25350
rect 13821 25162 13833 25338
rect 13867 25162 13879 25338
rect 13821 25150 13879 25162
rect 13939 25338 13997 25350
rect 13939 25162 13951 25338
rect 13985 25162 13997 25338
rect 13939 25150 13997 25162
rect 14057 25338 14115 25350
rect 14057 25162 14069 25338
rect 14103 25162 14115 25338
rect 14057 25150 14115 25162
rect 14175 25338 14233 25350
rect 14175 25162 14187 25338
rect 14221 25162 14233 25338
rect 14175 25150 14233 25162
rect 14305 25162 14317 25538
rect 14351 25162 14363 25538
rect 14305 25150 14363 25162
rect 14423 25538 14481 25550
rect 14423 25162 14435 25538
rect 14469 25162 14481 25538
rect 14423 25150 14481 25162
rect 14541 25538 14599 25550
rect 14541 25162 14553 25538
rect 14587 25162 14599 25538
rect 14541 25150 14599 25162
rect 14659 25538 14717 25550
rect 14659 25162 14671 25538
rect 14705 25162 14717 25538
rect 14659 25150 14717 25162
rect 14777 25538 14835 25550
rect 14777 25162 14789 25538
rect 14823 25162 14835 25538
rect 14777 25150 14835 25162
rect 14895 25538 14953 25550
rect 14895 25162 14907 25538
rect 14941 25162 14953 25538
rect 14895 25150 14953 25162
rect 15013 25538 15071 25550
rect 15013 25162 15025 25538
rect 15059 25162 15071 25538
rect 16203 25538 16261 25550
rect 15013 25150 15071 25162
rect 15142 25338 15200 25350
rect 15142 25162 15154 25338
rect 15188 25162 15200 25338
rect 15142 25150 15200 25162
rect 15260 25338 15318 25350
rect 15260 25162 15272 25338
rect 15306 25162 15318 25338
rect 15260 25150 15318 25162
rect 15378 25338 15436 25350
rect 15378 25162 15390 25338
rect 15424 25162 15436 25338
rect 15378 25150 15436 25162
rect 15496 25338 15554 25350
rect 15496 25162 15508 25338
rect 15542 25162 15554 25338
rect 15496 25150 15554 25162
rect 15719 25338 15777 25350
rect 15719 25162 15731 25338
rect 15765 25162 15777 25338
rect 15719 25150 15777 25162
rect 15837 25338 15895 25350
rect 15837 25162 15849 25338
rect 15883 25162 15895 25338
rect 15837 25150 15895 25162
rect 15955 25338 16013 25350
rect 15955 25162 15967 25338
rect 16001 25162 16013 25338
rect 15955 25150 16013 25162
rect 16073 25338 16131 25350
rect 16073 25162 16085 25338
rect 16119 25162 16131 25338
rect 16073 25150 16131 25162
rect 16203 25162 16215 25538
rect 16249 25162 16261 25538
rect 16203 25150 16261 25162
rect 16321 25538 16379 25550
rect 16321 25162 16333 25538
rect 16367 25162 16379 25538
rect 16321 25150 16379 25162
rect 16439 25538 16497 25550
rect 16439 25162 16451 25538
rect 16485 25162 16497 25538
rect 16439 25150 16497 25162
rect 16557 25538 16615 25550
rect 16557 25162 16569 25538
rect 16603 25162 16615 25538
rect 16557 25150 16615 25162
rect 16675 25538 16733 25550
rect 16675 25162 16687 25538
rect 16721 25162 16733 25538
rect 16675 25150 16733 25162
rect 16793 25538 16851 25550
rect 16793 25162 16805 25538
rect 16839 25162 16851 25538
rect 16793 25150 16851 25162
rect 16911 25538 16969 25550
rect 16911 25162 16923 25538
rect 16957 25162 16969 25538
rect 20839 25533 20897 25545
rect 16911 25150 16969 25162
rect 17040 25338 17098 25350
rect 17040 25162 17052 25338
rect 17086 25162 17098 25338
rect 17040 25150 17098 25162
rect 17158 25338 17216 25350
rect 17158 25162 17170 25338
rect 17204 25162 17216 25338
rect 17158 25150 17216 25162
rect 17276 25338 17334 25350
rect 17276 25162 17288 25338
rect 17322 25162 17334 25338
rect 17276 25150 17334 25162
rect 17394 25338 17452 25350
rect 17394 25162 17406 25338
rect 17440 25162 17452 25338
rect 17394 25150 17452 25162
rect 9633 24848 9691 24860
rect 9633 24472 9645 24848
rect 9679 24472 9691 24848
rect 9633 24460 9691 24472
rect 9751 24848 9809 24860
rect 9751 24472 9763 24848
rect 9797 24472 9809 24848
rect 9751 24460 9809 24472
rect 9869 24848 9927 24860
rect 9869 24472 9881 24848
rect 9915 24472 9927 24848
rect 9869 24460 9927 24472
rect 9987 24848 10045 24860
rect 9987 24472 9999 24848
rect 10033 24472 10045 24848
rect 9987 24460 10045 24472
rect 10105 24848 10163 24860
rect 10105 24472 10117 24848
rect 10151 24472 10163 24848
rect 10105 24460 10163 24472
rect 10223 24848 10281 24860
rect 10223 24472 10235 24848
rect 10269 24472 10281 24848
rect 10223 24460 10281 24472
rect 10341 24848 10399 24860
rect 10341 24472 10353 24848
rect 10387 24472 10399 24848
rect 10341 24460 10399 24472
rect 12352 24351 12410 24363
rect 12352 24175 12364 24351
rect 12398 24175 12410 24351
rect 12352 24163 12410 24175
rect 12470 24351 12528 24363
rect 12470 24175 12482 24351
rect 12516 24175 12528 24351
rect 12470 24163 12528 24175
rect 12588 24351 12646 24363
rect 12588 24175 12600 24351
rect 12634 24175 12646 24351
rect 12588 24163 12646 24175
rect 12706 24351 12764 24363
rect 12706 24175 12718 24351
rect 12752 24175 12764 24351
rect 12706 24163 12764 24175
rect 12824 24351 12882 24363
rect 12824 24175 12836 24351
rect 12870 24175 12882 24351
rect 12824 24163 12882 24175
rect 12942 24351 13000 24363
rect 12942 24175 12954 24351
rect 12988 24175 13000 24351
rect 12942 24163 13000 24175
rect 13060 24351 13118 24363
rect 13060 24175 13072 24351
rect 13106 24175 13118 24351
rect 13060 24163 13118 24175
rect 13178 24351 13236 24363
rect 13178 24175 13190 24351
rect 13224 24175 13236 24351
rect 13178 24163 13236 24175
rect 13296 24351 13354 24363
rect 13296 24175 13308 24351
rect 13342 24175 13354 24351
rect 13296 24163 13354 24175
rect 13414 24351 13472 24363
rect 13414 24175 13426 24351
rect 13460 24175 13472 24351
rect 13414 24163 13472 24175
rect 14248 24845 14306 24857
rect 14248 24469 14260 24845
rect 14294 24469 14306 24845
rect 14248 24457 14306 24469
rect 14366 24845 14424 24857
rect 14366 24469 14378 24845
rect 14412 24469 14424 24845
rect 14366 24457 14424 24469
rect 14484 24845 14542 24857
rect 14484 24469 14496 24845
rect 14530 24469 14542 24845
rect 14484 24457 14542 24469
rect 14602 24845 14660 24857
rect 14602 24469 14614 24845
rect 14648 24469 14660 24845
rect 14602 24457 14660 24469
rect 14720 24845 14778 24857
rect 14720 24469 14732 24845
rect 14766 24469 14778 24845
rect 14720 24457 14778 24469
rect 14838 24845 14896 24857
rect 14838 24469 14850 24845
rect 14884 24469 14896 24845
rect 14838 24457 14896 24469
rect 14956 24845 15014 24857
rect 14956 24469 14968 24845
rect 15002 24469 15014 24845
rect 14956 24457 15014 24469
rect 20355 25333 20413 25345
rect 20355 25157 20367 25333
rect 20401 25157 20413 25333
rect 20355 25145 20413 25157
rect 20473 25333 20531 25345
rect 20473 25157 20485 25333
rect 20519 25157 20531 25333
rect 20473 25145 20531 25157
rect 20591 25333 20649 25345
rect 20591 25157 20603 25333
rect 20637 25157 20649 25333
rect 20591 25145 20649 25157
rect 20709 25333 20767 25345
rect 20709 25157 20721 25333
rect 20755 25157 20767 25333
rect 20709 25145 20767 25157
rect 20839 25157 20851 25533
rect 20885 25157 20897 25533
rect 20839 25145 20897 25157
rect 20957 25533 21015 25545
rect 20957 25157 20969 25533
rect 21003 25157 21015 25533
rect 20957 25145 21015 25157
rect 21075 25533 21133 25545
rect 21075 25157 21087 25533
rect 21121 25157 21133 25533
rect 21075 25145 21133 25157
rect 21193 25533 21251 25545
rect 21193 25157 21205 25533
rect 21239 25157 21251 25533
rect 21193 25145 21251 25157
rect 21311 25533 21369 25545
rect 21311 25157 21323 25533
rect 21357 25157 21369 25533
rect 21311 25145 21369 25157
rect 21429 25533 21487 25545
rect 21429 25157 21441 25533
rect 21475 25157 21487 25533
rect 21429 25145 21487 25157
rect 21547 25533 21605 25545
rect 21547 25157 21559 25533
rect 21593 25157 21605 25533
rect 22737 25533 22795 25545
rect 21547 25145 21605 25157
rect 21676 25333 21734 25345
rect 21676 25157 21688 25333
rect 21722 25157 21734 25333
rect 21676 25145 21734 25157
rect 21794 25333 21852 25345
rect 21794 25157 21806 25333
rect 21840 25157 21852 25333
rect 21794 25145 21852 25157
rect 21912 25333 21970 25345
rect 21912 25157 21924 25333
rect 21958 25157 21970 25333
rect 21912 25145 21970 25157
rect 22030 25333 22088 25345
rect 22030 25157 22042 25333
rect 22076 25157 22088 25333
rect 22030 25145 22088 25157
rect 22253 25333 22311 25345
rect 22253 25157 22265 25333
rect 22299 25157 22311 25333
rect 22253 25145 22311 25157
rect 22371 25333 22429 25345
rect 22371 25157 22383 25333
rect 22417 25157 22429 25333
rect 22371 25145 22429 25157
rect 22489 25333 22547 25345
rect 22489 25157 22501 25333
rect 22535 25157 22547 25333
rect 22489 25145 22547 25157
rect 22607 25333 22665 25345
rect 22607 25157 22619 25333
rect 22653 25157 22665 25333
rect 22607 25145 22665 25157
rect 22737 25157 22749 25533
rect 22783 25157 22795 25533
rect 22737 25145 22795 25157
rect 22855 25533 22913 25545
rect 22855 25157 22867 25533
rect 22901 25157 22913 25533
rect 22855 25145 22913 25157
rect 22973 25533 23031 25545
rect 22973 25157 22985 25533
rect 23019 25157 23031 25533
rect 22973 25145 23031 25157
rect 23091 25533 23149 25545
rect 23091 25157 23103 25533
rect 23137 25157 23149 25533
rect 23091 25145 23149 25157
rect 23209 25533 23267 25545
rect 23209 25157 23221 25533
rect 23255 25157 23267 25533
rect 23209 25145 23267 25157
rect 23327 25533 23385 25545
rect 23327 25157 23339 25533
rect 23373 25157 23385 25533
rect 23327 25145 23385 25157
rect 23445 25533 23503 25545
rect 23445 25157 23457 25533
rect 23491 25157 23503 25533
rect 27397 25537 27455 25549
rect 23445 25145 23503 25157
rect 23574 25333 23632 25345
rect 23574 25157 23586 25333
rect 23620 25157 23632 25333
rect 23574 25145 23632 25157
rect 23692 25333 23750 25345
rect 23692 25157 23704 25333
rect 23738 25157 23750 25333
rect 23692 25145 23750 25157
rect 23810 25333 23868 25345
rect 23810 25157 23822 25333
rect 23856 25157 23868 25333
rect 23810 25145 23868 25157
rect 23928 25333 23986 25345
rect 23928 25157 23940 25333
rect 23974 25157 23986 25333
rect 23928 25145 23986 25157
rect 16146 24845 16204 24857
rect 16146 24469 16158 24845
rect 16192 24469 16204 24845
rect 16146 24457 16204 24469
rect 16264 24845 16322 24857
rect 16264 24469 16276 24845
rect 16310 24469 16322 24845
rect 16264 24457 16322 24469
rect 16382 24845 16440 24857
rect 16382 24469 16394 24845
rect 16428 24469 16440 24845
rect 16382 24457 16440 24469
rect 16500 24845 16558 24857
rect 16500 24469 16512 24845
rect 16546 24469 16558 24845
rect 16500 24457 16558 24469
rect 16618 24845 16676 24857
rect 16618 24469 16630 24845
rect 16664 24469 16676 24845
rect 16618 24457 16676 24469
rect 16736 24845 16794 24857
rect 16736 24469 16748 24845
rect 16782 24469 16794 24845
rect 16736 24457 16794 24469
rect 16854 24845 16912 24857
rect 16854 24469 16866 24845
rect 16900 24469 16912 24845
rect 16854 24457 16912 24469
rect 18886 24346 18944 24358
rect 18886 24170 18898 24346
rect 18932 24170 18944 24346
rect 18886 24158 18944 24170
rect 19004 24346 19062 24358
rect 19004 24170 19016 24346
rect 19050 24170 19062 24346
rect 19004 24158 19062 24170
rect 19122 24346 19180 24358
rect 19122 24170 19134 24346
rect 19168 24170 19180 24346
rect 19122 24158 19180 24170
rect 19240 24346 19298 24358
rect 19240 24170 19252 24346
rect 19286 24170 19298 24346
rect 19240 24158 19298 24170
rect 19358 24346 19416 24358
rect 19358 24170 19370 24346
rect 19404 24170 19416 24346
rect 19358 24158 19416 24170
rect 19476 24346 19534 24358
rect 19476 24170 19488 24346
rect 19522 24170 19534 24346
rect 19476 24158 19534 24170
rect 19594 24346 19652 24358
rect 19594 24170 19606 24346
rect 19640 24170 19652 24346
rect 19594 24158 19652 24170
rect 19712 24346 19770 24358
rect 19712 24170 19724 24346
rect 19758 24170 19770 24346
rect 19712 24158 19770 24170
rect 19830 24346 19888 24358
rect 19830 24170 19842 24346
rect 19876 24170 19888 24346
rect 19830 24158 19888 24170
rect 19948 24346 20006 24358
rect 19948 24170 19960 24346
rect 19994 24170 20006 24346
rect 19948 24158 20006 24170
rect 20782 24840 20840 24852
rect 20782 24464 20794 24840
rect 20828 24464 20840 24840
rect 20782 24452 20840 24464
rect 20900 24840 20958 24852
rect 20900 24464 20912 24840
rect 20946 24464 20958 24840
rect 20900 24452 20958 24464
rect 21018 24840 21076 24852
rect 21018 24464 21030 24840
rect 21064 24464 21076 24840
rect 21018 24452 21076 24464
rect 21136 24840 21194 24852
rect 21136 24464 21148 24840
rect 21182 24464 21194 24840
rect 21136 24452 21194 24464
rect 21254 24840 21312 24852
rect 21254 24464 21266 24840
rect 21300 24464 21312 24840
rect 21254 24452 21312 24464
rect 21372 24840 21430 24852
rect 21372 24464 21384 24840
rect 21418 24464 21430 24840
rect 21372 24452 21430 24464
rect 21490 24840 21548 24852
rect 21490 24464 21502 24840
rect 21536 24464 21548 24840
rect 21490 24452 21548 24464
rect 26913 25337 26971 25349
rect 26913 25161 26925 25337
rect 26959 25161 26971 25337
rect 26913 25149 26971 25161
rect 27031 25337 27089 25349
rect 27031 25161 27043 25337
rect 27077 25161 27089 25337
rect 27031 25149 27089 25161
rect 27149 25337 27207 25349
rect 27149 25161 27161 25337
rect 27195 25161 27207 25337
rect 27149 25149 27207 25161
rect 27267 25337 27325 25349
rect 27267 25161 27279 25337
rect 27313 25161 27325 25337
rect 27267 25149 27325 25161
rect 27397 25161 27409 25537
rect 27443 25161 27455 25537
rect 27397 25149 27455 25161
rect 27515 25537 27573 25549
rect 27515 25161 27527 25537
rect 27561 25161 27573 25537
rect 27515 25149 27573 25161
rect 27633 25537 27691 25549
rect 27633 25161 27645 25537
rect 27679 25161 27691 25537
rect 27633 25149 27691 25161
rect 27751 25537 27809 25549
rect 27751 25161 27763 25537
rect 27797 25161 27809 25537
rect 27751 25149 27809 25161
rect 27869 25537 27927 25549
rect 27869 25161 27881 25537
rect 27915 25161 27927 25537
rect 27869 25149 27927 25161
rect 27987 25537 28045 25549
rect 27987 25161 27999 25537
rect 28033 25161 28045 25537
rect 27987 25149 28045 25161
rect 28105 25537 28163 25549
rect 28105 25161 28117 25537
rect 28151 25161 28163 25537
rect 29295 25537 29353 25549
rect 28105 25149 28163 25161
rect 28234 25337 28292 25349
rect 28234 25161 28246 25337
rect 28280 25161 28292 25337
rect 28234 25149 28292 25161
rect 28352 25337 28410 25349
rect 28352 25161 28364 25337
rect 28398 25161 28410 25337
rect 28352 25149 28410 25161
rect 28470 25337 28528 25349
rect 28470 25161 28482 25337
rect 28516 25161 28528 25337
rect 28470 25149 28528 25161
rect 28588 25337 28646 25349
rect 28588 25161 28600 25337
rect 28634 25161 28646 25337
rect 28588 25149 28646 25161
rect 28811 25337 28869 25349
rect 28811 25161 28823 25337
rect 28857 25161 28869 25337
rect 28811 25149 28869 25161
rect 28929 25337 28987 25349
rect 28929 25161 28941 25337
rect 28975 25161 28987 25337
rect 28929 25149 28987 25161
rect 29047 25337 29105 25349
rect 29047 25161 29059 25337
rect 29093 25161 29105 25337
rect 29047 25149 29105 25161
rect 29165 25337 29223 25349
rect 29165 25161 29177 25337
rect 29211 25161 29223 25337
rect 29165 25149 29223 25161
rect 29295 25161 29307 25537
rect 29341 25161 29353 25537
rect 29295 25149 29353 25161
rect 29413 25537 29471 25549
rect 29413 25161 29425 25537
rect 29459 25161 29471 25537
rect 29413 25149 29471 25161
rect 29531 25537 29589 25549
rect 29531 25161 29543 25537
rect 29577 25161 29589 25537
rect 29531 25149 29589 25161
rect 29649 25537 29707 25549
rect 29649 25161 29661 25537
rect 29695 25161 29707 25537
rect 29649 25149 29707 25161
rect 29767 25537 29825 25549
rect 29767 25161 29779 25537
rect 29813 25161 29825 25537
rect 29767 25149 29825 25161
rect 29885 25537 29943 25549
rect 29885 25161 29897 25537
rect 29931 25161 29943 25537
rect 29885 25149 29943 25161
rect 30003 25537 30061 25549
rect 30003 25161 30015 25537
rect 30049 25161 30061 25537
rect 30003 25149 30061 25161
rect 30132 25337 30190 25349
rect 30132 25161 30144 25337
rect 30178 25161 30190 25337
rect 30132 25149 30190 25161
rect 30250 25337 30308 25349
rect 30250 25161 30262 25337
rect 30296 25161 30308 25337
rect 30250 25149 30308 25161
rect 30368 25337 30426 25349
rect 30368 25161 30380 25337
rect 30414 25161 30426 25337
rect 30368 25149 30426 25161
rect 30486 25337 30544 25349
rect 30486 25161 30498 25337
rect 30532 25161 30544 25337
rect 30486 25149 30544 25161
rect 22680 24840 22738 24852
rect 22680 24464 22692 24840
rect 22726 24464 22738 24840
rect 22680 24452 22738 24464
rect 22798 24840 22856 24852
rect 22798 24464 22810 24840
rect 22844 24464 22856 24840
rect 22798 24452 22856 24464
rect 22916 24840 22974 24852
rect 22916 24464 22928 24840
rect 22962 24464 22974 24840
rect 22916 24452 22974 24464
rect 23034 24840 23092 24852
rect 23034 24464 23046 24840
rect 23080 24464 23092 24840
rect 23034 24452 23092 24464
rect 23152 24840 23210 24852
rect 23152 24464 23164 24840
rect 23198 24464 23210 24840
rect 23152 24452 23210 24464
rect 23270 24840 23328 24852
rect 23270 24464 23282 24840
rect 23316 24464 23328 24840
rect 23270 24452 23328 24464
rect 23388 24840 23446 24852
rect 23388 24464 23400 24840
rect 23434 24464 23446 24840
rect 23388 24452 23446 24464
rect 25444 24350 25502 24362
rect 25444 24174 25456 24350
rect 25490 24174 25502 24350
rect 25444 24162 25502 24174
rect 25562 24350 25620 24362
rect 25562 24174 25574 24350
rect 25608 24174 25620 24350
rect 25562 24162 25620 24174
rect 25680 24350 25738 24362
rect 25680 24174 25692 24350
rect 25726 24174 25738 24350
rect 25680 24162 25738 24174
rect 25798 24350 25856 24362
rect 25798 24174 25810 24350
rect 25844 24174 25856 24350
rect 25798 24162 25856 24174
rect 25916 24350 25974 24362
rect 25916 24174 25928 24350
rect 25962 24174 25974 24350
rect 25916 24162 25974 24174
rect 26034 24350 26092 24362
rect 26034 24174 26046 24350
rect 26080 24174 26092 24350
rect 26034 24162 26092 24174
rect 26152 24350 26210 24362
rect 26152 24174 26164 24350
rect 26198 24174 26210 24350
rect 26152 24162 26210 24174
rect 26270 24350 26328 24362
rect 26270 24174 26282 24350
rect 26316 24174 26328 24350
rect 26270 24162 26328 24174
rect 26388 24350 26446 24362
rect 26388 24174 26400 24350
rect 26434 24174 26446 24350
rect 26388 24162 26446 24174
rect 26506 24350 26564 24362
rect 26506 24174 26518 24350
rect 26552 24174 26564 24350
rect 26506 24162 26564 24174
rect 27340 24844 27398 24856
rect 27340 24468 27352 24844
rect 27386 24468 27398 24844
rect 27340 24456 27398 24468
rect 27458 24844 27516 24856
rect 27458 24468 27470 24844
rect 27504 24468 27516 24844
rect 27458 24456 27516 24468
rect 27576 24844 27634 24856
rect 27576 24468 27588 24844
rect 27622 24468 27634 24844
rect 27576 24456 27634 24468
rect 27694 24844 27752 24856
rect 27694 24468 27706 24844
rect 27740 24468 27752 24844
rect 27694 24456 27752 24468
rect 27812 24844 27870 24856
rect 27812 24468 27824 24844
rect 27858 24468 27870 24844
rect 27812 24456 27870 24468
rect 27930 24844 27988 24856
rect 27930 24468 27942 24844
rect 27976 24468 27988 24844
rect 27930 24456 27988 24468
rect 28048 24844 28106 24856
rect 28048 24468 28060 24844
rect 28094 24468 28106 24844
rect 28048 24456 28106 24468
rect 36955 25148 37155 25160
rect 36955 25114 36967 25148
rect 37143 25114 37155 25148
rect 36955 25102 37155 25114
rect 36955 25030 37155 25042
rect 36955 24996 36967 25030
rect 37143 24996 37155 25030
rect 36955 24984 37155 24996
rect 29238 24844 29296 24856
rect 29238 24468 29250 24844
rect 29284 24468 29296 24844
rect 29238 24456 29296 24468
rect 29356 24844 29414 24856
rect 29356 24468 29368 24844
rect 29402 24468 29414 24844
rect 29356 24456 29414 24468
rect 29474 24844 29532 24856
rect 29474 24468 29486 24844
rect 29520 24468 29532 24844
rect 29474 24456 29532 24468
rect 29592 24844 29650 24856
rect 29592 24468 29604 24844
rect 29638 24468 29650 24844
rect 29592 24456 29650 24468
rect 29710 24844 29768 24856
rect 29710 24468 29722 24844
rect 29756 24468 29768 24844
rect 29710 24456 29768 24468
rect 29828 24844 29886 24856
rect 29828 24468 29840 24844
rect 29874 24468 29886 24844
rect 29828 24456 29886 24468
rect 29946 24844 30004 24856
rect 29946 24468 29958 24844
rect 29992 24468 30004 24844
rect 29946 24456 30004 24468
rect 36955 24912 37155 24924
rect 36955 24878 36967 24912
rect 37143 24878 37155 24912
rect 36955 24866 37155 24878
rect 36955 24794 37155 24806
rect 36955 24760 36967 24794
rect 37143 24760 37155 24794
rect 36955 24719 37155 24760
rect 36755 24707 37155 24719
rect 36755 24673 36767 24707
rect 37143 24673 37155 24707
rect 36755 24661 37155 24673
rect 36755 24589 37155 24601
rect 36755 24555 36767 24589
rect 37143 24555 37155 24589
rect 36755 24543 37155 24555
rect 36755 24471 37155 24483
rect 36755 24437 36767 24471
rect 37143 24437 37155 24471
rect 36755 24425 37155 24437
rect 36755 24353 37155 24365
rect 36755 24319 36767 24353
rect 37143 24319 37155 24353
rect 36755 24307 37155 24319
rect 36755 24240 37155 24252
rect 36755 24206 36767 24240
rect 37143 24206 37155 24240
rect 36755 24194 37155 24206
rect 36755 24122 37155 24134
rect 36755 24088 36767 24122
rect 37143 24088 37155 24122
rect 36755 24076 37155 24088
rect 36755 24004 37155 24016
rect 36755 23970 36767 24004
rect 37143 23970 37155 24004
rect 36755 23958 37155 23970
rect 36755 23886 37155 23898
rect 36755 23852 36767 23886
rect 37143 23852 37155 23886
rect 36755 23840 37155 23852
rect 36755 23768 37155 23780
rect 36755 23734 36767 23768
rect 37143 23734 37155 23768
rect 36755 23722 37155 23734
rect 36755 23650 37155 23662
rect 36755 23616 36767 23650
rect 37143 23616 37155 23650
rect 36755 23604 37155 23616
rect 36755 23532 37155 23544
rect 36755 23498 36767 23532
rect 37143 23498 37155 23532
rect 36755 23486 37155 23498
rect 36755 23413 37155 23425
rect 36755 23379 36767 23413
rect 37143 23379 37155 23413
rect 36755 23367 37155 23379
rect 36755 23295 37155 23307
rect 36755 23261 36767 23295
rect 37143 23261 37155 23295
rect 36755 23249 37155 23261
rect 36755 23177 37155 23189
rect 36755 23143 36767 23177
rect 37143 23143 37155 23177
rect 36755 23131 37155 23143
rect 36755 23059 37155 23071
rect 36755 23025 36767 23059
rect 37143 23025 37155 23059
rect 36755 23013 37155 23025
rect 36955 22940 37155 22952
rect 36955 22906 36967 22940
rect 37143 22906 37155 22940
rect 36955 22894 37155 22906
rect 36955 22822 37155 22834
rect 36955 22788 36967 22822
rect 37143 22788 37155 22822
rect 36955 22776 37155 22788
rect 36955 22704 37155 22716
rect 36955 22670 36967 22704
rect 37143 22670 37155 22704
rect 36955 22658 37155 22670
rect 36955 22586 37155 22598
rect 36955 22552 36967 22586
rect 37143 22552 37155 22586
rect 36955 22540 37155 22552
rect 5841 22076 5899 22088
rect 5841 21700 5853 22076
rect 5887 21700 5899 22076
rect 5841 21688 5899 21700
rect 5959 22076 6017 22088
rect 5959 21700 5971 22076
rect 6005 21700 6017 22076
rect 5959 21688 6017 21700
rect 6077 22076 6135 22088
rect 6077 21700 6089 22076
rect 6123 21700 6135 22076
rect 6077 21688 6135 21700
rect 6195 22076 6253 22088
rect 6195 21700 6207 22076
rect 6241 21700 6253 22076
rect 6195 21688 6253 21700
rect 6313 22076 6371 22088
rect 6313 21700 6325 22076
rect 6359 21700 6371 22076
rect 6313 21688 6371 21700
rect 6431 22076 6489 22088
rect 6431 21700 6443 22076
rect 6477 21700 6489 22076
rect 6431 21688 6489 21700
rect 6549 22076 6607 22088
rect 6549 21700 6561 22076
rect 6595 21700 6607 22076
rect 6549 21688 6607 21700
rect 6983 22072 7041 22084
rect 6983 21696 6995 22072
rect 7029 21696 7041 22072
rect 6983 21684 7041 21696
rect 7101 22072 7159 22084
rect 7101 21696 7113 22072
rect 7147 21696 7159 22072
rect 7101 21684 7159 21696
rect 7219 22072 7277 22084
rect 7219 21696 7231 22072
rect 7265 21696 7277 22072
rect 7219 21684 7277 21696
rect 7337 22072 7395 22084
rect 7337 21696 7349 22072
rect 7383 21696 7395 22072
rect 7337 21684 7395 21696
rect 7455 22072 7513 22084
rect 7455 21696 7467 22072
rect 7501 21696 7513 22072
rect 7455 21684 7513 21696
rect 7573 22072 7631 22084
rect 7573 21696 7585 22072
rect 7619 21696 7631 22072
rect 7573 21684 7631 21696
rect 7691 22072 7749 22084
rect 7691 21696 7703 22072
rect 7737 21696 7749 22072
rect 12399 22072 12457 22084
rect 8954 22000 9012 22012
rect 8954 21824 8966 22000
rect 9000 21824 9012 22000
rect 8954 21812 9012 21824
rect 9072 22000 9130 22012
rect 9072 21824 9084 22000
rect 9118 21824 9130 22000
rect 9072 21812 9130 21824
rect 9190 22000 9248 22012
rect 9190 21824 9202 22000
rect 9236 21824 9248 22000
rect 9190 21812 9248 21824
rect 9308 22000 9366 22012
rect 9308 21824 9320 22000
rect 9354 21824 9366 22000
rect 9308 21812 9366 21824
rect 9426 22000 9484 22012
rect 9426 21824 9438 22000
rect 9472 21824 9484 22000
rect 9426 21812 9484 21824
rect 9544 22000 9602 22012
rect 9544 21824 9556 22000
rect 9590 21824 9602 22000
rect 9544 21812 9602 21824
rect 9662 22000 9720 22012
rect 9662 21824 9674 22000
rect 9708 21824 9720 22000
rect 9662 21812 9720 21824
rect 9780 22000 9838 22012
rect 9780 21824 9792 22000
rect 9826 21824 9838 22000
rect 9780 21812 9838 21824
rect 9898 22000 9956 22012
rect 9898 21824 9910 22000
rect 9944 21824 9956 22000
rect 9898 21812 9956 21824
rect 10016 22000 10074 22012
rect 10016 21824 10028 22000
rect 10062 21824 10074 22000
rect 10016 21812 10074 21824
rect 7691 21684 7749 21696
rect 12399 21696 12411 22072
rect 12445 21696 12457 22072
rect 12399 21684 12457 21696
rect 12517 22072 12575 22084
rect 12517 21696 12529 22072
rect 12563 21696 12575 22072
rect 12517 21684 12575 21696
rect 12635 22072 12693 22084
rect 12635 21696 12647 22072
rect 12681 21696 12693 22072
rect 12635 21684 12693 21696
rect 12753 22072 12811 22084
rect 12753 21696 12765 22072
rect 12799 21696 12811 22072
rect 12753 21684 12811 21696
rect 12871 22072 12929 22084
rect 12871 21696 12883 22072
rect 12917 21696 12929 22072
rect 12871 21684 12929 21696
rect 12989 22072 13047 22084
rect 12989 21696 13001 22072
rect 13035 21696 13047 22072
rect 12989 21684 13047 21696
rect 13107 22072 13165 22084
rect 13107 21696 13119 22072
rect 13153 21696 13165 22072
rect 13107 21684 13165 21696
rect 13541 22068 13599 22080
rect 13541 21692 13553 22068
rect 13587 21692 13599 22068
rect 5766 21293 5824 21305
rect 5766 21117 5778 21293
rect 5812 21117 5824 21293
rect 5766 21105 5824 21117
rect 5884 21293 5942 21305
rect 5884 21117 5896 21293
rect 5930 21117 5942 21293
rect 5884 21105 5942 21117
rect 6002 21293 6060 21305
rect 6002 21117 6014 21293
rect 6048 21117 6060 21293
rect 6002 21105 6060 21117
rect 6120 21293 6178 21305
rect 6120 21117 6132 21293
rect 6166 21117 6178 21293
rect 6120 21105 6178 21117
rect 6908 21289 6966 21301
rect 6908 21113 6920 21289
rect 6954 21113 6966 21289
rect 6908 21101 6966 21113
rect 7026 21289 7084 21301
rect 7026 21113 7038 21289
rect 7072 21113 7084 21289
rect 7026 21101 7084 21113
rect 7144 21289 7202 21301
rect 7144 21113 7156 21289
rect 7190 21113 7202 21289
rect 7144 21101 7202 21113
rect 7262 21289 7320 21301
rect 7262 21113 7274 21289
rect 7308 21113 7320 21289
rect 7262 21101 7320 21113
rect 13541 21680 13599 21692
rect 13659 22068 13717 22080
rect 13659 21692 13671 22068
rect 13705 21692 13717 22068
rect 13659 21680 13717 21692
rect 13777 22068 13835 22080
rect 13777 21692 13789 22068
rect 13823 21692 13835 22068
rect 13777 21680 13835 21692
rect 13895 22068 13953 22080
rect 13895 21692 13907 22068
rect 13941 21692 13953 22068
rect 13895 21680 13953 21692
rect 14013 22068 14071 22080
rect 14013 21692 14025 22068
rect 14059 21692 14071 22068
rect 14013 21680 14071 21692
rect 14131 22068 14189 22080
rect 14131 21692 14143 22068
rect 14177 21692 14189 22068
rect 14131 21680 14189 21692
rect 14249 22068 14307 22080
rect 18933 22077 18991 22089
rect 14249 21692 14261 22068
rect 14295 21692 14307 22068
rect 15512 21996 15570 22008
rect 15512 21820 15524 21996
rect 15558 21820 15570 21996
rect 15512 21808 15570 21820
rect 15630 21996 15688 22008
rect 15630 21820 15642 21996
rect 15676 21820 15688 21996
rect 15630 21808 15688 21820
rect 15748 21996 15806 22008
rect 15748 21820 15760 21996
rect 15794 21820 15806 21996
rect 15748 21808 15806 21820
rect 15866 21996 15924 22008
rect 15866 21820 15878 21996
rect 15912 21820 15924 21996
rect 15866 21808 15924 21820
rect 15984 21996 16042 22008
rect 15984 21820 15996 21996
rect 16030 21820 16042 21996
rect 15984 21808 16042 21820
rect 16102 21996 16160 22008
rect 16102 21820 16114 21996
rect 16148 21820 16160 21996
rect 16102 21808 16160 21820
rect 16220 21996 16278 22008
rect 16220 21820 16232 21996
rect 16266 21820 16278 21996
rect 16220 21808 16278 21820
rect 16338 21996 16396 22008
rect 16338 21820 16350 21996
rect 16384 21820 16396 21996
rect 16338 21808 16396 21820
rect 16456 21996 16514 22008
rect 16456 21820 16468 21996
rect 16502 21820 16514 21996
rect 16456 21808 16514 21820
rect 16574 21996 16632 22008
rect 16574 21820 16586 21996
rect 16620 21820 16632 21996
rect 16574 21808 16632 21820
rect 14249 21680 14307 21692
rect 18933 21701 18945 22077
rect 18979 21701 18991 22077
rect 18933 21689 18991 21701
rect 19051 22077 19109 22089
rect 19051 21701 19063 22077
rect 19097 21701 19109 22077
rect 19051 21689 19109 21701
rect 19169 22077 19227 22089
rect 19169 21701 19181 22077
rect 19215 21701 19227 22077
rect 19169 21689 19227 21701
rect 19287 22077 19345 22089
rect 19287 21701 19299 22077
rect 19333 21701 19345 22077
rect 19287 21689 19345 21701
rect 19405 22077 19463 22089
rect 19405 21701 19417 22077
rect 19451 21701 19463 22077
rect 19405 21689 19463 21701
rect 19523 22077 19581 22089
rect 19523 21701 19535 22077
rect 19569 21701 19581 22077
rect 19523 21689 19581 21701
rect 19641 22077 19699 22089
rect 19641 21701 19653 22077
rect 19687 21701 19699 22077
rect 19641 21689 19699 21701
rect 20075 22073 20133 22085
rect 20075 21697 20087 22073
rect 20121 21697 20133 22073
rect 12324 21289 12382 21301
rect 12324 21113 12336 21289
rect 12370 21113 12382 21289
rect 12324 21101 12382 21113
rect 12442 21289 12500 21301
rect 12442 21113 12454 21289
rect 12488 21113 12500 21289
rect 12442 21101 12500 21113
rect 12560 21289 12618 21301
rect 12560 21113 12572 21289
rect 12606 21113 12618 21289
rect 12560 21101 12618 21113
rect 12678 21289 12736 21301
rect 12678 21113 12690 21289
rect 12724 21113 12736 21289
rect 12678 21101 12736 21113
rect 13466 21285 13524 21297
rect 13466 21109 13478 21285
rect 13512 21109 13524 21285
rect 13466 21097 13524 21109
rect 13584 21285 13642 21297
rect 13584 21109 13596 21285
rect 13630 21109 13642 21285
rect 13584 21097 13642 21109
rect 13702 21285 13760 21297
rect 13702 21109 13714 21285
rect 13748 21109 13760 21285
rect 13702 21097 13760 21109
rect 13820 21285 13878 21297
rect 13820 21109 13832 21285
rect 13866 21109 13878 21285
rect 13820 21097 13878 21109
rect 20075 21685 20133 21697
rect 20193 22073 20251 22085
rect 20193 21697 20205 22073
rect 20239 21697 20251 22073
rect 20193 21685 20251 21697
rect 20311 22073 20369 22085
rect 20311 21697 20323 22073
rect 20357 21697 20369 22073
rect 20311 21685 20369 21697
rect 20429 22073 20487 22085
rect 20429 21697 20441 22073
rect 20475 21697 20487 22073
rect 20429 21685 20487 21697
rect 20547 22073 20605 22085
rect 20547 21697 20559 22073
rect 20593 21697 20605 22073
rect 20547 21685 20605 21697
rect 20665 22073 20723 22085
rect 20665 21697 20677 22073
rect 20711 21697 20723 22073
rect 20665 21685 20723 21697
rect 20783 22073 20841 22085
rect 20783 21697 20795 22073
rect 20829 21697 20841 22073
rect 25446 22080 25504 22092
rect 22046 22001 22104 22013
rect 22046 21825 22058 22001
rect 22092 21825 22104 22001
rect 22046 21813 22104 21825
rect 22164 22001 22222 22013
rect 22164 21825 22176 22001
rect 22210 21825 22222 22001
rect 22164 21813 22222 21825
rect 22282 22001 22340 22013
rect 22282 21825 22294 22001
rect 22328 21825 22340 22001
rect 22282 21813 22340 21825
rect 22400 22001 22458 22013
rect 22400 21825 22412 22001
rect 22446 21825 22458 22001
rect 22400 21813 22458 21825
rect 22518 22001 22576 22013
rect 22518 21825 22530 22001
rect 22564 21825 22576 22001
rect 22518 21813 22576 21825
rect 22636 22001 22694 22013
rect 22636 21825 22648 22001
rect 22682 21825 22694 22001
rect 22636 21813 22694 21825
rect 22754 22001 22812 22013
rect 22754 21825 22766 22001
rect 22800 21825 22812 22001
rect 22754 21813 22812 21825
rect 22872 22001 22930 22013
rect 22872 21825 22884 22001
rect 22918 21825 22930 22001
rect 22872 21813 22930 21825
rect 22990 22001 23048 22013
rect 22990 21825 23002 22001
rect 23036 21825 23048 22001
rect 22990 21813 23048 21825
rect 23108 22001 23166 22013
rect 23108 21825 23120 22001
rect 23154 21825 23166 22001
rect 23108 21813 23166 21825
rect 20783 21685 20841 21697
rect 25446 21704 25458 22080
rect 25492 21704 25504 22080
rect 25446 21692 25504 21704
rect 25564 22080 25622 22092
rect 25564 21704 25576 22080
rect 25610 21704 25622 22080
rect 25564 21692 25622 21704
rect 25682 22080 25740 22092
rect 25682 21704 25694 22080
rect 25728 21704 25740 22080
rect 25682 21692 25740 21704
rect 25800 22080 25858 22092
rect 25800 21704 25812 22080
rect 25846 21704 25858 22080
rect 25800 21692 25858 21704
rect 25918 22080 25976 22092
rect 25918 21704 25930 22080
rect 25964 21704 25976 22080
rect 25918 21692 25976 21704
rect 26036 22080 26094 22092
rect 26036 21704 26048 22080
rect 26082 21704 26094 22080
rect 26036 21692 26094 21704
rect 26154 22080 26212 22092
rect 26154 21704 26166 22080
rect 26200 21704 26212 22080
rect 26154 21692 26212 21704
rect 26588 22076 26646 22088
rect 26588 21700 26600 22076
rect 26634 21700 26646 22076
rect 18858 21294 18916 21306
rect 18858 21118 18870 21294
rect 18904 21118 18916 21294
rect 18858 21106 18916 21118
rect 18976 21294 19034 21306
rect 18976 21118 18988 21294
rect 19022 21118 19034 21294
rect 18976 21106 19034 21118
rect 19094 21294 19152 21306
rect 19094 21118 19106 21294
rect 19140 21118 19152 21294
rect 19094 21106 19152 21118
rect 19212 21294 19270 21306
rect 19212 21118 19224 21294
rect 19258 21118 19270 21294
rect 19212 21106 19270 21118
rect 20000 21290 20058 21302
rect 20000 21114 20012 21290
rect 20046 21114 20058 21290
rect 20000 21102 20058 21114
rect 20118 21290 20176 21302
rect 20118 21114 20130 21290
rect 20164 21114 20176 21290
rect 20118 21102 20176 21114
rect 20236 21290 20294 21302
rect 20236 21114 20248 21290
rect 20282 21114 20294 21290
rect 20236 21102 20294 21114
rect 20354 21290 20412 21302
rect 20354 21114 20366 21290
rect 20400 21114 20412 21290
rect 20354 21102 20412 21114
rect 26588 21688 26646 21700
rect 26706 22076 26764 22088
rect 26706 21700 26718 22076
rect 26752 21700 26764 22076
rect 26706 21688 26764 21700
rect 26824 22076 26882 22088
rect 26824 21700 26836 22076
rect 26870 21700 26882 22076
rect 26824 21688 26882 21700
rect 26942 22076 27000 22088
rect 26942 21700 26954 22076
rect 26988 21700 27000 22076
rect 26942 21688 27000 21700
rect 27060 22076 27118 22088
rect 27060 21700 27072 22076
rect 27106 21700 27118 22076
rect 27060 21688 27118 21700
rect 27178 22076 27236 22088
rect 27178 21700 27190 22076
rect 27224 21700 27236 22076
rect 27178 21688 27236 21700
rect 27296 22076 27354 22088
rect 27296 21700 27308 22076
rect 27342 21700 27354 22076
rect 28559 22004 28617 22016
rect 28559 21828 28571 22004
rect 28605 21828 28617 22004
rect 28559 21816 28617 21828
rect 28677 22004 28735 22016
rect 28677 21828 28689 22004
rect 28723 21828 28735 22004
rect 28677 21816 28735 21828
rect 28795 22004 28853 22016
rect 28795 21828 28807 22004
rect 28841 21828 28853 22004
rect 28795 21816 28853 21828
rect 28913 22004 28971 22016
rect 28913 21828 28925 22004
rect 28959 21828 28971 22004
rect 28913 21816 28971 21828
rect 29031 22004 29089 22016
rect 29031 21828 29043 22004
rect 29077 21828 29089 22004
rect 29031 21816 29089 21828
rect 29149 22004 29207 22016
rect 29149 21828 29161 22004
rect 29195 21828 29207 22004
rect 29149 21816 29207 21828
rect 29267 22004 29325 22016
rect 29267 21828 29279 22004
rect 29313 21828 29325 22004
rect 29267 21816 29325 21828
rect 29385 22004 29443 22016
rect 29385 21828 29397 22004
rect 29431 21828 29443 22004
rect 29385 21816 29443 21828
rect 29503 22004 29561 22016
rect 29503 21828 29515 22004
rect 29549 21828 29561 22004
rect 29503 21816 29561 21828
rect 29621 22004 29679 22016
rect 29621 21828 29633 22004
rect 29667 21828 29679 22004
rect 36955 22004 37155 22016
rect 36955 21970 36967 22004
rect 37143 21970 37155 22004
rect 36955 21958 37155 21970
rect 29621 21816 29679 21828
rect 36955 21886 37155 21898
rect 36955 21852 36967 21886
rect 37143 21852 37155 21886
rect 36955 21840 37155 21852
rect 27296 21688 27354 21700
rect 36955 21768 37155 21780
rect 36955 21734 36967 21768
rect 37143 21734 37155 21768
rect 36955 21722 37155 21734
rect 36955 21650 37155 21662
rect 36955 21616 36967 21650
rect 37143 21616 37155 21650
rect 25371 21297 25429 21309
rect 25371 21121 25383 21297
rect 25417 21121 25429 21297
rect 25371 21109 25429 21121
rect 25489 21297 25547 21309
rect 25489 21121 25501 21297
rect 25535 21121 25547 21297
rect 25489 21109 25547 21121
rect 25607 21297 25665 21309
rect 25607 21121 25619 21297
rect 25653 21121 25665 21297
rect 25607 21109 25665 21121
rect 25725 21297 25783 21309
rect 25725 21121 25737 21297
rect 25771 21121 25783 21297
rect 25725 21109 25783 21121
rect 26513 21293 26571 21305
rect 26513 21117 26525 21293
rect 26559 21117 26571 21293
rect 26513 21105 26571 21117
rect 26631 21293 26689 21305
rect 26631 21117 26643 21293
rect 26677 21117 26689 21293
rect 26631 21105 26689 21117
rect 26749 21293 26807 21305
rect 26749 21117 26761 21293
rect 26795 21117 26807 21293
rect 26749 21105 26807 21117
rect 26867 21293 26925 21305
rect 26867 21117 26879 21293
rect 26913 21117 26925 21293
rect 26867 21105 26925 21117
rect 36955 21575 37155 21616
rect 36755 21563 37155 21575
rect 36755 21529 36767 21563
rect 37143 21529 37155 21563
rect 36755 21517 37155 21529
rect 36755 21445 37155 21457
rect 36755 21411 36767 21445
rect 37143 21411 37155 21445
rect 36755 21399 37155 21411
rect 36755 21327 37155 21339
rect 36755 21293 36767 21327
rect 37143 21293 37155 21327
rect 36755 21281 37155 21293
rect 36755 21209 37155 21221
rect 36755 21175 36767 21209
rect 37143 21175 37155 21209
rect 36755 21163 37155 21175
rect 36755 21096 37155 21108
rect 36755 21062 36767 21096
rect 37143 21062 37155 21096
rect 36755 21050 37155 21062
rect 36755 20978 37155 20990
rect 36755 20944 36767 20978
rect 37143 20944 37155 20978
rect 36755 20932 37155 20944
rect 36755 20860 37155 20872
rect 36755 20826 36767 20860
rect 37143 20826 37155 20860
rect 36755 20814 37155 20826
rect 36755 20742 37155 20754
rect 36755 20708 36767 20742
rect 37143 20708 37155 20742
rect 36755 20696 37155 20708
rect 36755 20624 37155 20636
rect 36755 20590 36767 20624
rect 37143 20590 37155 20624
rect 36755 20578 37155 20590
rect 8940 20350 8998 20362
rect 8940 20174 8952 20350
rect 8986 20174 8998 20350
rect 8940 20162 8998 20174
rect 9058 20350 9116 20362
rect 9058 20174 9070 20350
rect 9104 20174 9116 20350
rect 9058 20162 9116 20174
rect 9176 20350 9234 20362
rect 9176 20174 9188 20350
rect 9222 20174 9234 20350
rect 9176 20162 9234 20174
rect 9294 20350 9352 20362
rect 9294 20174 9306 20350
rect 9340 20174 9352 20350
rect 9294 20162 9352 20174
rect 9412 20350 9470 20362
rect 9412 20174 9424 20350
rect 9458 20174 9470 20350
rect 9412 20162 9470 20174
rect 9530 20350 9588 20362
rect 9530 20174 9542 20350
rect 9576 20174 9588 20350
rect 9530 20162 9588 20174
rect 9648 20350 9706 20362
rect 9648 20174 9660 20350
rect 9694 20174 9706 20350
rect 9648 20162 9706 20174
rect 9766 20350 9824 20362
rect 9766 20174 9778 20350
rect 9812 20174 9824 20350
rect 9766 20162 9824 20174
rect 9884 20350 9942 20362
rect 9884 20174 9896 20350
rect 9930 20174 9942 20350
rect 9884 20162 9942 20174
rect 10002 20350 10060 20362
rect 10002 20174 10014 20350
rect 10048 20174 10060 20350
rect 15498 20346 15556 20358
rect 10002 20162 10060 20174
rect 15498 20170 15510 20346
rect 15544 20170 15556 20346
rect 15498 20158 15556 20170
rect 15616 20346 15674 20358
rect 15616 20170 15628 20346
rect 15662 20170 15674 20346
rect 15616 20158 15674 20170
rect 15734 20346 15792 20358
rect 15734 20170 15746 20346
rect 15780 20170 15792 20346
rect 15734 20158 15792 20170
rect 15852 20346 15910 20358
rect 15852 20170 15864 20346
rect 15898 20170 15910 20346
rect 15852 20158 15910 20170
rect 15970 20346 16028 20358
rect 15970 20170 15982 20346
rect 16016 20170 16028 20346
rect 15970 20158 16028 20170
rect 16088 20346 16146 20358
rect 16088 20170 16100 20346
rect 16134 20170 16146 20346
rect 16088 20158 16146 20170
rect 16206 20346 16264 20358
rect 16206 20170 16218 20346
rect 16252 20170 16264 20346
rect 16206 20158 16264 20170
rect 16324 20346 16382 20358
rect 16324 20170 16336 20346
rect 16370 20170 16382 20346
rect 16324 20158 16382 20170
rect 16442 20346 16500 20358
rect 16442 20170 16454 20346
rect 16488 20170 16500 20346
rect 16442 20158 16500 20170
rect 16560 20346 16618 20358
rect 16560 20170 16572 20346
rect 16606 20170 16618 20346
rect 22032 20351 22090 20363
rect 16560 20158 16618 20170
rect 22032 20175 22044 20351
rect 22078 20175 22090 20351
rect 22032 20163 22090 20175
rect 22150 20351 22208 20363
rect 22150 20175 22162 20351
rect 22196 20175 22208 20351
rect 22150 20163 22208 20175
rect 22268 20351 22326 20363
rect 22268 20175 22280 20351
rect 22314 20175 22326 20351
rect 22268 20163 22326 20175
rect 22386 20351 22444 20363
rect 22386 20175 22398 20351
rect 22432 20175 22444 20351
rect 22386 20163 22444 20175
rect 22504 20351 22562 20363
rect 22504 20175 22516 20351
rect 22550 20175 22562 20351
rect 22504 20163 22562 20175
rect 22622 20351 22680 20363
rect 22622 20175 22634 20351
rect 22668 20175 22680 20351
rect 22622 20163 22680 20175
rect 22740 20351 22798 20363
rect 22740 20175 22752 20351
rect 22786 20175 22798 20351
rect 22740 20163 22798 20175
rect 22858 20351 22916 20363
rect 22858 20175 22870 20351
rect 22904 20175 22916 20351
rect 22858 20163 22916 20175
rect 22976 20351 23034 20363
rect 22976 20175 22988 20351
rect 23022 20175 23034 20351
rect 22976 20163 23034 20175
rect 23094 20351 23152 20363
rect 23094 20175 23106 20351
rect 23140 20175 23152 20351
rect 36755 20506 37155 20518
rect 36755 20472 36767 20506
rect 37143 20472 37155 20506
rect 36755 20460 37155 20472
rect 36755 20388 37155 20400
rect 28545 20354 28603 20366
rect 23094 20163 23152 20175
rect 28545 20178 28557 20354
rect 28591 20178 28603 20354
rect 28545 20166 28603 20178
rect 28663 20354 28721 20366
rect 28663 20178 28675 20354
rect 28709 20178 28721 20354
rect 28663 20166 28721 20178
rect 28781 20354 28839 20366
rect 28781 20178 28793 20354
rect 28827 20178 28839 20354
rect 28781 20166 28839 20178
rect 28899 20354 28957 20366
rect 28899 20178 28911 20354
rect 28945 20178 28957 20354
rect 28899 20166 28957 20178
rect 29017 20354 29075 20366
rect 29017 20178 29029 20354
rect 29063 20178 29075 20354
rect 29017 20166 29075 20178
rect 29135 20354 29193 20366
rect 29135 20178 29147 20354
rect 29181 20178 29193 20354
rect 29135 20166 29193 20178
rect 29253 20354 29311 20366
rect 29253 20178 29265 20354
rect 29299 20178 29311 20354
rect 29253 20166 29311 20178
rect 29371 20354 29429 20366
rect 29371 20178 29383 20354
rect 29417 20178 29429 20354
rect 29371 20166 29429 20178
rect 29489 20354 29547 20366
rect 29489 20178 29501 20354
rect 29535 20178 29547 20354
rect 29489 20166 29547 20178
rect 29607 20354 29665 20366
rect 29607 20178 29619 20354
rect 29653 20178 29665 20354
rect 36755 20354 36767 20388
rect 37143 20354 37155 20388
rect 36755 20342 37155 20354
rect 36755 20269 37155 20281
rect 36755 20235 36767 20269
rect 37143 20235 37155 20269
rect 36755 20223 37155 20235
rect 29607 20166 29665 20178
rect 5448 19933 5506 19945
rect 4965 19733 5023 19745
rect 4965 19557 4977 19733
rect 5011 19557 5023 19733
rect 4965 19545 5023 19557
rect 5083 19733 5141 19745
rect 5083 19557 5095 19733
rect 5129 19557 5141 19733
rect 5083 19545 5141 19557
rect 5201 19733 5259 19745
rect 5201 19557 5213 19733
rect 5247 19557 5259 19733
rect 5201 19545 5259 19557
rect 5319 19733 5377 19745
rect 5319 19557 5331 19733
rect 5365 19557 5377 19733
rect 5319 19545 5377 19557
rect 5448 19557 5460 19933
rect 5494 19557 5506 19933
rect 5448 19545 5506 19557
rect 5566 19933 5624 19945
rect 5566 19557 5578 19933
rect 5612 19557 5624 19933
rect 5566 19545 5624 19557
rect 5684 19933 5742 19945
rect 5684 19557 5696 19933
rect 5730 19557 5742 19933
rect 5684 19545 5742 19557
rect 5802 19933 5860 19945
rect 5802 19557 5814 19933
rect 5848 19557 5860 19933
rect 5802 19545 5860 19557
rect 5920 19933 5978 19945
rect 5920 19557 5932 19933
rect 5966 19557 5978 19933
rect 5920 19545 5978 19557
rect 6038 19933 6096 19945
rect 6038 19557 6050 19933
rect 6084 19557 6096 19933
rect 6038 19545 6096 19557
rect 6156 19933 6214 19945
rect 6156 19557 6168 19933
rect 6202 19557 6214 19933
rect 7346 19933 7404 19945
rect 6156 19545 6214 19557
rect 6286 19733 6344 19745
rect 6286 19557 6298 19733
rect 6332 19557 6344 19733
rect 6286 19545 6344 19557
rect 6404 19733 6462 19745
rect 6404 19557 6416 19733
rect 6450 19557 6462 19733
rect 6404 19545 6462 19557
rect 6522 19733 6580 19745
rect 6522 19557 6534 19733
rect 6568 19557 6580 19733
rect 6522 19545 6580 19557
rect 6640 19733 6698 19745
rect 6640 19557 6652 19733
rect 6686 19557 6698 19733
rect 6640 19545 6698 19557
rect 6863 19733 6921 19745
rect 6863 19557 6875 19733
rect 6909 19557 6921 19733
rect 6863 19545 6921 19557
rect 6981 19733 7039 19745
rect 6981 19557 6993 19733
rect 7027 19557 7039 19733
rect 6981 19545 7039 19557
rect 7099 19733 7157 19745
rect 7099 19557 7111 19733
rect 7145 19557 7157 19733
rect 7099 19545 7157 19557
rect 7217 19733 7275 19745
rect 7217 19557 7229 19733
rect 7263 19557 7275 19733
rect 7217 19545 7275 19557
rect 7346 19557 7358 19933
rect 7392 19557 7404 19933
rect 7346 19545 7404 19557
rect 7464 19933 7522 19945
rect 7464 19557 7476 19933
rect 7510 19557 7522 19933
rect 7464 19545 7522 19557
rect 7582 19933 7640 19945
rect 7582 19557 7594 19933
rect 7628 19557 7640 19933
rect 7582 19545 7640 19557
rect 7700 19933 7758 19945
rect 7700 19557 7712 19933
rect 7746 19557 7758 19933
rect 7700 19545 7758 19557
rect 7818 19933 7876 19945
rect 7818 19557 7830 19933
rect 7864 19557 7876 19933
rect 7818 19545 7876 19557
rect 7936 19933 7994 19945
rect 7936 19557 7948 19933
rect 7982 19557 7994 19933
rect 7936 19545 7994 19557
rect 8054 19933 8112 19945
rect 8054 19557 8066 19933
rect 8100 19557 8112 19933
rect 12006 19929 12064 19941
rect 8054 19545 8112 19557
rect 8184 19733 8242 19745
rect 8184 19557 8196 19733
rect 8230 19557 8242 19733
rect 8184 19545 8242 19557
rect 8302 19733 8360 19745
rect 8302 19557 8314 19733
rect 8348 19557 8360 19733
rect 8302 19545 8360 19557
rect 8420 19733 8478 19745
rect 8420 19557 8432 19733
rect 8466 19557 8478 19733
rect 8420 19545 8478 19557
rect 8538 19733 8596 19745
rect 8538 19557 8550 19733
rect 8584 19557 8596 19733
rect 8538 19545 8596 19557
rect 5505 19240 5563 19252
rect 5505 18864 5517 19240
rect 5551 18864 5563 19240
rect 5505 18852 5563 18864
rect 5623 19240 5681 19252
rect 5623 18864 5635 19240
rect 5669 18864 5681 19240
rect 5623 18852 5681 18864
rect 5741 19240 5799 19252
rect 5741 18864 5753 19240
rect 5787 18864 5799 19240
rect 5741 18852 5799 18864
rect 5859 19240 5917 19252
rect 5859 18864 5871 19240
rect 5905 18864 5917 19240
rect 5859 18852 5917 18864
rect 5977 19240 6035 19252
rect 5977 18864 5989 19240
rect 6023 18864 6035 19240
rect 5977 18852 6035 18864
rect 6095 19240 6153 19252
rect 6095 18864 6107 19240
rect 6141 18864 6153 19240
rect 6095 18852 6153 18864
rect 6213 19240 6271 19252
rect 6213 18864 6225 19240
rect 6259 18864 6271 19240
rect 6213 18852 6271 18864
rect 11523 19729 11581 19741
rect 11523 19553 11535 19729
rect 11569 19553 11581 19729
rect 11523 19541 11581 19553
rect 11641 19729 11699 19741
rect 11641 19553 11653 19729
rect 11687 19553 11699 19729
rect 11641 19541 11699 19553
rect 11759 19729 11817 19741
rect 11759 19553 11771 19729
rect 11805 19553 11817 19729
rect 11759 19541 11817 19553
rect 11877 19729 11935 19741
rect 11877 19553 11889 19729
rect 11923 19553 11935 19729
rect 11877 19541 11935 19553
rect 12006 19553 12018 19929
rect 12052 19553 12064 19929
rect 12006 19541 12064 19553
rect 12124 19929 12182 19941
rect 12124 19553 12136 19929
rect 12170 19553 12182 19929
rect 12124 19541 12182 19553
rect 12242 19929 12300 19941
rect 12242 19553 12254 19929
rect 12288 19553 12300 19929
rect 12242 19541 12300 19553
rect 12360 19929 12418 19941
rect 12360 19553 12372 19929
rect 12406 19553 12418 19929
rect 12360 19541 12418 19553
rect 12478 19929 12536 19941
rect 12478 19553 12490 19929
rect 12524 19553 12536 19929
rect 12478 19541 12536 19553
rect 12596 19929 12654 19941
rect 12596 19553 12608 19929
rect 12642 19553 12654 19929
rect 12596 19541 12654 19553
rect 12714 19929 12772 19941
rect 12714 19553 12726 19929
rect 12760 19553 12772 19929
rect 13904 19929 13962 19941
rect 12714 19541 12772 19553
rect 12844 19729 12902 19741
rect 12844 19553 12856 19729
rect 12890 19553 12902 19729
rect 12844 19541 12902 19553
rect 12962 19729 13020 19741
rect 12962 19553 12974 19729
rect 13008 19553 13020 19729
rect 12962 19541 13020 19553
rect 13080 19729 13138 19741
rect 13080 19553 13092 19729
rect 13126 19553 13138 19729
rect 13080 19541 13138 19553
rect 13198 19729 13256 19741
rect 13198 19553 13210 19729
rect 13244 19553 13256 19729
rect 13198 19541 13256 19553
rect 13421 19729 13479 19741
rect 13421 19553 13433 19729
rect 13467 19553 13479 19729
rect 13421 19541 13479 19553
rect 13539 19729 13597 19741
rect 13539 19553 13551 19729
rect 13585 19553 13597 19729
rect 13539 19541 13597 19553
rect 13657 19729 13715 19741
rect 13657 19553 13669 19729
rect 13703 19553 13715 19729
rect 13657 19541 13715 19553
rect 13775 19729 13833 19741
rect 13775 19553 13787 19729
rect 13821 19553 13833 19729
rect 13775 19541 13833 19553
rect 13904 19553 13916 19929
rect 13950 19553 13962 19929
rect 13904 19541 13962 19553
rect 14022 19929 14080 19941
rect 14022 19553 14034 19929
rect 14068 19553 14080 19929
rect 14022 19541 14080 19553
rect 14140 19929 14198 19941
rect 14140 19553 14152 19929
rect 14186 19553 14198 19929
rect 14140 19541 14198 19553
rect 14258 19929 14316 19941
rect 14258 19553 14270 19929
rect 14304 19553 14316 19929
rect 14258 19541 14316 19553
rect 14376 19929 14434 19941
rect 14376 19553 14388 19929
rect 14422 19553 14434 19929
rect 14376 19541 14434 19553
rect 14494 19929 14552 19941
rect 14494 19553 14506 19929
rect 14540 19553 14552 19929
rect 14494 19541 14552 19553
rect 14612 19929 14670 19941
rect 14612 19553 14624 19929
rect 14658 19553 14670 19929
rect 18540 19934 18598 19946
rect 14612 19541 14670 19553
rect 14742 19729 14800 19741
rect 14742 19553 14754 19729
rect 14788 19553 14800 19729
rect 14742 19541 14800 19553
rect 14860 19729 14918 19741
rect 14860 19553 14872 19729
rect 14906 19553 14918 19729
rect 14860 19541 14918 19553
rect 14978 19729 15036 19741
rect 14978 19553 14990 19729
rect 15024 19553 15036 19729
rect 14978 19541 15036 19553
rect 15096 19729 15154 19741
rect 15096 19553 15108 19729
rect 15142 19553 15154 19729
rect 15096 19541 15154 19553
rect 7403 19240 7461 19252
rect 7403 18864 7415 19240
rect 7449 18864 7461 19240
rect 7403 18852 7461 18864
rect 7521 19240 7579 19252
rect 7521 18864 7533 19240
rect 7567 18864 7579 19240
rect 7521 18852 7579 18864
rect 7639 19240 7697 19252
rect 7639 18864 7651 19240
rect 7685 18864 7697 19240
rect 7639 18852 7697 18864
rect 7757 19240 7815 19252
rect 7757 18864 7769 19240
rect 7803 18864 7815 19240
rect 7757 18852 7815 18864
rect 7875 19240 7933 19252
rect 7875 18864 7887 19240
rect 7921 18864 7933 19240
rect 7875 18852 7933 18864
rect 7993 19240 8051 19252
rect 7993 18864 8005 19240
rect 8039 18864 8051 19240
rect 7993 18852 8051 18864
rect 8111 19240 8169 19252
rect 8111 18864 8123 19240
rect 8157 18864 8169 19240
rect 8111 18852 8169 18864
rect 8945 18746 9003 18758
rect 8945 18570 8957 18746
rect 8991 18570 9003 18746
rect 8945 18558 9003 18570
rect 9063 18746 9121 18758
rect 9063 18570 9075 18746
rect 9109 18570 9121 18746
rect 9063 18558 9121 18570
rect 9181 18746 9239 18758
rect 9181 18570 9193 18746
rect 9227 18570 9239 18746
rect 9181 18558 9239 18570
rect 9299 18746 9357 18758
rect 9299 18570 9311 18746
rect 9345 18570 9357 18746
rect 9299 18558 9357 18570
rect 9417 18746 9475 18758
rect 9417 18570 9429 18746
rect 9463 18570 9475 18746
rect 9417 18558 9475 18570
rect 9535 18746 9593 18758
rect 9535 18570 9547 18746
rect 9581 18570 9593 18746
rect 9535 18558 9593 18570
rect 9653 18746 9711 18758
rect 9653 18570 9665 18746
rect 9699 18570 9711 18746
rect 9653 18558 9711 18570
rect 9771 18746 9829 18758
rect 9771 18570 9783 18746
rect 9817 18570 9829 18746
rect 9771 18558 9829 18570
rect 9889 18746 9947 18758
rect 9889 18570 9901 18746
rect 9935 18570 9947 18746
rect 9889 18558 9947 18570
rect 10007 18746 10065 18758
rect 10007 18570 10019 18746
rect 10053 18570 10065 18746
rect 10007 18558 10065 18570
rect 12063 19236 12121 19248
rect 12063 18860 12075 19236
rect 12109 18860 12121 19236
rect 12063 18848 12121 18860
rect 12181 19236 12239 19248
rect 12181 18860 12193 19236
rect 12227 18860 12239 19236
rect 12181 18848 12239 18860
rect 12299 19236 12357 19248
rect 12299 18860 12311 19236
rect 12345 18860 12357 19236
rect 12299 18848 12357 18860
rect 12417 19236 12475 19248
rect 12417 18860 12429 19236
rect 12463 18860 12475 19236
rect 12417 18848 12475 18860
rect 12535 19236 12593 19248
rect 12535 18860 12547 19236
rect 12581 18860 12593 19236
rect 12535 18848 12593 18860
rect 12653 19236 12711 19248
rect 12653 18860 12665 19236
rect 12699 18860 12711 19236
rect 12653 18848 12711 18860
rect 12771 19236 12829 19248
rect 12771 18860 12783 19236
rect 12817 18860 12829 19236
rect 12771 18848 12829 18860
rect 18057 19734 18115 19746
rect 18057 19558 18069 19734
rect 18103 19558 18115 19734
rect 18057 19546 18115 19558
rect 18175 19734 18233 19746
rect 18175 19558 18187 19734
rect 18221 19558 18233 19734
rect 18175 19546 18233 19558
rect 18293 19734 18351 19746
rect 18293 19558 18305 19734
rect 18339 19558 18351 19734
rect 18293 19546 18351 19558
rect 18411 19734 18469 19746
rect 18411 19558 18423 19734
rect 18457 19558 18469 19734
rect 18411 19546 18469 19558
rect 18540 19558 18552 19934
rect 18586 19558 18598 19934
rect 18540 19546 18598 19558
rect 18658 19934 18716 19946
rect 18658 19558 18670 19934
rect 18704 19558 18716 19934
rect 18658 19546 18716 19558
rect 18776 19934 18834 19946
rect 18776 19558 18788 19934
rect 18822 19558 18834 19934
rect 18776 19546 18834 19558
rect 18894 19934 18952 19946
rect 18894 19558 18906 19934
rect 18940 19558 18952 19934
rect 18894 19546 18952 19558
rect 19012 19934 19070 19946
rect 19012 19558 19024 19934
rect 19058 19558 19070 19934
rect 19012 19546 19070 19558
rect 19130 19934 19188 19946
rect 19130 19558 19142 19934
rect 19176 19558 19188 19934
rect 19130 19546 19188 19558
rect 19248 19934 19306 19946
rect 19248 19558 19260 19934
rect 19294 19558 19306 19934
rect 20438 19934 20496 19946
rect 19248 19546 19306 19558
rect 19378 19734 19436 19746
rect 19378 19558 19390 19734
rect 19424 19558 19436 19734
rect 19378 19546 19436 19558
rect 19496 19734 19554 19746
rect 19496 19558 19508 19734
rect 19542 19558 19554 19734
rect 19496 19546 19554 19558
rect 19614 19734 19672 19746
rect 19614 19558 19626 19734
rect 19660 19558 19672 19734
rect 19614 19546 19672 19558
rect 19732 19734 19790 19746
rect 19732 19558 19744 19734
rect 19778 19558 19790 19734
rect 19732 19546 19790 19558
rect 19955 19734 20013 19746
rect 19955 19558 19967 19734
rect 20001 19558 20013 19734
rect 19955 19546 20013 19558
rect 20073 19734 20131 19746
rect 20073 19558 20085 19734
rect 20119 19558 20131 19734
rect 20073 19546 20131 19558
rect 20191 19734 20249 19746
rect 20191 19558 20203 19734
rect 20237 19558 20249 19734
rect 20191 19546 20249 19558
rect 20309 19734 20367 19746
rect 20309 19558 20321 19734
rect 20355 19558 20367 19734
rect 20309 19546 20367 19558
rect 20438 19558 20450 19934
rect 20484 19558 20496 19934
rect 20438 19546 20496 19558
rect 20556 19934 20614 19946
rect 20556 19558 20568 19934
rect 20602 19558 20614 19934
rect 20556 19546 20614 19558
rect 20674 19934 20732 19946
rect 20674 19558 20686 19934
rect 20720 19558 20732 19934
rect 20674 19546 20732 19558
rect 20792 19934 20850 19946
rect 20792 19558 20804 19934
rect 20838 19558 20850 19934
rect 20792 19546 20850 19558
rect 20910 19934 20968 19946
rect 20910 19558 20922 19934
rect 20956 19558 20968 19934
rect 20910 19546 20968 19558
rect 21028 19934 21086 19946
rect 21028 19558 21040 19934
rect 21074 19558 21086 19934
rect 21028 19546 21086 19558
rect 21146 19934 21204 19946
rect 21146 19558 21158 19934
rect 21192 19558 21204 19934
rect 25053 19937 25111 19949
rect 21146 19546 21204 19558
rect 21276 19734 21334 19746
rect 21276 19558 21288 19734
rect 21322 19558 21334 19734
rect 21276 19546 21334 19558
rect 21394 19734 21452 19746
rect 21394 19558 21406 19734
rect 21440 19558 21452 19734
rect 21394 19546 21452 19558
rect 21512 19734 21570 19746
rect 21512 19558 21524 19734
rect 21558 19558 21570 19734
rect 21512 19546 21570 19558
rect 21630 19734 21688 19746
rect 21630 19558 21642 19734
rect 21676 19558 21688 19734
rect 21630 19546 21688 19558
rect 13961 19236 14019 19248
rect 13961 18860 13973 19236
rect 14007 18860 14019 19236
rect 13961 18848 14019 18860
rect 14079 19236 14137 19248
rect 14079 18860 14091 19236
rect 14125 18860 14137 19236
rect 14079 18848 14137 18860
rect 14197 19236 14255 19248
rect 14197 18860 14209 19236
rect 14243 18860 14255 19236
rect 14197 18848 14255 18860
rect 14315 19236 14373 19248
rect 14315 18860 14327 19236
rect 14361 18860 14373 19236
rect 14315 18848 14373 18860
rect 14433 19236 14491 19248
rect 14433 18860 14445 19236
rect 14479 18860 14491 19236
rect 14433 18848 14491 18860
rect 14551 19236 14609 19248
rect 14551 18860 14563 19236
rect 14597 18860 14609 19236
rect 14551 18848 14609 18860
rect 14669 19236 14727 19248
rect 14669 18860 14681 19236
rect 14715 18860 14727 19236
rect 14669 18848 14727 18860
rect 15503 18742 15561 18754
rect 15503 18566 15515 18742
rect 15549 18566 15561 18742
rect 15503 18554 15561 18566
rect 15621 18742 15679 18754
rect 15621 18566 15633 18742
rect 15667 18566 15679 18742
rect 15621 18554 15679 18566
rect 15739 18742 15797 18754
rect 15739 18566 15751 18742
rect 15785 18566 15797 18742
rect 15739 18554 15797 18566
rect 15857 18742 15915 18754
rect 15857 18566 15869 18742
rect 15903 18566 15915 18742
rect 15857 18554 15915 18566
rect 15975 18742 16033 18754
rect 15975 18566 15987 18742
rect 16021 18566 16033 18742
rect 15975 18554 16033 18566
rect 16093 18742 16151 18754
rect 16093 18566 16105 18742
rect 16139 18566 16151 18742
rect 16093 18554 16151 18566
rect 16211 18742 16269 18754
rect 16211 18566 16223 18742
rect 16257 18566 16269 18742
rect 16211 18554 16269 18566
rect 16329 18742 16387 18754
rect 16329 18566 16341 18742
rect 16375 18566 16387 18742
rect 16329 18554 16387 18566
rect 16447 18742 16505 18754
rect 16447 18566 16459 18742
rect 16493 18566 16505 18742
rect 16447 18554 16505 18566
rect 16565 18742 16623 18754
rect 16565 18566 16577 18742
rect 16611 18566 16623 18742
rect 16565 18554 16623 18566
rect 18597 19241 18655 19253
rect 18597 18865 18609 19241
rect 18643 18865 18655 19241
rect 18597 18853 18655 18865
rect 18715 19241 18773 19253
rect 18715 18865 18727 19241
rect 18761 18865 18773 19241
rect 18715 18853 18773 18865
rect 18833 19241 18891 19253
rect 18833 18865 18845 19241
rect 18879 18865 18891 19241
rect 18833 18853 18891 18865
rect 18951 19241 19009 19253
rect 18951 18865 18963 19241
rect 18997 18865 19009 19241
rect 18951 18853 19009 18865
rect 19069 19241 19127 19253
rect 19069 18865 19081 19241
rect 19115 18865 19127 19241
rect 19069 18853 19127 18865
rect 19187 19241 19245 19253
rect 19187 18865 19199 19241
rect 19233 18865 19245 19241
rect 19187 18853 19245 18865
rect 19305 19241 19363 19253
rect 19305 18865 19317 19241
rect 19351 18865 19363 19241
rect 19305 18853 19363 18865
rect 24570 19737 24628 19749
rect 24570 19561 24582 19737
rect 24616 19561 24628 19737
rect 24570 19549 24628 19561
rect 24688 19737 24746 19749
rect 24688 19561 24700 19737
rect 24734 19561 24746 19737
rect 24688 19549 24746 19561
rect 24806 19737 24864 19749
rect 24806 19561 24818 19737
rect 24852 19561 24864 19737
rect 24806 19549 24864 19561
rect 24924 19737 24982 19749
rect 24924 19561 24936 19737
rect 24970 19561 24982 19737
rect 24924 19549 24982 19561
rect 25053 19561 25065 19937
rect 25099 19561 25111 19937
rect 25053 19549 25111 19561
rect 25171 19937 25229 19949
rect 25171 19561 25183 19937
rect 25217 19561 25229 19937
rect 25171 19549 25229 19561
rect 25289 19937 25347 19949
rect 25289 19561 25301 19937
rect 25335 19561 25347 19937
rect 25289 19549 25347 19561
rect 25407 19937 25465 19949
rect 25407 19561 25419 19937
rect 25453 19561 25465 19937
rect 25407 19549 25465 19561
rect 25525 19937 25583 19949
rect 25525 19561 25537 19937
rect 25571 19561 25583 19937
rect 25525 19549 25583 19561
rect 25643 19937 25701 19949
rect 25643 19561 25655 19937
rect 25689 19561 25701 19937
rect 25643 19549 25701 19561
rect 25761 19937 25819 19949
rect 25761 19561 25773 19937
rect 25807 19561 25819 19937
rect 26951 19937 27009 19949
rect 25761 19549 25819 19561
rect 25891 19737 25949 19749
rect 25891 19561 25903 19737
rect 25937 19561 25949 19737
rect 25891 19549 25949 19561
rect 26009 19737 26067 19749
rect 26009 19561 26021 19737
rect 26055 19561 26067 19737
rect 26009 19549 26067 19561
rect 26127 19737 26185 19749
rect 26127 19561 26139 19737
rect 26173 19561 26185 19737
rect 26127 19549 26185 19561
rect 26245 19737 26303 19749
rect 26245 19561 26257 19737
rect 26291 19561 26303 19737
rect 26245 19549 26303 19561
rect 26468 19737 26526 19749
rect 26468 19561 26480 19737
rect 26514 19561 26526 19737
rect 26468 19549 26526 19561
rect 26586 19737 26644 19749
rect 26586 19561 26598 19737
rect 26632 19561 26644 19737
rect 26586 19549 26644 19561
rect 26704 19737 26762 19749
rect 26704 19561 26716 19737
rect 26750 19561 26762 19737
rect 26704 19549 26762 19561
rect 26822 19737 26880 19749
rect 26822 19561 26834 19737
rect 26868 19561 26880 19737
rect 26822 19549 26880 19561
rect 26951 19561 26963 19937
rect 26997 19561 27009 19937
rect 26951 19549 27009 19561
rect 27069 19937 27127 19949
rect 27069 19561 27081 19937
rect 27115 19561 27127 19937
rect 27069 19549 27127 19561
rect 27187 19937 27245 19949
rect 27187 19561 27199 19937
rect 27233 19561 27245 19937
rect 27187 19549 27245 19561
rect 27305 19937 27363 19949
rect 27305 19561 27317 19937
rect 27351 19561 27363 19937
rect 27305 19549 27363 19561
rect 27423 19937 27481 19949
rect 27423 19561 27435 19937
rect 27469 19561 27481 19937
rect 27423 19549 27481 19561
rect 27541 19937 27599 19949
rect 27541 19561 27553 19937
rect 27587 19561 27599 19937
rect 27541 19549 27599 19561
rect 27659 19937 27717 19949
rect 27659 19561 27671 19937
rect 27705 19561 27717 19937
rect 36755 20151 37155 20163
rect 36755 20117 36767 20151
rect 37143 20117 37155 20151
rect 36755 20105 37155 20117
rect 36755 20033 37155 20045
rect 36755 19999 36767 20033
rect 37143 19999 37155 20033
rect 36755 19987 37155 19999
rect 27659 19549 27717 19561
rect 27789 19737 27847 19749
rect 27789 19561 27801 19737
rect 27835 19561 27847 19737
rect 27789 19549 27847 19561
rect 27907 19737 27965 19749
rect 27907 19561 27919 19737
rect 27953 19561 27965 19737
rect 27907 19549 27965 19561
rect 28025 19737 28083 19749
rect 28025 19561 28037 19737
rect 28071 19561 28083 19737
rect 28025 19549 28083 19561
rect 28143 19737 28201 19749
rect 28143 19561 28155 19737
rect 28189 19561 28201 19737
rect 28143 19549 28201 19561
rect 20495 19241 20553 19253
rect 20495 18865 20507 19241
rect 20541 18865 20553 19241
rect 20495 18853 20553 18865
rect 20613 19241 20671 19253
rect 20613 18865 20625 19241
rect 20659 18865 20671 19241
rect 20613 18853 20671 18865
rect 20731 19241 20789 19253
rect 20731 18865 20743 19241
rect 20777 18865 20789 19241
rect 20731 18853 20789 18865
rect 20849 19241 20907 19253
rect 20849 18865 20861 19241
rect 20895 18865 20907 19241
rect 20849 18853 20907 18865
rect 20967 19241 21025 19253
rect 20967 18865 20979 19241
rect 21013 18865 21025 19241
rect 20967 18853 21025 18865
rect 21085 19241 21143 19253
rect 21085 18865 21097 19241
rect 21131 18865 21143 19241
rect 21085 18853 21143 18865
rect 21203 19241 21261 19253
rect 21203 18865 21215 19241
rect 21249 18865 21261 19241
rect 21203 18853 21261 18865
rect 22037 18747 22095 18759
rect 22037 18571 22049 18747
rect 22083 18571 22095 18747
rect 22037 18559 22095 18571
rect 22155 18747 22213 18759
rect 22155 18571 22167 18747
rect 22201 18571 22213 18747
rect 22155 18559 22213 18571
rect 22273 18747 22331 18759
rect 22273 18571 22285 18747
rect 22319 18571 22331 18747
rect 22273 18559 22331 18571
rect 22391 18747 22449 18759
rect 22391 18571 22403 18747
rect 22437 18571 22449 18747
rect 22391 18559 22449 18571
rect 22509 18747 22567 18759
rect 22509 18571 22521 18747
rect 22555 18571 22567 18747
rect 22509 18559 22567 18571
rect 22627 18747 22685 18759
rect 22627 18571 22639 18747
rect 22673 18571 22685 18747
rect 22627 18559 22685 18571
rect 22745 18747 22803 18759
rect 22745 18571 22757 18747
rect 22791 18571 22803 18747
rect 22745 18559 22803 18571
rect 22863 18747 22921 18759
rect 22863 18571 22875 18747
rect 22909 18571 22921 18747
rect 22863 18559 22921 18571
rect 22981 18747 23039 18759
rect 22981 18571 22993 18747
rect 23027 18571 23039 18747
rect 22981 18559 23039 18571
rect 23099 18747 23157 18759
rect 23099 18571 23111 18747
rect 23145 18571 23157 18747
rect 23099 18559 23157 18571
rect 25110 19244 25168 19256
rect 25110 18868 25122 19244
rect 25156 18868 25168 19244
rect 25110 18856 25168 18868
rect 25228 19244 25286 19256
rect 25228 18868 25240 19244
rect 25274 18868 25286 19244
rect 25228 18856 25286 18868
rect 25346 19244 25404 19256
rect 25346 18868 25358 19244
rect 25392 18868 25404 19244
rect 25346 18856 25404 18868
rect 25464 19244 25522 19256
rect 25464 18868 25476 19244
rect 25510 18868 25522 19244
rect 25464 18856 25522 18868
rect 25582 19244 25640 19256
rect 25582 18868 25594 19244
rect 25628 18868 25640 19244
rect 25582 18856 25640 18868
rect 25700 19244 25758 19256
rect 25700 18868 25712 19244
rect 25746 18868 25758 19244
rect 25700 18856 25758 18868
rect 25818 19244 25876 19256
rect 25818 18868 25830 19244
rect 25864 18868 25876 19244
rect 25818 18856 25876 18868
rect 36755 19915 37155 19927
rect 36755 19881 36767 19915
rect 37143 19881 37155 19915
rect 36755 19869 37155 19881
rect 36955 19796 37155 19808
rect 36955 19762 36967 19796
rect 37143 19762 37155 19796
rect 36955 19750 37155 19762
rect 36955 19678 37155 19690
rect 36955 19644 36967 19678
rect 37143 19644 37155 19678
rect 36955 19632 37155 19644
rect 36955 19560 37155 19572
rect 36955 19526 36967 19560
rect 37143 19526 37155 19560
rect 36955 19514 37155 19526
rect 36955 19442 37155 19454
rect 36955 19408 36967 19442
rect 37143 19408 37155 19442
rect 36955 19396 37155 19408
rect 27008 19244 27066 19256
rect 27008 18868 27020 19244
rect 27054 18868 27066 19244
rect 27008 18856 27066 18868
rect 27126 19244 27184 19256
rect 27126 18868 27138 19244
rect 27172 18868 27184 19244
rect 27126 18856 27184 18868
rect 27244 19244 27302 19256
rect 27244 18868 27256 19244
rect 27290 18868 27302 19244
rect 27244 18856 27302 18868
rect 27362 19244 27420 19256
rect 27362 18868 27374 19244
rect 27408 18868 27420 19244
rect 27362 18856 27420 18868
rect 27480 19244 27538 19256
rect 27480 18868 27492 19244
rect 27526 18868 27538 19244
rect 27480 18856 27538 18868
rect 27598 19244 27656 19256
rect 27598 18868 27610 19244
rect 27644 18868 27656 19244
rect 27598 18856 27656 18868
rect 27716 19244 27774 19256
rect 27716 18868 27728 19244
rect 27762 18868 27774 19244
rect 27716 18856 27774 18868
rect 36951 18872 37151 18884
rect 36951 18838 36963 18872
rect 37139 18838 37151 18872
rect 36951 18826 37151 18838
rect 28550 18750 28608 18762
rect 28550 18574 28562 18750
rect 28596 18574 28608 18750
rect 28550 18562 28608 18574
rect 28668 18750 28726 18762
rect 28668 18574 28680 18750
rect 28714 18574 28726 18750
rect 28668 18562 28726 18574
rect 28786 18750 28844 18762
rect 28786 18574 28798 18750
rect 28832 18574 28844 18750
rect 28786 18562 28844 18574
rect 28904 18750 28962 18762
rect 28904 18574 28916 18750
rect 28950 18574 28962 18750
rect 28904 18562 28962 18574
rect 29022 18750 29080 18762
rect 29022 18574 29034 18750
rect 29068 18574 29080 18750
rect 29022 18562 29080 18574
rect 29140 18750 29198 18762
rect 29140 18574 29152 18750
rect 29186 18574 29198 18750
rect 29140 18562 29198 18574
rect 29258 18750 29316 18762
rect 29258 18574 29270 18750
rect 29304 18574 29316 18750
rect 29258 18562 29316 18574
rect 29376 18750 29434 18762
rect 29376 18574 29388 18750
rect 29422 18574 29434 18750
rect 29376 18562 29434 18574
rect 29494 18750 29552 18762
rect 29494 18574 29506 18750
rect 29540 18574 29552 18750
rect 29494 18562 29552 18574
rect 29612 18750 29670 18762
rect 29612 18574 29624 18750
rect 29658 18574 29670 18750
rect 29612 18562 29670 18574
rect 36951 18754 37151 18766
rect 36951 18720 36963 18754
rect 37139 18720 37151 18754
rect 36951 18708 37151 18720
rect 36951 18636 37151 18648
rect 36951 18602 36963 18636
rect 37139 18602 37151 18636
rect 36951 18590 37151 18602
rect 36951 18518 37151 18530
rect 36951 18484 36963 18518
rect 37139 18484 37151 18518
rect 36951 18443 37151 18484
rect 36751 18431 37151 18443
rect 36751 18397 36763 18431
rect 37139 18397 37151 18431
rect 36751 18385 37151 18397
rect 36751 18313 37151 18325
rect 36751 18279 36763 18313
rect 37139 18279 37151 18313
rect 36751 18267 37151 18279
rect 36751 18195 37151 18207
rect 36751 18161 36763 18195
rect 37139 18161 37151 18195
rect 36751 18149 37151 18161
rect 36751 18077 37151 18089
rect 36751 18043 36763 18077
rect 37139 18043 37151 18077
rect 36751 18031 37151 18043
rect 36751 17964 37151 17976
rect 36751 17930 36763 17964
rect 37139 17930 37151 17964
rect 36751 17918 37151 17930
rect 36751 17846 37151 17858
rect 36751 17812 36763 17846
rect 37139 17812 37151 17846
rect 36751 17800 37151 17812
rect 36751 17728 37151 17740
rect 36751 17694 36763 17728
rect 37139 17694 37151 17728
rect 36751 17682 37151 17694
rect 36751 17610 37151 17622
rect 36751 17576 36763 17610
rect 37139 17576 37151 17610
rect 36751 17564 37151 17576
rect 36751 17492 37151 17504
rect 36751 17458 36763 17492
rect 37139 17458 37151 17492
rect 36751 17446 37151 17458
rect 36751 17374 37151 17386
rect 36751 17340 36763 17374
rect 37139 17340 37151 17374
rect 36751 17328 37151 17340
rect 36751 17256 37151 17268
rect 36751 17222 36763 17256
rect 37139 17222 37151 17256
rect 36751 17210 37151 17222
rect 36751 17137 37151 17149
rect 36751 17103 36763 17137
rect 37139 17103 37151 17137
rect 36751 17091 37151 17103
rect 36751 17019 37151 17031
rect 36751 16985 36763 17019
rect 37139 16985 37151 17019
rect 36751 16973 37151 16985
rect 36751 16901 37151 16913
rect 36751 16867 36763 16901
rect 37139 16867 37151 16901
rect 36751 16855 37151 16867
rect 36751 16783 37151 16795
rect 36751 16749 36763 16783
rect 37139 16749 37151 16783
rect 36751 16737 37151 16749
rect 36951 16664 37151 16676
rect 36951 16630 36963 16664
rect 37139 16630 37151 16664
rect 36951 16618 37151 16630
rect 36951 16546 37151 16558
rect 36951 16512 36963 16546
rect 37139 16512 37151 16546
rect 36951 16500 37151 16512
rect 36951 16428 37151 16440
rect 36951 16394 36963 16428
rect 37139 16394 37151 16428
rect 36951 16382 37151 16394
rect 36951 16310 37151 16322
rect 36951 16276 36963 16310
rect 37139 16276 37151 16310
rect -3604 16255 -3404 16267
rect 36951 16264 37151 16276
rect -3604 16221 -3592 16255
rect -3416 16221 -3404 16255
rect -3604 16209 -3404 16221
rect -3604 16137 -3404 16149
rect -3604 16103 -3592 16137
rect -3416 16103 -3404 16137
rect -3604 16091 -3404 16103
rect -3604 16019 -3404 16031
rect -3604 15985 -3592 16019
rect -3416 15985 -3404 16019
rect -3604 15973 -3404 15985
rect -3604 15901 -3404 15913
rect -3604 15867 -3592 15901
rect -3416 15867 -3404 15901
rect -3604 15855 -3404 15867
rect -3804 15771 -3404 15783
rect -3804 15737 -3792 15771
rect -3416 15737 -3404 15771
rect -3804 15725 -3404 15737
rect -3111 15828 -2711 15840
rect -3111 15794 -3099 15828
rect -2723 15794 -2711 15828
rect -3111 15782 -2711 15794
rect -3804 15653 -3404 15665
rect -3804 15619 -3792 15653
rect -3416 15619 -3404 15653
rect -3804 15607 -3404 15619
rect -3111 15710 -2711 15722
rect -3111 15676 -3099 15710
rect -2723 15676 -2711 15710
rect -3111 15664 -2711 15676
rect 36951 15728 37151 15740
rect 36951 15694 36963 15728
rect 37139 15694 37151 15728
rect 36951 15682 37151 15694
rect -3804 15535 -3404 15547
rect -3804 15501 -3792 15535
rect -3416 15501 -3404 15535
rect -3804 15489 -3404 15501
rect -3111 15592 -2711 15604
rect -3111 15558 -3099 15592
rect -2723 15558 -2711 15592
rect -3111 15546 -2711 15558
rect 36951 15610 37151 15622
rect 36951 15576 36963 15610
rect 37139 15576 37151 15610
rect 36951 15564 37151 15576
rect -3111 15474 -2711 15486
rect -3111 15440 -3099 15474
rect -2723 15440 -2711 15474
rect -3804 15417 -3404 15429
rect -3111 15428 -2711 15440
rect -3804 15383 -3792 15417
rect -3416 15383 -3404 15417
rect -3804 15371 -3404 15383
rect -3804 15299 -3404 15311
rect -3804 15265 -3792 15299
rect -3416 15265 -3404 15299
rect -3804 15253 -3404 15265
rect -3804 15181 -3404 15193
rect -3804 15147 -3792 15181
rect -3416 15147 -3404 15181
rect -3804 15135 -3404 15147
rect -3111 15356 -2711 15368
rect -3111 15322 -3099 15356
rect -2723 15322 -2711 15356
rect -3111 15310 -2711 15322
rect 36951 15492 37151 15504
rect 36951 15458 36963 15492
rect 37139 15458 37151 15492
rect 36951 15446 37151 15458
rect -3111 15238 -2711 15250
rect -3111 15204 -3099 15238
rect -2723 15204 -2711 15238
rect -3111 15192 -2711 15204
rect 7800 15224 7858 15236
rect -3804 15063 -3404 15075
rect -3804 15029 -3792 15063
rect -3416 15029 -3404 15063
rect -3804 15017 -3404 15029
rect -3604 14934 -3404 14946
rect -3604 14900 -3592 14934
rect -3416 14900 -3404 14934
rect -3604 14888 -3404 14900
rect -3111 15120 -2711 15132
rect -3111 15086 -3099 15120
rect -2723 15086 -2711 15120
rect -3111 15074 -2711 15086
rect 7800 15048 7812 15224
rect 7846 15048 7858 15224
rect 7800 15036 7858 15048
rect 7918 15224 7976 15236
rect 7918 15048 7930 15224
rect 7964 15048 7976 15224
rect 7918 15036 7976 15048
rect 8036 15224 8094 15236
rect 8036 15048 8048 15224
rect 8082 15048 8094 15224
rect 8036 15036 8094 15048
rect 8154 15224 8212 15236
rect 8154 15048 8166 15224
rect 8200 15048 8212 15224
rect 8154 15036 8212 15048
rect 8272 15224 8330 15236
rect 8272 15048 8284 15224
rect 8318 15048 8330 15224
rect 8272 15036 8330 15048
rect 8390 15224 8448 15236
rect 8390 15048 8402 15224
rect 8436 15048 8448 15224
rect 8390 15036 8448 15048
rect 8508 15224 8566 15236
rect 8508 15048 8520 15224
rect 8554 15048 8566 15224
rect 8508 15036 8566 15048
rect 8626 15224 8684 15236
rect 8626 15048 8638 15224
rect 8672 15048 8684 15224
rect 8626 15036 8684 15048
rect 8744 15224 8802 15236
rect 8744 15048 8756 15224
rect 8790 15048 8802 15224
rect 8744 15036 8802 15048
rect 8862 15224 8920 15236
rect 21003 15244 21061 15256
rect 8862 15048 8874 15224
rect 8908 15048 8920 15224
rect 8862 15036 8920 15048
rect 14349 15223 14407 15235
rect 14349 15047 14361 15223
rect 14395 15047 14407 15223
rect -3604 14816 -3404 14828
rect -3604 14782 -3592 14816
rect -3416 14782 -3404 14816
rect 14349 15035 14407 15047
rect 14467 15223 14525 15235
rect 14467 15047 14479 15223
rect 14513 15047 14525 15223
rect 14467 15035 14525 15047
rect 14585 15223 14643 15235
rect 14585 15047 14597 15223
rect 14631 15047 14643 15223
rect 14585 15035 14643 15047
rect 14703 15223 14761 15235
rect 14703 15047 14715 15223
rect 14749 15047 14761 15223
rect 14703 15035 14761 15047
rect 14821 15223 14879 15235
rect 14821 15047 14833 15223
rect 14867 15047 14879 15223
rect 14821 15035 14879 15047
rect 14939 15223 14997 15235
rect 14939 15047 14951 15223
rect 14985 15047 14997 15223
rect 14939 15035 14997 15047
rect 15057 15223 15115 15235
rect 15057 15047 15069 15223
rect 15103 15047 15115 15223
rect 15057 15035 15115 15047
rect 15175 15223 15233 15235
rect 15175 15047 15187 15223
rect 15221 15047 15233 15223
rect 15175 15035 15233 15047
rect 15293 15223 15351 15235
rect 15293 15047 15305 15223
rect 15339 15047 15351 15223
rect 15293 15035 15351 15047
rect 15411 15223 15469 15235
rect 15411 15047 15423 15223
rect 15457 15047 15469 15223
rect 21003 15068 21015 15244
rect 21049 15068 21061 15244
rect 21003 15056 21061 15068
rect 21121 15244 21179 15256
rect 21121 15068 21133 15244
rect 21167 15068 21179 15244
rect 21121 15056 21179 15068
rect 21239 15244 21297 15256
rect 21239 15068 21251 15244
rect 21285 15068 21297 15244
rect 21239 15056 21297 15068
rect 21357 15244 21415 15256
rect 21357 15068 21369 15244
rect 21403 15068 21415 15244
rect 21357 15056 21415 15068
rect 21475 15244 21533 15256
rect 21475 15068 21487 15244
rect 21521 15068 21533 15244
rect 21475 15056 21533 15068
rect 21593 15244 21651 15256
rect 21593 15068 21605 15244
rect 21639 15068 21651 15244
rect 21593 15056 21651 15068
rect 21711 15244 21769 15256
rect 21711 15068 21723 15244
rect 21757 15068 21769 15244
rect 21711 15056 21769 15068
rect 21829 15244 21887 15256
rect 21829 15068 21841 15244
rect 21875 15068 21887 15244
rect 21829 15056 21887 15068
rect 21947 15244 22005 15256
rect 21947 15068 21959 15244
rect 21993 15068 22005 15244
rect 21947 15056 22005 15068
rect 22065 15244 22123 15256
rect 22065 15068 22077 15244
rect 22111 15068 22123 15244
rect 36951 15374 37151 15386
rect 36951 15340 36963 15374
rect 37139 15340 37151 15374
rect 36951 15299 37151 15340
rect 36751 15287 37151 15299
rect 36751 15253 36763 15287
rect 37139 15253 37151 15287
rect 36751 15241 37151 15253
rect 36751 15169 37151 15181
rect 36751 15135 36763 15169
rect 37139 15135 37151 15169
rect 36751 15123 37151 15135
rect 22065 15056 22123 15068
rect 29656 15077 29714 15089
rect 15411 15035 15469 15047
rect -3604 14770 -3404 14782
rect -3604 14698 -3404 14710
rect -3604 14664 -3592 14698
rect -3416 14664 -3404 14698
rect -3604 14652 -3404 14664
rect -3604 14580 -3404 14592
rect -3604 14546 -3592 14580
rect -3416 14546 -3404 14580
rect -3604 14534 -3404 14546
rect 29656 14901 29668 15077
rect 29702 14901 29714 15077
rect 29656 14889 29714 14901
rect 29774 15077 29832 15089
rect 29774 14901 29786 15077
rect 29820 14901 29832 15077
rect 29774 14889 29832 14901
rect 29892 15077 29950 15089
rect 29892 14901 29904 15077
rect 29938 14901 29950 15077
rect 29892 14889 29950 14901
rect 30010 15077 30068 15089
rect 30010 14901 30022 15077
rect 30056 14901 30068 15077
rect 30010 14889 30068 14901
rect 30128 15077 30186 15089
rect 30128 14901 30140 15077
rect 30174 14901 30186 15077
rect 30128 14889 30186 14901
rect 30246 15077 30304 15089
rect 30246 14901 30258 15077
rect 30292 14901 30304 15077
rect 30246 14889 30304 14901
rect 30364 15077 30422 15089
rect 30364 14901 30376 15077
rect 30410 14901 30422 15077
rect 30364 14889 30422 14901
rect 30482 15077 30540 15089
rect 30482 14901 30494 15077
rect 30528 14901 30540 15077
rect 30482 14889 30540 14901
rect 30600 15077 30658 15089
rect 30600 14901 30612 15077
rect 30646 14901 30658 15077
rect 30600 14889 30658 14901
rect 30718 15077 30776 15089
rect 30718 14901 30730 15077
rect 30764 14901 30776 15077
rect 36751 15051 37151 15063
rect 36751 15017 36763 15051
rect 37139 15017 37151 15051
rect 36751 15005 37151 15017
rect 30718 14889 30776 14901
rect 31948 14872 32006 14884
rect 31464 14672 31522 14684
rect -3606 14187 -3406 14199
rect -3606 14153 -3594 14187
rect -3418 14153 -3406 14187
rect -3606 14141 -3406 14153
rect 31464 14496 31476 14672
rect 31510 14496 31522 14672
rect 31464 14484 31522 14496
rect 31582 14672 31640 14684
rect 31582 14496 31594 14672
rect 31628 14496 31640 14672
rect 31582 14484 31640 14496
rect 31700 14672 31758 14684
rect 31700 14496 31712 14672
rect 31746 14496 31758 14672
rect 31700 14484 31758 14496
rect 31818 14672 31876 14684
rect 31818 14496 31830 14672
rect 31864 14496 31876 14672
rect 31818 14484 31876 14496
rect 31948 14496 31960 14872
rect 31994 14496 32006 14872
rect 31948 14484 32006 14496
rect 32066 14872 32124 14884
rect 32066 14496 32078 14872
rect 32112 14496 32124 14872
rect 32066 14484 32124 14496
rect 32184 14872 32242 14884
rect 32184 14496 32196 14872
rect 32230 14496 32242 14872
rect 32184 14484 32242 14496
rect 32302 14872 32360 14884
rect 32302 14496 32314 14872
rect 32348 14496 32360 14872
rect 32302 14484 32360 14496
rect 32420 14872 32478 14884
rect 32420 14496 32432 14872
rect 32466 14496 32478 14872
rect 32420 14484 32478 14496
rect 32538 14872 32596 14884
rect 32538 14496 32550 14872
rect 32584 14496 32596 14872
rect 32538 14484 32596 14496
rect 32656 14872 32714 14884
rect 32656 14496 32668 14872
rect 32702 14496 32714 14872
rect 36751 14933 37151 14945
rect 36751 14899 36763 14933
rect 37139 14899 37151 14933
rect 36751 14887 37151 14899
rect 36751 14820 37151 14832
rect 36751 14786 36763 14820
rect 37139 14786 37151 14820
rect 36751 14774 37151 14786
rect 32656 14484 32714 14496
rect 32785 14672 32843 14684
rect 32785 14496 32797 14672
rect 32831 14496 32843 14672
rect 32785 14484 32843 14496
rect 32903 14672 32961 14684
rect 32903 14496 32915 14672
rect 32949 14496 32961 14672
rect 32903 14484 32961 14496
rect 33021 14672 33079 14684
rect 33021 14496 33033 14672
rect 33067 14496 33079 14672
rect 33021 14484 33079 14496
rect 33139 14672 33197 14684
rect 33139 14496 33151 14672
rect 33185 14496 33197 14672
rect 33139 14484 33197 14496
rect 33257 14669 33315 14681
rect 33257 14493 33269 14669
rect 33303 14493 33315 14669
rect 33257 14481 33315 14493
rect 33375 14669 33433 14681
rect 33375 14493 33387 14669
rect 33421 14493 33433 14669
rect 33375 14481 33433 14493
rect 33493 14669 33551 14681
rect 33493 14493 33505 14669
rect 33539 14493 33551 14669
rect 33493 14481 33551 14493
rect 33611 14669 33669 14681
rect 33611 14493 33623 14669
rect 33657 14493 33669 14669
rect 33611 14481 33669 14493
rect 33729 14669 33787 14681
rect 33729 14493 33741 14669
rect 33775 14493 33787 14669
rect 33729 14481 33787 14493
rect 33847 14669 33905 14681
rect 33847 14493 33859 14669
rect 33893 14493 33905 14669
rect 33847 14481 33905 14493
rect 33965 14669 34023 14681
rect 33965 14493 33977 14669
rect 34011 14493 34023 14669
rect 33965 14481 34023 14493
rect 34083 14669 34141 14681
rect 34083 14493 34095 14669
rect 34129 14493 34141 14669
rect 34083 14481 34141 14493
rect 34201 14669 34259 14681
rect 34201 14493 34213 14669
rect 34247 14493 34259 14669
rect 34201 14481 34259 14493
rect 34319 14669 34377 14681
rect 34319 14493 34331 14669
rect 34365 14493 34377 14669
rect 36751 14702 37151 14714
rect 36751 14668 36763 14702
rect 37139 14668 37151 14702
rect 36751 14656 37151 14668
rect 34319 14481 34377 14493
rect -3606 14069 -3406 14081
rect -3606 14035 -3594 14069
rect -3418 14035 -3406 14069
rect -3606 14023 -3406 14035
rect 31891 14179 31949 14191
rect -3606 13951 -3406 13963
rect -3606 13917 -3594 13951
rect -3418 13917 -3406 13951
rect -3606 13905 -3406 13917
rect -3606 13833 -3406 13845
rect -3606 13799 -3594 13833
rect -3418 13799 -3406 13833
rect -3606 13787 -3406 13799
rect -3806 13703 -3406 13715
rect -3806 13669 -3794 13703
rect -3418 13669 -3406 13703
rect -3806 13657 -3406 13669
rect -3113 13760 -2713 13772
rect -3113 13726 -3101 13760
rect -2725 13726 -2713 13760
rect -3113 13714 -2713 13726
rect -3806 13585 -3406 13597
rect -3806 13551 -3794 13585
rect -3418 13551 -3406 13585
rect -3806 13539 -3406 13551
rect -3113 13642 -2713 13654
rect -3113 13608 -3101 13642
rect -2725 13608 -2713 13642
rect -3113 13596 -2713 13608
rect -3806 13467 -3406 13479
rect -3806 13433 -3794 13467
rect -3418 13433 -3406 13467
rect -3806 13421 -3406 13433
rect -3113 13524 -2713 13536
rect -3113 13490 -3101 13524
rect -2725 13490 -2713 13524
rect -3113 13478 -2713 13490
rect -3113 13406 -2713 13418
rect -3113 13372 -3101 13406
rect -2725 13372 -2713 13406
rect -3806 13349 -3406 13361
rect -3113 13360 -2713 13372
rect -3806 13315 -3794 13349
rect -3418 13315 -3406 13349
rect -3806 13303 -3406 13315
rect -3806 13231 -3406 13243
rect -3806 13197 -3794 13231
rect -3418 13197 -3406 13231
rect -3806 13185 -3406 13197
rect -3806 13113 -3406 13125
rect -3806 13079 -3794 13113
rect -3418 13079 -3406 13113
rect -3806 13067 -3406 13079
rect -3113 13288 -2713 13300
rect -3113 13254 -3101 13288
rect -2725 13254 -2713 13288
rect -3113 13242 -2713 13254
rect 1136 13324 1194 13336
rect -3113 13170 -2713 13182
rect -3113 13136 -3101 13170
rect -2725 13136 -2713 13170
rect -3113 13124 -2713 13136
rect 1136 13148 1148 13324
rect 1182 13148 1194 13324
rect 1136 13136 1194 13148
rect 1254 13324 1312 13336
rect 1254 13148 1266 13324
rect 1300 13148 1312 13324
rect 1254 13136 1312 13148
rect 1372 13324 1430 13336
rect 1372 13148 1384 13324
rect 1418 13148 1430 13324
rect 1372 13136 1430 13148
rect 1490 13324 1548 13336
rect 1490 13148 1502 13324
rect 1536 13148 1548 13324
rect 1490 13136 1548 13148
rect 1608 13324 1666 13336
rect 1608 13148 1620 13324
rect 1654 13148 1666 13324
rect 1608 13136 1666 13148
rect 1726 13324 1784 13336
rect 1726 13148 1738 13324
rect 1772 13148 1784 13324
rect 1726 13136 1784 13148
rect 1844 13324 1902 13336
rect 1844 13148 1856 13324
rect 1890 13148 1902 13324
rect 1844 13136 1902 13148
rect 1962 13324 2020 13336
rect 1962 13148 1974 13324
rect 2008 13148 2020 13324
rect 1962 13136 2020 13148
rect 2080 13324 2138 13336
rect 2080 13148 2092 13324
rect 2126 13148 2138 13324
rect 2080 13136 2138 13148
rect 2198 13324 2256 13336
rect 2198 13148 2210 13324
rect 2244 13148 2256 13324
rect 31891 13803 31903 14179
rect 31937 13803 31949 14179
rect 31891 13791 31949 13803
rect 32009 14179 32067 14191
rect 32009 13803 32021 14179
rect 32055 13803 32067 14179
rect 32009 13791 32067 13803
rect 32127 14179 32185 14191
rect 32127 13803 32139 14179
rect 32173 13803 32185 14179
rect 32127 13791 32185 13803
rect 32245 14179 32303 14191
rect 32245 13803 32257 14179
rect 32291 13803 32303 14179
rect 32245 13791 32303 13803
rect 32363 14179 32421 14191
rect 32363 13803 32375 14179
rect 32409 13803 32421 14179
rect 32363 13791 32421 13803
rect 32481 14179 32539 14191
rect 32481 13803 32493 14179
rect 32527 13803 32539 14179
rect 32481 13791 32539 13803
rect 32599 14179 32657 14191
rect 32599 13803 32611 14179
rect 32645 13803 32657 14179
rect 32599 13791 32657 13803
rect 36751 14584 37151 14596
rect 36751 14550 36763 14584
rect 37139 14550 37151 14584
rect 36751 14538 37151 14550
rect 36751 14466 37151 14478
rect 36751 14432 36763 14466
rect 37139 14432 37151 14466
rect 36751 14420 37151 14432
rect 36751 14348 37151 14360
rect 36751 14314 36763 14348
rect 37139 14314 37151 14348
rect 36751 14302 37151 14314
rect 36751 14230 37151 14242
rect 36751 14196 36763 14230
rect 37139 14196 37151 14230
rect 36751 14184 37151 14196
rect 36751 14112 37151 14124
rect 36751 14078 36763 14112
rect 37139 14078 37151 14112
rect 36751 14066 37151 14078
rect 36751 13993 37151 14005
rect 36751 13959 36763 13993
rect 37139 13959 37151 13993
rect 36751 13947 37151 13959
rect 36751 13875 37151 13887
rect 36751 13841 36763 13875
rect 37139 13841 37151 13875
rect 36751 13829 37151 13841
rect 36751 13757 37151 13769
rect 36751 13723 36763 13757
rect 37139 13723 37151 13757
rect 36751 13711 37151 13723
rect 36751 13639 37151 13651
rect 36751 13605 36763 13639
rect 37139 13605 37151 13639
rect 36751 13593 37151 13605
rect 36951 13520 37151 13532
rect 36951 13486 36963 13520
rect 37139 13486 37151 13520
rect 36951 13474 37151 13486
rect 12900 13217 12958 13229
rect 2198 13136 2256 13148
rect 10575 13145 10633 13157
rect -3806 12995 -3406 13007
rect -3806 12961 -3794 12995
rect -3418 12961 -3406 12995
rect -3806 12949 -3406 12961
rect -3606 12866 -3406 12878
rect -3606 12832 -3594 12866
rect -3418 12832 -3406 12866
rect -3606 12820 -3406 12832
rect -3113 13052 -2713 13064
rect -3113 13018 -3101 13052
rect -2725 13018 -2713 13052
rect -3113 13006 -2713 13018
rect 6351 13129 6409 13141
rect 4026 13057 4084 13069
rect -3606 12748 -3406 12760
rect -3606 12714 -3594 12748
rect -3418 12714 -3406 12748
rect -3606 12702 -3406 12714
rect -3606 12630 -3406 12642
rect -3606 12596 -3594 12630
rect -3418 12596 -3406 12630
rect -3606 12584 -3406 12596
rect -3606 12512 -3406 12524
rect -3606 12478 -3594 12512
rect -3418 12478 -3406 12512
rect 4026 12881 4038 13057
rect 4072 12881 4084 13057
rect 4026 12869 4084 12881
rect 4144 13057 4202 13069
rect 4144 12881 4156 13057
rect 4190 12881 4202 13057
rect 4144 12869 4202 12881
rect 4262 13057 4320 13069
rect 4262 12881 4274 13057
rect 4308 12881 4320 13057
rect 4262 12869 4320 12881
rect 4380 13057 4438 13069
rect 4380 12881 4392 13057
rect 4426 12881 4438 13057
rect 4380 12869 4438 12881
rect 4498 13057 4556 13069
rect 4498 12881 4510 13057
rect 4544 12881 4556 13057
rect 4498 12869 4556 12881
rect 4616 13057 4674 13069
rect 4616 12881 4628 13057
rect 4662 12881 4674 13057
rect 4616 12869 4674 12881
rect 4734 13057 4792 13069
rect 4734 12881 4746 13057
rect 4780 12881 4792 13057
rect 4734 12869 4792 12881
rect 4852 13057 4910 13069
rect 4852 12881 4864 13057
rect 4898 12881 4910 13057
rect 4852 12869 4910 12881
rect 4970 13057 5028 13069
rect 4970 12881 4982 13057
rect 5016 12881 5028 13057
rect 4970 12869 5028 12881
rect 5088 13057 5146 13069
rect 5088 12881 5100 13057
rect 5134 12881 5146 13057
rect 5088 12869 5146 12881
rect 6351 12753 6363 13129
rect 6397 12753 6409 13129
rect 6351 12741 6409 12753
rect 6469 13129 6527 13141
rect 6469 12753 6481 13129
rect 6515 12753 6527 13129
rect 6469 12741 6527 12753
rect 6587 13129 6645 13141
rect 6587 12753 6599 13129
rect 6633 12753 6645 13129
rect 6587 12741 6645 12753
rect 6705 13129 6763 13141
rect 6705 12753 6717 13129
rect 6751 12753 6763 13129
rect 6705 12741 6763 12753
rect 6823 13129 6881 13141
rect 6823 12753 6835 13129
rect 6869 12753 6881 13129
rect 6823 12741 6881 12753
rect 6941 13129 6999 13141
rect 6941 12753 6953 13129
rect 6987 12753 6999 13129
rect 6941 12741 6999 12753
rect 7059 13129 7117 13141
rect 7059 12753 7071 13129
rect 7105 12753 7117 13129
rect 7059 12741 7117 12753
rect 7493 13133 7551 13145
rect 7493 12757 7505 13133
rect 7539 12757 7551 13133
rect 7493 12745 7551 12757
rect 7611 13133 7669 13145
rect 7611 12757 7623 13133
rect 7657 12757 7669 13133
rect 7611 12745 7669 12757
rect 7729 13133 7787 13145
rect 7729 12757 7741 13133
rect 7775 12757 7787 13133
rect 7729 12745 7787 12757
rect 7847 13133 7905 13145
rect 7847 12757 7859 13133
rect 7893 12757 7905 13133
rect 7847 12745 7905 12757
rect 7965 13133 8023 13145
rect 7965 12757 7977 13133
rect 8011 12757 8023 13133
rect 7965 12745 8023 12757
rect 8083 13133 8141 13145
rect 8083 12757 8095 13133
rect 8129 12757 8141 13133
rect 8083 12745 8141 12757
rect 8201 13133 8259 13145
rect 8201 12757 8213 13133
rect 8247 12757 8259 13133
rect 10575 12969 10587 13145
rect 10621 12969 10633 13145
rect 10575 12957 10633 12969
rect 10693 13145 10751 13157
rect 10693 12969 10705 13145
rect 10739 12969 10751 13145
rect 10693 12957 10751 12969
rect 10811 13145 10869 13157
rect 10811 12969 10823 13145
rect 10857 12969 10869 13145
rect 10811 12957 10869 12969
rect 10929 13145 10987 13157
rect 10929 12969 10941 13145
rect 10975 12969 10987 13145
rect 10929 12957 10987 12969
rect 11047 13145 11105 13157
rect 11047 12969 11059 13145
rect 11093 12969 11105 13145
rect 11047 12957 11105 12969
rect 11165 13145 11223 13157
rect 11165 12969 11177 13145
rect 11211 12969 11223 13145
rect 11165 12957 11223 12969
rect 11283 13145 11341 13157
rect 11283 12969 11295 13145
rect 11329 12969 11341 13145
rect 11283 12957 11341 12969
rect 11401 13145 11459 13157
rect 11401 12969 11413 13145
rect 11447 12969 11459 13145
rect 11401 12957 11459 12969
rect 11519 13145 11577 13157
rect 11519 12969 11531 13145
rect 11565 12969 11577 13145
rect 11519 12957 11577 12969
rect 11637 13145 11695 13157
rect 11637 12969 11649 13145
rect 11683 12969 11695 13145
rect 11637 12957 11695 12969
rect 8201 12745 8259 12757
rect -3606 12466 -3406 12478
rect 12900 12841 12912 13217
rect 12946 12841 12958 13217
rect 12900 12829 12958 12841
rect 13018 13217 13076 13229
rect 13018 12841 13030 13217
rect 13064 12841 13076 13217
rect 13018 12829 13076 12841
rect 13136 13217 13194 13229
rect 13136 12841 13148 13217
rect 13182 12841 13194 13217
rect 13136 12829 13194 12841
rect 13254 13217 13312 13229
rect 13254 12841 13266 13217
rect 13300 12841 13312 13217
rect 13254 12829 13312 12841
rect 13372 13217 13430 13229
rect 13372 12841 13384 13217
rect 13418 12841 13430 13217
rect 13372 12829 13430 12841
rect 13490 13217 13548 13229
rect 13490 12841 13502 13217
rect 13536 12841 13548 13217
rect 13490 12829 13548 12841
rect 13608 13217 13666 13229
rect 13608 12841 13620 13217
rect 13654 12841 13666 13217
rect 13608 12829 13666 12841
rect 14042 13221 14100 13233
rect 14042 12845 14054 13221
rect 14088 12845 14100 13221
rect 14042 12833 14100 12845
rect 14160 13221 14218 13233
rect 14160 12845 14172 13221
rect 14206 12845 14218 13221
rect 14160 12833 14218 12845
rect 14278 13221 14336 13233
rect 14278 12845 14290 13221
rect 14324 12845 14336 13221
rect 14278 12833 14336 12845
rect 14396 13221 14454 13233
rect 14396 12845 14408 13221
rect 14442 12845 14454 13221
rect 14396 12833 14454 12845
rect 14514 13221 14572 13233
rect 14514 12845 14526 13221
rect 14560 12845 14572 13221
rect 14514 12833 14572 12845
rect 14632 13221 14690 13233
rect 14632 12845 14644 13221
rect 14678 12845 14690 13221
rect 14632 12833 14690 12845
rect 14750 13221 14808 13233
rect 14750 12845 14762 13221
rect 14796 12845 14808 13221
rect 26179 13217 26237 13229
rect 19554 13149 19612 13161
rect 17229 13077 17287 13089
rect 17229 12901 17241 13077
rect 17275 12901 17287 13077
rect 17229 12889 17287 12901
rect 17347 13077 17405 13089
rect 17347 12901 17359 13077
rect 17393 12901 17405 13077
rect 17347 12889 17405 12901
rect 17465 13077 17523 13089
rect 17465 12901 17477 13077
rect 17511 12901 17523 13077
rect 17465 12889 17523 12901
rect 17583 13077 17641 13089
rect 17583 12901 17595 13077
rect 17629 12901 17641 13077
rect 17583 12889 17641 12901
rect 17701 13077 17759 13089
rect 17701 12901 17713 13077
rect 17747 12901 17759 13077
rect 17701 12889 17759 12901
rect 17819 13077 17877 13089
rect 17819 12901 17831 13077
rect 17865 12901 17877 13077
rect 17819 12889 17877 12901
rect 17937 13077 17995 13089
rect 17937 12901 17949 13077
rect 17983 12901 17995 13077
rect 17937 12889 17995 12901
rect 18055 13077 18113 13089
rect 18055 12901 18067 13077
rect 18101 12901 18113 13077
rect 18055 12889 18113 12901
rect 18173 13077 18231 13089
rect 18173 12901 18185 13077
rect 18219 12901 18231 13077
rect 18173 12889 18231 12901
rect 18291 13077 18349 13089
rect 18291 12901 18303 13077
rect 18337 12901 18349 13077
rect 18291 12889 18349 12901
rect 14750 12833 14808 12845
rect 6780 12346 6838 12358
rect 6780 12170 6792 12346
rect 6826 12170 6838 12346
rect 6780 12158 6838 12170
rect 6898 12346 6956 12358
rect 6898 12170 6910 12346
rect 6944 12170 6956 12346
rect 6898 12158 6956 12170
rect 7016 12346 7074 12358
rect 7016 12170 7028 12346
rect 7062 12170 7074 12346
rect 7016 12158 7074 12170
rect 7134 12346 7192 12358
rect 7134 12170 7146 12346
rect 7180 12170 7192 12346
rect 7134 12158 7192 12170
rect 7922 12350 7980 12362
rect 7922 12174 7934 12350
rect 7968 12174 7980 12350
rect 7922 12162 7980 12174
rect 8040 12350 8098 12362
rect 8040 12174 8052 12350
rect 8086 12174 8098 12350
rect 8040 12162 8098 12174
rect 8158 12350 8216 12362
rect 8158 12174 8170 12350
rect 8204 12174 8216 12350
rect 8158 12162 8216 12174
rect 8276 12350 8334 12362
rect 8276 12174 8288 12350
rect 8322 12174 8334 12350
rect 19554 12773 19566 13149
rect 19600 12773 19612 13149
rect 19554 12761 19612 12773
rect 19672 13149 19730 13161
rect 19672 12773 19684 13149
rect 19718 12773 19730 13149
rect 19672 12761 19730 12773
rect 19790 13149 19848 13161
rect 19790 12773 19802 13149
rect 19836 12773 19848 13149
rect 19790 12761 19848 12773
rect 19908 13149 19966 13161
rect 19908 12773 19920 13149
rect 19954 12773 19966 13149
rect 19908 12761 19966 12773
rect 20026 13149 20084 13161
rect 20026 12773 20038 13149
rect 20072 12773 20084 13149
rect 20026 12761 20084 12773
rect 20144 13149 20202 13161
rect 20144 12773 20156 13149
rect 20190 12773 20202 13149
rect 20144 12761 20202 12773
rect 20262 13149 20320 13161
rect 20262 12773 20274 13149
rect 20308 12773 20320 13149
rect 20262 12761 20320 12773
rect 20696 13153 20754 13165
rect 20696 12777 20708 13153
rect 20742 12777 20754 13153
rect 20696 12765 20754 12777
rect 20814 13153 20872 13165
rect 20814 12777 20826 13153
rect 20860 12777 20872 13153
rect 20814 12765 20872 12777
rect 20932 13153 20990 13165
rect 20932 12777 20944 13153
rect 20978 12777 20990 13153
rect 20932 12765 20990 12777
rect 21050 13153 21108 13165
rect 21050 12777 21062 13153
rect 21096 12777 21108 13153
rect 21050 12765 21108 12777
rect 21168 13153 21226 13165
rect 21168 12777 21180 13153
rect 21214 12777 21226 13153
rect 21168 12765 21226 12777
rect 21286 13153 21344 13165
rect 21286 12777 21298 13153
rect 21332 12777 21344 13153
rect 21286 12765 21344 12777
rect 21404 13153 21462 13165
rect 21404 12777 21416 13153
rect 21450 12777 21462 13153
rect 23854 13145 23912 13157
rect 23854 12969 23866 13145
rect 23900 12969 23912 13145
rect 23854 12957 23912 12969
rect 23972 13145 24030 13157
rect 23972 12969 23984 13145
rect 24018 12969 24030 13145
rect 23972 12957 24030 12969
rect 24090 13145 24148 13157
rect 24090 12969 24102 13145
rect 24136 12969 24148 13145
rect 24090 12957 24148 12969
rect 24208 13145 24266 13157
rect 24208 12969 24220 13145
rect 24254 12969 24266 13145
rect 24208 12957 24266 12969
rect 24326 13145 24384 13157
rect 24326 12969 24338 13145
rect 24372 12969 24384 13145
rect 24326 12957 24384 12969
rect 24444 13145 24502 13157
rect 24444 12969 24456 13145
rect 24490 12969 24502 13145
rect 24444 12957 24502 12969
rect 24562 13145 24620 13157
rect 24562 12969 24574 13145
rect 24608 12969 24620 13145
rect 24562 12957 24620 12969
rect 24680 13145 24738 13157
rect 24680 12969 24692 13145
rect 24726 12969 24738 13145
rect 24680 12957 24738 12969
rect 24798 13145 24856 13157
rect 24798 12969 24810 13145
rect 24844 12969 24856 13145
rect 24798 12957 24856 12969
rect 24916 13145 24974 13157
rect 24916 12969 24928 13145
rect 24962 12969 24974 13145
rect 24916 12957 24974 12969
rect 21404 12765 21462 12777
rect 13329 12434 13387 12446
rect 13329 12258 13341 12434
rect 13375 12258 13387 12434
rect 13329 12246 13387 12258
rect 13447 12434 13505 12446
rect 13447 12258 13459 12434
rect 13493 12258 13505 12434
rect 13447 12246 13505 12258
rect 13565 12434 13623 12446
rect 13565 12258 13577 12434
rect 13611 12258 13623 12434
rect 13565 12246 13623 12258
rect 13683 12434 13741 12446
rect 13683 12258 13695 12434
rect 13729 12258 13741 12434
rect 13683 12246 13741 12258
rect 14471 12438 14529 12450
rect 14471 12262 14483 12438
rect 14517 12262 14529 12438
rect 14471 12250 14529 12262
rect 14589 12438 14647 12450
rect 14589 12262 14601 12438
rect 14635 12262 14647 12438
rect 14589 12250 14647 12262
rect 14707 12438 14765 12450
rect 14707 12262 14719 12438
rect 14753 12262 14765 12438
rect 14707 12250 14765 12262
rect 14825 12438 14883 12450
rect 14825 12262 14837 12438
rect 14871 12262 14883 12438
rect 14825 12250 14883 12262
rect 26179 12841 26191 13217
rect 26225 12841 26237 13217
rect 26179 12829 26237 12841
rect 26297 13217 26355 13229
rect 26297 12841 26309 13217
rect 26343 12841 26355 13217
rect 26297 12829 26355 12841
rect 26415 13217 26473 13229
rect 26415 12841 26427 13217
rect 26461 12841 26473 13217
rect 26415 12829 26473 12841
rect 26533 13217 26591 13229
rect 26533 12841 26545 13217
rect 26579 12841 26591 13217
rect 26533 12829 26591 12841
rect 26651 13217 26709 13229
rect 26651 12841 26663 13217
rect 26697 12841 26709 13217
rect 26651 12829 26709 12841
rect 26769 13217 26827 13229
rect 26769 12841 26781 13217
rect 26815 12841 26827 13217
rect 26769 12829 26827 12841
rect 26887 13217 26945 13229
rect 26887 12841 26899 13217
rect 26933 12841 26945 13217
rect 26887 12829 26945 12841
rect 27321 13221 27379 13233
rect 27321 12845 27333 13221
rect 27367 12845 27379 13221
rect 27321 12833 27379 12845
rect 27439 13221 27497 13233
rect 27439 12845 27451 13221
rect 27485 12845 27497 13221
rect 27439 12833 27497 12845
rect 27557 13221 27615 13233
rect 27557 12845 27569 13221
rect 27603 12845 27615 13221
rect 27557 12833 27615 12845
rect 27675 13221 27733 13233
rect 27675 12845 27687 13221
rect 27721 12845 27733 13221
rect 27675 12833 27733 12845
rect 27793 13221 27851 13233
rect 27793 12845 27805 13221
rect 27839 12845 27851 13221
rect 27793 12833 27851 12845
rect 27911 13221 27969 13233
rect 27911 12845 27923 13221
rect 27957 12845 27969 13221
rect 27911 12833 27969 12845
rect 28029 13221 28087 13233
rect 28029 12845 28041 13221
rect 28075 12845 28087 13221
rect 36951 13402 37151 13414
rect 36951 13368 36963 13402
rect 37139 13368 37151 13402
rect 36951 13356 37151 13368
rect 36951 13284 37151 13296
rect 36951 13250 36963 13284
rect 37139 13250 37151 13284
rect 36951 13238 37151 13250
rect 36951 13166 37151 13178
rect 36951 13132 36963 13166
rect 37139 13132 37151 13166
rect 36951 13120 37151 13132
rect 28029 12833 28087 12845
rect 8276 12162 8334 12174
rect 19983 12366 20041 12378
rect 19983 12190 19995 12366
rect 20029 12190 20041 12366
rect 19983 12178 20041 12190
rect 20101 12366 20159 12378
rect 20101 12190 20113 12366
rect 20147 12190 20159 12366
rect 20101 12178 20159 12190
rect 20219 12366 20277 12378
rect 20219 12190 20231 12366
rect 20265 12190 20277 12366
rect 20219 12178 20277 12190
rect 20337 12366 20395 12378
rect 20337 12190 20349 12366
rect 20383 12190 20395 12366
rect 20337 12178 20395 12190
rect 21125 12370 21183 12382
rect 21125 12194 21137 12370
rect 21171 12194 21183 12370
rect 21125 12182 21183 12194
rect 21243 12370 21301 12382
rect 21243 12194 21255 12370
rect 21289 12194 21301 12370
rect 21243 12182 21301 12194
rect 21361 12370 21419 12382
rect 21361 12194 21373 12370
rect 21407 12194 21419 12370
rect 21361 12182 21419 12194
rect 21479 12370 21537 12382
rect 21479 12194 21491 12370
rect 21525 12194 21537 12370
rect 36955 12526 37155 12538
rect 29651 12506 29709 12518
rect 26608 12434 26666 12446
rect 26608 12258 26620 12434
rect 26654 12258 26666 12434
rect 26608 12246 26666 12258
rect 26726 12434 26784 12446
rect 26726 12258 26738 12434
rect 26772 12258 26784 12434
rect 26726 12246 26784 12258
rect 26844 12434 26902 12446
rect 26844 12258 26856 12434
rect 26890 12258 26902 12434
rect 26844 12246 26902 12258
rect 26962 12434 27020 12446
rect 26962 12258 26974 12434
rect 27008 12258 27020 12434
rect 26962 12246 27020 12258
rect 27750 12438 27808 12450
rect 27750 12262 27762 12438
rect 27796 12262 27808 12438
rect 27750 12250 27808 12262
rect 27868 12438 27926 12450
rect 27868 12262 27880 12438
rect 27914 12262 27926 12438
rect 27868 12250 27926 12262
rect 27986 12438 28044 12450
rect 27986 12262 27998 12438
rect 28032 12262 28044 12438
rect 27986 12250 28044 12262
rect 28104 12438 28162 12450
rect 28104 12262 28116 12438
rect 28150 12262 28162 12438
rect 29651 12330 29663 12506
rect 29697 12330 29709 12506
rect 29651 12318 29709 12330
rect 29769 12506 29827 12518
rect 29769 12330 29781 12506
rect 29815 12330 29827 12506
rect 29769 12318 29827 12330
rect 29887 12506 29945 12518
rect 29887 12330 29899 12506
rect 29933 12330 29945 12506
rect 29887 12318 29945 12330
rect 30005 12506 30063 12518
rect 30005 12330 30017 12506
rect 30051 12330 30063 12506
rect 30005 12318 30063 12330
rect 30123 12506 30181 12518
rect 30123 12330 30135 12506
rect 30169 12330 30181 12506
rect 30123 12318 30181 12330
rect 30241 12506 30299 12518
rect 30241 12330 30253 12506
rect 30287 12330 30299 12506
rect 30241 12318 30299 12330
rect 30359 12506 30417 12518
rect 30359 12330 30371 12506
rect 30405 12330 30417 12506
rect 30359 12318 30417 12330
rect 30477 12506 30535 12518
rect 30477 12330 30489 12506
rect 30523 12330 30535 12506
rect 30477 12318 30535 12330
rect 30595 12506 30653 12518
rect 30595 12330 30607 12506
rect 30641 12330 30653 12506
rect 30595 12318 30653 12330
rect 30713 12506 30771 12518
rect 30713 12330 30725 12506
rect 30759 12330 30771 12506
rect 36955 12492 36967 12526
rect 37143 12492 37155 12526
rect 36955 12480 37155 12492
rect 30713 12318 30771 12330
rect 36955 12408 37155 12420
rect 36955 12374 36967 12408
rect 37143 12374 37155 12408
rect 36955 12362 37155 12374
rect 28104 12250 28162 12262
rect 21479 12182 21537 12194
rect -3604 12118 -3404 12130
rect -3604 12084 -3592 12118
rect -3416 12084 -3404 12118
rect -3604 12072 -3404 12084
rect -3604 12000 -3404 12012
rect -3604 11966 -3592 12000
rect -3416 11966 -3404 12000
rect -3604 11954 -3404 11966
rect 36955 12290 37155 12302
rect 36955 12256 36967 12290
rect 37143 12256 37155 12290
rect 36955 12244 37155 12256
rect 36955 12172 37155 12184
rect 36955 12138 36967 12172
rect 37143 12138 37155 12172
rect 36955 12097 37155 12138
rect 36755 12085 37155 12097
rect -3604 11882 -3404 11894
rect -3604 11848 -3592 11882
rect -3416 11848 -3404 11882
rect -3604 11836 -3404 11848
rect -3604 11764 -3404 11776
rect -3604 11730 -3592 11764
rect -3416 11730 -3404 11764
rect -3604 11718 -3404 11730
rect -3804 11634 -3404 11646
rect -3804 11600 -3792 11634
rect -3416 11600 -3404 11634
rect -3804 11588 -3404 11600
rect -3111 11691 -2711 11703
rect -3111 11657 -3099 11691
rect -2723 11657 -2711 11691
rect -3111 11645 -2711 11657
rect -3804 11516 -3404 11528
rect -3804 11482 -3792 11516
rect -3416 11482 -3404 11516
rect -3804 11470 -3404 11482
rect -3111 11573 -2711 11585
rect -3111 11539 -3099 11573
rect -2723 11539 -2711 11573
rect -3111 11527 -2711 11539
rect 36755 12051 36767 12085
rect 37143 12051 37155 12085
rect 36755 12039 37155 12051
rect 36755 11967 37155 11979
rect 36755 11933 36767 11967
rect 37143 11933 37155 11967
rect 36755 11921 37155 11933
rect 36755 11849 37155 11861
rect 36755 11815 36767 11849
rect 37143 11815 37155 11849
rect 36755 11803 37155 11815
rect 36755 11731 37155 11743
rect 36755 11697 36767 11731
rect 37143 11697 37155 11731
rect 36755 11685 37155 11697
rect -3804 11398 -3404 11410
rect -3804 11364 -3792 11398
rect -3416 11364 -3404 11398
rect -3804 11352 -3404 11364
rect -3111 11455 -2711 11467
rect -3111 11421 -3099 11455
rect -2723 11421 -2711 11455
rect -3111 11409 -2711 11421
rect -3111 11337 -2711 11349
rect -3111 11303 -3099 11337
rect -2723 11303 -2711 11337
rect -3804 11280 -3404 11292
rect -3111 11291 -2711 11303
rect -3804 11246 -3792 11280
rect -3416 11246 -3404 11280
rect -3804 11234 -3404 11246
rect -3804 11162 -3404 11174
rect -3804 11128 -3792 11162
rect -3416 11128 -3404 11162
rect -3804 11116 -3404 11128
rect -3804 11044 -3404 11056
rect -3804 11010 -3792 11044
rect -3416 11010 -3404 11044
rect -3804 10998 -3404 11010
rect -3111 11219 -2711 11231
rect -3111 11185 -3099 11219
rect -2723 11185 -2711 11219
rect -3111 11173 -2711 11185
rect 4040 11407 4098 11419
rect 4040 11231 4052 11407
rect 4086 11231 4098 11407
rect 4040 11219 4098 11231
rect 4158 11407 4216 11419
rect 4158 11231 4170 11407
rect 4204 11231 4216 11407
rect 4158 11219 4216 11231
rect 4276 11407 4334 11419
rect 4276 11231 4288 11407
rect 4322 11231 4334 11407
rect 4276 11219 4334 11231
rect 4394 11407 4452 11419
rect 4394 11231 4406 11407
rect 4440 11231 4452 11407
rect 4394 11219 4452 11231
rect 4512 11407 4570 11419
rect 4512 11231 4524 11407
rect 4558 11231 4570 11407
rect 4512 11219 4570 11231
rect 4630 11407 4688 11419
rect 4630 11231 4642 11407
rect 4676 11231 4688 11407
rect 4630 11219 4688 11231
rect 4748 11407 4806 11419
rect 4748 11231 4760 11407
rect 4794 11231 4806 11407
rect 4748 11219 4806 11231
rect 4866 11407 4924 11419
rect 4866 11231 4878 11407
rect 4912 11231 4924 11407
rect 4866 11219 4924 11231
rect 4984 11407 5042 11419
rect 4984 11231 4996 11407
rect 5030 11231 5042 11407
rect 4984 11219 5042 11231
rect 5102 11407 5160 11419
rect 5102 11231 5114 11407
rect 5148 11231 5160 11407
rect 10589 11495 10647 11507
rect 10589 11319 10601 11495
rect 10635 11319 10647 11495
rect 10589 11307 10647 11319
rect 10707 11495 10765 11507
rect 10707 11319 10719 11495
rect 10753 11319 10765 11495
rect 10707 11307 10765 11319
rect 10825 11495 10883 11507
rect 10825 11319 10837 11495
rect 10871 11319 10883 11495
rect 10825 11307 10883 11319
rect 10943 11495 11001 11507
rect 10943 11319 10955 11495
rect 10989 11319 11001 11495
rect 10943 11307 11001 11319
rect 11061 11495 11119 11507
rect 11061 11319 11073 11495
rect 11107 11319 11119 11495
rect 11061 11307 11119 11319
rect 11179 11495 11237 11507
rect 11179 11319 11191 11495
rect 11225 11319 11237 11495
rect 11179 11307 11237 11319
rect 11297 11495 11355 11507
rect 11297 11319 11309 11495
rect 11343 11319 11355 11495
rect 11297 11307 11355 11319
rect 11415 11495 11473 11507
rect 11415 11319 11427 11495
rect 11461 11319 11473 11495
rect 11415 11307 11473 11319
rect 11533 11495 11591 11507
rect 11533 11319 11545 11495
rect 11579 11319 11591 11495
rect 11533 11307 11591 11319
rect 11651 11495 11709 11507
rect 11651 11319 11663 11495
rect 11697 11319 11709 11495
rect 36755 11618 37155 11630
rect 36755 11584 36767 11618
rect 37143 11584 37155 11618
rect 36755 11572 37155 11584
rect 17243 11427 17301 11439
rect 11651 11307 11709 11319
rect 5102 11219 5160 11231
rect -3111 11101 -2711 11113
rect -3111 11067 -3099 11101
rect -2723 11067 -2711 11101
rect -3111 11055 -2711 11067
rect -3804 10926 -3404 10938
rect -3804 10892 -3792 10926
rect -3416 10892 -3404 10926
rect -3804 10880 -3404 10892
rect -3604 10797 -3404 10809
rect -3604 10763 -3592 10797
rect -3416 10763 -3404 10797
rect -3604 10751 -3404 10763
rect -3111 10983 -2711 10995
rect -3111 10949 -3099 10983
rect -2723 10949 -2711 10983
rect 17243 11251 17255 11427
rect 17289 11251 17301 11427
rect 17243 11239 17301 11251
rect 17361 11427 17419 11439
rect 17361 11251 17373 11427
rect 17407 11251 17419 11427
rect 17361 11239 17419 11251
rect 17479 11427 17537 11439
rect 17479 11251 17491 11427
rect 17525 11251 17537 11427
rect 17479 11239 17537 11251
rect 17597 11427 17655 11439
rect 17597 11251 17609 11427
rect 17643 11251 17655 11427
rect 17597 11239 17655 11251
rect 17715 11427 17773 11439
rect 17715 11251 17727 11427
rect 17761 11251 17773 11427
rect 17715 11239 17773 11251
rect 17833 11427 17891 11439
rect 17833 11251 17845 11427
rect 17879 11251 17891 11427
rect 17833 11239 17891 11251
rect 17951 11427 18009 11439
rect 17951 11251 17963 11427
rect 17997 11251 18009 11427
rect 17951 11239 18009 11251
rect 18069 11427 18127 11439
rect 18069 11251 18081 11427
rect 18115 11251 18127 11427
rect 18069 11239 18127 11251
rect 18187 11427 18245 11439
rect 18187 11251 18199 11427
rect 18233 11251 18245 11427
rect 18187 11239 18245 11251
rect 18305 11427 18363 11439
rect 18305 11251 18317 11427
rect 18351 11251 18363 11427
rect 23868 11495 23926 11507
rect 23868 11319 23880 11495
rect 23914 11319 23926 11495
rect 23868 11307 23926 11319
rect 23986 11495 24044 11507
rect 23986 11319 23998 11495
rect 24032 11319 24044 11495
rect 23986 11307 24044 11319
rect 24104 11495 24162 11507
rect 24104 11319 24116 11495
rect 24150 11319 24162 11495
rect 24104 11307 24162 11319
rect 24222 11495 24280 11507
rect 24222 11319 24234 11495
rect 24268 11319 24280 11495
rect 24222 11307 24280 11319
rect 24340 11495 24398 11507
rect 24340 11319 24352 11495
rect 24386 11319 24398 11495
rect 24340 11307 24398 11319
rect 24458 11495 24516 11507
rect 24458 11319 24470 11495
rect 24504 11319 24516 11495
rect 24458 11307 24516 11319
rect 24576 11495 24634 11507
rect 24576 11319 24588 11495
rect 24622 11319 24634 11495
rect 24576 11307 24634 11319
rect 24694 11495 24752 11507
rect 24694 11319 24706 11495
rect 24740 11319 24752 11495
rect 24694 11307 24752 11319
rect 24812 11495 24870 11507
rect 24812 11319 24824 11495
rect 24858 11319 24870 11495
rect 24812 11307 24870 11319
rect 24930 11495 24988 11507
rect 24930 11319 24942 11495
rect 24976 11319 24988 11495
rect 36755 11500 37155 11512
rect 36755 11466 36767 11500
rect 37143 11466 37155 11500
rect 36755 11454 37155 11466
rect 24930 11307 24988 11319
rect 18305 11239 18363 11251
rect 12537 11078 12595 11090
rect 5988 10990 6046 11002
rect -3111 10937 -2711 10949
rect 1128 10739 1186 10751
rect -3604 10679 -3404 10691
rect -3604 10645 -3592 10679
rect -3416 10645 -3404 10679
rect -3604 10633 -3404 10645
rect -3604 10561 -3404 10573
rect -3604 10527 -3592 10561
rect -3416 10527 -3404 10561
rect 1128 10563 1140 10739
rect 1174 10563 1186 10739
rect 1128 10551 1186 10563
rect 1246 10739 1304 10751
rect 1246 10563 1258 10739
rect 1292 10563 1304 10739
rect 1246 10551 1304 10563
rect 1364 10739 1422 10751
rect 1364 10563 1376 10739
rect 1410 10563 1422 10739
rect 1364 10551 1422 10563
rect 1482 10739 1540 10751
rect 1482 10563 1494 10739
rect 1528 10563 1540 10739
rect 1482 10551 1540 10563
rect 1600 10739 1658 10751
rect 1600 10563 1612 10739
rect 1646 10563 1658 10739
rect 1600 10551 1658 10563
rect 1718 10739 1776 10751
rect 1718 10563 1730 10739
rect 1764 10563 1776 10739
rect 1718 10551 1776 10563
rect 1836 10739 1894 10751
rect 1836 10563 1848 10739
rect 1882 10563 1894 10739
rect 1836 10551 1894 10563
rect 1954 10739 2012 10751
rect 1954 10563 1966 10739
rect 2000 10563 2012 10739
rect 1954 10551 2012 10563
rect 2072 10739 2130 10751
rect 2072 10563 2084 10739
rect 2118 10563 2130 10739
rect 2072 10551 2130 10563
rect 2190 10739 2248 10751
rect 2190 10563 2202 10739
rect 2236 10563 2248 10739
rect 5504 10790 5562 10802
rect 2190 10551 2248 10563
rect -3604 10515 -3404 10527
rect -3604 10443 -3404 10455
rect -3604 10409 -3592 10443
rect -3416 10409 -3404 10443
rect -3604 10397 -3404 10409
rect 5504 10614 5516 10790
rect 5550 10614 5562 10790
rect 5504 10602 5562 10614
rect 5622 10790 5680 10802
rect 5622 10614 5634 10790
rect 5668 10614 5680 10790
rect 5622 10602 5680 10614
rect 5740 10790 5798 10802
rect 5740 10614 5752 10790
rect 5786 10614 5798 10790
rect 5740 10602 5798 10614
rect 5858 10790 5916 10802
rect 5858 10614 5870 10790
rect 5904 10614 5916 10790
rect 5858 10602 5916 10614
rect 5988 10614 6000 10990
rect 6034 10614 6046 10990
rect 5988 10602 6046 10614
rect 6106 10990 6164 11002
rect 6106 10614 6118 10990
rect 6152 10614 6164 10990
rect 6106 10602 6164 10614
rect 6224 10990 6282 11002
rect 6224 10614 6236 10990
rect 6270 10614 6282 10990
rect 6224 10602 6282 10614
rect 6342 10990 6400 11002
rect 6342 10614 6354 10990
rect 6388 10614 6400 10990
rect 6342 10602 6400 10614
rect 6460 10990 6518 11002
rect 6460 10614 6472 10990
rect 6506 10614 6518 10990
rect 6460 10602 6518 10614
rect 6578 10990 6636 11002
rect 6578 10614 6590 10990
rect 6624 10614 6636 10990
rect 6578 10602 6636 10614
rect 6696 10990 6754 11002
rect 6696 10614 6708 10990
rect 6742 10614 6754 10990
rect 7886 10990 7944 11002
rect 6696 10602 6754 10614
rect 6825 10790 6883 10802
rect 6825 10614 6837 10790
rect 6871 10614 6883 10790
rect 6825 10602 6883 10614
rect 6943 10790 7001 10802
rect 6943 10614 6955 10790
rect 6989 10614 7001 10790
rect 6943 10602 7001 10614
rect 7061 10790 7119 10802
rect 7061 10614 7073 10790
rect 7107 10614 7119 10790
rect 7061 10602 7119 10614
rect 7179 10790 7237 10802
rect 7179 10614 7191 10790
rect 7225 10614 7237 10790
rect 7179 10602 7237 10614
rect 7402 10790 7460 10802
rect 7402 10614 7414 10790
rect 7448 10614 7460 10790
rect 7402 10602 7460 10614
rect 7520 10790 7578 10802
rect 7520 10614 7532 10790
rect 7566 10614 7578 10790
rect 7520 10602 7578 10614
rect 7638 10790 7696 10802
rect 7638 10614 7650 10790
rect 7684 10614 7696 10790
rect 7638 10602 7696 10614
rect 7756 10790 7814 10802
rect 7756 10614 7768 10790
rect 7802 10614 7814 10790
rect 7756 10602 7814 10614
rect 7886 10614 7898 10990
rect 7932 10614 7944 10990
rect 7886 10602 7944 10614
rect 8004 10990 8062 11002
rect 8004 10614 8016 10990
rect 8050 10614 8062 10990
rect 8004 10602 8062 10614
rect 8122 10990 8180 11002
rect 8122 10614 8134 10990
rect 8168 10614 8180 10990
rect 8122 10602 8180 10614
rect 8240 10990 8298 11002
rect 8240 10614 8252 10990
rect 8286 10614 8298 10990
rect 8240 10602 8298 10614
rect 8358 10990 8416 11002
rect 8358 10614 8370 10990
rect 8404 10614 8416 10990
rect 8358 10602 8416 10614
rect 8476 10990 8534 11002
rect 8476 10614 8488 10990
rect 8522 10614 8534 10990
rect 8476 10602 8534 10614
rect 8594 10990 8652 11002
rect 8594 10614 8606 10990
rect 8640 10614 8652 10990
rect 8594 10602 8652 10614
rect 8723 10790 8781 10802
rect 8723 10614 8735 10790
rect 8769 10614 8781 10790
rect 8723 10602 8781 10614
rect 8841 10790 8899 10802
rect 8841 10614 8853 10790
rect 8887 10614 8899 10790
rect 8841 10602 8899 10614
rect 8959 10790 9017 10802
rect 8959 10614 8971 10790
rect 9005 10614 9017 10790
rect 8959 10602 9017 10614
rect 9077 10790 9135 10802
rect 9077 10614 9089 10790
rect 9123 10614 9135 10790
rect 12053 10878 12111 10890
rect 9077 10602 9135 10614
rect -3606 10050 -3406 10062
rect -3606 10016 -3594 10050
rect -3418 10016 -3406 10050
rect -3606 10004 -3406 10016
rect -3606 9932 -3406 9944
rect -3606 9898 -3594 9932
rect -3418 9898 -3406 9932
rect -3606 9886 -3406 9898
rect -3606 9814 -3406 9826
rect -3606 9780 -3594 9814
rect -3418 9780 -3406 9814
rect -3606 9768 -3406 9780
rect 4035 9803 4093 9815
rect -3606 9696 -3406 9708
rect -3606 9662 -3594 9696
rect -3418 9662 -3406 9696
rect -3606 9650 -3406 9662
rect -3806 9566 -3406 9578
rect -3806 9532 -3794 9566
rect -3418 9532 -3406 9566
rect -3806 9520 -3406 9532
rect -3113 9623 -2713 9635
rect -3113 9589 -3101 9623
rect -2725 9589 -2713 9623
rect 4035 9627 4047 9803
rect 4081 9627 4093 9803
rect 4035 9615 4093 9627
rect 4153 9803 4211 9815
rect 4153 9627 4165 9803
rect 4199 9627 4211 9803
rect 4153 9615 4211 9627
rect 4271 9803 4329 9815
rect 4271 9627 4283 9803
rect 4317 9627 4329 9803
rect 4271 9615 4329 9627
rect 4389 9803 4447 9815
rect 4389 9627 4401 9803
rect 4435 9627 4447 9803
rect 4389 9615 4447 9627
rect 4507 9803 4565 9815
rect 4507 9627 4519 9803
rect 4553 9627 4565 9803
rect 4507 9615 4565 9627
rect 4625 9803 4683 9815
rect 4625 9627 4637 9803
rect 4671 9627 4683 9803
rect 4625 9615 4683 9627
rect 4743 9803 4801 9815
rect 4743 9627 4755 9803
rect 4789 9627 4801 9803
rect 4743 9615 4801 9627
rect 4861 9803 4919 9815
rect 4861 9627 4873 9803
rect 4907 9627 4919 9803
rect 4861 9615 4919 9627
rect 4979 9803 5037 9815
rect 4979 9627 4991 9803
rect 5025 9627 5037 9803
rect 4979 9615 5037 9627
rect 5097 9803 5155 9815
rect 5097 9627 5109 9803
rect 5143 9627 5155 9803
rect 5097 9615 5155 9627
rect 5931 10297 5989 10309
rect 5931 9921 5943 10297
rect 5977 9921 5989 10297
rect 5931 9909 5989 9921
rect 6049 10297 6107 10309
rect 6049 9921 6061 10297
rect 6095 9921 6107 10297
rect 6049 9909 6107 9921
rect 6167 10297 6225 10309
rect 6167 9921 6179 10297
rect 6213 9921 6225 10297
rect 6167 9909 6225 9921
rect 6285 10297 6343 10309
rect 6285 9921 6297 10297
rect 6331 9921 6343 10297
rect 6285 9909 6343 9921
rect 6403 10297 6461 10309
rect 6403 9921 6415 10297
rect 6449 9921 6461 10297
rect 6403 9909 6461 9921
rect 6521 10297 6579 10309
rect 6521 9921 6533 10297
rect 6567 9921 6579 10297
rect 6521 9909 6579 9921
rect 6639 10297 6697 10309
rect 6639 9921 6651 10297
rect 6685 9921 6697 10297
rect 6639 9909 6697 9921
rect -3113 9577 -2713 9589
rect -3806 9448 -3406 9460
rect -3806 9414 -3794 9448
rect -3418 9414 -3406 9448
rect -3806 9402 -3406 9414
rect -3113 9505 -2713 9517
rect -3113 9471 -3101 9505
rect -2725 9471 -2713 9505
rect -3113 9459 -2713 9471
rect -3806 9330 -3406 9342
rect -3806 9296 -3794 9330
rect -3418 9296 -3406 9330
rect -3806 9284 -3406 9296
rect -3113 9387 -2713 9399
rect -3113 9353 -3101 9387
rect -2725 9353 -2713 9387
rect -3113 9341 -2713 9353
rect 12053 10702 12065 10878
rect 12099 10702 12111 10878
rect 12053 10690 12111 10702
rect 12171 10878 12229 10890
rect 12171 10702 12183 10878
rect 12217 10702 12229 10878
rect 12171 10690 12229 10702
rect 12289 10878 12347 10890
rect 12289 10702 12301 10878
rect 12335 10702 12347 10878
rect 12289 10690 12347 10702
rect 12407 10878 12465 10890
rect 12407 10702 12419 10878
rect 12453 10702 12465 10878
rect 12407 10690 12465 10702
rect 12537 10702 12549 11078
rect 12583 10702 12595 11078
rect 12537 10690 12595 10702
rect 12655 11078 12713 11090
rect 12655 10702 12667 11078
rect 12701 10702 12713 11078
rect 12655 10690 12713 10702
rect 12773 11078 12831 11090
rect 12773 10702 12785 11078
rect 12819 10702 12831 11078
rect 12773 10690 12831 10702
rect 12891 11078 12949 11090
rect 12891 10702 12903 11078
rect 12937 10702 12949 11078
rect 12891 10690 12949 10702
rect 13009 11078 13067 11090
rect 13009 10702 13021 11078
rect 13055 10702 13067 11078
rect 13009 10690 13067 10702
rect 13127 11078 13185 11090
rect 13127 10702 13139 11078
rect 13173 10702 13185 11078
rect 13127 10690 13185 10702
rect 13245 11078 13303 11090
rect 13245 10702 13257 11078
rect 13291 10702 13303 11078
rect 14435 11078 14493 11090
rect 13245 10690 13303 10702
rect 13374 10878 13432 10890
rect 13374 10702 13386 10878
rect 13420 10702 13432 10878
rect 13374 10690 13432 10702
rect 13492 10878 13550 10890
rect 13492 10702 13504 10878
rect 13538 10702 13550 10878
rect 13492 10690 13550 10702
rect 13610 10878 13668 10890
rect 13610 10702 13622 10878
rect 13656 10702 13668 10878
rect 13610 10690 13668 10702
rect 13728 10878 13786 10890
rect 13728 10702 13740 10878
rect 13774 10702 13786 10878
rect 13728 10690 13786 10702
rect 13951 10878 14009 10890
rect 13951 10702 13963 10878
rect 13997 10702 14009 10878
rect 13951 10690 14009 10702
rect 14069 10878 14127 10890
rect 14069 10702 14081 10878
rect 14115 10702 14127 10878
rect 14069 10690 14127 10702
rect 14187 10878 14245 10890
rect 14187 10702 14199 10878
rect 14233 10702 14245 10878
rect 14187 10690 14245 10702
rect 14305 10878 14363 10890
rect 14305 10702 14317 10878
rect 14351 10702 14363 10878
rect 14305 10690 14363 10702
rect 14435 10702 14447 11078
rect 14481 10702 14493 11078
rect 14435 10690 14493 10702
rect 14553 11078 14611 11090
rect 14553 10702 14565 11078
rect 14599 10702 14611 11078
rect 14553 10690 14611 10702
rect 14671 11078 14729 11090
rect 14671 10702 14683 11078
rect 14717 10702 14729 11078
rect 14671 10690 14729 10702
rect 14789 11078 14847 11090
rect 14789 10702 14801 11078
rect 14835 10702 14847 11078
rect 14789 10690 14847 10702
rect 14907 11078 14965 11090
rect 14907 10702 14919 11078
rect 14953 10702 14965 11078
rect 14907 10690 14965 10702
rect 15025 11078 15083 11090
rect 15025 10702 15037 11078
rect 15071 10702 15083 11078
rect 15025 10690 15083 10702
rect 15143 11078 15201 11090
rect 15143 10702 15155 11078
rect 15189 10702 15201 11078
rect 36755 11382 37155 11394
rect 36755 11348 36767 11382
rect 37143 11348 37155 11382
rect 36755 11336 37155 11348
rect 36755 11264 37155 11276
rect 36755 11230 36767 11264
rect 37143 11230 37155 11264
rect 36755 11218 37155 11230
rect 36755 11146 37155 11158
rect 36755 11112 36767 11146
rect 37143 11112 37155 11146
rect 36755 11100 37155 11112
rect 25816 11078 25874 11090
rect 19191 11010 19249 11022
rect 15143 10690 15201 10702
rect 15272 10878 15330 10890
rect 15272 10702 15284 10878
rect 15318 10702 15330 10878
rect 15272 10690 15330 10702
rect 15390 10878 15448 10890
rect 15390 10702 15402 10878
rect 15436 10702 15448 10878
rect 15390 10690 15448 10702
rect 15508 10878 15566 10890
rect 15508 10702 15520 10878
rect 15554 10702 15566 10878
rect 15508 10690 15566 10702
rect 15626 10878 15684 10890
rect 15626 10702 15638 10878
rect 15672 10702 15684 10878
rect 15626 10690 15684 10702
rect 7829 10297 7887 10309
rect 7829 9921 7841 10297
rect 7875 9921 7887 10297
rect 7829 9909 7887 9921
rect 7947 10297 8005 10309
rect 7947 9921 7959 10297
rect 7993 9921 8005 10297
rect 7947 9909 8005 9921
rect 8065 10297 8123 10309
rect 8065 9921 8077 10297
rect 8111 9921 8123 10297
rect 8065 9909 8123 9921
rect 8183 10297 8241 10309
rect 8183 9921 8195 10297
rect 8229 9921 8241 10297
rect 8183 9909 8241 9921
rect 8301 10297 8359 10309
rect 8301 9921 8313 10297
rect 8347 9921 8359 10297
rect 8301 9909 8359 9921
rect 8419 10297 8477 10309
rect 8419 9921 8431 10297
rect 8465 9921 8477 10297
rect 8419 9909 8477 9921
rect 8537 10297 8595 10309
rect 8537 9921 8549 10297
rect 8583 9921 8595 10297
rect 8537 9909 8595 9921
rect 10584 9891 10642 9903
rect 10584 9715 10596 9891
rect 10630 9715 10642 9891
rect 10584 9703 10642 9715
rect 10702 9891 10760 9903
rect 10702 9715 10714 9891
rect 10748 9715 10760 9891
rect 10702 9703 10760 9715
rect 10820 9891 10878 9903
rect 10820 9715 10832 9891
rect 10866 9715 10878 9891
rect 10820 9703 10878 9715
rect 10938 9891 10996 9903
rect 10938 9715 10950 9891
rect 10984 9715 10996 9891
rect 10938 9703 10996 9715
rect 11056 9891 11114 9903
rect 11056 9715 11068 9891
rect 11102 9715 11114 9891
rect 11056 9703 11114 9715
rect 11174 9891 11232 9903
rect 11174 9715 11186 9891
rect 11220 9715 11232 9891
rect 11174 9703 11232 9715
rect 11292 9891 11350 9903
rect 11292 9715 11304 9891
rect 11338 9715 11350 9891
rect 11292 9703 11350 9715
rect 11410 9891 11468 9903
rect 11410 9715 11422 9891
rect 11456 9715 11468 9891
rect 11410 9703 11468 9715
rect 11528 9891 11586 9903
rect 11528 9715 11540 9891
rect 11574 9715 11586 9891
rect 11528 9703 11586 9715
rect 11646 9891 11704 9903
rect 11646 9715 11658 9891
rect 11692 9715 11704 9891
rect 11646 9703 11704 9715
rect 12480 10385 12538 10397
rect 12480 10009 12492 10385
rect 12526 10009 12538 10385
rect 12480 9997 12538 10009
rect 12598 10385 12656 10397
rect 12598 10009 12610 10385
rect 12644 10009 12656 10385
rect 12598 9997 12656 10009
rect 12716 10385 12774 10397
rect 12716 10009 12728 10385
rect 12762 10009 12774 10385
rect 12716 9997 12774 10009
rect 12834 10385 12892 10397
rect 12834 10009 12846 10385
rect 12880 10009 12892 10385
rect 12834 9997 12892 10009
rect 12952 10385 13010 10397
rect 12952 10009 12964 10385
rect 12998 10009 13010 10385
rect 12952 9997 13010 10009
rect 13070 10385 13128 10397
rect 13070 10009 13082 10385
rect 13116 10009 13128 10385
rect 13070 9997 13128 10009
rect 13188 10385 13246 10397
rect 13188 10009 13200 10385
rect 13234 10009 13246 10385
rect 13188 9997 13246 10009
rect -3113 9269 -2713 9281
rect -3113 9235 -3101 9269
rect -2725 9235 -2713 9269
rect -3806 9212 -3406 9224
rect -3113 9223 -2713 9235
rect -3806 9178 -3794 9212
rect -3418 9178 -3406 9212
rect -3806 9166 -3406 9178
rect -3806 9094 -3406 9106
rect -3806 9060 -3794 9094
rect -3418 9060 -3406 9094
rect -3806 9048 -3406 9060
rect -3806 8976 -3406 8988
rect -3806 8942 -3794 8976
rect -3418 8942 -3406 8976
rect -3806 8930 -3406 8942
rect -3113 9151 -2713 9163
rect -3113 9117 -3101 9151
rect -2725 9117 -2713 9151
rect -3113 9105 -2713 9117
rect -3113 9033 -2713 9045
rect -3113 8999 -3101 9033
rect -2725 8999 -2713 9033
rect -3113 8987 -2713 8999
rect 18707 10810 18765 10822
rect 18707 10634 18719 10810
rect 18753 10634 18765 10810
rect 18707 10622 18765 10634
rect 18825 10810 18883 10822
rect 18825 10634 18837 10810
rect 18871 10634 18883 10810
rect 18825 10622 18883 10634
rect 18943 10810 19001 10822
rect 18943 10634 18955 10810
rect 18989 10634 19001 10810
rect 18943 10622 19001 10634
rect 19061 10810 19119 10822
rect 19061 10634 19073 10810
rect 19107 10634 19119 10810
rect 19061 10622 19119 10634
rect 19191 10634 19203 11010
rect 19237 10634 19249 11010
rect 19191 10622 19249 10634
rect 19309 11010 19367 11022
rect 19309 10634 19321 11010
rect 19355 10634 19367 11010
rect 19309 10622 19367 10634
rect 19427 11010 19485 11022
rect 19427 10634 19439 11010
rect 19473 10634 19485 11010
rect 19427 10622 19485 10634
rect 19545 11010 19603 11022
rect 19545 10634 19557 11010
rect 19591 10634 19603 11010
rect 19545 10622 19603 10634
rect 19663 11010 19721 11022
rect 19663 10634 19675 11010
rect 19709 10634 19721 11010
rect 19663 10622 19721 10634
rect 19781 11010 19839 11022
rect 19781 10634 19793 11010
rect 19827 10634 19839 11010
rect 19781 10622 19839 10634
rect 19899 11010 19957 11022
rect 19899 10634 19911 11010
rect 19945 10634 19957 11010
rect 21089 11010 21147 11022
rect 19899 10622 19957 10634
rect 20028 10810 20086 10822
rect 20028 10634 20040 10810
rect 20074 10634 20086 10810
rect 20028 10622 20086 10634
rect 20146 10810 20204 10822
rect 20146 10634 20158 10810
rect 20192 10634 20204 10810
rect 20146 10622 20204 10634
rect 20264 10810 20322 10822
rect 20264 10634 20276 10810
rect 20310 10634 20322 10810
rect 20264 10622 20322 10634
rect 20382 10810 20440 10822
rect 20382 10634 20394 10810
rect 20428 10634 20440 10810
rect 20382 10622 20440 10634
rect 20605 10810 20663 10822
rect 20605 10634 20617 10810
rect 20651 10634 20663 10810
rect 20605 10622 20663 10634
rect 20723 10810 20781 10822
rect 20723 10634 20735 10810
rect 20769 10634 20781 10810
rect 20723 10622 20781 10634
rect 20841 10810 20899 10822
rect 20841 10634 20853 10810
rect 20887 10634 20899 10810
rect 20841 10622 20899 10634
rect 20959 10810 21017 10822
rect 20959 10634 20971 10810
rect 21005 10634 21017 10810
rect 20959 10622 21017 10634
rect 21089 10634 21101 11010
rect 21135 10634 21147 11010
rect 21089 10622 21147 10634
rect 21207 11010 21265 11022
rect 21207 10634 21219 11010
rect 21253 10634 21265 11010
rect 21207 10622 21265 10634
rect 21325 11010 21383 11022
rect 21325 10634 21337 11010
rect 21371 10634 21383 11010
rect 21325 10622 21383 10634
rect 21443 11010 21501 11022
rect 21443 10634 21455 11010
rect 21489 10634 21501 11010
rect 21443 10622 21501 10634
rect 21561 11010 21619 11022
rect 21561 10634 21573 11010
rect 21607 10634 21619 11010
rect 21561 10622 21619 10634
rect 21679 11010 21737 11022
rect 21679 10634 21691 11010
rect 21725 10634 21737 11010
rect 21679 10622 21737 10634
rect 21797 11010 21855 11022
rect 21797 10634 21809 11010
rect 21843 10634 21855 11010
rect 21797 10622 21855 10634
rect 21926 10810 21984 10822
rect 21926 10634 21938 10810
rect 21972 10634 21984 10810
rect 21926 10622 21984 10634
rect 22044 10810 22102 10822
rect 22044 10634 22056 10810
rect 22090 10634 22102 10810
rect 22044 10622 22102 10634
rect 22162 10810 22220 10822
rect 22162 10634 22174 10810
rect 22208 10634 22220 10810
rect 22162 10622 22220 10634
rect 22280 10810 22338 10822
rect 22280 10634 22292 10810
rect 22326 10634 22338 10810
rect 25332 10878 25390 10890
rect 22280 10622 22338 10634
rect 14378 10385 14436 10397
rect 14378 10009 14390 10385
rect 14424 10009 14436 10385
rect 14378 9997 14436 10009
rect 14496 10385 14554 10397
rect 14496 10009 14508 10385
rect 14542 10009 14554 10385
rect 14496 9997 14554 10009
rect 14614 10385 14672 10397
rect 14614 10009 14626 10385
rect 14660 10009 14672 10385
rect 14614 9997 14672 10009
rect 14732 10385 14790 10397
rect 14732 10009 14744 10385
rect 14778 10009 14790 10385
rect 14732 9997 14790 10009
rect 14850 10385 14908 10397
rect 14850 10009 14862 10385
rect 14896 10009 14908 10385
rect 14850 9997 14908 10009
rect 14968 10385 15026 10397
rect 14968 10009 14980 10385
rect 15014 10009 15026 10385
rect 14968 9997 15026 10009
rect 15086 10385 15144 10397
rect 15086 10009 15098 10385
rect 15132 10009 15144 10385
rect 15086 9997 15144 10009
rect 17238 9823 17296 9835
rect 17238 9647 17250 9823
rect 17284 9647 17296 9823
rect 17238 9635 17296 9647
rect 17356 9823 17414 9835
rect 17356 9647 17368 9823
rect 17402 9647 17414 9823
rect 17356 9635 17414 9647
rect 17474 9823 17532 9835
rect 17474 9647 17486 9823
rect 17520 9647 17532 9823
rect 17474 9635 17532 9647
rect 17592 9823 17650 9835
rect 17592 9647 17604 9823
rect 17638 9647 17650 9823
rect 17592 9635 17650 9647
rect 17710 9823 17768 9835
rect 17710 9647 17722 9823
rect 17756 9647 17768 9823
rect 17710 9635 17768 9647
rect 17828 9823 17886 9835
rect 17828 9647 17840 9823
rect 17874 9647 17886 9823
rect 17828 9635 17886 9647
rect 17946 9823 18004 9835
rect 17946 9647 17958 9823
rect 17992 9647 18004 9823
rect 17946 9635 18004 9647
rect 18064 9823 18122 9835
rect 18064 9647 18076 9823
rect 18110 9647 18122 9823
rect 18064 9635 18122 9647
rect 18182 9823 18240 9835
rect 18182 9647 18194 9823
rect 18228 9647 18240 9823
rect 18182 9635 18240 9647
rect 18300 9823 18358 9835
rect 18300 9647 18312 9823
rect 18346 9647 18358 9823
rect 18300 9635 18358 9647
rect 19134 10317 19192 10329
rect 19134 9941 19146 10317
rect 19180 9941 19192 10317
rect 19134 9929 19192 9941
rect 19252 10317 19310 10329
rect 19252 9941 19264 10317
rect 19298 9941 19310 10317
rect 19252 9929 19310 9941
rect 19370 10317 19428 10329
rect 19370 9941 19382 10317
rect 19416 9941 19428 10317
rect 19370 9929 19428 9941
rect 19488 10317 19546 10329
rect 19488 9941 19500 10317
rect 19534 9941 19546 10317
rect 19488 9929 19546 9941
rect 19606 10317 19664 10329
rect 19606 9941 19618 10317
rect 19652 9941 19664 10317
rect 19606 9929 19664 9941
rect 19724 10317 19782 10329
rect 19724 9941 19736 10317
rect 19770 9941 19782 10317
rect 19724 9929 19782 9941
rect 19842 10317 19900 10329
rect 19842 9941 19854 10317
rect 19888 9941 19900 10317
rect 19842 9929 19900 9941
rect 25332 10702 25344 10878
rect 25378 10702 25390 10878
rect 25332 10690 25390 10702
rect 25450 10878 25508 10890
rect 25450 10702 25462 10878
rect 25496 10702 25508 10878
rect 25450 10690 25508 10702
rect 25568 10878 25626 10890
rect 25568 10702 25580 10878
rect 25614 10702 25626 10878
rect 25568 10690 25626 10702
rect 25686 10878 25744 10890
rect 25686 10702 25698 10878
rect 25732 10702 25744 10878
rect 25686 10690 25744 10702
rect 25816 10702 25828 11078
rect 25862 10702 25874 11078
rect 25816 10690 25874 10702
rect 25934 11078 25992 11090
rect 25934 10702 25946 11078
rect 25980 10702 25992 11078
rect 25934 10690 25992 10702
rect 26052 11078 26110 11090
rect 26052 10702 26064 11078
rect 26098 10702 26110 11078
rect 26052 10690 26110 10702
rect 26170 11078 26228 11090
rect 26170 10702 26182 11078
rect 26216 10702 26228 11078
rect 26170 10690 26228 10702
rect 26288 11078 26346 11090
rect 26288 10702 26300 11078
rect 26334 10702 26346 11078
rect 26288 10690 26346 10702
rect 26406 11078 26464 11090
rect 26406 10702 26418 11078
rect 26452 10702 26464 11078
rect 26406 10690 26464 10702
rect 26524 11078 26582 11090
rect 26524 10702 26536 11078
rect 26570 10702 26582 11078
rect 27714 11078 27772 11090
rect 26524 10690 26582 10702
rect 26653 10878 26711 10890
rect 26653 10702 26665 10878
rect 26699 10702 26711 10878
rect 26653 10690 26711 10702
rect 26771 10878 26829 10890
rect 26771 10702 26783 10878
rect 26817 10702 26829 10878
rect 26771 10690 26829 10702
rect 26889 10878 26947 10890
rect 26889 10702 26901 10878
rect 26935 10702 26947 10878
rect 26889 10690 26947 10702
rect 27007 10878 27065 10890
rect 27007 10702 27019 10878
rect 27053 10702 27065 10878
rect 27007 10690 27065 10702
rect 27230 10878 27288 10890
rect 27230 10702 27242 10878
rect 27276 10702 27288 10878
rect 27230 10690 27288 10702
rect 27348 10878 27406 10890
rect 27348 10702 27360 10878
rect 27394 10702 27406 10878
rect 27348 10690 27406 10702
rect 27466 10878 27524 10890
rect 27466 10702 27478 10878
rect 27512 10702 27524 10878
rect 27466 10690 27524 10702
rect 27584 10878 27642 10890
rect 27584 10702 27596 10878
rect 27630 10702 27642 10878
rect 27584 10690 27642 10702
rect 27714 10702 27726 11078
rect 27760 10702 27772 11078
rect 27714 10690 27772 10702
rect 27832 11078 27890 11090
rect 27832 10702 27844 11078
rect 27878 10702 27890 11078
rect 27832 10690 27890 10702
rect 27950 11078 28008 11090
rect 27950 10702 27962 11078
rect 27996 10702 28008 11078
rect 27950 10690 28008 10702
rect 28068 11078 28126 11090
rect 28068 10702 28080 11078
rect 28114 10702 28126 11078
rect 28068 10690 28126 10702
rect 28186 11078 28244 11090
rect 28186 10702 28198 11078
rect 28232 10702 28244 11078
rect 28186 10690 28244 10702
rect 28304 11078 28362 11090
rect 28304 10702 28316 11078
rect 28350 10702 28362 11078
rect 28304 10690 28362 10702
rect 28422 11078 28480 11090
rect 28422 10702 28434 11078
rect 28468 10702 28480 11078
rect 36755 11028 37155 11040
rect 36755 10994 36767 11028
rect 37143 10994 37155 11028
rect 36755 10982 37155 10994
rect 36755 10910 37155 10922
rect 28422 10690 28480 10702
rect 28551 10878 28609 10890
rect 28551 10702 28563 10878
rect 28597 10702 28609 10878
rect 28551 10690 28609 10702
rect 28669 10878 28727 10890
rect 28669 10702 28681 10878
rect 28715 10702 28727 10878
rect 28669 10690 28727 10702
rect 28787 10878 28845 10890
rect 28787 10702 28799 10878
rect 28833 10702 28845 10878
rect 28787 10690 28845 10702
rect 28905 10878 28963 10890
rect 28905 10702 28917 10878
rect 28951 10702 28963 10878
rect 36755 10876 36767 10910
rect 37143 10876 37155 10910
rect 36755 10864 37155 10876
rect 28905 10690 28963 10702
rect 31950 10781 32008 10793
rect 21032 10317 21090 10329
rect 21032 9941 21044 10317
rect 21078 9941 21090 10317
rect 21032 9929 21090 9941
rect 21150 10317 21208 10329
rect 21150 9941 21162 10317
rect 21196 9941 21208 10317
rect 21150 9929 21208 9941
rect 21268 10317 21326 10329
rect 21268 9941 21280 10317
rect 21314 9941 21326 10317
rect 21268 9929 21326 9941
rect 21386 10317 21444 10329
rect 21386 9941 21398 10317
rect 21432 9941 21444 10317
rect 21386 9929 21444 9941
rect 21504 10317 21562 10329
rect 21504 9941 21516 10317
rect 21550 9941 21562 10317
rect 21504 9929 21562 9941
rect 21622 10317 21680 10329
rect 21622 9941 21634 10317
rect 21668 9941 21680 10317
rect 21622 9929 21680 9941
rect 21740 10317 21798 10329
rect 21740 9941 21752 10317
rect 21786 9941 21798 10317
rect 21740 9929 21798 9941
rect 23863 9891 23921 9903
rect 23863 9715 23875 9891
rect 23909 9715 23921 9891
rect 23863 9703 23921 9715
rect 23981 9891 24039 9903
rect 23981 9715 23993 9891
rect 24027 9715 24039 9891
rect 23981 9703 24039 9715
rect 24099 9891 24157 9903
rect 24099 9715 24111 9891
rect 24145 9715 24157 9891
rect 24099 9703 24157 9715
rect 24217 9891 24275 9903
rect 24217 9715 24229 9891
rect 24263 9715 24275 9891
rect 24217 9703 24275 9715
rect 24335 9891 24393 9903
rect 24335 9715 24347 9891
rect 24381 9715 24393 9891
rect 24335 9703 24393 9715
rect 24453 9891 24511 9903
rect 24453 9715 24465 9891
rect 24499 9715 24511 9891
rect 24453 9703 24511 9715
rect 24571 9891 24629 9903
rect 24571 9715 24583 9891
rect 24617 9715 24629 9891
rect 24571 9703 24629 9715
rect 24689 9891 24747 9903
rect 24689 9715 24701 9891
rect 24735 9715 24747 9891
rect 24689 9703 24747 9715
rect 24807 9891 24865 9903
rect 24807 9715 24819 9891
rect 24853 9715 24865 9891
rect 24807 9703 24865 9715
rect 24925 9891 24983 9903
rect 24925 9715 24937 9891
rect 24971 9715 24983 9891
rect 24925 9703 24983 9715
rect 25759 10385 25817 10397
rect 25759 10009 25771 10385
rect 25805 10009 25817 10385
rect 25759 9997 25817 10009
rect 25877 10385 25935 10397
rect 25877 10009 25889 10385
rect 25923 10009 25935 10385
rect 25877 9997 25935 10009
rect 25995 10385 26053 10397
rect 25995 10009 26007 10385
rect 26041 10009 26053 10385
rect 25995 9997 26053 10009
rect 26113 10385 26171 10397
rect 26113 10009 26125 10385
rect 26159 10009 26171 10385
rect 26113 9997 26171 10009
rect 26231 10385 26289 10397
rect 26231 10009 26243 10385
rect 26277 10009 26289 10385
rect 26231 9997 26289 10009
rect 26349 10385 26407 10397
rect 26349 10009 26361 10385
rect 26395 10009 26407 10385
rect 26349 9997 26407 10009
rect 26467 10385 26525 10397
rect 26467 10009 26479 10385
rect 26513 10009 26525 10385
rect 26467 9997 26525 10009
rect -3806 8858 -3406 8870
rect -3806 8824 -3794 8858
rect -3418 8824 -3406 8858
rect -3806 8812 -3406 8824
rect -3606 8729 -3406 8741
rect -3606 8695 -3594 8729
rect -3418 8695 -3406 8729
rect -3606 8683 -3406 8695
rect -3113 8915 -2713 8927
rect -3113 8881 -3101 8915
rect -2725 8881 -2713 8915
rect 31466 10581 31524 10593
rect 27657 10385 27715 10397
rect 27657 10009 27669 10385
rect 27703 10009 27715 10385
rect 27657 9997 27715 10009
rect 27775 10385 27833 10397
rect 27775 10009 27787 10385
rect 27821 10009 27833 10385
rect 27775 9997 27833 10009
rect 27893 10385 27951 10397
rect 27893 10009 27905 10385
rect 27939 10009 27951 10385
rect 27893 9997 27951 10009
rect 28011 10385 28069 10397
rect 28011 10009 28023 10385
rect 28057 10009 28069 10385
rect 28011 9997 28069 10009
rect 28129 10385 28187 10397
rect 28129 10009 28141 10385
rect 28175 10009 28187 10385
rect 28129 9997 28187 10009
rect 28247 10385 28305 10397
rect 28247 10009 28259 10385
rect 28293 10009 28305 10385
rect 28247 9997 28305 10009
rect 28365 10385 28423 10397
rect 28365 10009 28377 10385
rect 28411 10009 28423 10385
rect 28365 9997 28423 10009
rect 31466 10405 31478 10581
rect 31512 10405 31524 10581
rect 31466 10393 31524 10405
rect 31584 10581 31642 10593
rect 31584 10405 31596 10581
rect 31630 10405 31642 10581
rect 31584 10393 31642 10405
rect 31702 10581 31760 10593
rect 31702 10405 31714 10581
rect 31748 10405 31760 10581
rect 31702 10393 31760 10405
rect 31820 10581 31878 10593
rect 31820 10405 31832 10581
rect 31866 10405 31878 10581
rect 31820 10393 31878 10405
rect 31950 10405 31962 10781
rect 31996 10405 32008 10781
rect 31950 10393 32008 10405
rect 32068 10781 32126 10793
rect 32068 10405 32080 10781
rect 32114 10405 32126 10781
rect 32068 10393 32126 10405
rect 32186 10781 32244 10793
rect 32186 10405 32198 10781
rect 32232 10405 32244 10781
rect 32186 10393 32244 10405
rect 32304 10781 32362 10793
rect 32304 10405 32316 10781
rect 32350 10405 32362 10781
rect 32304 10393 32362 10405
rect 32422 10781 32480 10793
rect 32422 10405 32434 10781
rect 32468 10405 32480 10781
rect 32422 10393 32480 10405
rect 32540 10781 32598 10793
rect 32540 10405 32552 10781
rect 32586 10405 32598 10781
rect 32540 10393 32598 10405
rect 32658 10781 32716 10793
rect 32658 10405 32670 10781
rect 32704 10405 32716 10781
rect 36755 10791 37155 10803
rect 36755 10757 36767 10791
rect 37143 10757 37155 10791
rect 36755 10745 37155 10757
rect 32658 10393 32716 10405
rect 32787 10581 32845 10593
rect 32787 10405 32799 10581
rect 32833 10405 32845 10581
rect 32787 10393 32845 10405
rect 32905 10581 32963 10593
rect 32905 10405 32917 10581
rect 32951 10405 32963 10581
rect 32905 10393 32963 10405
rect 33023 10581 33081 10593
rect 33023 10405 33035 10581
rect 33069 10405 33081 10581
rect 33023 10393 33081 10405
rect 33141 10581 33199 10593
rect 36755 10673 37155 10685
rect 36755 10639 36767 10673
rect 37143 10639 37155 10673
rect 36755 10627 37155 10639
rect 33141 10405 33153 10581
rect 33187 10405 33199 10581
rect 33141 10393 33199 10405
rect 33259 10578 33317 10590
rect 33259 10402 33271 10578
rect 33305 10402 33317 10578
rect 33259 10390 33317 10402
rect 33377 10578 33435 10590
rect 33377 10402 33389 10578
rect 33423 10402 33435 10578
rect 33377 10390 33435 10402
rect 33495 10578 33553 10590
rect 33495 10402 33507 10578
rect 33541 10402 33553 10578
rect 33495 10390 33553 10402
rect 33613 10578 33671 10590
rect 33613 10402 33625 10578
rect 33659 10402 33671 10578
rect 33613 10390 33671 10402
rect 33731 10578 33789 10590
rect 33731 10402 33743 10578
rect 33777 10402 33789 10578
rect 33731 10390 33789 10402
rect 33849 10578 33907 10590
rect 33849 10402 33861 10578
rect 33895 10402 33907 10578
rect 33849 10390 33907 10402
rect 33967 10578 34025 10590
rect 33967 10402 33979 10578
rect 34013 10402 34025 10578
rect 33967 10390 34025 10402
rect 34085 10578 34143 10590
rect 34085 10402 34097 10578
rect 34131 10402 34143 10578
rect 34085 10390 34143 10402
rect 34203 10578 34261 10590
rect 34203 10402 34215 10578
rect 34249 10402 34261 10578
rect 34203 10390 34261 10402
rect 34321 10578 34379 10590
rect 34321 10402 34333 10578
rect 34367 10402 34379 10578
rect 36755 10555 37155 10567
rect 36755 10521 36767 10555
rect 37143 10521 37155 10555
rect 36755 10509 37155 10521
rect 34321 10390 34379 10402
rect 36755 10437 37155 10449
rect 36755 10403 36767 10437
rect 37143 10403 37155 10437
rect 36755 10391 37155 10403
rect 31893 10088 31951 10100
rect 29651 9473 29709 9485
rect 29651 9297 29663 9473
rect 29697 9297 29709 9473
rect 29651 9285 29709 9297
rect 29769 9473 29827 9485
rect 29769 9297 29781 9473
rect 29815 9297 29827 9473
rect 29769 9285 29827 9297
rect 29887 9473 29945 9485
rect 29887 9297 29899 9473
rect 29933 9297 29945 9473
rect 29887 9285 29945 9297
rect 30005 9473 30063 9485
rect 30005 9297 30017 9473
rect 30051 9297 30063 9473
rect 30005 9285 30063 9297
rect 30123 9473 30181 9485
rect 30123 9297 30135 9473
rect 30169 9297 30181 9473
rect 30123 9285 30181 9297
rect 30241 9473 30299 9485
rect 30241 9297 30253 9473
rect 30287 9297 30299 9473
rect 30241 9285 30299 9297
rect 30359 9473 30417 9485
rect 30359 9297 30371 9473
rect 30405 9297 30417 9473
rect 30359 9285 30417 9297
rect 30477 9473 30535 9485
rect 30477 9297 30489 9473
rect 30523 9297 30535 9473
rect 30477 9285 30535 9297
rect 30595 9473 30653 9485
rect 30595 9297 30607 9473
rect 30641 9297 30653 9473
rect 30595 9285 30653 9297
rect 30713 9473 30771 9485
rect 30713 9297 30725 9473
rect 30759 9297 30771 9473
rect 31893 9712 31905 10088
rect 31939 9712 31951 10088
rect 31893 9700 31951 9712
rect 32011 10088 32069 10100
rect 32011 9712 32023 10088
rect 32057 9712 32069 10088
rect 32011 9700 32069 9712
rect 32129 10088 32187 10100
rect 32129 9712 32141 10088
rect 32175 9712 32187 10088
rect 32129 9700 32187 9712
rect 32247 10088 32305 10100
rect 32247 9712 32259 10088
rect 32293 9712 32305 10088
rect 32247 9700 32305 9712
rect 32365 10088 32423 10100
rect 32365 9712 32377 10088
rect 32411 9712 32423 10088
rect 32365 9700 32423 9712
rect 32483 10088 32541 10100
rect 32483 9712 32495 10088
rect 32529 9712 32541 10088
rect 32483 9700 32541 9712
rect 32601 10088 32659 10100
rect 32601 9712 32613 10088
rect 32647 9712 32659 10088
rect 32601 9700 32659 9712
rect 36955 10318 37155 10330
rect 36955 10284 36967 10318
rect 37143 10284 37155 10318
rect 36955 10272 37155 10284
rect 36955 10200 37155 10212
rect 36955 10166 36967 10200
rect 37143 10166 37155 10200
rect 36955 10154 37155 10166
rect 36955 10082 37155 10094
rect 36955 10048 36967 10082
rect 37143 10048 37155 10082
rect 36955 10036 37155 10048
rect 36955 9964 37155 9976
rect 36955 9930 36967 9964
rect 37143 9930 37155 9964
rect 36955 9918 37155 9930
rect 36955 9382 37155 9394
rect 30713 9285 30771 9297
rect -3113 8869 -2713 8881
rect -3606 8611 -3406 8623
rect -3606 8577 -3594 8611
rect -3418 8577 -3406 8611
rect 36955 9348 36967 9382
rect 37143 9348 37155 9382
rect 36955 9336 37155 9348
rect 36955 9264 37155 9276
rect 36955 9230 36967 9264
rect 37143 9230 37155 9264
rect 36955 9218 37155 9230
rect 36955 9146 37155 9158
rect 36955 9112 36967 9146
rect 37143 9112 37155 9146
rect 36955 9100 37155 9112
rect 36955 9028 37155 9040
rect 36955 8994 36967 9028
rect 37143 8994 37155 9028
rect 36955 8953 37155 8994
rect 36755 8941 37155 8953
rect 36755 8907 36767 8941
rect 37143 8907 37155 8941
rect 36755 8895 37155 8907
rect 36755 8823 37155 8835
rect 36755 8789 36767 8823
rect 37143 8789 37155 8823
rect 36755 8777 37155 8789
rect 36755 8705 37155 8717
rect 36755 8671 36767 8705
rect 37143 8671 37155 8705
rect 36755 8659 37155 8671
rect -3606 8565 -3406 8577
rect 36755 8587 37155 8599
rect 36755 8553 36767 8587
rect 37143 8553 37155 8587
rect 36755 8541 37155 8553
rect -3606 8493 -3406 8505
rect -3606 8459 -3594 8493
rect -3418 8459 -3406 8493
rect -3606 8447 -3406 8459
rect 36755 8474 37155 8486
rect 36755 8440 36767 8474
rect 37143 8440 37155 8474
rect 36755 8428 37155 8440
rect -3606 8375 -3406 8387
rect -3606 8341 -3594 8375
rect -3418 8341 -3406 8375
rect -3606 8329 -3406 8341
rect 36755 8356 37155 8368
rect 36755 8322 36767 8356
rect 37143 8322 37155 8356
rect 36755 8310 37155 8322
rect 36755 8238 37155 8250
rect 36755 8204 36767 8238
rect 37143 8204 37155 8238
rect 36755 8192 37155 8204
rect 36755 8120 37155 8132
rect 36755 8086 36767 8120
rect 37143 8086 37155 8120
rect 36755 8074 37155 8086
rect -3606 7981 -3406 7993
rect -3606 7947 -3594 7981
rect -3418 7947 -3406 7981
rect -3606 7935 -3406 7947
rect -3606 7863 -3406 7875
rect -3606 7829 -3594 7863
rect -3418 7829 -3406 7863
rect -3606 7817 -3406 7829
rect 36755 8002 37155 8014
rect 36755 7968 36767 8002
rect 37143 7968 37155 8002
rect 36755 7956 37155 7968
rect 36755 7884 37155 7896
rect 36755 7850 36767 7884
rect 37143 7850 37155 7884
rect 36755 7838 37155 7850
rect -3606 7745 -3406 7757
rect -3606 7711 -3594 7745
rect -3418 7711 -3406 7745
rect -3606 7699 -3406 7711
rect -3606 7627 -3406 7639
rect -3606 7593 -3594 7627
rect -3418 7593 -3406 7627
rect -3606 7581 -3406 7593
rect -3806 7497 -3406 7509
rect -3806 7463 -3794 7497
rect -3418 7463 -3406 7497
rect -3806 7451 -3406 7463
rect -3113 7554 -2713 7566
rect -3113 7520 -3101 7554
rect -2725 7520 -2713 7554
rect -3113 7508 -2713 7520
rect -3806 7379 -3406 7391
rect -3806 7345 -3794 7379
rect -3418 7345 -3406 7379
rect -3806 7333 -3406 7345
rect -3113 7436 -2713 7448
rect -3113 7402 -3101 7436
rect -2725 7402 -2713 7436
rect -3113 7390 -2713 7402
rect 1109 7461 1167 7473
rect -3806 7261 -3406 7273
rect -3806 7227 -3794 7261
rect -3418 7227 -3406 7261
rect -3806 7215 -3406 7227
rect -3113 7318 -2713 7330
rect -3113 7284 -3101 7318
rect -2725 7284 -2713 7318
rect -3113 7272 -2713 7284
rect 1109 7285 1121 7461
rect 1155 7285 1167 7461
rect 1109 7273 1167 7285
rect 1227 7461 1285 7473
rect 1227 7285 1239 7461
rect 1273 7285 1285 7461
rect 1227 7273 1285 7285
rect 1345 7461 1403 7473
rect 1345 7285 1357 7461
rect 1391 7285 1403 7461
rect 1345 7273 1403 7285
rect 1463 7461 1521 7473
rect 1463 7285 1475 7461
rect 1509 7285 1521 7461
rect 1463 7273 1521 7285
rect 1581 7461 1639 7473
rect 1581 7285 1593 7461
rect 1627 7285 1639 7461
rect 1581 7273 1639 7285
rect 1699 7461 1757 7473
rect 1699 7285 1711 7461
rect 1745 7285 1757 7461
rect 1699 7273 1757 7285
rect 1817 7461 1875 7473
rect 1817 7285 1829 7461
rect 1863 7285 1875 7461
rect 1817 7273 1875 7285
rect 1935 7461 1993 7473
rect 1935 7285 1947 7461
rect 1981 7285 1993 7461
rect 1935 7273 1993 7285
rect 2053 7461 2111 7473
rect 2053 7285 2065 7461
rect 2099 7285 2111 7461
rect 2053 7273 2111 7285
rect 2171 7461 2229 7473
rect 2171 7285 2183 7461
rect 2217 7285 2229 7461
rect 6343 7349 6401 7361
rect 2171 7273 2229 7285
rect 4018 7277 4076 7289
rect -3113 7200 -2713 7212
rect -3113 7166 -3101 7200
rect -2725 7166 -2713 7200
rect -3806 7143 -3406 7155
rect -3113 7154 -2713 7166
rect -3806 7109 -3794 7143
rect -3418 7109 -3406 7143
rect -3806 7097 -3406 7109
rect -3806 7025 -3406 7037
rect -3806 6991 -3794 7025
rect -3418 6991 -3406 7025
rect -3806 6979 -3406 6991
rect -3806 6907 -3406 6919
rect -3806 6873 -3794 6907
rect -3418 6873 -3406 6907
rect -3806 6861 -3406 6873
rect -3113 7082 -2713 7094
rect -3113 7048 -3101 7082
rect -2725 7048 -2713 7082
rect -3113 7036 -2713 7048
rect 4018 7101 4030 7277
rect 4064 7101 4076 7277
rect 4018 7089 4076 7101
rect 4136 7277 4194 7289
rect 4136 7101 4148 7277
rect 4182 7101 4194 7277
rect 4136 7089 4194 7101
rect 4254 7277 4312 7289
rect 4254 7101 4266 7277
rect 4300 7101 4312 7277
rect 4254 7089 4312 7101
rect 4372 7277 4430 7289
rect 4372 7101 4384 7277
rect 4418 7101 4430 7277
rect 4372 7089 4430 7101
rect 4490 7277 4548 7289
rect 4490 7101 4502 7277
rect 4536 7101 4548 7277
rect 4490 7089 4548 7101
rect 4608 7277 4666 7289
rect 4608 7101 4620 7277
rect 4654 7101 4666 7277
rect 4608 7089 4666 7101
rect 4726 7277 4784 7289
rect 4726 7101 4738 7277
rect 4772 7101 4784 7277
rect 4726 7089 4784 7101
rect 4844 7277 4902 7289
rect 4844 7101 4856 7277
rect 4890 7101 4902 7277
rect 4844 7089 4902 7101
rect 4962 7277 5020 7289
rect 4962 7101 4974 7277
rect 5008 7101 5020 7277
rect 4962 7089 5020 7101
rect 5080 7277 5138 7289
rect 5080 7101 5092 7277
rect 5126 7101 5138 7277
rect 5080 7089 5138 7101
rect -3113 6964 -2713 6976
rect -3113 6930 -3101 6964
rect -2725 6930 -2713 6964
rect -3113 6918 -2713 6930
rect -3806 6789 -3406 6801
rect -3806 6755 -3794 6789
rect -3418 6755 -3406 6789
rect -3806 6743 -3406 6755
rect -3606 6660 -3406 6672
rect -3606 6626 -3594 6660
rect -3418 6626 -3406 6660
rect -3606 6614 -3406 6626
rect -3113 6846 -2713 6858
rect -3113 6812 -3101 6846
rect -2725 6812 -2713 6846
rect -3113 6800 -2713 6812
rect 6343 6973 6355 7349
rect 6389 6973 6401 7349
rect 6343 6961 6401 6973
rect 6461 7349 6519 7361
rect 6461 6973 6473 7349
rect 6507 6973 6519 7349
rect 6461 6961 6519 6973
rect 6579 7349 6637 7361
rect 6579 6973 6591 7349
rect 6625 6973 6637 7349
rect 6579 6961 6637 6973
rect 6697 7349 6755 7361
rect 6697 6973 6709 7349
rect 6743 6973 6755 7349
rect 6697 6961 6755 6973
rect 6815 7349 6873 7361
rect 6815 6973 6827 7349
rect 6861 6973 6873 7349
rect 6815 6961 6873 6973
rect 6933 7349 6991 7361
rect 6933 6973 6945 7349
rect 6979 6973 6991 7349
rect 6933 6961 6991 6973
rect 7051 7349 7109 7361
rect 7051 6973 7063 7349
rect 7097 6973 7109 7349
rect 7051 6961 7109 6973
rect 7485 7353 7543 7365
rect 7485 6977 7497 7353
rect 7531 6977 7543 7353
rect 7485 6965 7543 6977
rect 7603 7353 7661 7365
rect 7603 6977 7615 7353
rect 7649 6977 7661 7353
rect 7603 6965 7661 6977
rect 7721 7353 7779 7365
rect 7721 6977 7733 7353
rect 7767 6977 7779 7353
rect 7721 6965 7779 6977
rect 7839 7353 7897 7365
rect 7839 6977 7851 7353
rect 7885 6977 7897 7353
rect 7839 6965 7897 6977
rect 7957 7353 8015 7365
rect 7957 6977 7969 7353
rect 8003 6977 8015 7353
rect 7957 6965 8015 6977
rect 8075 7353 8133 7365
rect 8075 6977 8087 7353
rect 8121 6977 8133 7353
rect 8075 6965 8133 6977
rect 8193 7353 8251 7365
rect 36755 7766 37155 7778
rect 36755 7732 36767 7766
rect 37143 7732 37155 7766
rect 36755 7720 37155 7732
rect 36755 7647 37155 7659
rect 36755 7613 36767 7647
rect 37143 7613 37155 7647
rect 36755 7601 37155 7613
rect 29722 7553 29780 7565
rect 8193 6977 8205 7353
rect 8239 6977 8251 7353
rect 12894 7347 12952 7359
rect 10569 7275 10627 7287
rect 10569 7099 10581 7275
rect 10615 7099 10627 7275
rect 10569 7087 10627 7099
rect 10687 7275 10745 7287
rect 10687 7099 10699 7275
rect 10733 7099 10745 7275
rect 10687 7087 10745 7099
rect 10805 7275 10863 7287
rect 10805 7099 10817 7275
rect 10851 7099 10863 7275
rect 10805 7087 10863 7099
rect 10923 7275 10981 7287
rect 10923 7099 10935 7275
rect 10969 7099 10981 7275
rect 10923 7087 10981 7099
rect 11041 7275 11099 7287
rect 11041 7099 11053 7275
rect 11087 7099 11099 7275
rect 11041 7087 11099 7099
rect 11159 7275 11217 7287
rect 11159 7099 11171 7275
rect 11205 7099 11217 7275
rect 11159 7087 11217 7099
rect 11277 7275 11335 7287
rect 11277 7099 11289 7275
rect 11323 7099 11335 7275
rect 11277 7087 11335 7099
rect 11395 7275 11453 7287
rect 11395 7099 11407 7275
rect 11441 7099 11453 7275
rect 11395 7087 11453 7099
rect 11513 7275 11571 7287
rect 11513 7099 11525 7275
rect 11559 7099 11571 7275
rect 11513 7087 11571 7099
rect 11631 7275 11689 7287
rect 11631 7099 11643 7275
rect 11677 7099 11689 7275
rect 11631 7087 11689 7099
rect 8193 6965 8251 6977
rect -3606 6542 -3406 6554
rect -3606 6508 -3594 6542
rect -3418 6508 -3406 6542
rect -3606 6496 -3406 6508
rect -3606 6424 -3406 6436
rect -3606 6390 -3594 6424
rect -3418 6390 -3406 6424
rect 12894 6971 12906 7347
rect 12940 6971 12952 7347
rect 12894 6959 12952 6971
rect 13012 7347 13070 7359
rect 13012 6971 13024 7347
rect 13058 6971 13070 7347
rect 13012 6959 13070 6971
rect 13130 7347 13188 7359
rect 13130 6971 13142 7347
rect 13176 6971 13188 7347
rect 13130 6959 13188 6971
rect 13248 7347 13306 7359
rect 13248 6971 13260 7347
rect 13294 6971 13306 7347
rect 13248 6959 13306 6971
rect 13366 7347 13424 7359
rect 13366 6971 13378 7347
rect 13412 6971 13424 7347
rect 13366 6959 13424 6971
rect 13484 7347 13542 7359
rect 13484 6971 13496 7347
rect 13530 6971 13542 7347
rect 13484 6959 13542 6971
rect 13602 7347 13660 7359
rect 13602 6971 13614 7347
rect 13648 6971 13660 7347
rect 13602 6959 13660 6971
rect 14036 7351 14094 7363
rect 14036 6975 14048 7351
rect 14082 6975 14094 7351
rect 14036 6963 14094 6975
rect 14154 7351 14212 7363
rect 14154 6975 14166 7351
rect 14200 6975 14212 7351
rect 14154 6963 14212 6975
rect 14272 7351 14330 7363
rect 14272 6975 14284 7351
rect 14318 6975 14330 7351
rect 14272 6963 14330 6975
rect 14390 7351 14448 7363
rect 14390 6975 14402 7351
rect 14436 6975 14448 7351
rect 14390 6963 14448 6975
rect 14508 7351 14566 7363
rect 14508 6975 14520 7351
rect 14554 6975 14566 7351
rect 14508 6963 14566 6975
rect 14626 7351 14684 7363
rect 14626 6975 14638 7351
rect 14672 6975 14684 7351
rect 14626 6963 14684 6975
rect 14744 7351 14802 7363
rect 14744 6975 14756 7351
rect 14790 6975 14802 7351
rect 19549 7348 19607 7360
rect 17224 7276 17282 7288
rect 17224 7100 17236 7276
rect 17270 7100 17282 7276
rect 17224 7088 17282 7100
rect 17342 7276 17400 7288
rect 17342 7100 17354 7276
rect 17388 7100 17400 7276
rect 17342 7088 17400 7100
rect 17460 7276 17518 7288
rect 17460 7100 17472 7276
rect 17506 7100 17518 7276
rect 17460 7088 17518 7100
rect 17578 7276 17636 7288
rect 17578 7100 17590 7276
rect 17624 7100 17636 7276
rect 17578 7088 17636 7100
rect 17696 7276 17754 7288
rect 17696 7100 17708 7276
rect 17742 7100 17754 7276
rect 17696 7088 17754 7100
rect 17814 7276 17872 7288
rect 17814 7100 17826 7276
rect 17860 7100 17872 7276
rect 17814 7088 17872 7100
rect 17932 7276 17990 7288
rect 17932 7100 17944 7276
rect 17978 7100 17990 7276
rect 17932 7088 17990 7100
rect 18050 7276 18108 7288
rect 18050 7100 18062 7276
rect 18096 7100 18108 7276
rect 18050 7088 18108 7100
rect 18168 7276 18226 7288
rect 18168 7100 18180 7276
rect 18214 7100 18226 7276
rect 18168 7088 18226 7100
rect 18286 7276 18344 7288
rect 18286 7100 18298 7276
rect 18332 7100 18344 7276
rect 18286 7088 18344 7100
rect 14744 6963 14802 6975
rect -3606 6378 -3406 6390
rect 6772 6566 6830 6578
rect 6772 6390 6784 6566
rect 6818 6390 6830 6566
rect 6772 6378 6830 6390
rect 6890 6566 6948 6578
rect 6890 6390 6902 6566
rect 6936 6390 6948 6566
rect 6890 6378 6948 6390
rect 7008 6566 7066 6578
rect 7008 6390 7020 6566
rect 7054 6390 7066 6566
rect 7008 6378 7066 6390
rect 7126 6566 7184 6578
rect 7126 6390 7138 6566
rect 7172 6390 7184 6566
rect 7126 6378 7184 6390
rect 7914 6570 7972 6582
rect 7914 6394 7926 6570
rect 7960 6394 7972 6570
rect 7914 6382 7972 6394
rect 8032 6570 8090 6582
rect 8032 6394 8044 6570
rect 8078 6394 8090 6570
rect 8032 6382 8090 6394
rect 8150 6570 8208 6582
rect 8150 6394 8162 6570
rect 8196 6394 8208 6570
rect 8150 6382 8208 6394
rect 8268 6570 8326 6582
rect 8268 6394 8280 6570
rect 8314 6394 8326 6570
rect 19549 6972 19561 7348
rect 19595 6972 19607 7348
rect 19549 6960 19607 6972
rect 19667 7348 19725 7360
rect 19667 6972 19679 7348
rect 19713 6972 19725 7348
rect 19667 6960 19725 6972
rect 19785 7348 19843 7360
rect 19785 6972 19797 7348
rect 19831 6972 19843 7348
rect 19785 6960 19843 6972
rect 19903 7348 19961 7360
rect 19903 6972 19915 7348
rect 19949 6972 19961 7348
rect 19903 6960 19961 6972
rect 20021 7348 20079 7360
rect 20021 6972 20033 7348
rect 20067 6972 20079 7348
rect 20021 6960 20079 6972
rect 20139 7348 20197 7360
rect 20139 6972 20151 7348
rect 20185 6972 20197 7348
rect 20139 6960 20197 6972
rect 20257 7348 20315 7360
rect 20257 6972 20269 7348
rect 20303 6972 20315 7348
rect 20257 6960 20315 6972
rect 20691 7352 20749 7364
rect 20691 6976 20703 7352
rect 20737 6976 20749 7352
rect 20691 6964 20749 6976
rect 20809 7352 20867 7364
rect 20809 6976 20821 7352
rect 20855 6976 20867 7352
rect 20809 6964 20867 6976
rect 20927 7352 20985 7364
rect 20927 6976 20939 7352
rect 20973 6976 20985 7352
rect 20927 6964 20985 6976
rect 21045 7352 21103 7364
rect 21045 6976 21057 7352
rect 21091 6976 21103 7352
rect 21045 6964 21103 6976
rect 21163 7352 21221 7364
rect 21163 6976 21175 7352
rect 21209 6976 21221 7352
rect 21163 6964 21221 6976
rect 21281 7352 21339 7364
rect 21281 6976 21293 7352
rect 21327 6976 21339 7352
rect 21281 6964 21339 6976
rect 21399 7352 21457 7364
rect 29722 7377 29734 7553
rect 29768 7377 29780 7553
rect 29722 7365 29780 7377
rect 29840 7553 29898 7565
rect 29840 7377 29852 7553
rect 29886 7377 29898 7553
rect 29840 7365 29898 7377
rect 29958 7553 30016 7565
rect 29958 7377 29970 7553
rect 30004 7377 30016 7553
rect 29958 7365 30016 7377
rect 30076 7553 30134 7565
rect 30076 7377 30088 7553
rect 30122 7377 30134 7553
rect 30076 7365 30134 7377
rect 30194 7553 30252 7565
rect 30194 7377 30206 7553
rect 30240 7377 30252 7553
rect 30194 7365 30252 7377
rect 30312 7553 30370 7565
rect 30312 7377 30324 7553
rect 30358 7377 30370 7553
rect 30312 7365 30370 7377
rect 30430 7553 30488 7565
rect 30430 7377 30442 7553
rect 30476 7377 30488 7553
rect 30430 7365 30488 7377
rect 30548 7553 30606 7565
rect 30548 7377 30560 7553
rect 30594 7377 30606 7553
rect 30548 7365 30606 7377
rect 30666 7553 30724 7565
rect 30666 7377 30678 7553
rect 30712 7377 30724 7553
rect 30666 7365 30724 7377
rect 30784 7553 30842 7565
rect 30784 7377 30796 7553
rect 30830 7377 30842 7553
rect 30784 7365 30842 7377
rect 36755 7529 37155 7541
rect 36755 7495 36767 7529
rect 37143 7495 37155 7529
rect 36755 7483 37155 7495
rect 36755 7411 37155 7423
rect 36755 7377 36767 7411
rect 37143 7377 37155 7411
rect 36755 7365 37155 7377
rect 21399 6976 21411 7352
rect 21445 6976 21457 7352
rect 26171 7349 26229 7361
rect 23846 7277 23904 7289
rect 23846 7101 23858 7277
rect 23892 7101 23904 7277
rect 23846 7089 23904 7101
rect 23964 7277 24022 7289
rect 23964 7101 23976 7277
rect 24010 7101 24022 7277
rect 23964 7089 24022 7101
rect 24082 7277 24140 7289
rect 24082 7101 24094 7277
rect 24128 7101 24140 7277
rect 24082 7089 24140 7101
rect 24200 7277 24258 7289
rect 24200 7101 24212 7277
rect 24246 7101 24258 7277
rect 24200 7089 24258 7101
rect 24318 7277 24376 7289
rect 24318 7101 24330 7277
rect 24364 7101 24376 7277
rect 24318 7089 24376 7101
rect 24436 7277 24494 7289
rect 24436 7101 24448 7277
rect 24482 7101 24494 7277
rect 24436 7089 24494 7101
rect 24554 7277 24612 7289
rect 24554 7101 24566 7277
rect 24600 7101 24612 7277
rect 24554 7089 24612 7101
rect 24672 7277 24730 7289
rect 24672 7101 24684 7277
rect 24718 7101 24730 7277
rect 24672 7089 24730 7101
rect 24790 7277 24848 7289
rect 24790 7101 24802 7277
rect 24836 7101 24848 7277
rect 24790 7089 24848 7101
rect 24908 7277 24966 7289
rect 24908 7101 24920 7277
rect 24954 7101 24966 7277
rect 24908 7089 24966 7101
rect 21399 6964 21457 6976
rect 8268 6382 8326 6394
rect -3606 6306 -3406 6318
rect -3606 6272 -3594 6306
rect -3418 6272 -3406 6306
rect 13323 6564 13381 6576
rect 13323 6388 13335 6564
rect 13369 6388 13381 6564
rect 13323 6376 13381 6388
rect 13441 6564 13499 6576
rect 13441 6388 13453 6564
rect 13487 6388 13499 6564
rect 13441 6376 13499 6388
rect 13559 6564 13617 6576
rect 13559 6388 13571 6564
rect 13605 6388 13617 6564
rect 13559 6376 13617 6388
rect 13677 6564 13735 6576
rect 13677 6388 13689 6564
rect 13723 6388 13735 6564
rect 13677 6376 13735 6388
rect 14465 6568 14523 6580
rect 14465 6392 14477 6568
rect 14511 6392 14523 6568
rect 14465 6380 14523 6392
rect 14583 6568 14641 6580
rect 14583 6392 14595 6568
rect 14629 6392 14641 6568
rect 14583 6380 14641 6392
rect 14701 6568 14759 6580
rect 14701 6392 14713 6568
rect 14747 6392 14759 6568
rect 14701 6380 14759 6392
rect 14819 6568 14877 6580
rect 14819 6392 14831 6568
rect 14865 6392 14877 6568
rect 26171 6973 26183 7349
rect 26217 6973 26229 7349
rect 26171 6961 26229 6973
rect 26289 7349 26347 7361
rect 26289 6973 26301 7349
rect 26335 6973 26347 7349
rect 26289 6961 26347 6973
rect 26407 7349 26465 7361
rect 26407 6973 26419 7349
rect 26453 6973 26465 7349
rect 26407 6961 26465 6973
rect 26525 7349 26583 7361
rect 26525 6973 26537 7349
rect 26571 6973 26583 7349
rect 26525 6961 26583 6973
rect 26643 7349 26701 7361
rect 26643 6973 26655 7349
rect 26689 6973 26701 7349
rect 26643 6961 26701 6973
rect 26761 7349 26819 7361
rect 26761 6973 26773 7349
rect 26807 6973 26819 7349
rect 26761 6961 26819 6973
rect 26879 7349 26937 7361
rect 26879 6973 26891 7349
rect 26925 6973 26937 7349
rect 26879 6961 26937 6973
rect 27313 7353 27371 7365
rect 27313 6977 27325 7353
rect 27359 6977 27371 7353
rect 27313 6965 27371 6977
rect 27431 7353 27489 7365
rect 27431 6977 27443 7353
rect 27477 6977 27489 7353
rect 27431 6965 27489 6977
rect 27549 7353 27607 7365
rect 27549 6977 27561 7353
rect 27595 6977 27607 7353
rect 27549 6965 27607 6977
rect 27667 7353 27725 7365
rect 27667 6977 27679 7353
rect 27713 6977 27725 7353
rect 27667 6965 27725 6977
rect 27785 7353 27843 7365
rect 27785 6977 27797 7353
rect 27831 6977 27843 7353
rect 27785 6965 27843 6977
rect 27903 7353 27961 7365
rect 27903 6977 27915 7353
rect 27949 6977 27961 7353
rect 27903 6965 27961 6977
rect 28021 7353 28079 7365
rect 28021 6977 28033 7353
rect 28067 6977 28079 7353
rect 31950 7286 32008 7298
rect 28021 6965 28079 6977
rect 14819 6380 14877 6392
rect 19978 6565 20036 6577
rect 19978 6389 19990 6565
rect 20024 6389 20036 6565
rect 19978 6377 20036 6389
rect 20096 6565 20154 6577
rect 20096 6389 20108 6565
rect 20142 6389 20154 6565
rect 20096 6377 20154 6389
rect 20214 6565 20272 6577
rect 20214 6389 20226 6565
rect 20260 6389 20272 6565
rect 20214 6377 20272 6389
rect 20332 6565 20390 6577
rect 20332 6389 20344 6565
rect 20378 6389 20390 6565
rect 20332 6377 20390 6389
rect 21120 6569 21178 6581
rect 21120 6393 21132 6569
rect 21166 6393 21178 6569
rect 21120 6381 21178 6393
rect 21238 6569 21296 6581
rect 21238 6393 21250 6569
rect 21284 6393 21296 6569
rect 21238 6381 21296 6393
rect 21356 6569 21414 6581
rect 21356 6393 21368 6569
rect 21402 6393 21414 6569
rect 21356 6381 21414 6393
rect 21474 6569 21532 6581
rect 21474 6393 21486 6569
rect 21520 6393 21532 6569
rect 31466 7086 31524 7098
rect 31466 6910 31478 7086
rect 31512 6910 31524 7086
rect 31466 6898 31524 6910
rect 31584 7086 31642 7098
rect 31584 6910 31596 7086
rect 31630 6910 31642 7086
rect 31584 6898 31642 6910
rect 31702 7086 31760 7098
rect 31702 6910 31714 7086
rect 31748 6910 31760 7086
rect 31702 6898 31760 6910
rect 31820 7086 31878 7098
rect 31820 6910 31832 7086
rect 31866 6910 31878 7086
rect 31820 6898 31878 6910
rect 31950 6910 31962 7286
rect 31996 6910 32008 7286
rect 31950 6898 32008 6910
rect 32068 7286 32126 7298
rect 32068 6910 32080 7286
rect 32114 6910 32126 7286
rect 32068 6898 32126 6910
rect 32186 7286 32244 7298
rect 32186 6910 32198 7286
rect 32232 6910 32244 7286
rect 32186 6898 32244 6910
rect 32304 7286 32362 7298
rect 32304 6910 32316 7286
rect 32350 6910 32362 7286
rect 32304 6898 32362 6910
rect 32422 7286 32480 7298
rect 32422 6910 32434 7286
rect 32468 6910 32480 7286
rect 32422 6898 32480 6910
rect 32540 7286 32598 7298
rect 32540 6910 32552 7286
rect 32586 6910 32598 7286
rect 32540 6898 32598 6910
rect 32658 7286 32716 7298
rect 32658 6910 32670 7286
rect 32704 6910 32716 7286
rect 36755 7293 37155 7305
rect 36755 7259 36767 7293
rect 37143 7259 37155 7293
rect 36755 7247 37155 7259
rect 36955 7174 37155 7186
rect 32658 6898 32716 6910
rect 32787 7086 32845 7098
rect 32787 6910 32799 7086
rect 32833 6910 32845 7086
rect 32787 6898 32845 6910
rect 32905 7086 32963 7098
rect 32905 6910 32917 7086
rect 32951 6910 32963 7086
rect 32905 6898 32963 6910
rect 33023 7086 33081 7098
rect 33023 6910 33035 7086
rect 33069 6910 33081 7086
rect 33023 6898 33081 6910
rect 33141 7086 33199 7098
rect 36955 7140 36967 7174
rect 37143 7140 37155 7174
rect 36955 7128 37155 7140
rect 33141 6910 33153 7086
rect 33187 6910 33199 7086
rect 33141 6898 33199 6910
rect 33259 7083 33317 7095
rect 33259 6907 33271 7083
rect 33305 6907 33317 7083
rect 33259 6895 33317 6907
rect 33377 7083 33435 7095
rect 33377 6907 33389 7083
rect 33423 6907 33435 7083
rect 33377 6895 33435 6907
rect 33495 7083 33553 7095
rect 33495 6907 33507 7083
rect 33541 6907 33553 7083
rect 33495 6895 33553 6907
rect 33613 7083 33671 7095
rect 33613 6907 33625 7083
rect 33659 6907 33671 7083
rect 33613 6895 33671 6907
rect 33731 7083 33789 7095
rect 33731 6907 33743 7083
rect 33777 6907 33789 7083
rect 33731 6895 33789 6907
rect 33849 7083 33907 7095
rect 33849 6907 33861 7083
rect 33895 6907 33907 7083
rect 33849 6895 33907 6907
rect 33967 7083 34025 7095
rect 33967 6907 33979 7083
rect 34013 6907 34025 7083
rect 33967 6895 34025 6907
rect 34085 7083 34143 7095
rect 34085 6907 34097 7083
rect 34131 6907 34143 7083
rect 34085 6895 34143 6907
rect 34203 7083 34261 7095
rect 34203 6907 34215 7083
rect 34249 6907 34261 7083
rect 34203 6895 34261 6907
rect 34321 7083 34379 7095
rect 34321 6907 34333 7083
rect 34367 6907 34379 7083
rect 34321 6895 34379 6907
rect 36955 7056 37155 7068
rect 36955 7022 36967 7056
rect 37143 7022 37155 7056
rect 36955 7010 37155 7022
rect 21474 6381 21532 6393
rect 26600 6566 26658 6578
rect 26600 6390 26612 6566
rect 26646 6390 26658 6566
rect 26600 6378 26658 6390
rect 26718 6566 26776 6578
rect 26718 6390 26730 6566
rect 26764 6390 26776 6566
rect 26718 6378 26776 6390
rect 26836 6566 26894 6578
rect 26836 6390 26848 6566
rect 26882 6390 26894 6566
rect 26836 6378 26894 6390
rect 26954 6566 27012 6578
rect 26954 6390 26966 6566
rect 27000 6390 27012 6566
rect 26954 6378 27012 6390
rect 27742 6570 27800 6582
rect 27742 6394 27754 6570
rect 27788 6394 27800 6570
rect 27742 6382 27800 6394
rect 27860 6570 27918 6582
rect 27860 6394 27872 6570
rect 27906 6394 27918 6570
rect 27860 6382 27918 6394
rect 27978 6570 28036 6582
rect 27978 6394 27990 6570
rect 28024 6394 28036 6570
rect 27978 6382 28036 6394
rect 28096 6570 28154 6582
rect 28096 6394 28108 6570
rect 28142 6394 28154 6570
rect 31893 6593 31951 6605
rect 28096 6382 28154 6394
rect -3606 6260 -3406 6272
rect -3608 5913 -3408 5925
rect -3608 5879 -3596 5913
rect -3420 5879 -3408 5913
rect -3608 5867 -3408 5879
rect -3608 5795 -3408 5807
rect -3608 5761 -3596 5795
rect -3420 5761 -3408 5795
rect -3608 5749 -3408 5761
rect 31893 6217 31905 6593
rect 31939 6217 31951 6593
rect 31893 6205 31951 6217
rect 32011 6593 32069 6605
rect 32011 6217 32023 6593
rect 32057 6217 32069 6593
rect 32011 6205 32069 6217
rect 32129 6593 32187 6605
rect 32129 6217 32141 6593
rect 32175 6217 32187 6593
rect 32129 6205 32187 6217
rect 32247 6593 32305 6605
rect 32247 6217 32259 6593
rect 32293 6217 32305 6593
rect 32247 6205 32305 6217
rect 32365 6593 32423 6605
rect 32365 6217 32377 6593
rect 32411 6217 32423 6593
rect 32365 6205 32423 6217
rect 32483 6593 32541 6605
rect 32483 6217 32495 6593
rect 32529 6217 32541 6593
rect 32483 6205 32541 6217
rect 32601 6593 32659 6605
rect 32601 6217 32613 6593
rect 32647 6217 32659 6593
rect 32601 6205 32659 6217
rect 36955 6938 37155 6950
rect 36955 6904 36967 6938
rect 37143 6904 37155 6938
rect 36955 6892 37155 6904
rect 36955 6820 37155 6832
rect 36955 6786 36967 6820
rect 37143 6786 37155 6820
rect 36955 6774 37155 6786
rect 36951 6250 37151 6262
rect 36951 6216 36963 6250
rect 37139 6216 37151 6250
rect 36951 6204 37151 6216
rect 36951 6132 37151 6144
rect 36951 6098 36963 6132
rect 37139 6098 37151 6132
rect 36951 6086 37151 6098
rect 36951 6014 37151 6026
rect 36951 5980 36963 6014
rect 37139 5980 37151 6014
rect 36951 5968 37151 5980
rect 36951 5896 37151 5908
rect -3608 5677 -3408 5689
rect -3608 5643 -3596 5677
rect -3420 5643 -3408 5677
rect -3608 5631 -3408 5643
rect 4032 5627 4090 5639
rect -3608 5559 -3408 5571
rect -3608 5525 -3596 5559
rect -3420 5525 -3408 5559
rect -3608 5513 -3408 5525
rect -3808 5429 -3408 5441
rect -3808 5395 -3796 5429
rect -3420 5395 -3408 5429
rect -3808 5383 -3408 5395
rect -3115 5486 -2715 5498
rect -3115 5452 -3103 5486
rect -2727 5452 -2715 5486
rect -3115 5440 -2715 5452
rect 4032 5451 4044 5627
rect 4078 5451 4090 5627
rect 4032 5439 4090 5451
rect 4150 5627 4208 5639
rect 4150 5451 4162 5627
rect 4196 5451 4208 5627
rect 4150 5439 4208 5451
rect 4268 5627 4326 5639
rect 4268 5451 4280 5627
rect 4314 5451 4326 5627
rect 4268 5439 4326 5451
rect 4386 5627 4444 5639
rect 4386 5451 4398 5627
rect 4432 5451 4444 5627
rect 4386 5439 4444 5451
rect 4504 5627 4562 5639
rect 4504 5451 4516 5627
rect 4550 5451 4562 5627
rect 4504 5439 4562 5451
rect 4622 5627 4680 5639
rect 4622 5451 4634 5627
rect 4668 5451 4680 5627
rect 4622 5439 4680 5451
rect 4740 5627 4798 5639
rect 4740 5451 4752 5627
rect 4786 5451 4798 5627
rect 4740 5439 4798 5451
rect 4858 5627 4916 5639
rect 4858 5451 4870 5627
rect 4904 5451 4916 5627
rect 4858 5439 4916 5451
rect 4976 5627 5034 5639
rect 4976 5451 4988 5627
rect 5022 5451 5034 5627
rect 4976 5439 5034 5451
rect 5094 5627 5152 5639
rect 5094 5451 5106 5627
rect 5140 5451 5152 5627
rect 10583 5625 10641 5637
rect 5094 5439 5152 5451
rect 10583 5449 10595 5625
rect 10629 5449 10641 5625
rect -3808 5311 -3408 5323
rect -3808 5277 -3796 5311
rect -3420 5277 -3408 5311
rect -3808 5265 -3408 5277
rect -3115 5368 -2715 5380
rect -3115 5334 -3103 5368
rect -2727 5334 -2715 5368
rect -3115 5322 -2715 5334
rect -3808 5193 -3408 5205
rect -3808 5159 -3796 5193
rect -3420 5159 -3408 5193
rect -3808 5147 -3408 5159
rect -3115 5250 -2715 5262
rect -3115 5216 -3103 5250
rect -2727 5216 -2715 5250
rect -3115 5204 -2715 5216
rect 10583 5437 10641 5449
rect 10701 5625 10759 5637
rect 10701 5449 10713 5625
rect 10747 5449 10759 5625
rect 10701 5437 10759 5449
rect 10819 5625 10877 5637
rect 10819 5449 10831 5625
rect 10865 5449 10877 5625
rect 10819 5437 10877 5449
rect 10937 5625 10995 5637
rect 10937 5449 10949 5625
rect 10983 5449 10995 5625
rect 10937 5437 10995 5449
rect 11055 5625 11113 5637
rect 11055 5449 11067 5625
rect 11101 5449 11113 5625
rect 11055 5437 11113 5449
rect 11173 5625 11231 5637
rect 11173 5449 11185 5625
rect 11219 5449 11231 5625
rect 11173 5437 11231 5449
rect 11291 5625 11349 5637
rect 11291 5449 11303 5625
rect 11337 5449 11349 5625
rect 11291 5437 11349 5449
rect 11409 5625 11467 5637
rect 11409 5449 11421 5625
rect 11455 5449 11467 5625
rect 11409 5437 11467 5449
rect 11527 5625 11585 5637
rect 11527 5449 11539 5625
rect 11573 5449 11585 5625
rect 11527 5437 11585 5449
rect 11645 5625 11703 5637
rect 11645 5449 11657 5625
rect 11691 5449 11703 5625
rect 17238 5626 17296 5638
rect 11645 5437 11703 5449
rect 17238 5450 17250 5626
rect 17284 5450 17296 5626
rect 17238 5438 17296 5450
rect 17356 5626 17414 5638
rect 17356 5450 17368 5626
rect 17402 5450 17414 5626
rect 17356 5438 17414 5450
rect 17474 5626 17532 5638
rect 17474 5450 17486 5626
rect 17520 5450 17532 5626
rect 17474 5438 17532 5450
rect 17592 5626 17650 5638
rect 17592 5450 17604 5626
rect 17638 5450 17650 5626
rect 17592 5438 17650 5450
rect 17710 5626 17768 5638
rect 17710 5450 17722 5626
rect 17756 5450 17768 5626
rect 17710 5438 17768 5450
rect 17828 5626 17886 5638
rect 17828 5450 17840 5626
rect 17874 5450 17886 5626
rect 17828 5438 17886 5450
rect 17946 5626 18004 5638
rect 17946 5450 17958 5626
rect 17992 5450 18004 5626
rect 17946 5438 18004 5450
rect 18064 5626 18122 5638
rect 18064 5450 18076 5626
rect 18110 5450 18122 5626
rect 18064 5438 18122 5450
rect 18182 5626 18240 5638
rect 18182 5450 18194 5626
rect 18228 5450 18240 5626
rect 18182 5438 18240 5450
rect 18300 5626 18358 5638
rect 18300 5450 18312 5626
rect 18346 5450 18358 5626
rect 23860 5627 23918 5639
rect 18300 5438 18358 5450
rect 23860 5451 23872 5627
rect 23906 5451 23918 5627
rect 23860 5439 23918 5451
rect 23978 5627 24036 5639
rect 23978 5451 23990 5627
rect 24024 5451 24036 5627
rect 23978 5439 24036 5451
rect 24096 5627 24154 5639
rect 24096 5451 24108 5627
rect 24142 5451 24154 5627
rect 24096 5439 24154 5451
rect 24214 5627 24272 5639
rect 24214 5451 24226 5627
rect 24260 5451 24272 5627
rect 24214 5439 24272 5451
rect 24332 5627 24390 5639
rect 24332 5451 24344 5627
rect 24378 5451 24390 5627
rect 24332 5439 24390 5451
rect 24450 5627 24508 5639
rect 24450 5451 24462 5627
rect 24496 5451 24508 5627
rect 24450 5439 24508 5451
rect 24568 5627 24626 5639
rect 24568 5451 24580 5627
rect 24614 5451 24626 5627
rect 24568 5439 24626 5451
rect 24686 5627 24744 5639
rect 24686 5451 24698 5627
rect 24732 5451 24744 5627
rect 24686 5439 24744 5451
rect 24804 5627 24862 5639
rect 24804 5451 24816 5627
rect 24850 5451 24862 5627
rect 24804 5439 24862 5451
rect 24922 5627 24980 5639
rect 24922 5451 24934 5627
rect 24968 5451 24980 5627
rect 36951 5862 36963 5896
rect 37139 5862 37151 5896
rect 36951 5821 37151 5862
rect 36751 5809 37151 5821
rect 36751 5775 36763 5809
rect 37139 5775 37151 5809
rect 36751 5763 37151 5775
rect 36751 5691 37151 5703
rect 36751 5657 36763 5691
rect 37139 5657 37151 5691
rect 36751 5645 37151 5657
rect 36751 5573 37151 5585
rect 36751 5539 36763 5573
rect 37139 5539 37151 5573
rect 36751 5527 37151 5539
rect 24922 5439 24980 5451
rect 36751 5455 37151 5467
rect 5980 5210 6038 5222
rect -3115 5132 -2715 5144
rect -3115 5098 -3103 5132
rect -2727 5098 -2715 5132
rect -3808 5075 -3408 5087
rect -3115 5086 -2715 5098
rect -3808 5041 -3796 5075
rect -3420 5041 -3408 5075
rect -3808 5029 -3408 5041
rect -3808 4957 -3408 4969
rect -3808 4923 -3796 4957
rect -3420 4923 -3408 4957
rect -3808 4911 -3408 4923
rect -3808 4839 -3408 4851
rect -3808 4805 -3796 4839
rect -3420 4805 -3408 4839
rect -3808 4793 -3408 4805
rect -3115 5014 -2715 5026
rect -3115 4980 -3103 5014
rect -2727 4980 -2715 5014
rect -3115 4968 -2715 4980
rect -3115 4896 -2715 4908
rect -3115 4862 -3103 4896
rect -2727 4862 -2715 4896
rect -3115 4850 -2715 4862
rect -3808 4721 -3408 4733
rect -3808 4687 -3796 4721
rect -3420 4687 -3408 4721
rect -3808 4675 -3408 4687
rect -3608 4592 -3408 4604
rect -3608 4558 -3596 4592
rect -3420 4558 -3408 4592
rect -3608 4546 -3408 4558
rect -3115 4778 -2715 4790
rect -3115 4744 -3103 4778
rect -2727 4744 -2715 4778
rect 5496 5010 5554 5022
rect -3115 4732 -2715 4744
rect 5496 4834 5508 5010
rect 5542 4834 5554 5010
rect 5496 4822 5554 4834
rect 5614 5010 5672 5022
rect 5614 4834 5626 5010
rect 5660 4834 5672 5010
rect 5614 4822 5672 4834
rect 5732 5010 5790 5022
rect 5732 4834 5744 5010
rect 5778 4834 5790 5010
rect 5732 4822 5790 4834
rect 5850 5010 5908 5022
rect 5850 4834 5862 5010
rect 5896 4834 5908 5010
rect 5850 4822 5908 4834
rect 5980 4834 5992 5210
rect 6026 4834 6038 5210
rect 5980 4822 6038 4834
rect 6098 5210 6156 5222
rect 6098 4834 6110 5210
rect 6144 4834 6156 5210
rect 6098 4822 6156 4834
rect 6216 5210 6274 5222
rect 6216 4834 6228 5210
rect 6262 4834 6274 5210
rect 6216 4822 6274 4834
rect 6334 5210 6392 5222
rect 6334 4834 6346 5210
rect 6380 4834 6392 5210
rect 6334 4822 6392 4834
rect 6452 5210 6510 5222
rect 6452 4834 6464 5210
rect 6498 4834 6510 5210
rect 6452 4822 6510 4834
rect 6570 5210 6628 5222
rect 6570 4834 6582 5210
rect 6616 4834 6628 5210
rect 6570 4822 6628 4834
rect 6688 5210 6746 5222
rect 6688 4834 6700 5210
rect 6734 4834 6746 5210
rect 7878 5210 7936 5222
rect 6688 4822 6746 4834
rect 6817 5010 6875 5022
rect 6817 4834 6829 5010
rect 6863 4834 6875 5010
rect 6817 4822 6875 4834
rect 6935 5010 6993 5022
rect 6935 4834 6947 5010
rect 6981 4834 6993 5010
rect 6935 4822 6993 4834
rect 7053 5010 7111 5022
rect 7053 4834 7065 5010
rect 7099 4834 7111 5010
rect 7053 4822 7111 4834
rect 7171 5010 7229 5022
rect 7171 4834 7183 5010
rect 7217 4834 7229 5010
rect 7171 4822 7229 4834
rect 7394 5010 7452 5022
rect 7394 4834 7406 5010
rect 7440 4834 7452 5010
rect 7394 4822 7452 4834
rect 7512 5010 7570 5022
rect 7512 4834 7524 5010
rect 7558 4834 7570 5010
rect 7512 4822 7570 4834
rect 7630 5010 7688 5022
rect 7630 4834 7642 5010
rect 7676 4834 7688 5010
rect 7630 4822 7688 4834
rect 7748 5010 7806 5022
rect 7748 4834 7760 5010
rect 7794 4834 7806 5010
rect 7748 4822 7806 4834
rect 7878 4834 7890 5210
rect 7924 4834 7936 5210
rect 7878 4822 7936 4834
rect 7996 5210 8054 5222
rect 7996 4834 8008 5210
rect 8042 4834 8054 5210
rect 7996 4822 8054 4834
rect 8114 5210 8172 5222
rect 8114 4834 8126 5210
rect 8160 4834 8172 5210
rect 8114 4822 8172 4834
rect 8232 5210 8290 5222
rect 8232 4834 8244 5210
rect 8278 4834 8290 5210
rect 8232 4822 8290 4834
rect 8350 5210 8408 5222
rect 8350 4834 8362 5210
rect 8396 4834 8408 5210
rect 8350 4822 8408 4834
rect 8468 5210 8526 5222
rect 8468 4834 8480 5210
rect 8514 4834 8526 5210
rect 8468 4822 8526 4834
rect 8586 5210 8644 5222
rect 8586 4834 8598 5210
rect 8632 4834 8644 5210
rect 12531 5208 12589 5220
rect 8586 4822 8644 4834
rect 8715 5010 8773 5022
rect 8715 4834 8727 5010
rect 8761 4834 8773 5010
rect 8715 4822 8773 4834
rect 8833 5010 8891 5022
rect 8833 4834 8845 5010
rect 8879 4834 8891 5010
rect 8833 4822 8891 4834
rect 8951 5010 9009 5022
rect 8951 4834 8963 5010
rect 8997 4834 9009 5010
rect 8951 4822 9009 4834
rect 9069 5010 9127 5022
rect 9069 4834 9081 5010
rect 9115 4834 9127 5010
rect 9069 4822 9127 4834
rect 1125 4701 1183 4713
rect -3608 4474 -3408 4486
rect -3608 4440 -3596 4474
rect -3420 4440 -3408 4474
rect 1125 4525 1137 4701
rect 1171 4525 1183 4701
rect 1125 4513 1183 4525
rect 1243 4701 1301 4713
rect 1243 4525 1255 4701
rect 1289 4525 1301 4701
rect 1243 4513 1301 4525
rect 1361 4701 1419 4713
rect 1361 4525 1373 4701
rect 1407 4525 1419 4701
rect 1361 4513 1419 4525
rect 1479 4701 1537 4713
rect 1479 4525 1491 4701
rect 1525 4525 1537 4701
rect 1479 4513 1537 4525
rect 1597 4701 1655 4713
rect 1597 4525 1609 4701
rect 1643 4525 1655 4701
rect 1597 4513 1655 4525
rect 1715 4701 1773 4713
rect 1715 4525 1727 4701
rect 1761 4525 1773 4701
rect 1715 4513 1773 4525
rect 1833 4701 1891 4713
rect 1833 4525 1845 4701
rect 1879 4525 1891 4701
rect 1833 4513 1891 4525
rect 1951 4701 2009 4713
rect 1951 4525 1963 4701
rect 1997 4525 2009 4701
rect 1951 4513 2009 4525
rect 2069 4701 2127 4713
rect 2069 4525 2081 4701
rect 2115 4525 2127 4701
rect 2069 4513 2127 4525
rect 2187 4701 2245 4713
rect 2187 4525 2199 4701
rect 2233 4525 2245 4701
rect 2187 4513 2245 4525
rect -3608 4428 -3408 4440
rect -3608 4356 -3408 4368
rect -3608 4322 -3596 4356
rect -3420 4322 -3408 4356
rect -3608 4310 -3408 4322
rect -3608 4238 -3408 4250
rect -3608 4204 -3596 4238
rect -3420 4204 -3408 4238
rect -3608 4192 -3408 4204
rect 4027 4023 4085 4035
rect -3606 3844 -3406 3856
rect -3606 3810 -3594 3844
rect -3418 3810 -3406 3844
rect -3606 3798 -3406 3810
rect -3606 3726 -3406 3738
rect -3606 3692 -3594 3726
rect -3418 3692 -3406 3726
rect -3606 3680 -3406 3692
rect 4027 3847 4039 4023
rect 4073 3847 4085 4023
rect 4027 3835 4085 3847
rect 4145 4023 4203 4035
rect 4145 3847 4157 4023
rect 4191 3847 4203 4023
rect 4145 3835 4203 3847
rect 4263 4023 4321 4035
rect 4263 3847 4275 4023
rect 4309 3847 4321 4023
rect 4263 3835 4321 3847
rect 4381 4023 4439 4035
rect 4381 3847 4393 4023
rect 4427 3847 4439 4023
rect 4381 3835 4439 3847
rect 4499 4023 4557 4035
rect 4499 3847 4511 4023
rect 4545 3847 4557 4023
rect 4499 3835 4557 3847
rect 4617 4023 4675 4035
rect 4617 3847 4629 4023
rect 4663 3847 4675 4023
rect 4617 3835 4675 3847
rect 4735 4023 4793 4035
rect 4735 3847 4747 4023
rect 4781 3847 4793 4023
rect 4735 3835 4793 3847
rect 4853 4023 4911 4035
rect 4853 3847 4865 4023
rect 4899 3847 4911 4023
rect 4853 3835 4911 3847
rect 4971 4023 5029 4035
rect 4971 3847 4983 4023
rect 5017 3847 5029 4023
rect 4971 3835 5029 3847
rect 5089 4023 5147 4035
rect 5089 3847 5101 4023
rect 5135 3847 5147 4023
rect 5089 3835 5147 3847
rect 5923 4517 5981 4529
rect 5923 4141 5935 4517
rect 5969 4141 5981 4517
rect 5923 4129 5981 4141
rect 6041 4517 6099 4529
rect 6041 4141 6053 4517
rect 6087 4141 6099 4517
rect 6041 4129 6099 4141
rect 6159 4517 6217 4529
rect 6159 4141 6171 4517
rect 6205 4141 6217 4517
rect 6159 4129 6217 4141
rect 6277 4517 6335 4529
rect 6277 4141 6289 4517
rect 6323 4141 6335 4517
rect 6277 4129 6335 4141
rect 6395 4517 6453 4529
rect 6395 4141 6407 4517
rect 6441 4141 6453 4517
rect 6395 4129 6453 4141
rect 6513 4517 6571 4529
rect 6513 4141 6525 4517
rect 6559 4141 6571 4517
rect 6513 4129 6571 4141
rect 6631 4517 6689 4529
rect 6631 4141 6643 4517
rect 6677 4141 6689 4517
rect 6631 4129 6689 4141
rect -3606 3608 -3406 3620
rect -3606 3574 -3594 3608
rect -3418 3574 -3406 3608
rect -3606 3562 -3406 3574
rect 12047 5008 12105 5020
rect 12047 4832 12059 5008
rect 12093 4832 12105 5008
rect 12047 4820 12105 4832
rect 12165 5008 12223 5020
rect 12165 4832 12177 5008
rect 12211 4832 12223 5008
rect 12165 4820 12223 4832
rect 12283 5008 12341 5020
rect 12283 4832 12295 5008
rect 12329 4832 12341 5008
rect 12283 4820 12341 4832
rect 12401 5008 12459 5020
rect 12401 4832 12413 5008
rect 12447 4832 12459 5008
rect 12401 4820 12459 4832
rect 12531 4832 12543 5208
rect 12577 4832 12589 5208
rect 12531 4820 12589 4832
rect 12649 5208 12707 5220
rect 12649 4832 12661 5208
rect 12695 4832 12707 5208
rect 12649 4820 12707 4832
rect 12767 5208 12825 5220
rect 12767 4832 12779 5208
rect 12813 4832 12825 5208
rect 12767 4820 12825 4832
rect 12885 5208 12943 5220
rect 12885 4832 12897 5208
rect 12931 4832 12943 5208
rect 12885 4820 12943 4832
rect 13003 5208 13061 5220
rect 13003 4832 13015 5208
rect 13049 4832 13061 5208
rect 13003 4820 13061 4832
rect 13121 5208 13179 5220
rect 13121 4832 13133 5208
rect 13167 4832 13179 5208
rect 13121 4820 13179 4832
rect 13239 5208 13297 5220
rect 13239 4832 13251 5208
rect 13285 4832 13297 5208
rect 14429 5208 14487 5220
rect 13239 4820 13297 4832
rect 13368 5008 13426 5020
rect 13368 4832 13380 5008
rect 13414 4832 13426 5008
rect 13368 4820 13426 4832
rect 13486 5008 13544 5020
rect 13486 4832 13498 5008
rect 13532 4832 13544 5008
rect 13486 4820 13544 4832
rect 13604 5008 13662 5020
rect 13604 4832 13616 5008
rect 13650 4832 13662 5008
rect 13604 4820 13662 4832
rect 13722 5008 13780 5020
rect 13722 4832 13734 5008
rect 13768 4832 13780 5008
rect 13722 4820 13780 4832
rect 13945 5008 14003 5020
rect 13945 4832 13957 5008
rect 13991 4832 14003 5008
rect 13945 4820 14003 4832
rect 14063 5008 14121 5020
rect 14063 4832 14075 5008
rect 14109 4832 14121 5008
rect 14063 4820 14121 4832
rect 14181 5008 14239 5020
rect 14181 4832 14193 5008
rect 14227 4832 14239 5008
rect 14181 4820 14239 4832
rect 14299 5008 14357 5020
rect 14299 4832 14311 5008
rect 14345 4832 14357 5008
rect 14299 4820 14357 4832
rect 14429 4832 14441 5208
rect 14475 4832 14487 5208
rect 14429 4820 14487 4832
rect 14547 5208 14605 5220
rect 14547 4832 14559 5208
rect 14593 4832 14605 5208
rect 14547 4820 14605 4832
rect 14665 5208 14723 5220
rect 14665 4832 14677 5208
rect 14711 4832 14723 5208
rect 14665 4820 14723 4832
rect 14783 5208 14841 5220
rect 14783 4832 14795 5208
rect 14829 4832 14841 5208
rect 14783 4820 14841 4832
rect 14901 5208 14959 5220
rect 14901 4832 14913 5208
rect 14947 4832 14959 5208
rect 14901 4820 14959 4832
rect 15019 5208 15077 5220
rect 15019 4832 15031 5208
rect 15065 4832 15077 5208
rect 15019 4820 15077 4832
rect 15137 5208 15195 5220
rect 15137 4832 15149 5208
rect 15183 4832 15195 5208
rect 19186 5209 19244 5221
rect 15137 4820 15195 4832
rect 15266 5008 15324 5020
rect 15266 4832 15278 5008
rect 15312 4832 15324 5008
rect 15266 4820 15324 4832
rect 15384 5008 15442 5020
rect 15384 4832 15396 5008
rect 15430 4832 15442 5008
rect 15384 4820 15442 4832
rect 15502 5008 15560 5020
rect 15502 4832 15514 5008
rect 15548 4832 15560 5008
rect 15502 4820 15560 4832
rect 15620 5008 15678 5020
rect 15620 4832 15632 5008
rect 15666 4832 15678 5008
rect 15620 4820 15678 4832
rect 7821 4517 7879 4529
rect 7821 4141 7833 4517
rect 7867 4141 7879 4517
rect 7821 4129 7879 4141
rect 7939 4517 7997 4529
rect 7939 4141 7951 4517
rect 7985 4141 7997 4517
rect 7939 4129 7997 4141
rect 8057 4517 8115 4529
rect 8057 4141 8069 4517
rect 8103 4141 8115 4517
rect 8057 4129 8115 4141
rect 8175 4517 8233 4529
rect 8175 4141 8187 4517
rect 8221 4141 8233 4517
rect 8175 4129 8233 4141
rect 8293 4517 8351 4529
rect 8293 4141 8305 4517
rect 8339 4141 8351 4517
rect 8293 4129 8351 4141
rect 8411 4517 8469 4529
rect 8411 4141 8423 4517
rect 8457 4141 8469 4517
rect 8411 4129 8469 4141
rect 8529 4517 8587 4529
rect 8529 4141 8541 4517
rect 8575 4141 8587 4517
rect 8529 4129 8587 4141
rect 10578 4021 10636 4033
rect 10578 3845 10590 4021
rect 10624 3845 10636 4021
rect 10578 3833 10636 3845
rect 10696 4021 10754 4033
rect 10696 3845 10708 4021
rect 10742 3845 10754 4021
rect 10696 3833 10754 3845
rect 10814 4021 10872 4033
rect 10814 3845 10826 4021
rect 10860 3845 10872 4021
rect 10814 3833 10872 3845
rect 10932 4021 10990 4033
rect 10932 3845 10944 4021
rect 10978 3845 10990 4021
rect 10932 3833 10990 3845
rect 11050 4021 11108 4033
rect 11050 3845 11062 4021
rect 11096 3845 11108 4021
rect 11050 3833 11108 3845
rect 11168 4021 11226 4033
rect 11168 3845 11180 4021
rect 11214 3845 11226 4021
rect 11168 3833 11226 3845
rect 11286 4021 11344 4033
rect 11286 3845 11298 4021
rect 11332 3845 11344 4021
rect 11286 3833 11344 3845
rect 11404 4021 11462 4033
rect 11404 3845 11416 4021
rect 11450 3845 11462 4021
rect 11404 3833 11462 3845
rect 11522 4021 11580 4033
rect 11522 3845 11534 4021
rect 11568 3845 11580 4021
rect 11522 3833 11580 3845
rect 11640 4021 11698 4033
rect 11640 3845 11652 4021
rect 11686 3845 11698 4021
rect 11640 3833 11698 3845
rect 12474 4515 12532 4527
rect 12474 4139 12486 4515
rect 12520 4139 12532 4515
rect 12474 4127 12532 4139
rect 12592 4515 12650 4527
rect 12592 4139 12604 4515
rect 12638 4139 12650 4515
rect 12592 4127 12650 4139
rect 12710 4515 12768 4527
rect 12710 4139 12722 4515
rect 12756 4139 12768 4515
rect 12710 4127 12768 4139
rect 12828 4515 12886 4527
rect 12828 4139 12840 4515
rect 12874 4139 12886 4515
rect 12828 4127 12886 4139
rect 12946 4515 13004 4527
rect 12946 4139 12958 4515
rect 12992 4139 13004 4515
rect 12946 4127 13004 4139
rect 13064 4515 13122 4527
rect 13064 4139 13076 4515
rect 13110 4139 13122 4515
rect 13064 4127 13122 4139
rect 13182 4515 13240 4527
rect 13182 4139 13194 4515
rect 13228 4139 13240 4515
rect 13182 4127 13240 4139
rect -3606 3490 -3406 3502
rect -3606 3456 -3594 3490
rect -3418 3456 -3406 3490
rect -3606 3444 -3406 3456
rect -3806 3360 -3406 3372
rect -3806 3326 -3794 3360
rect -3418 3326 -3406 3360
rect -3806 3314 -3406 3326
rect -3113 3417 -2713 3429
rect -3113 3383 -3101 3417
rect -2725 3383 -2713 3417
rect -3113 3371 -2713 3383
rect -3806 3242 -3406 3254
rect -3806 3208 -3794 3242
rect -3418 3208 -3406 3242
rect -3806 3196 -3406 3208
rect -3113 3299 -2713 3311
rect -3113 3265 -3101 3299
rect -2725 3265 -2713 3299
rect -3113 3253 -2713 3265
rect 18702 5009 18760 5021
rect 18702 4833 18714 5009
rect 18748 4833 18760 5009
rect 18702 4821 18760 4833
rect 18820 5009 18878 5021
rect 18820 4833 18832 5009
rect 18866 4833 18878 5009
rect 18820 4821 18878 4833
rect 18938 5009 18996 5021
rect 18938 4833 18950 5009
rect 18984 4833 18996 5009
rect 18938 4821 18996 4833
rect 19056 5009 19114 5021
rect 19056 4833 19068 5009
rect 19102 4833 19114 5009
rect 19056 4821 19114 4833
rect 19186 4833 19198 5209
rect 19232 4833 19244 5209
rect 19186 4821 19244 4833
rect 19304 5209 19362 5221
rect 19304 4833 19316 5209
rect 19350 4833 19362 5209
rect 19304 4821 19362 4833
rect 19422 5209 19480 5221
rect 19422 4833 19434 5209
rect 19468 4833 19480 5209
rect 19422 4821 19480 4833
rect 19540 5209 19598 5221
rect 19540 4833 19552 5209
rect 19586 4833 19598 5209
rect 19540 4821 19598 4833
rect 19658 5209 19716 5221
rect 19658 4833 19670 5209
rect 19704 4833 19716 5209
rect 19658 4821 19716 4833
rect 19776 5209 19834 5221
rect 19776 4833 19788 5209
rect 19822 4833 19834 5209
rect 19776 4821 19834 4833
rect 19894 5209 19952 5221
rect 19894 4833 19906 5209
rect 19940 4833 19952 5209
rect 21084 5209 21142 5221
rect 19894 4821 19952 4833
rect 20023 5009 20081 5021
rect 20023 4833 20035 5009
rect 20069 4833 20081 5009
rect 20023 4821 20081 4833
rect 20141 5009 20199 5021
rect 20141 4833 20153 5009
rect 20187 4833 20199 5009
rect 20141 4821 20199 4833
rect 20259 5009 20317 5021
rect 20259 4833 20271 5009
rect 20305 4833 20317 5009
rect 20259 4821 20317 4833
rect 20377 5009 20435 5021
rect 20377 4833 20389 5009
rect 20423 4833 20435 5009
rect 20377 4821 20435 4833
rect 20600 5009 20658 5021
rect 20600 4833 20612 5009
rect 20646 4833 20658 5009
rect 20600 4821 20658 4833
rect 20718 5009 20776 5021
rect 20718 4833 20730 5009
rect 20764 4833 20776 5009
rect 20718 4821 20776 4833
rect 20836 5009 20894 5021
rect 20836 4833 20848 5009
rect 20882 4833 20894 5009
rect 20836 4821 20894 4833
rect 20954 5009 21012 5021
rect 20954 4833 20966 5009
rect 21000 4833 21012 5009
rect 20954 4821 21012 4833
rect 21084 4833 21096 5209
rect 21130 4833 21142 5209
rect 21084 4821 21142 4833
rect 21202 5209 21260 5221
rect 21202 4833 21214 5209
rect 21248 4833 21260 5209
rect 21202 4821 21260 4833
rect 21320 5209 21378 5221
rect 21320 4833 21332 5209
rect 21366 4833 21378 5209
rect 21320 4821 21378 4833
rect 21438 5209 21496 5221
rect 21438 4833 21450 5209
rect 21484 4833 21496 5209
rect 21438 4821 21496 4833
rect 21556 5209 21614 5221
rect 21556 4833 21568 5209
rect 21602 4833 21614 5209
rect 21556 4821 21614 4833
rect 21674 5209 21732 5221
rect 21674 4833 21686 5209
rect 21720 4833 21732 5209
rect 21674 4821 21732 4833
rect 21792 5209 21850 5221
rect 21792 4833 21804 5209
rect 21838 4833 21850 5209
rect 36751 5421 36763 5455
rect 37139 5421 37151 5455
rect 36751 5409 37151 5421
rect 36751 5342 37151 5354
rect 25808 5210 25866 5222
rect 21792 4821 21850 4833
rect 21921 5009 21979 5021
rect 21921 4833 21933 5009
rect 21967 4833 21979 5009
rect 21921 4821 21979 4833
rect 22039 5009 22097 5021
rect 22039 4833 22051 5009
rect 22085 4833 22097 5009
rect 22039 4821 22097 4833
rect 22157 5009 22215 5021
rect 22157 4833 22169 5009
rect 22203 4833 22215 5009
rect 22157 4821 22215 4833
rect 22275 5009 22333 5021
rect 22275 4833 22287 5009
rect 22321 4833 22333 5009
rect 22275 4821 22333 4833
rect 14372 4515 14430 4527
rect 14372 4139 14384 4515
rect 14418 4139 14430 4515
rect 14372 4127 14430 4139
rect 14490 4515 14548 4527
rect 14490 4139 14502 4515
rect 14536 4139 14548 4515
rect 14490 4127 14548 4139
rect 14608 4515 14666 4527
rect 14608 4139 14620 4515
rect 14654 4139 14666 4515
rect 14608 4127 14666 4139
rect 14726 4515 14784 4527
rect 14726 4139 14738 4515
rect 14772 4139 14784 4515
rect 14726 4127 14784 4139
rect 14844 4515 14902 4527
rect 14844 4139 14856 4515
rect 14890 4139 14902 4515
rect 14844 4127 14902 4139
rect 14962 4515 15020 4527
rect 14962 4139 14974 4515
rect 15008 4139 15020 4515
rect 14962 4127 15020 4139
rect 15080 4515 15138 4527
rect 15080 4139 15092 4515
rect 15126 4139 15138 4515
rect 15080 4127 15138 4139
rect 17233 4022 17291 4034
rect 17233 3846 17245 4022
rect 17279 3846 17291 4022
rect 17233 3834 17291 3846
rect 17351 4022 17409 4034
rect 17351 3846 17363 4022
rect 17397 3846 17409 4022
rect 17351 3834 17409 3846
rect 17469 4022 17527 4034
rect 17469 3846 17481 4022
rect 17515 3846 17527 4022
rect 17469 3834 17527 3846
rect 17587 4022 17645 4034
rect 17587 3846 17599 4022
rect 17633 3846 17645 4022
rect 17587 3834 17645 3846
rect 17705 4022 17763 4034
rect 17705 3846 17717 4022
rect 17751 3846 17763 4022
rect 17705 3834 17763 3846
rect 17823 4022 17881 4034
rect 17823 3846 17835 4022
rect 17869 3846 17881 4022
rect 17823 3834 17881 3846
rect 17941 4022 17999 4034
rect 17941 3846 17953 4022
rect 17987 3846 17999 4022
rect 17941 3834 17999 3846
rect 18059 4022 18117 4034
rect 18059 3846 18071 4022
rect 18105 3846 18117 4022
rect 18059 3834 18117 3846
rect 18177 4022 18235 4034
rect 18177 3846 18189 4022
rect 18223 3846 18235 4022
rect 18177 3834 18235 3846
rect 18295 4022 18353 4034
rect 18295 3846 18307 4022
rect 18341 3846 18353 4022
rect 18295 3834 18353 3846
rect 19129 4516 19187 4528
rect 19129 4140 19141 4516
rect 19175 4140 19187 4516
rect 19129 4128 19187 4140
rect 19247 4516 19305 4528
rect 19247 4140 19259 4516
rect 19293 4140 19305 4516
rect 19247 4128 19305 4140
rect 19365 4516 19423 4528
rect 19365 4140 19377 4516
rect 19411 4140 19423 4516
rect 19365 4128 19423 4140
rect 19483 4516 19541 4528
rect 19483 4140 19495 4516
rect 19529 4140 19541 4516
rect 19483 4128 19541 4140
rect 19601 4516 19659 4528
rect 19601 4140 19613 4516
rect 19647 4140 19659 4516
rect 19601 4128 19659 4140
rect 19719 4516 19777 4528
rect 19719 4140 19731 4516
rect 19765 4140 19777 4516
rect 19719 4128 19777 4140
rect 19837 4516 19895 4528
rect 19837 4140 19849 4516
rect 19883 4140 19895 4516
rect 19837 4128 19895 4140
rect -3806 3124 -3406 3136
rect -3806 3090 -3794 3124
rect -3418 3090 -3406 3124
rect -3806 3078 -3406 3090
rect -3113 3181 -2713 3193
rect -3113 3147 -3101 3181
rect -2725 3147 -2713 3181
rect -3113 3135 -2713 3147
rect 25324 5010 25382 5022
rect 25324 4834 25336 5010
rect 25370 4834 25382 5010
rect 25324 4822 25382 4834
rect 25442 5010 25500 5022
rect 25442 4834 25454 5010
rect 25488 4834 25500 5010
rect 25442 4822 25500 4834
rect 25560 5010 25618 5022
rect 25560 4834 25572 5010
rect 25606 4834 25618 5010
rect 25560 4822 25618 4834
rect 25678 5010 25736 5022
rect 25678 4834 25690 5010
rect 25724 4834 25736 5010
rect 25678 4822 25736 4834
rect 25808 4834 25820 5210
rect 25854 4834 25866 5210
rect 25808 4822 25866 4834
rect 25926 5210 25984 5222
rect 25926 4834 25938 5210
rect 25972 4834 25984 5210
rect 25926 4822 25984 4834
rect 26044 5210 26102 5222
rect 26044 4834 26056 5210
rect 26090 4834 26102 5210
rect 26044 4822 26102 4834
rect 26162 5210 26220 5222
rect 26162 4834 26174 5210
rect 26208 4834 26220 5210
rect 26162 4822 26220 4834
rect 26280 5210 26338 5222
rect 26280 4834 26292 5210
rect 26326 4834 26338 5210
rect 26280 4822 26338 4834
rect 26398 5210 26456 5222
rect 26398 4834 26410 5210
rect 26444 4834 26456 5210
rect 26398 4822 26456 4834
rect 26516 5210 26574 5222
rect 26516 4834 26528 5210
rect 26562 4834 26574 5210
rect 27706 5210 27764 5222
rect 26516 4822 26574 4834
rect 26645 5010 26703 5022
rect 26645 4834 26657 5010
rect 26691 4834 26703 5010
rect 26645 4822 26703 4834
rect 26763 5010 26821 5022
rect 26763 4834 26775 5010
rect 26809 4834 26821 5010
rect 26763 4822 26821 4834
rect 26881 5010 26939 5022
rect 26881 4834 26893 5010
rect 26927 4834 26939 5010
rect 26881 4822 26939 4834
rect 26999 5010 27057 5022
rect 26999 4834 27011 5010
rect 27045 4834 27057 5010
rect 26999 4822 27057 4834
rect 27222 5010 27280 5022
rect 27222 4834 27234 5010
rect 27268 4834 27280 5010
rect 27222 4822 27280 4834
rect 27340 5010 27398 5022
rect 27340 4834 27352 5010
rect 27386 4834 27398 5010
rect 27340 4822 27398 4834
rect 27458 5010 27516 5022
rect 27458 4834 27470 5010
rect 27504 4834 27516 5010
rect 27458 4822 27516 4834
rect 27576 5010 27634 5022
rect 27576 4834 27588 5010
rect 27622 4834 27634 5010
rect 27576 4822 27634 4834
rect 27706 4834 27718 5210
rect 27752 4834 27764 5210
rect 27706 4822 27764 4834
rect 27824 5210 27882 5222
rect 27824 4834 27836 5210
rect 27870 4834 27882 5210
rect 27824 4822 27882 4834
rect 27942 5210 28000 5222
rect 27942 4834 27954 5210
rect 27988 4834 28000 5210
rect 27942 4822 28000 4834
rect 28060 5210 28118 5222
rect 28060 4834 28072 5210
rect 28106 4834 28118 5210
rect 28060 4822 28118 4834
rect 28178 5210 28236 5222
rect 28178 4834 28190 5210
rect 28224 4834 28236 5210
rect 28178 4822 28236 4834
rect 28296 5210 28354 5222
rect 28296 4834 28308 5210
rect 28342 4834 28354 5210
rect 28296 4822 28354 4834
rect 28414 5210 28472 5222
rect 28414 4834 28426 5210
rect 28460 4834 28472 5210
rect 36751 5308 36763 5342
rect 37139 5308 37151 5342
rect 36751 5296 37151 5308
rect 36751 5224 37151 5236
rect 36751 5190 36763 5224
rect 37139 5190 37151 5224
rect 36751 5178 37151 5190
rect 28414 4822 28472 4834
rect 28543 5010 28601 5022
rect 28543 4834 28555 5010
rect 28589 4834 28601 5010
rect 28543 4822 28601 4834
rect 28661 5010 28719 5022
rect 28661 4834 28673 5010
rect 28707 4834 28719 5010
rect 28661 4822 28719 4834
rect 28779 5010 28837 5022
rect 28779 4834 28791 5010
rect 28825 4834 28837 5010
rect 28779 4822 28837 4834
rect 28897 5010 28955 5022
rect 28897 4834 28909 5010
rect 28943 4834 28955 5010
rect 28897 4822 28955 4834
rect 36751 5106 37151 5118
rect 36751 5072 36763 5106
rect 37139 5072 37151 5106
rect 36751 5060 37151 5072
rect 36751 4988 37151 5000
rect 36751 4954 36763 4988
rect 37139 4954 37151 4988
rect 36751 4942 37151 4954
rect 21027 4516 21085 4528
rect 21027 4140 21039 4516
rect 21073 4140 21085 4516
rect 21027 4128 21085 4140
rect 21145 4516 21203 4528
rect 21145 4140 21157 4516
rect 21191 4140 21203 4516
rect 21145 4128 21203 4140
rect 21263 4516 21321 4528
rect 21263 4140 21275 4516
rect 21309 4140 21321 4516
rect 21263 4128 21321 4140
rect 21381 4516 21439 4528
rect 21381 4140 21393 4516
rect 21427 4140 21439 4516
rect 21381 4128 21439 4140
rect 21499 4516 21557 4528
rect 21499 4140 21511 4516
rect 21545 4140 21557 4516
rect 21499 4128 21557 4140
rect 21617 4516 21675 4528
rect 21617 4140 21629 4516
rect 21663 4140 21675 4516
rect 21617 4128 21675 4140
rect 21735 4516 21793 4528
rect 21735 4140 21747 4516
rect 21781 4140 21793 4516
rect 21735 4128 21793 4140
rect 23855 4023 23913 4035
rect 23855 3847 23867 4023
rect 23901 3847 23913 4023
rect 23855 3835 23913 3847
rect 23973 4023 24031 4035
rect 23973 3847 23985 4023
rect 24019 3847 24031 4023
rect 23973 3835 24031 3847
rect 24091 4023 24149 4035
rect 24091 3847 24103 4023
rect 24137 3847 24149 4023
rect 24091 3835 24149 3847
rect 24209 4023 24267 4035
rect 24209 3847 24221 4023
rect 24255 3847 24267 4023
rect 24209 3835 24267 3847
rect 24327 4023 24385 4035
rect 24327 3847 24339 4023
rect 24373 3847 24385 4023
rect 24327 3835 24385 3847
rect 24445 4023 24503 4035
rect 24445 3847 24457 4023
rect 24491 3847 24503 4023
rect 24445 3835 24503 3847
rect 24563 4023 24621 4035
rect 24563 3847 24575 4023
rect 24609 3847 24621 4023
rect 24563 3835 24621 3847
rect 24681 4023 24739 4035
rect 24681 3847 24693 4023
rect 24727 3847 24739 4023
rect 24681 3835 24739 3847
rect 24799 4023 24857 4035
rect 24799 3847 24811 4023
rect 24845 3847 24857 4023
rect 24799 3835 24857 3847
rect 24917 4023 24975 4035
rect 24917 3847 24929 4023
rect 24963 3847 24975 4023
rect 24917 3835 24975 3847
rect 25751 4517 25809 4529
rect 25751 4141 25763 4517
rect 25797 4141 25809 4517
rect 25751 4129 25809 4141
rect 25869 4517 25927 4529
rect 25869 4141 25881 4517
rect 25915 4141 25927 4517
rect 25869 4129 25927 4141
rect 25987 4517 26045 4529
rect 25987 4141 25999 4517
rect 26033 4141 26045 4517
rect 25987 4129 26045 4141
rect 26105 4517 26163 4529
rect 26105 4141 26117 4517
rect 26151 4141 26163 4517
rect 26105 4129 26163 4141
rect 26223 4517 26281 4529
rect 26223 4141 26235 4517
rect 26269 4141 26281 4517
rect 26223 4129 26281 4141
rect 26341 4517 26399 4529
rect 26341 4141 26353 4517
rect 26387 4141 26399 4517
rect 26341 4129 26399 4141
rect 26459 4517 26517 4529
rect 26459 4141 26471 4517
rect 26505 4141 26517 4517
rect 26459 4129 26517 4141
rect -3113 3063 -2713 3075
rect -3113 3029 -3101 3063
rect -2725 3029 -2713 3063
rect -3806 3006 -3406 3018
rect -3113 3017 -2713 3029
rect -3806 2972 -3794 3006
rect -3418 2972 -3406 3006
rect -3806 2960 -3406 2972
rect -3806 2888 -3406 2900
rect -3806 2854 -3794 2888
rect -3418 2854 -3406 2888
rect -3806 2842 -3406 2854
rect -3806 2770 -3406 2782
rect -3806 2736 -3794 2770
rect -3418 2736 -3406 2770
rect -3806 2724 -3406 2736
rect -3113 2945 -2713 2957
rect -3113 2911 -3101 2945
rect -2725 2911 -2713 2945
rect -3113 2899 -2713 2911
rect 36751 4870 37151 4882
rect 36751 4836 36763 4870
rect 37139 4836 37151 4870
rect 36751 4824 37151 4836
rect 36751 4752 37151 4764
rect 36751 4718 36763 4752
rect 37139 4718 37151 4752
rect 36751 4706 37151 4718
rect 36751 4634 37151 4646
rect 36751 4600 36763 4634
rect 37139 4600 37151 4634
rect 36751 4588 37151 4600
rect 27649 4517 27707 4529
rect 27649 4141 27661 4517
rect 27695 4141 27707 4517
rect 27649 4129 27707 4141
rect 27767 4517 27825 4529
rect 27767 4141 27779 4517
rect 27813 4141 27825 4517
rect 27767 4129 27825 4141
rect 27885 4517 27943 4529
rect 27885 4141 27897 4517
rect 27931 4141 27943 4517
rect 27885 4129 27943 4141
rect 28003 4517 28061 4529
rect 28003 4141 28015 4517
rect 28049 4141 28061 4517
rect 28003 4129 28061 4141
rect 28121 4517 28179 4529
rect 28121 4141 28133 4517
rect 28167 4141 28179 4517
rect 28121 4129 28179 4141
rect 28239 4517 28297 4529
rect 28239 4141 28251 4517
rect 28285 4141 28297 4517
rect 28239 4129 28297 4141
rect 28357 4517 28415 4529
rect 28357 4141 28369 4517
rect 28403 4141 28415 4517
rect 28357 4129 28415 4141
rect 36751 4515 37151 4527
rect 29719 4483 29777 4495
rect 29719 4307 29731 4483
rect 29765 4307 29777 4483
rect 29719 4295 29777 4307
rect 29837 4483 29895 4495
rect 29837 4307 29849 4483
rect 29883 4307 29895 4483
rect 29837 4295 29895 4307
rect 29955 4483 30013 4495
rect 29955 4307 29967 4483
rect 30001 4307 30013 4483
rect 29955 4295 30013 4307
rect 30073 4483 30131 4495
rect 30073 4307 30085 4483
rect 30119 4307 30131 4483
rect 30073 4295 30131 4307
rect 30191 4483 30249 4495
rect 30191 4307 30203 4483
rect 30237 4307 30249 4483
rect 30191 4295 30249 4307
rect 30309 4483 30367 4495
rect 30309 4307 30321 4483
rect 30355 4307 30367 4483
rect 30309 4295 30367 4307
rect 30427 4483 30485 4495
rect 30427 4307 30439 4483
rect 30473 4307 30485 4483
rect 30427 4295 30485 4307
rect 30545 4483 30603 4495
rect 30545 4307 30557 4483
rect 30591 4307 30603 4483
rect 30545 4295 30603 4307
rect 30663 4483 30721 4495
rect 30663 4307 30675 4483
rect 30709 4307 30721 4483
rect 30663 4295 30721 4307
rect 30781 4483 30839 4495
rect 30781 4307 30793 4483
rect 30827 4307 30839 4483
rect 36751 4481 36763 4515
rect 37139 4481 37151 4515
rect 36751 4469 37151 4481
rect 30781 4295 30839 4307
rect 36751 4397 37151 4409
rect 36751 4363 36763 4397
rect 37139 4363 37151 4397
rect 36751 4351 37151 4363
rect 36751 4279 37151 4291
rect 36751 4245 36763 4279
rect 37139 4245 37151 4279
rect 36751 4233 37151 4245
rect 36751 4161 37151 4173
rect 36751 4127 36763 4161
rect 37139 4127 37151 4161
rect 36751 4115 37151 4127
rect 36951 4042 37151 4054
rect 36951 4008 36963 4042
rect 37139 4008 37151 4042
rect 36951 3996 37151 4008
rect 36951 3924 37151 3936
rect 36951 3890 36963 3924
rect 37139 3890 37151 3924
rect 36951 3878 37151 3890
rect 36951 3806 37151 3818
rect 36951 3772 36963 3806
rect 37139 3772 37151 3806
rect 36951 3760 37151 3772
rect 36951 3688 37151 3700
rect 36951 3654 36963 3688
rect 37139 3654 37151 3688
rect 36951 3642 37151 3654
rect 36951 3106 37151 3118
rect 36951 3072 36963 3106
rect 37139 3072 37151 3106
rect 36951 3060 37151 3072
rect 31950 2938 32008 2950
rect -3113 2827 -2713 2839
rect -3113 2793 -3101 2827
rect -2725 2793 -2713 2827
rect -3113 2781 -2713 2793
rect -3806 2652 -3406 2664
rect -3806 2618 -3794 2652
rect -3418 2618 -3406 2652
rect -3806 2606 -3406 2618
rect -3606 2523 -3406 2535
rect -3606 2489 -3594 2523
rect -3418 2489 -3406 2523
rect -3606 2477 -3406 2489
rect -3113 2709 -2713 2721
rect -3113 2675 -3101 2709
rect -2725 2675 -2713 2709
rect 31466 2738 31524 2750
rect -3113 2663 -2713 2675
rect 31466 2562 31478 2738
rect 31512 2562 31524 2738
rect 31466 2550 31524 2562
rect 31584 2738 31642 2750
rect 31584 2562 31596 2738
rect 31630 2562 31642 2738
rect 31584 2550 31642 2562
rect 31702 2738 31760 2750
rect 31702 2562 31714 2738
rect 31748 2562 31760 2738
rect 31702 2550 31760 2562
rect 31820 2738 31878 2750
rect 31820 2562 31832 2738
rect 31866 2562 31878 2738
rect 31820 2550 31878 2562
rect 31950 2562 31962 2938
rect 31996 2562 32008 2938
rect 31950 2550 32008 2562
rect 32068 2938 32126 2950
rect 32068 2562 32080 2938
rect 32114 2562 32126 2938
rect 32068 2550 32126 2562
rect 32186 2938 32244 2950
rect 32186 2562 32198 2938
rect 32232 2562 32244 2938
rect 32186 2550 32244 2562
rect 32304 2938 32362 2950
rect 32304 2562 32316 2938
rect 32350 2562 32362 2938
rect 32304 2550 32362 2562
rect 32422 2938 32480 2950
rect 32422 2562 32434 2938
rect 32468 2562 32480 2938
rect 32422 2550 32480 2562
rect 32540 2938 32598 2950
rect 32540 2562 32552 2938
rect 32586 2562 32598 2938
rect 32540 2550 32598 2562
rect 32658 2938 32716 2950
rect 32658 2562 32670 2938
rect 32704 2562 32716 2938
rect 36951 2988 37151 3000
rect 36951 2954 36963 2988
rect 37139 2954 37151 2988
rect 36951 2942 37151 2954
rect 36951 2870 37151 2882
rect 36951 2836 36963 2870
rect 37139 2836 37151 2870
rect 36951 2824 37151 2836
rect 32658 2550 32716 2562
rect 32787 2738 32845 2750
rect 32787 2562 32799 2738
rect 32833 2562 32845 2738
rect 32787 2550 32845 2562
rect 32905 2738 32963 2750
rect 32905 2562 32917 2738
rect 32951 2562 32963 2738
rect 32905 2550 32963 2562
rect 33023 2738 33081 2750
rect 33023 2562 33035 2738
rect 33069 2562 33081 2738
rect 33023 2550 33081 2562
rect 33141 2738 33199 2750
rect 36951 2752 37151 2764
rect 33141 2562 33153 2738
rect 33187 2562 33199 2738
rect 33141 2550 33199 2562
rect 33259 2735 33317 2747
rect 33259 2559 33271 2735
rect 33305 2559 33317 2735
rect -3606 2405 -3406 2417
rect -3606 2371 -3594 2405
rect -3418 2371 -3406 2405
rect -3606 2359 -3406 2371
rect -3606 2287 -3406 2299
rect -3606 2253 -3594 2287
rect -3418 2253 -3406 2287
rect 33259 2547 33317 2559
rect 33377 2735 33435 2747
rect 33377 2559 33389 2735
rect 33423 2559 33435 2735
rect 33377 2547 33435 2559
rect 33495 2735 33553 2747
rect 33495 2559 33507 2735
rect 33541 2559 33553 2735
rect 33495 2547 33553 2559
rect 33613 2735 33671 2747
rect 33613 2559 33625 2735
rect 33659 2559 33671 2735
rect 33613 2547 33671 2559
rect 33731 2735 33789 2747
rect 33731 2559 33743 2735
rect 33777 2559 33789 2735
rect 33731 2547 33789 2559
rect 33849 2735 33907 2747
rect 33849 2559 33861 2735
rect 33895 2559 33907 2735
rect 33849 2547 33907 2559
rect 33967 2735 34025 2747
rect 33967 2559 33979 2735
rect 34013 2559 34025 2735
rect 33967 2547 34025 2559
rect 34085 2735 34143 2747
rect 34085 2559 34097 2735
rect 34131 2559 34143 2735
rect 34085 2547 34143 2559
rect 34203 2735 34261 2747
rect 34203 2559 34215 2735
rect 34249 2559 34261 2735
rect 34203 2547 34261 2559
rect 34321 2735 34379 2747
rect 34321 2559 34333 2735
rect 34367 2559 34379 2735
rect 36951 2718 36963 2752
rect 37139 2718 37151 2752
rect 36951 2677 37151 2718
rect 36751 2665 37151 2677
rect 36751 2631 36763 2665
rect 37139 2631 37151 2665
rect 36751 2619 37151 2631
rect 34321 2547 34379 2559
rect -3606 2241 -3406 2253
rect -3606 2169 -3406 2181
rect 31893 2245 31951 2257
rect -3606 2135 -3594 2169
rect -3418 2135 -3406 2169
rect -3606 2123 -3406 2135
rect -3608 1776 -3408 1788
rect -3608 1742 -3596 1776
rect -3420 1742 -3408 1776
rect -3608 1730 -3408 1742
rect -3608 1658 -3408 1670
rect -3608 1624 -3596 1658
rect -3420 1624 -3408 1658
rect -3608 1612 -3408 1624
rect -3608 1540 -3408 1552
rect -3608 1506 -3596 1540
rect -3420 1506 -3408 1540
rect -3608 1494 -3408 1506
rect 29726 1638 29784 1650
rect 7835 1520 7893 1532
rect -3608 1422 -3408 1434
rect -3608 1388 -3596 1422
rect -3420 1388 -3408 1422
rect -3608 1376 -3408 1388
rect -3808 1292 -3408 1304
rect -3808 1258 -3796 1292
rect -3420 1258 -3408 1292
rect -3808 1246 -3408 1258
rect -3115 1349 -2715 1361
rect -3115 1315 -3103 1349
rect -2727 1315 -2715 1349
rect 7835 1344 7847 1520
rect 7881 1344 7893 1520
rect -3115 1303 -2715 1315
rect 7835 1332 7893 1344
rect 7953 1520 8011 1532
rect 7953 1344 7965 1520
rect 7999 1344 8011 1520
rect 7953 1332 8011 1344
rect 8071 1520 8129 1532
rect 8071 1344 8083 1520
rect 8117 1344 8129 1520
rect 8071 1332 8129 1344
rect 8189 1520 8247 1532
rect 8189 1344 8201 1520
rect 8235 1344 8247 1520
rect 8189 1332 8247 1344
rect 8307 1520 8365 1532
rect 8307 1344 8319 1520
rect 8353 1344 8365 1520
rect 8307 1332 8365 1344
rect 8425 1520 8483 1532
rect 8425 1344 8437 1520
rect 8471 1344 8483 1520
rect 8425 1332 8483 1344
rect 8543 1520 8601 1532
rect 8543 1344 8555 1520
rect 8589 1344 8601 1520
rect 8543 1332 8601 1344
rect 8661 1520 8719 1532
rect 8661 1344 8673 1520
rect 8707 1344 8719 1520
rect 8661 1332 8719 1344
rect 8779 1520 8837 1532
rect 8779 1344 8791 1520
rect 8825 1344 8837 1520
rect 8779 1332 8837 1344
rect 8897 1520 8955 1532
rect 8897 1344 8909 1520
rect 8943 1344 8955 1520
rect 8897 1332 8955 1344
rect 14389 1525 14447 1537
rect 14389 1349 14401 1525
rect 14435 1349 14447 1525
rect 14389 1337 14447 1349
rect 14507 1525 14565 1537
rect 14507 1349 14519 1525
rect 14553 1349 14565 1525
rect 14507 1337 14565 1349
rect 14625 1525 14683 1537
rect 14625 1349 14637 1525
rect 14671 1349 14683 1525
rect 14625 1337 14683 1349
rect 14743 1525 14801 1537
rect 14743 1349 14755 1525
rect 14789 1349 14801 1525
rect 14743 1337 14801 1349
rect 14861 1525 14919 1537
rect 14861 1349 14873 1525
rect 14907 1349 14919 1525
rect 14861 1337 14919 1349
rect 14979 1525 15037 1537
rect 14979 1349 14991 1525
rect 15025 1349 15037 1525
rect 14979 1337 15037 1349
rect 15097 1525 15155 1537
rect 15097 1349 15109 1525
rect 15143 1349 15155 1525
rect 15097 1337 15155 1349
rect 15215 1525 15273 1537
rect 15215 1349 15227 1525
rect 15261 1349 15273 1525
rect 15215 1337 15273 1349
rect 15333 1525 15391 1537
rect 15333 1349 15345 1525
rect 15379 1349 15391 1525
rect 15333 1337 15391 1349
rect 15451 1525 15509 1537
rect 15451 1349 15463 1525
rect 15497 1349 15509 1525
rect 15451 1337 15509 1349
rect 21038 1513 21096 1525
rect 21038 1337 21050 1513
rect 21084 1337 21096 1513
rect 21038 1325 21096 1337
rect 21156 1513 21214 1525
rect 21156 1337 21168 1513
rect 21202 1337 21214 1513
rect 21156 1325 21214 1337
rect 21274 1513 21332 1525
rect 21274 1337 21286 1513
rect 21320 1337 21332 1513
rect 21274 1325 21332 1337
rect 21392 1513 21450 1525
rect 21392 1337 21404 1513
rect 21438 1337 21450 1513
rect 21392 1325 21450 1337
rect 21510 1513 21568 1525
rect 21510 1337 21522 1513
rect 21556 1337 21568 1513
rect 21510 1325 21568 1337
rect 21628 1513 21686 1525
rect 21628 1337 21640 1513
rect 21674 1337 21686 1513
rect 21628 1325 21686 1337
rect 21746 1513 21804 1525
rect 21746 1337 21758 1513
rect 21792 1337 21804 1513
rect 21746 1325 21804 1337
rect 21864 1513 21922 1525
rect 21864 1337 21876 1513
rect 21910 1337 21922 1513
rect 21864 1325 21922 1337
rect 21982 1513 22040 1525
rect 21982 1337 21994 1513
rect 22028 1337 22040 1513
rect 21982 1325 22040 1337
rect 22100 1513 22158 1525
rect 22100 1337 22112 1513
rect 22146 1337 22158 1513
rect 29726 1462 29738 1638
rect 29772 1462 29784 1638
rect 29726 1450 29784 1462
rect 29844 1638 29902 1650
rect 29844 1462 29856 1638
rect 29890 1462 29902 1638
rect 29844 1450 29902 1462
rect 29962 1638 30020 1650
rect 29962 1462 29974 1638
rect 30008 1462 30020 1638
rect 29962 1450 30020 1462
rect 30080 1638 30138 1650
rect 30080 1462 30092 1638
rect 30126 1462 30138 1638
rect 30080 1450 30138 1462
rect 30198 1638 30256 1650
rect 30198 1462 30210 1638
rect 30244 1462 30256 1638
rect 30198 1450 30256 1462
rect 30316 1638 30374 1650
rect 30316 1462 30328 1638
rect 30362 1462 30374 1638
rect 30316 1450 30374 1462
rect 30434 1638 30492 1650
rect 30434 1462 30446 1638
rect 30480 1462 30492 1638
rect 30434 1450 30492 1462
rect 30552 1638 30610 1650
rect 30552 1462 30564 1638
rect 30598 1462 30610 1638
rect 30552 1450 30610 1462
rect 30670 1638 30728 1650
rect 30670 1462 30682 1638
rect 30716 1462 30728 1638
rect 30670 1450 30728 1462
rect 30788 1638 30846 1650
rect 30788 1462 30800 1638
rect 30834 1462 30846 1638
rect 31893 1869 31905 2245
rect 31939 1869 31951 2245
rect 31893 1857 31951 1869
rect 32011 2245 32069 2257
rect 32011 1869 32023 2245
rect 32057 1869 32069 2245
rect 32011 1857 32069 1869
rect 32129 2245 32187 2257
rect 32129 1869 32141 2245
rect 32175 1869 32187 2245
rect 32129 1857 32187 1869
rect 32247 2245 32305 2257
rect 32247 1869 32259 2245
rect 32293 1869 32305 2245
rect 32247 1857 32305 1869
rect 32365 2245 32423 2257
rect 32365 1869 32377 2245
rect 32411 1869 32423 2245
rect 32365 1857 32423 1869
rect 32483 2245 32541 2257
rect 32483 1869 32495 2245
rect 32529 1869 32541 2245
rect 32483 1857 32541 1869
rect 32601 2245 32659 2257
rect 32601 1869 32613 2245
rect 32647 1869 32659 2245
rect 32601 1857 32659 1869
rect 36751 2547 37151 2559
rect 36751 2513 36763 2547
rect 37139 2513 37151 2547
rect 36751 2501 37151 2513
rect 36751 2429 37151 2441
rect 36751 2395 36763 2429
rect 37139 2395 37151 2429
rect 36751 2383 37151 2395
rect 36751 2311 37151 2323
rect 36751 2277 36763 2311
rect 37139 2277 37151 2311
rect 36751 2265 37151 2277
rect 36751 2198 37151 2210
rect 36751 2164 36763 2198
rect 37139 2164 37151 2198
rect 36751 2152 37151 2164
rect 36751 2080 37151 2092
rect 36751 2046 36763 2080
rect 37139 2046 37151 2080
rect 36751 2034 37151 2046
rect 36751 1962 37151 1974
rect 36751 1928 36763 1962
rect 37139 1928 37151 1962
rect 36751 1916 37151 1928
rect 36751 1844 37151 1856
rect 36751 1810 36763 1844
rect 37139 1810 37151 1844
rect 36751 1798 37151 1810
rect 36751 1726 37151 1738
rect 36751 1692 36763 1726
rect 37139 1692 37151 1726
rect 36751 1680 37151 1692
rect 36751 1608 37151 1620
rect 36751 1574 36763 1608
rect 37139 1574 37151 1608
rect 36751 1562 37151 1574
rect 30788 1450 30846 1462
rect 22100 1325 22158 1337
rect -3808 1174 -3408 1186
rect -3808 1140 -3796 1174
rect -3420 1140 -3408 1174
rect -3808 1128 -3408 1140
rect -3115 1231 -2715 1243
rect -3115 1197 -3103 1231
rect -2727 1197 -2715 1231
rect -3115 1185 -2715 1197
rect -3808 1056 -3408 1068
rect -3808 1022 -3796 1056
rect -3420 1022 -3408 1056
rect -3808 1010 -3408 1022
rect -3115 1113 -2715 1125
rect -3115 1079 -3103 1113
rect -2727 1079 -2715 1113
rect -3115 1067 -2715 1079
rect -3115 995 -2715 1007
rect -3115 961 -3103 995
rect -2727 961 -2715 995
rect -3808 938 -3408 950
rect -3115 949 -2715 961
rect -3808 904 -3796 938
rect -3420 904 -3408 938
rect -3808 892 -3408 904
rect -3808 820 -3408 832
rect -3808 786 -3796 820
rect -3420 786 -3408 820
rect -3808 774 -3408 786
rect -3808 702 -3408 714
rect -3808 668 -3796 702
rect -3420 668 -3408 702
rect -3808 656 -3408 668
rect -3115 877 -2715 889
rect -3115 843 -3103 877
rect -2727 843 -2715 877
rect -3115 831 -2715 843
rect 36751 1490 37151 1502
rect 36751 1456 36763 1490
rect 37139 1456 37151 1490
rect 36751 1444 37151 1456
rect 36751 1371 37151 1383
rect 36751 1337 36763 1371
rect 37139 1337 37151 1371
rect 36751 1325 37151 1337
rect 36751 1253 37151 1265
rect 36751 1219 36763 1253
rect 37139 1219 37151 1253
rect 36751 1207 37151 1219
rect 36751 1135 37151 1147
rect 36751 1101 36763 1135
rect 37139 1101 37151 1135
rect 36751 1089 37151 1101
rect 36751 1017 37151 1029
rect 36751 983 36763 1017
rect 37139 983 37151 1017
rect 36751 971 37151 983
rect 36951 898 37151 910
rect 36951 864 36963 898
rect 37139 864 37151 898
rect 36951 852 37151 864
rect -3115 759 -2715 771
rect -3115 725 -3103 759
rect -2727 725 -2715 759
rect -3115 713 -2715 725
rect 36951 780 37151 792
rect 36951 746 36963 780
rect 37139 746 37151 780
rect 36951 734 37151 746
rect -3808 584 -3408 596
rect -3808 550 -3796 584
rect -3420 550 -3408 584
rect -3808 538 -3408 550
rect -3608 455 -3408 467
rect -3608 421 -3596 455
rect -3420 421 -3408 455
rect -3608 409 -3408 421
rect -3115 641 -2715 653
rect -3115 607 -3103 641
rect -2727 607 -2715 641
rect -3115 595 -2715 607
rect 36951 662 37151 674
rect 36951 628 36963 662
rect 37139 628 37151 662
rect 36951 616 37151 628
rect 36951 544 37151 556
rect 36951 510 36963 544
rect 37139 510 37151 544
rect 36951 498 37151 510
rect -3608 337 -3408 349
rect -3608 303 -3596 337
rect -3420 303 -3408 337
rect -3608 291 -3408 303
rect -3608 219 -3408 231
rect -3608 185 -3596 219
rect -3420 185 -3408 219
rect -3608 173 -3408 185
rect -3608 101 -3408 113
rect -3608 67 -3596 101
rect -3420 67 -3408 101
rect -3608 55 -3408 67
<< ndiffc >>
rect 6079 26795 6113 27171
rect 6197 26795 6231 27171
rect 6315 26795 6349 27171
rect 6432 26995 6466 27171
rect 6550 26995 6584 27171
rect 8077 26721 8111 26897
rect 8195 26721 8229 26897
rect 8313 26721 8347 26897
rect 8431 26721 8465 26897
rect 9219 26725 9253 26901
rect 9337 26725 9371 26901
rect 9455 26725 9489 26901
rect 9573 26725 9607 26901
rect 12592 26792 12626 27168
rect 12710 26792 12744 27168
rect 12828 26792 12862 27168
rect 12945 26992 12979 27168
rect 13063 26992 13097 27168
rect 14590 26718 14624 26894
rect 14708 26718 14742 26894
rect 14826 26718 14860 26894
rect 14944 26718 14978 26894
rect 15732 26722 15766 26898
rect 15850 26722 15884 26898
rect 15968 26722 16002 26898
rect 16086 26722 16120 26898
rect 19126 26787 19160 27163
rect 19244 26787 19278 27163
rect 19362 26787 19396 27163
rect 19479 26987 19513 27163
rect 19597 26987 19631 27163
rect 21124 26713 21158 26889
rect 21242 26713 21276 26889
rect 21360 26713 21394 26889
rect 21478 26713 21512 26889
rect 22266 26717 22300 26893
rect 22384 26717 22418 26893
rect 22502 26717 22536 26893
rect 22620 26717 22654 26893
rect 25684 26791 25718 27167
rect 25802 26791 25836 27167
rect 25920 26791 25954 27167
rect 26037 26991 26071 27167
rect 26155 26991 26189 27167
rect 27682 26717 27716 26893
rect 27800 26717 27834 26893
rect 27918 26717 27952 26893
rect 28036 26717 28070 26893
rect 28824 26721 28858 26897
rect 28942 26721 28976 26897
rect 29060 26721 29094 26897
rect 29178 26721 29212 26897
rect 6093 25145 6127 25521
rect 6211 25145 6245 25521
rect 6329 25145 6363 25521
rect 6446 25345 6480 25521
rect 6564 25345 6598 25521
rect 12606 25142 12640 25518
rect 12724 25142 12758 25518
rect 12842 25142 12876 25518
rect 12959 25342 12993 25518
rect 13077 25342 13111 25518
rect 7445 23940 7479 24116
rect 6088 23541 6122 23917
rect 6206 23541 6240 23917
rect 6324 23541 6358 23917
rect 6441 23741 6475 23917
rect 7563 23940 7597 24116
rect 6559 23741 6593 23917
rect 7865 23740 7899 24116
rect 7983 23740 8017 24116
rect 8101 23740 8135 24116
rect 8219 23740 8253 24116
rect 8337 23740 8371 24116
rect 8743 23940 8777 24116
rect 8861 23940 8895 24116
rect 9343 23940 9377 24116
rect 9461 23940 9495 24116
rect 9763 23740 9797 24116
rect 9881 23740 9915 24116
rect 9999 23740 10033 24116
rect 10117 23740 10151 24116
rect 10235 23740 10269 24116
rect 10641 23940 10675 24116
rect 10759 23940 10793 24116
rect 19140 25137 19174 25513
rect 19258 25137 19292 25513
rect 19376 25137 19410 25513
rect 19493 25337 19527 25513
rect 19611 25337 19645 25513
rect 13958 23937 13992 24113
rect 12601 23538 12635 23914
rect 12719 23538 12753 23914
rect 12837 23538 12871 23914
rect 12954 23738 12988 23914
rect 14076 23937 14110 24113
rect 13072 23738 13106 23914
rect 14378 23737 14412 24113
rect 14496 23737 14530 24113
rect 14614 23737 14648 24113
rect 14732 23737 14766 24113
rect 14850 23737 14884 24113
rect 15256 23937 15290 24113
rect 15374 23937 15408 24113
rect 15856 23937 15890 24113
rect 15974 23937 16008 24113
rect 16276 23737 16310 24113
rect 16394 23737 16428 24113
rect 16512 23737 16546 24113
rect 16630 23737 16664 24113
rect 16748 23737 16782 24113
rect 17154 23937 17188 24113
rect 17272 23937 17306 24113
rect 25698 25141 25732 25517
rect 25816 25141 25850 25517
rect 25934 25141 25968 25517
rect 26051 25341 26085 25517
rect 26169 25341 26203 25517
rect 20492 23932 20526 24108
rect 19135 23533 19169 23909
rect 19253 23533 19287 23909
rect 19371 23533 19405 23909
rect 19488 23733 19522 23909
rect 20610 23932 20644 24108
rect 19606 23733 19640 23909
rect 20912 23732 20946 24108
rect 21030 23732 21064 24108
rect 21148 23732 21182 24108
rect 21266 23732 21300 24108
rect 21384 23732 21418 24108
rect 21790 23932 21824 24108
rect 21908 23932 21942 24108
rect 22390 23932 22424 24108
rect 22508 23932 22542 24108
rect 22810 23732 22844 24108
rect 22928 23732 22962 24108
rect 23046 23732 23080 24108
rect 23164 23732 23198 24108
rect 23282 23732 23316 24108
rect 23688 23932 23722 24108
rect 23806 23932 23840 24108
rect 27050 23936 27084 24112
rect 25693 23537 25727 23913
rect 25811 23537 25845 23913
rect 25929 23537 25963 23913
rect 26046 23737 26080 23913
rect 27168 23936 27202 24112
rect 26164 23737 26198 23913
rect 27470 23736 27504 24112
rect 27588 23736 27622 24112
rect 27706 23736 27740 24112
rect 27824 23736 27858 24112
rect 27942 23736 27976 24112
rect 28348 23936 28382 24112
rect 28466 23936 28500 24112
rect 28948 23936 28982 24112
rect 29066 23936 29100 24112
rect 29368 23736 29402 24112
rect 29486 23736 29520 24112
rect 29604 23736 29638 24112
rect 29722 23736 29756 24112
rect 29840 23736 29874 24112
rect 30246 23936 30280 24112
rect 30364 23936 30398 24112
rect 38100 24280 38276 24314
rect 38100 24162 38276 24196
rect 38100 24088 38476 24122
rect 38100 23970 38476 24004
rect 38100 23852 38476 23886
rect 38100 23734 38476 23768
rect 38100 23616 38476 23650
rect 38100 23538 38276 23572
rect 38100 23420 38276 23454
rect 6297 21117 6331 21293
rect 6415 21117 6449 21293
rect 6533 21117 6567 21293
rect 9320 21387 9354 21563
rect 9438 21387 9472 21563
rect 6651 21117 6685 21293
rect 7439 21113 7473 21289
rect 7557 21113 7591 21289
rect 7675 21113 7709 21289
rect 7793 21113 7827 21289
rect 9555 21187 9589 21563
rect 9673 21187 9707 21563
rect 9791 21187 9825 21563
rect 12855 21113 12889 21289
rect 12973 21113 13007 21289
rect 13091 21113 13125 21289
rect 15878 21383 15912 21559
rect 15996 21383 16030 21559
rect 13209 21113 13243 21289
rect 13997 21109 14031 21285
rect 14115 21109 14149 21285
rect 14233 21109 14267 21285
rect 14351 21109 14385 21285
rect 16113 21183 16147 21559
rect 16231 21183 16265 21559
rect 16349 21183 16383 21559
rect 19389 21118 19423 21294
rect 19507 21118 19541 21294
rect 19625 21118 19659 21294
rect 22412 21388 22446 21564
rect 22530 21388 22564 21564
rect 19743 21118 19777 21294
rect 20531 21114 20565 21290
rect 20649 21114 20683 21290
rect 20767 21114 20801 21290
rect 20885 21114 20919 21290
rect 22647 21188 22681 21564
rect 22765 21188 22799 21564
rect 22883 21188 22917 21564
rect 25902 21121 25936 21297
rect 26020 21121 26054 21297
rect 26138 21121 26172 21297
rect 28925 21391 28959 21567
rect 29043 21391 29077 21567
rect 26256 21121 26290 21297
rect 27044 21117 27078 21293
rect 27162 21117 27196 21293
rect 27280 21117 27314 21293
rect 27398 21117 27432 21293
rect 29160 21191 29194 21567
rect 29278 21191 29312 21567
rect 29396 21191 29430 21567
rect 38100 21136 38276 21170
rect 38100 21018 38276 21052
rect 38100 20944 38476 20978
rect 38100 20826 38476 20860
rect 38100 20708 38476 20742
rect 38100 20590 38476 20624
rect 9306 19737 9340 19913
rect 9424 19737 9458 19913
rect 9541 19537 9575 19913
rect 9659 19537 9693 19913
rect 9777 19537 9811 19913
rect 15864 19733 15898 19909
rect 15982 19733 16016 19909
rect 5111 18332 5145 18508
rect 5229 18332 5263 18508
rect 5635 18132 5669 18508
rect 5753 18132 5787 18508
rect 5871 18132 5905 18508
rect 5989 18132 6023 18508
rect 6107 18132 6141 18508
rect 6409 18332 6443 18508
rect 6527 18332 6561 18508
rect 7009 18332 7043 18508
rect 7127 18332 7161 18508
rect 7533 18132 7567 18508
rect 7651 18132 7685 18508
rect 7769 18132 7803 18508
rect 7887 18132 7921 18508
rect 8005 18132 8039 18508
rect 8307 18332 8341 18508
rect 8425 18332 8459 18508
rect 16099 19533 16133 19909
rect 16217 19533 16251 19909
rect 16335 19533 16369 19909
rect 22398 19738 22432 19914
rect 22516 19738 22550 19914
rect 11669 18328 11703 18504
rect 9311 18133 9345 18309
rect 9429 18133 9463 18309
rect 9546 17933 9580 18309
rect 9664 17933 9698 18309
rect 11787 18328 11821 18504
rect 9782 17933 9816 18309
rect 12193 18128 12227 18504
rect 12311 18128 12345 18504
rect 12429 18128 12463 18504
rect 12547 18128 12581 18504
rect 12665 18128 12699 18504
rect 12967 18328 13001 18504
rect 13085 18328 13119 18504
rect 13567 18328 13601 18504
rect 13685 18328 13719 18504
rect 14091 18128 14125 18504
rect 14209 18128 14243 18504
rect 14327 18128 14361 18504
rect 14445 18128 14479 18504
rect 14563 18128 14597 18504
rect 14865 18328 14899 18504
rect 14983 18328 15017 18504
rect 22633 19538 22667 19914
rect 22751 19538 22785 19914
rect 22869 19538 22903 19914
rect 38100 20472 38476 20506
rect 38100 20394 38276 20428
rect 28911 19741 28945 19917
rect 29029 19741 29063 19917
rect 18203 18333 18237 18509
rect 18321 18333 18355 18509
rect 15869 18129 15903 18305
rect 15987 18129 16021 18305
rect 16104 17929 16138 18305
rect 16222 17929 16256 18305
rect 16340 17929 16374 18305
rect 18727 18133 18761 18509
rect 18845 18133 18879 18509
rect 18963 18133 18997 18509
rect 19081 18133 19115 18509
rect 19199 18133 19233 18509
rect 19501 18333 19535 18509
rect 19619 18333 19653 18509
rect 20101 18333 20135 18509
rect 20219 18333 20253 18509
rect 20625 18133 20659 18509
rect 20743 18133 20777 18509
rect 20861 18133 20895 18509
rect 20979 18133 21013 18509
rect 21097 18133 21131 18509
rect 21399 18333 21433 18509
rect 21517 18333 21551 18509
rect 29146 19541 29180 19917
rect 29264 19541 29298 19917
rect 29382 19541 29416 19917
rect 38100 20276 38276 20310
rect 24716 18336 24750 18512
rect 24834 18336 24868 18512
rect 22403 18134 22437 18310
rect 22521 18134 22555 18310
rect 22638 17934 22672 18310
rect 22756 17934 22790 18310
rect 22874 17934 22908 18310
rect 25240 18136 25274 18512
rect 25358 18136 25392 18512
rect 25476 18136 25510 18512
rect 25594 18136 25628 18512
rect 25712 18136 25746 18512
rect 26014 18336 26048 18512
rect 26132 18336 26166 18512
rect 26614 18336 26648 18512
rect 26732 18336 26766 18512
rect 27138 18136 27172 18512
rect 27256 18136 27290 18512
rect 27374 18136 27408 18512
rect 27492 18136 27526 18512
rect 27610 18136 27644 18512
rect 27912 18336 27946 18512
rect 28030 18336 28064 18512
rect 28916 18137 28950 18313
rect 29034 18137 29068 18313
rect 29151 17937 29185 18313
rect 29269 17937 29303 18313
rect 29387 17937 29421 18313
rect 38096 18004 38272 18038
rect 38096 17886 38272 17920
rect 38096 17812 38472 17846
rect 38096 17694 38472 17728
rect 38096 17576 38472 17610
rect 38096 17458 38472 17492
rect 38096 17340 38472 17374
rect 38096 17262 38272 17296
rect 38096 17144 38272 17178
rect -2367 16096 -2191 16130
rect -2367 15978 -2191 16012
rect -2367 15676 -1991 15710
rect -2367 15558 -1991 15592
rect -2367 15440 -1991 15474
rect -2367 15322 -1991 15356
rect -2367 15204 -1991 15238
rect -2367 14798 -2191 14832
rect -2367 14680 -2191 14714
rect 8049 14411 8083 14787
rect 8167 14411 8201 14787
rect 8285 14411 8319 14787
rect 8402 14611 8436 14787
rect 8520 14611 8554 14787
rect 14598 14410 14632 14786
rect 14716 14410 14750 14786
rect 14834 14410 14868 14786
rect 14951 14610 14985 14786
rect 15069 14610 15103 14786
rect 21252 14431 21286 14807
rect 21370 14431 21404 14807
rect 21488 14431 21522 14807
rect 21605 14631 21639 14807
rect 21723 14631 21757 14807
rect 29905 14264 29939 14640
rect 30023 14264 30057 14640
rect 30141 14264 30175 14640
rect 30258 14464 30292 14640
rect 30376 14464 30410 14640
rect 38096 14860 38272 14894
rect 38096 14742 38272 14776
rect 38096 14668 38472 14702
rect -2369 14028 -2193 14062
rect -2369 13910 -2193 13944
rect -2369 13608 -1993 13642
rect -2369 13490 -1993 13524
rect -2369 13372 -1993 13406
rect -2369 13254 -1993 13288
rect -2369 13136 -1993 13170
rect 38096 14550 38472 14584
rect 38096 14432 38472 14466
rect 38096 14314 38472 14348
rect 33506 13856 33540 14232
rect 33624 13856 33658 14232
rect 33742 13856 33776 14232
rect 33859 14056 33893 14232
rect 33977 14056 34011 14232
rect 38096 14196 38472 14230
rect 38096 14118 38272 14152
rect -2369 12730 -2193 12764
rect -2369 12612 -2193 12646
rect 1385 12511 1419 12887
rect 1503 12511 1537 12887
rect 1621 12511 1655 12887
rect 1738 12711 1772 12887
rect 1856 12711 1890 12887
rect 4275 12244 4309 12620
rect 4393 12244 4427 12620
rect 4511 12244 4545 12620
rect 4628 12444 4662 12620
rect 4746 12444 4780 12620
rect 31601 13271 31635 13447
rect 31719 13271 31753 13447
rect 6273 12170 6307 12346
rect 6391 12170 6425 12346
rect 6509 12170 6543 12346
rect 6627 12170 6661 12346
rect 7415 12174 7449 12350
rect 7533 12174 7567 12350
rect 7651 12174 7685 12350
rect 7769 12174 7803 12350
rect 10824 12332 10858 12708
rect 10942 12332 10976 12708
rect 11060 12332 11094 12708
rect 11177 12532 11211 12708
rect 11295 12532 11329 12708
rect 12822 12258 12856 12434
rect 12940 12258 12974 12434
rect 13058 12258 13092 12434
rect 13176 12258 13210 12434
rect 13964 12262 13998 12438
rect 14082 12262 14116 12438
rect 14200 12262 14234 12438
rect 14318 12262 14352 12438
rect 17478 12264 17512 12640
rect 17596 12264 17630 12640
rect 17714 12264 17748 12640
rect 17831 12464 17865 12640
rect 17949 12464 17983 12640
rect 32021 13071 32055 13447
rect 32139 13071 32173 13447
rect 32257 13071 32291 13447
rect 32375 13071 32409 13447
rect 32493 13071 32527 13447
rect 32899 13271 32933 13447
rect 33017 13271 33051 13447
rect 38096 14000 38272 14034
rect 19476 12190 19510 12366
rect 19594 12190 19628 12366
rect 19712 12190 19746 12366
rect 19830 12190 19864 12366
rect 20618 12194 20652 12370
rect 20736 12194 20770 12370
rect 20854 12194 20888 12370
rect 20972 12194 21006 12370
rect 24103 12332 24137 12708
rect 24221 12332 24255 12708
rect 24339 12332 24373 12708
rect 24456 12532 24490 12708
rect 24574 12532 24608 12708
rect 26101 12258 26135 12434
rect 26219 12258 26253 12434
rect 26337 12258 26371 12434
rect 26455 12258 26489 12434
rect 27243 12262 27277 12438
rect 27361 12262 27395 12438
rect 27479 12262 27513 12438
rect 27597 12262 27631 12438
rect -2367 11959 -2191 11993
rect -2367 11841 -2191 11875
rect 29900 11693 29934 12069
rect 30018 11693 30052 12069
rect 30136 11693 30170 12069
rect 30253 11893 30287 12069
rect 30371 11893 30405 12069
rect -2367 11539 -1991 11573
rect -2367 11421 -1991 11455
rect -2367 11303 -1991 11337
rect -2367 11185 -1991 11219
rect -2367 11067 -1991 11101
rect 38100 11658 38276 11692
rect 38100 11540 38276 11574
rect 38100 11466 38476 11500
rect -2367 10661 -2191 10695
rect -2367 10543 -2191 10577
rect 4289 10594 4323 10970
rect 4407 10594 4441 10970
rect 4525 10594 4559 10970
rect 4642 10794 4676 10970
rect 4760 10794 4794 10970
rect 10838 10682 10872 11058
rect 10956 10682 10990 11058
rect 11074 10682 11108 11058
rect 11191 10882 11225 11058
rect 11309 10882 11343 11058
rect -2369 9891 -2193 9925
rect 1377 9926 1411 10302
rect 1495 9926 1529 10302
rect 1613 9926 1647 10302
rect 1730 10126 1764 10302
rect 1848 10126 1882 10302
rect -2369 9773 -2193 9807
rect -2369 9471 -1993 9505
rect -2369 9353 -1993 9387
rect 38100 11348 38476 11382
rect 38100 11230 38476 11264
rect 38100 11112 38476 11146
rect 5641 9389 5675 9565
rect -2369 9235 -1993 9269
rect -2369 9117 -1993 9151
rect -2369 8999 -1993 9033
rect 4284 8990 4318 9366
rect 4402 8990 4436 9366
rect 4520 8990 4554 9366
rect 4637 9190 4671 9366
rect 5759 9389 5793 9565
rect 4755 9190 4789 9366
rect 6061 9189 6095 9565
rect 6179 9189 6213 9565
rect 6297 9189 6331 9565
rect 6415 9189 6449 9565
rect 6533 9189 6567 9565
rect 6939 9389 6973 9565
rect 7057 9389 7091 9565
rect 7539 9389 7573 9565
rect 7657 9389 7691 9565
rect 7959 9189 7993 9565
rect 8077 9189 8111 9565
rect 8195 9189 8229 9565
rect 8313 9189 8347 9565
rect 8431 9189 8465 9565
rect 8837 9389 8871 9565
rect 8955 9389 8989 9565
rect 17492 10614 17526 10990
rect 17610 10614 17644 10990
rect 17728 10614 17762 10990
rect 17845 10814 17879 10990
rect 17963 10814 17997 10990
rect 24117 10682 24151 11058
rect 24235 10682 24269 11058
rect 24353 10682 24387 11058
rect 24470 10882 24504 11058
rect 24588 10882 24622 11058
rect 12190 9477 12224 9653
rect 10833 9078 10867 9454
rect 10951 9078 10985 9454
rect 11069 9078 11103 9454
rect 11186 9278 11220 9454
rect 12308 9477 12342 9653
rect 11304 9278 11338 9454
rect 12610 9277 12644 9653
rect 12728 9277 12762 9653
rect 12846 9277 12880 9653
rect 12964 9277 12998 9653
rect 13082 9277 13116 9653
rect 13488 9477 13522 9653
rect 13606 9477 13640 9653
rect 14088 9477 14122 9653
rect 14206 9477 14240 9653
rect 14508 9277 14542 9653
rect 14626 9277 14660 9653
rect 14744 9277 14778 9653
rect 14862 9277 14896 9653
rect 14980 9277 15014 9653
rect 15386 9477 15420 9653
rect 15504 9477 15538 9653
rect 18844 9409 18878 9585
rect 17487 9010 17521 9386
rect 17605 9010 17639 9386
rect 17723 9010 17757 9386
rect 17840 9210 17874 9386
rect 18962 9409 18996 9585
rect 17958 9210 17992 9386
rect 19264 9209 19298 9585
rect 19382 9209 19416 9585
rect 19500 9209 19534 9585
rect 19618 9209 19652 9585
rect 19736 9209 19770 9585
rect 20142 9409 20176 9585
rect 20260 9409 20294 9585
rect 20742 9409 20776 9585
rect 20860 9409 20894 9585
rect 21162 9209 21196 9585
rect 21280 9209 21314 9585
rect 21398 9209 21432 9585
rect 21516 9209 21550 9585
rect 21634 9209 21668 9585
rect 22040 9409 22074 9585
rect 22158 9409 22192 9585
rect 38100 10994 38476 11028
rect 38100 10916 38276 10950
rect 25469 9477 25503 9653
rect 24112 9078 24146 9454
rect 24230 9078 24264 9454
rect 24348 9078 24382 9454
rect 24465 9278 24499 9454
rect 25587 9477 25621 9653
rect 24583 9278 24617 9454
rect 25889 9277 25923 9653
rect 26007 9277 26041 9653
rect 26125 9277 26159 9653
rect 26243 9277 26277 9653
rect 26361 9277 26395 9653
rect 26767 9477 26801 9653
rect 26885 9477 26919 9653
rect 27367 9477 27401 9653
rect 27485 9477 27519 9653
rect 27787 9277 27821 9653
rect 27905 9277 27939 9653
rect 28023 9277 28057 9653
rect 28141 9277 28175 9653
rect 28259 9277 28293 9653
rect 28665 9477 28699 9653
rect 28783 9477 28817 9653
rect 33508 9765 33542 10141
rect 33626 9765 33660 10141
rect 33744 9765 33778 10141
rect 33861 9965 33895 10141
rect 33979 9965 34013 10141
rect 38100 10798 38276 10832
rect 31603 9180 31637 9356
rect 31721 9180 31755 9356
rect 29900 8660 29934 9036
rect 30018 8660 30052 9036
rect 30136 8660 30170 9036
rect 30253 8860 30287 9036
rect 30371 8860 30405 9036
rect 32023 8980 32057 9356
rect 32141 8980 32175 9356
rect 32259 8980 32293 9356
rect 32377 8980 32411 9356
rect 32495 8980 32529 9356
rect 32901 9180 32935 9356
rect 33019 9180 33053 9356
rect -2369 8593 -2193 8627
rect -2369 8475 -2193 8509
rect 38100 8514 38276 8548
rect 38100 8396 38276 8430
rect 38100 8322 38476 8356
rect 38100 8204 38476 8238
rect 38100 8086 38476 8120
rect 38100 7968 38476 8002
rect -2369 7822 -2193 7856
rect -2369 7704 -2193 7738
rect -2369 7402 -1993 7436
rect -2369 7284 -1993 7318
rect -2369 7166 -1993 7200
rect -2369 7048 -1993 7082
rect -2369 6930 -1993 6964
rect 1358 6648 1392 7024
rect 1476 6648 1510 7024
rect 1594 6648 1628 7024
rect 1711 6848 1745 7024
rect 1829 6848 1863 7024
rect -2369 6524 -2193 6558
rect -2369 6406 -2193 6440
rect 4267 6464 4301 6840
rect 4385 6464 4419 6840
rect 4503 6464 4537 6840
rect 4620 6664 4654 6840
rect 4738 6664 4772 6840
rect 6265 6390 6299 6566
rect 6383 6390 6417 6566
rect 6501 6390 6535 6566
rect 6619 6390 6653 6566
rect 7407 6394 7441 6570
rect 7525 6394 7559 6570
rect 7643 6394 7677 6570
rect 7761 6394 7795 6570
rect 10818 6462 10852 6838
rect 10936 6462 10970 6838
rect 11054 6462 11088 6838
rect 11171 6662 11205 6838
rect 11289 6662 11323 6838
rect 38100 7850 38476 7884
rect 38100 7772 38276 7806
rect 12816 6388 12850 6564
rect 12934 6388 12968 6564
rect 13052 6388 13086 6564
rect 13170 6388 13204 6564
rect 13958 6392 13992 6568
rect 14076 6392 14110 6568
rect 14194 6392 14228 6568
rect 14312 6392 14346 6568
rect 17473 6463 17507 6839
rect 17591 6463 17625 6839
rect 17709 6463 17743 6839
rect 17826 6663 17860 6839
rect 17944 6663 17978 6839
rect 19471 6389 19505 6565
rect 19589 6389 19623 6565
rect 19707 6389 19741 6565
rect 19825 6389 19859 6565
rect 20613 6393 20647 6569
rect 20731 6393 20765 6569
rect 20849 6393 20883 6569
rect 20967 6393 21001 6569
rect 24095 6464 24129 6840
rect 24213 6464 24247 6840
rect 24331 6464 24365 6840
rect 24448 6664 24482 6840
rect 24566 6664 24600 6840
rect 29971 6740 30005 7116
rect 30089 6740 30123 7116
rect 30207 6740 30241 7116
rect 30324 6940 30358 7116
rect 30442 6940 30476 7116
rect 26093 6390 26127 6566
rect 26211 6390 26245 6566
rect 26329 6390 26363 6566
rect 26447 6390 26481 6566
rect 27235 6394 27269 6570
rect 27353 6394 27387 6570
rect 27471 6394 27505 6570
rect 27589 6394 27623 6570
rect 38100 7654 38276 7688
rect 33508 6270 33542 6646
rect 33626 6270 33660 6646
rect 33744 6270 33778 6646
rect 33861 6470 33895 6646
rect 33979 6470 34013 6646
rect -2371 5754 -2195 5788
rect -2371 5636 -2195 5670
rect -2371 5334 -1995 5368
rect -2371 5216 -1995 5250
rect 31603 5685 31637 5861
rect 31721 5685 31755 5861
rect 32023 5485 32057 5861
rect 32141 5485 32175 5861
rect 32259 5485 32293 5861
rect 32377 5485 32411 5861
rect 32495 5485 32529 5861
rect 32901 5685 32935 5861
rect 33019 5685 33053 5861
rect -2371 5098 -1995 5132
rect -2371 4980 -1995 5014
rect -2371 4862 -1995 4896
rect 4281 4814 4315 5190
rect 4399 4814 4433 5190
rect 4517 4814 4551 5190
rect 4634 5014 4668 5190
rect 4752 5014 4786 5190
rect -2371 4456 -2195 4490
rect -2371 4338 -2195 4372
rect 1374 3888 1408 4264
rect 1492 3888 1526 4264
rect 1610 3888 1644 4264
rect 1727 4088 1761 4264
rect 1845 4088 1879 4264
rect -2369 3685 -2193 3719
rect -2369 3567 -2193 3601
rect 10832 4812 10866 5188
rect 10950 4812 10984 5188
rect 11068 4812 11102 5188
rect 11185 5012 11219 5188
rect 11303 5012 11337 5188
rect 5633 3609 5667 3785
rect -2369 3265 -1993 3299
rect 4276 3210 4310 3586
rect 4394 3210 4428 3586
rect 4512 3210 4546 3586
rect 4629 3410 4663 3586
rect 5751 3609 5785 3785
rect 4747 3410 4781 3586
rect 6053 3409 6087 3785
rect 6171 3409 6205 3785
rect 6289 3409 6323 3785
rect 6407 3409 6441 3785
rect 6525 3409 6559 3785
rect 6931 3609 6965 3785
rect 7049 3609 7083 3785
rect 7531 3609 7565 3785
rect 7649 3609 7683 3785
rect 7951 3409 7985 3785
rect 8069 3409 8103 3785
rect 8187 3409 8221 3785
rect 8305 3409 8339 3785
rect 8423 3409 8457 3785
rect 8829 3609 8863 3785
rect 8947 3609 8981 3785
rect 17487 4813 17521 5189
rect 17605 4813 17639 5189
rect 17723 4813 17757 5189
rect 17840 5013 17874 5189
rect 17958 5013 17992 5189
rect 12184 3607 12218 3783
rect -2369 3147 -1993 3181
rect 10827 3208 10861 3584
rect 10945 3208 10979 3584
rect 11063 3208 11097 3584
rect 11180 3408 11214 3584
rect 12302 3607 12336 3783
rect 11298 3408 11332 3584
rect 12604 3407 12638 3783
rect 12722 3407 12756 3783
rect 12840 3407 12874 3783
rect 12958 3407 12992 3783
rect 13076 3407 13110 3783
rect 13482 3607 13516 3783
rect 13600 3607 13634 3783
rect 14082 3607 14116 3783
rect 14200 3607 14234 3783
rect 14502 3407 14536 3783
rect 14620 3407 14654 3783
rect 14738 3407 14772 3783
rect 14856 3407 14890 3783
rect 14974 3407 15008 3783
rect 15380 3607 15414 3783
rect 15498 3607 15532 3783
rect 24109 4814 24143 5190
rect 24227 4814 24261 5190
rect 24345 4814 24379 5190
rect 24462 5014 24496 5190
rect 24580 5014 24614 5190
rect 38096 5382 38272 5416
rect 38096 5264 38272 5298
rect 38096 5190 38472 5224
rect 38096 5072 38472 5106
rect 18839 3608 18873 3784
rect -2369 3029 -1993 3063
rect -2369 2911 -1993 2945
rect 17482 3209 17516 3585
rect 17600 3209 17634 3585
rect 17718 3209 17752 3585
rect 17835 3409 17869 3585
rect 18957 3608 18991 3784
rect 17953 3409 17987 3585
rect 19259 3408 19293 3784
rect 19377 3408 19411 3784
rect 19495 3408 19529 3784
rect 19613 3408 19647 3784
rect 19731 3408 19765 3784
rect 20137 3608 20171 3784
rect 20255 3608 20289 3784
rect 20737 3608 20771 3784
rect 20855 3608 20889 3784
rect 21157 3408 21191 3784
rect 21275 3408 21309 3784
rect 21393 3408 21427 3784
rect 21511 3408 21545 3784
rect 21629 3408 21663 3784
rect 22035 3608 22069 3784
rect 22153 3608 22187 3784
rect 38096 4954 38472 4988
rect 38096 4836 38472 4870
rect 38096 4718 38472 4752
rect 38096 4640 38272 4674
rect 25461 3609 25495 3785
rect 24104 3210 24138 3586
rect 24222 3210 24256 3586
rect 24340 3210 24374 3586
rect 24457 3410 24491 3586
rect 25579 3609 25613 3785
rect 24575 3410 24609 3586
rect 25881 3409 25915 3785
rect 25999 3409 26033 3785
rect 26117 3409 26151 3785
rect 26235 3409 26269 3785
rect 26353 3409 26387 3785
rect 26759 3609 26793 3785
rect 26877 3609 26911 3785
rect 27359 3609 27393 3785
rect 27477 3609 27511 3785
rect 27779 3409 27813 3785
rect 27897 3409 27931 3785
rect 28015 3409 28049 3785
rect 28133 3409 28167 3785
rect 28251 3409 28285 3785
rect 28657 3609 28691 3785
rect 28775 3609 28809 3785
rect 29968 3670 30002 4046
rect 30086 3670 30120 4046
rect 30204 3670 30238 4046
rect 30321 3870 30355 4046
rect 30439 3870 30473 4046
rect 38096 4522 38272 4556
rect -2369 2793 -1993 2827
rect -2369 2387 -2193 2421
rect -2369 2269 -2193 2303
rect 8084 1781 8118 2157
rect 8202 1781 8236 2157
rect 8320 1781 8354 2157
rect 8437 1781 8471 1957
rect 8555 1781 8589 1957
rect 14638 1786 14672 2162
rect 14756 1786 14790 2162
rect 14874 1786 14908 2162
rect 14991 1786 15025 1962
rect 15109 1786 15143 1962
rect 21287 1774 21321 2150
rect -2371 1617 -2195 1651
rect -2371 1499 -2195 1533
rect 21405 1774 21439 2150
rect 21523 1774 21557 2150
rect 21640 1774 21674 1950
rect 21758 1774 21792 1950
rect 33508 1922 33542 2298
rect 33626 1922 33660 2298
rect 33744 1922 33778 2298
rect 33861 2122 33895 2298
rect 33979 2122 34013 2298
rect 38096 2238 38272 2272
rect 38096 2120 38272 2154
rect 38096 2046 38472 2080
rect 38096 1928 38472 1962
rect 38096 1810 38472 1844
rect 38096 1692 38472 1726
rect -2371 1197 -1995 1231
rect 31603 1337 31637 1513
rect 31721 1337 31755 1513
rect -2371 1079 -1995 1113
rect -2371 961 -1995 995
rect -2371 843 -1995 877
rect 29975 825 30009 1201
rect 30093 825 30127 1201
rect 30211 825 30245 1201
rect 30328 1025 30362 1201
rect 30446 1025 30480 1201
rect 32023 1137 32057 1513
rect 32141 1137 32175 1513
rect 32259 1137 32293 1513
rect 32377 1137 32411 1513
rect 32495 1137 32529 1513
rect 32901 1337 32935 1513
rect 33019 1337 33053 1513
rect 38096 1574 38472 1608
rect 38096 1496 38272 1530
rect -2371 725 -1995 759
rect 38096 1378 38272 1412
rect -2371 319 -2195 353
rect -2371 201 -2195 235
<< pdiffc >>
rect 5842 27432 5876 27608
rect 5960 27432 5994 27608
rect 6078 27432 6112 27608
rect 6196 27432 6230 27608
rect 6314 27432 6348 27608
rect 6432 27432 6466 27608
rect 6550 27432 6584 27608
rect 6668 27432 6702 27608
rect 6786 27432 6820 27608
rect 6904 27432 6938 27608
rect 8167 27304 8201 27680
rect 8285 27304 8319 27680
rect 8403 27304 8437 27680
rect 8521 27304 8555 27680
rect 8639 27304 8673 27680
rect 8757 27304 8791 27680
rect 8875 27304 8909 27680
rect 9309 27308 9343 27684
rect 9427 27308 9461 27684
rect 9545 27308 9579 27684
rect 9663 27308 9697 27684
rect 9781 27308 9815 27684
rect 9899 27308 9933 27684
rect 10017 27308 10051 27684
rect 12355 27429 12389 27605
rect 12473 27429 12507 27605
rect 12591 27429 12625 27605
rect 12709 27429 12743 27605
rect 12827 27429 12861 27605
rect 12945 27429 12979 27605
rect 13063 27429 13097 27605
rect 13181 27429 13215 27605
rect 13299 27429 13333 27605
rect 13417 27429 13451 27605
rect 14680 27301 14714 27677
rect 14798 27301 14832 27677
rect 14916 27301 14950 27677
rect 15034 27301 15068 27677
rect 15152 27301 15186 27677
rect 15270 27301 15304 27677
rect 15388 27301 15422 27677
rect 15822 27305 15856 27681
rect 15940 27305 15974 27681
rect 16058 27305 16092 27681
rect 16176 27305 16210 27681
rect 16294 27305 16328 27681
rect 16412 27305 16446 27681
rect 16530 27305 16564 27681
rect 18889 27424 18923 27600
rect 19007 27424 19041 27600
rect 19125 27424 19159 27600
rect 19243 27424 19277 27600
rect 19361 27424 19395 27600
rect 19479 27424 19513 27600
rect 19597 27424 19631 27600
rect 19715 27424 19749 27600
rect 19833 27424 19867 27600
rect 19951 27424 19985 27600
rect 8596 26721 8630 26897
rect 8714 26721 8748 26897
rect 8832 26721 8866 26897
rect 8950 26721 8984 26897
rect 9738 26725 9772 26901
rect 9856 26725 9890 26901
rect 9974 26725 10008 26901
rect 10092 26725 10126 26901
rect 21214 27296 21248 27672
rect 21332 27296 21366 27672
rect 21450 27296 21484 27672
rect 21568 27296 21602 27672
rect 21686 27296 21720 27672
rect 21804 27296 21838 27672
rect 21922 27296 21956 27672
rect 22356 27300 22390 27676
rect 22474 27300 22508 27676
rect 22592 27300 22626 27676
rect 22710 27300 22744 27676
rect 22828 27300 22862 27676
rect 22946 27300 22980 27676
rect 23064 27300 23098 27676
rect 25447 27428 25481 27604
rect 25565 27428 25599 27604
rect 25683 27428 25717 27604
rect 25801 27428 25835 27604
rect 25919 27428 25953 27604
rect 26037 27428 26071 27604
rect 26155 27428 26189 27604
rect 26273 27428 26307 27604
rect 26391 27428 26425 27604
rect 26509 27428 26543 27604
rect 15109 26718 15143 26894
rect 15227 26718 15261 26894
rect 15345 26718 15379 26894
rect 15463 26718 15497 26894
rect 16251 26722 16285 26898
rect 16369 26722 16403 26898
rect 16487 26722 16521 26898
rect 16605 26722 16639 26898
rect 27772 27300 27806 27676
rect 27890 27300 27924 27676
rect 28008 27300 28042 27676
rect 28126 27300 28160 27676
rect 28244 27300 28278 27676
rect 28362 27300 28396 27676
rect 28480 27300 28514 27676
rect 28914 27304 28948 27680
rect 29032 27304 29066 27680
rect 29150 27304 29184 27680
rect 29268 27304 29302 27680
rect 29386 27304 29420 27680
rect 29504 27304 29538 27680
rect 29622 27304 29656 27680
rect 21643 26713 21677 26889
rect 21761 26713 21795 26889
rect 21879 26713 21913 26889
rect 21997 26713 22031 26889
rect 22785 26717 22819 26893
rect 22903 26717 22937 26893
rect 23021 26717 23055 26893
rect 23139 26717 23173 26893
rect 28201 26717 28235 26893
rect 28319 26717 28353 26893
rect 28437 26717 28471 26893
rect 28555 26717 28589 26893
rect 29343 26721 29377 26897
rect 29461 26721 29495 26897
rect 29579 26721 29613 26897
rect 29697 26721 29731 26897
rect 5856 25782 5890 25958
rect 5974 25782 6008 25958
rect 6092 25782 6126 25958
rect 6210 25782 6244 25958
rect 6328 25782 6362 25958
rect 6446 25782 6480 25958
rect 6564 25782 6598 25958
rect 6682 25782 6716 25958
rect 6800 25782 6834 25958
rect 6918 25782 6952 25958
rect 12369 25779 12403 25955
rect 12487 25779 12521 25955
rect 12605 25779 12639 25955
rect 12723 25779 12757 25955
rect 12841 25779 12875 25955
rect 12959 25779 12993 25955
rect 13077 25779 13111 25955
rect 13195 25779 13229 25955
rect 13313 25779 13347 25955
rect 13431 25779 13465 25955
rect 18903 25774 18937 25950
rect 7320 25165 7354 25341
rect 7438 25165 7472 25341
rect 7556 25165 7590 25341
rect 7674 25165 7708 25341
rect 7804 25165 7838 25541
rect 7922 25165 7956 25541
rect 8040 25165 8074 25541
rect 8158 25165 8192 25541
rect 8276 25165 8310 25541
rect 8394 25165 8428 25541
rect 8512 25165 8546 25541
rect 8641 25165 8675 25341
rect 8759 25165 8793 25341
rect 8877 25165 8911 25341
rect 8995 25165 9029 25341
rect 9218 25165 9252 25341
rect 9336 25165 9370 25341
rect 9454 25165 9488 25341
rect 9572 25165 9606 25341
rect 9702 25165 9736 25541
rect 9820 25165 9854 25541
rect 9938 25165 9972 25541
rect 10056 25165 10090 25541
rect 10174 25165 10208 25541
rect 10292 25165 10326 25541
rect 10410 25165 10444 25541
rect 19021 25774 19055 25950
rect 19139 25774 19173 25950
rect 19257 25774 19291 25950
rect 19375 25774 19409 25950
rect 19493 25774 19527 25950
rect 19611 25774 19645 25950
rect 19729 25774 19763 25950
rect 19847 25774 19881 25950
rect 19965 25774 19999 25950
rect 25461 25778 25495 25954
rect 25579 25778 25613 25954
rect 25697 25778 25731 25954
rect 25815 25778 25849 25954
rect 25933 25778 25967 25954
rect 26051 25778 26085 25954
rect 26169 25778 26203 25954
rect 26287 25778 26321 25954
rect 26405 25778 26439 25954
rect 26523 25778 26557 25954
rect 10539 25165 10573 25341
rect 10657 25165 10691 25341
rect 10775 25165 10809 25341
rect 10893 25165 10927 25341
rect 5851 24178 5885 24354
rect 5969 24178 6003 24354
rect 6087 24178 6121 24354
rect 6205 24178 6239 24354
rect 6323 24178 6357 24354
rect 6441 24178 6475 24354
rect 6559 24178 6593 24354
rect 6677 24178 6711 24354
rect 6795 24178 6829 24354
rect 6913 24178 6947 24354
rect 7747 24472 7781 24848
rect 7865 24472 7899 24848
rect 7983 24472 8017 24848
rect 8101 24472 8135 24848
rect 8219 24472 8253 24848
rect 8337 24472 8371 24848
rect 8455 24472 8489 24848
rect 13833 25162 13867 25338
rect 13951 25162 13985 25338
rect 14069 25162 14103 25338
rect 14187 25162 14221 25338
rect 14317 25162 14351 25538
rect 14435 25162 14469 25538
rect 14553 25162 14587 25538
rect 14671 25162 14705 25538
rect 14789 25162 14823 25538
rect 14907 25162 14941 25538
rect 15025 25162 15059 25538
rect 15154 25162 15188 25338
rect 15272 25162 15306 25338
rect 15390 25162 15424 25338
rect 15508 25162 15542 25338
rect 15731 25162 15765 25338
rect 15849 25162 15883 25338
rect 15967 25162 16001 25338
rect 16085 25162 16119 25338
rect 16215 25162 16249 25538
rect 16333 25162 16367 25538
rect 16451 25162 16485 25538
rect 16569 25162 16603 25538
rect 16687 25162 16721 25538
rect 16805 25162 16839 25538
rect 16923 25162 16957 25538
rect 17052 25162 17086 25338
rect 17170 25162 17204 25338
rect 17288 25162 17322 25338
rect 17406 25162 17440 25338
rect 9645 24472 9679 24848
rect 9763 24472 9797 24848
rect 9881 24472 9915 24848
rect 9999 24472 10033 24848
rect 10117 24472 10151 24848
rect 10235 24472 10269 24848
rect 10353 24472 10387 24848
rect 12364 24175 12398 24351
rect 12482 24175 12516 24351
rect 12600 24175 12634 24351
rect 12718 24175 12752 24351
rect 12836 24175 12870 24351
rect 12954 24175 12988 24351
rect 13072 24175 13106 24351
rect 13190 24175 13224 24351
rect 13308 24175 13342 24351
rect 13426 24175 13460 24351
rect 14260 24469 14294 24845
rect 14378 24469 14412 24845
rect 14496 24469 14530 24845
rect 14614 24469 14648 24845
rect 14732 24469 14766 24845
rect 14850 24469 14884 24845
rect 14968 24469 15002 24845
rect 20367 25157 20401 25333
rect 20485 25157 20519 25333
rect 20603 25157 20637 25333
rect 20721 25157 20755 25333
rect 20851 25157 20885 25533
rect 20969 25157 21003 25533
rect 21087 25157 21121 25533
rect 21205 25157 21239 25533
rect 21323 25157 21357 25533
rect 21441 25157 21475 25533
rect 21559 25157 21593 25533
rect 21688 25157 21722 25333
rect 21806 25157 21840 25333
rect 21924 25157 21958 25333
rect 22042 25157 22076 25333
rect 22265 25157 22299 25333
rect 22383 25157 22417 25333
rect 22501 25157 22535 25333
rect 22619 25157 22653 25333
rect 22749 25157 22783 25533
rect 22867 25157 22901 25533
rect 22985 25157 23019 25533
rect 23103 25157 23137 25533
rect 23221 25157 23255 25533
rect 23339 25157 23373 25533
rect 23457 25157 23491 25533
rect 23586 25157 23620 25333
rect 23704 25157 23738 25333
rect 23822 25157 23856 25333
rect 23940 25157 23974 25333
rect 16158 24469 16192 24845
rect 16276 24469 16310 24845
rect 16394 24469 16428 24845
rect 16512 24469 16546 24845
rect 16630 24469 16664 24845
rect 16748 24469 16782 24845
rect 16866 24469 16900 24845
rect 18898 24170 18932 24346
rect 19016 24170 19050 24346
rect 19134 24170 19168 24346
rect 19252 24170 19286 24346
rect 19370 24170 19404 24346
rect 19488 24170 19522 24346
rect 19606 24170 19640 24346
rect 19724 24170 19758 24346
rect 19842 24170 19876 24346
rect 19960 24170 19994 24346
rect 20794 24464 20828 24840
rect 20912 24464 20946 24840
rect 21030 24464 21064 24840
rect 21148 24464 21182 24840
rect 21266 24464 21300 24840
rect 21384 24464 21418 24840
rect 21502 24464 21536 24840
rect 26925 25161 26959 25337
rect 27043 25161 27077 25337
rect 27161 25161 27195 25337
rect 27279 25161 27313 25337
rect 27409 25161 27443 25537
rect 27527 25161 27561 25537
rect 27645 25161 27679 25537
rect 27763 25161 27797 25537
rect 27881 25161 27915 25537
rect 27999 25161 28033 25537
rect 28117 25161 28151 25537
rect 28246 25161 28280 25337
rect 28364 25161 28398 25337
rect 28482 25161 28516 25337
rect 28600 25161 28634 25337
rect 28823 25161 28857 25337
rect 28941 25161 28975 25337
rect 29059 25161 29093 25337
rect 29177 25161 29211 25337
rect 29307 25161 29341 25537
rect 29425 25161 29459 25537
rect 29543 25161 29577 25537
rect 29661 25161 29695 25537
rect 29779 25161 29813 25537
rect 29897 25161 29931 25537
rect 30015 25161 30049 25537
rect 30144 25161 30178 25337
rect 30262 25161 30296 25337
rect 30380 25161 30414 25337
rect 30498 25161 30532 25337
rect 22692 24464 22726 24840
rect 22810 24464 22844 24840
rect 22928 24464 22962 24840
rect 23046 24464 23080 24840
rect 23164 24464 23198 24840
rect 23282 24464 23316 24840
rect 23400 24464 23434 24840
rect 25456 24174 25490 24350
rect 25574 24174 25608 24350
rect 25692 24174 25726 24350
rect 25810 24174 25844 24350
rect 25928 24174 25962 24350
rect 26046 24174 26080 24350
rect 26164 24174 26198 24350
rect 26282 24174 26316 24350
rect 26400 24174 26434 24350
rect 26518 24174 26552 24350
rect 27352 24468 27386 24844
rect 27470 24468 27504 24844
rect 27588 24468 27622 24844
rect 27706 24468 27740 24844
rect 27824 24468 27858 24844
rect 27942 24468 27976 24844
rect 28060 24468 28094 24844
rect 36967 25114 37143 25148
rect 36967 24996 37143 25030
rect 29250 24468 29284 24844
rect 29368 24468 29402 24844
rect 29486 24468 29520 24844
rect 29604 24468 29638 24844
rect 29722 24468 29756 24844
rect 29840 24468 29874 24844
rect 29958 24468 29992 24844
rect 36967 24878 37143 24912
rect 36967 24760 37143 24794
rect 36767 24673 37143 24707
rect 36767 24555 37143 24589
rect 36767 24437 37143 24471
rect 36767 24319 37143 24353
rect 36767 24206 37143 24240
rect 36767 24088 37143 24122
rect 36767 23970 37143 24004
rect 36767 23852 37143 23886
rect 36767 23734 37143 23768
rect 36767 23616 37143 23650
rect 36767 23498 37143 23532
rect 36767 23379 37143 23413
rect 36767 23261 37143 23295
rect 36767 23143 37143 23177
rect 36767 23025 37143 23059
rect 36967 22906 37143 22940
rect 36967 22788 37143 22822
rect 36967 22670 37143 22704
rect 36967 22552 37143 22586
rect 5853 21700 5887 22076
rect 5971 21700 6005 22076
rect 6089 21700 6123 22076
rect 6207 21700 6241 22076
rect 6325 21700 6359 22076
rect 6443 21700 6477 22076
rect 6561 21700 6595 22076
rect 6995 21696 7029 22072
rect 7113 21696 7147 22072
rect 7231 21696 7265 22072
rect 7349 21696 7383 22072
rect 7467 21696 7501 22072
rect 7585 21696 7619 22072
rect 7703 21696 7737 22072
rect 8966 21824 9000 22000
rect 9084 21824 9118 22000
rect 9202 21824 9236 22000
rect 9320 21824 9354 22000
rect 9438 21824 9472 22000
rect 9556 21824 9590 22000
rect 9674 21824 9708 22000
rect 9792 21824 9826 22000
rect 9910 21824 9944 22000
rect 10028 21824 10062 22000
rect 12411 21696 12445 22072
rect 12529 21696 12563 22072
rect 12647 21696 12681 22072
rect 12765 21696 12799 22072
rect 12883 21696 12917 22072
rect 13001 21696 13035 22072
rect 13119 21696 13153 22072
rect 13553 21692 13587 22068
rect 5778 21117 5812 21293
rect 5896 21117 5930 21293
rect 6014 21117 6048 21293
rect 6132 21117 6166 21293
rect 6920 21113 6954 21289
rect 7038 21113 7072 21289
rect 7156 21113 7190 21289
rect 7274 21113 7308 21289
rect 13671 21692 13705 22068
rect 13789 21692 13823 22068
rect 13907 21692 13941 22068
rect 14025 21692 14059 22068
rect 14143 21692 14177 22068
rect 14261 21692 14295 22068
rect 15524 21820 15558 21996
rect 15642 21820 15676 21996
rect 15760 21820 15794 21996
rect 15878 21820 15912 21996
rect 15996 21820 16030 21996
rect 16114 21820 16148 21996
rect 16232 21820 16266 21996
rect 16350 21820 16384 21996
rect 16468 21820 16502 21996
rect 16586 21820 16620 21996
rect 18945 21701 18979 22077
rect 19063 21701 19097 22077
rect 19181 21701 19215 22077
rect 19299 21701 19333 22077
rect 19417 21701 19451 22077
rect 19535 21701 19569 22077
rect 19653 21701 19687 22077
rect 20087 21697 20121 22073
rect 12336 21113 12370 21289
rect 12454 21113 12488 21289
rect 12572 21113 12606 21289
rect 12690 21113 12724 21289
rect 13478 21109 13512 21285
rect 13596 21109 13630 21285
rect 13714 21109 13748 21285
rect 13832 21109 13866 21285
rect 20205 21697 20239 22073
rect 20323 21697 20357 22073
rect 20441 21697 20475 22073
rect 20559 21697 20593 22073
rect 20677 21697 20711 22073
rect 20795 21697 20829 22073
rect 22058 21825 22092 22001
rect 22176 21825 22210 22001
rect 22294 21825 22328 22001
rect 22412 21825 22446 22001
rect 22530 21825 22564 22001
rect 22648 21825 22682 22001
rect 22766 21825 22800 22001
rect 22884 21825 22918 22001
rect 23002 21825 23036 22001
rect 23120 21825 23154 22001
rect 25458 21704 25492 22080
rect 25576 21704 25610 22080
rect 25694 21704 25728 22080
rect 25812 21704 25846 22080
rect 25930 21704 25964 22080
rect 26048 21704 26082 22080
rect 26166 21704 26200 22080
rect 26600 21700 26634 22076
rect 18870 21118 18904 21294
rect 18988 21118 19022 21294
rect 19106 21118 19140 21294
rect 19224 21118 19258 21294
rect 20012 21114 20046 21290
rect 20130 21114 20164 21290
rect 20248 21114 20282 21290
rect 20366 21114 20400 21290
rect 26718 21700 26752 22076
rect 26836 21700 26870 22076
rect 26954 21700 26988 22076
rect 27072 21700 27106 22076
rect 27190 21700 27224 22076
rect 27308 21700 27342 22076
rect 28571 21828 28605 22004
rect 28689 21828 28723 22004
rect 28807 21828 28841 22004
rect 28925 21828 28959 22004
rect 29043 21828 29077 22004
rect 29161 21828 29195 22004
rect 29279 21828 29313 22004
rect 29397 21828 29431 22004
rect 29515 21828 29549 22004
rect 29633 21828 29667 22004
rect 36967 21970 37143 22004
rect 36967 21852 37143 21886
rect 36967 21734 37143 21768
rect 36967 21616 37143 21650
rect 25383 21121 25417 21297
rect 25501 21121 25535 21297
rect 25619 21121 25653 21297
rect 25737 21121 25771 21297
rect 26525 21117 26559 21293
rect 26643 21117 26677 21293
rect 26761 21117 26795 21293
rect 26879 21117 26913 21293
rect 36767 21529 37143 21563
rect 36767 21411 37143 21445
rect 36767 21293 37143 21327
rect 36767 21175 37143 21209
rect 36767 21062 37143 21096
rect 36767 20944 37143 20978
rect 36767 20826 37143 20860
rect 36767 20708 37143 20742
rect 36767 20590 37143 20624
rect 8952 20174 8986 20350
rect 9070 20174 9104 20350
rect 9188 20174 9222 20350
rect 9306 20174 9340 20350
rect 9424 20174 9458 20350
rect 9542 20174 9576 20350
rect 9660 20174 9694 20350
rect 9778 20174 9812 20350
rect 9896 20174 9930 20350
rect 10014 20174 10048 20350
rect 15510 20170 15544 20346
rect 15628 20170 15662 20346
rect 15746 20170 15780 20346
rect 15864 20170 15898 20346
rect 15982 20170 16016 20346
rect 16100 20170 16134 20346
rect 16218 20170 16252 20346
rect 16336 20170 16370 20346
rect 16454 20170 16488 20346
rect 16572 20170 16606 20346
rect 22044 20175 22078 20351
rect 22162 20175 22196 20351
rect 22280 20175 22314 20351
rect 22398 20175 22432 20351
rect 22516 20175 22550 20351
rect 22634 20175 22668 20351
rect 22752 20175 22786 20351
rect 22870 20175 22904 20351
rect 22988 20175 23022 20351
rect 23106 20175 23140 20351
rect 36767 20472 37143 20506
rect 28557 20178 28591 20354
rect 28675 20178 28709 20354
rect 28793 20178 28827 20354
rect 28911 20178 28945 20354
rect 29029 20178 29063 20354
rect 29147 20178 29181 20354
rect 29265 20178 29299 20354
rect 29383 20178 29417 20354
rect 29501 20178 29535 20354
rect 29619 20178 29653 20354
rect 36767 20354 37143 20388
rect 36767 20235 37143 20269
rect 4977 19557 5011 19733
rect 5095 19557 5129 19733
rect 5213 19557 5247 19733
rect 5331 19557 5365 19733
rect 5460 19557 5494 19933
rect 5578 19557 5612 19933
rect 5696 19557 5730 19933
rect 5814 19557 5848 19933
rect 5932 19557 5966 19933
rect 6050 19557 6084 19933
rect 6168 19557 6202 19933
rect 6298 19557 6332 19733
rect 6416 19557 6450 19733
rect 6534 19557 6568 19733
rect 6652 19557 6686 19733
rect 6875 19557 6909 19733
rect 6993 19557 7027 19733
rect 7111 19557 7145 19733
rect 7229 19557 7263 19733
rect 7358 19557 7392 19933
rect 7476 19557 7510 19933
rect 7594 19557 7628 19933
rect 7712 19557 7746 19933
rect 7830 19557 7864 19933
rect 7948 19557 7982 19933
rect 8066 19557 8100 19933
rect 8196 19557 8230 19733
rect 8314 19557 8348 19733
rect 8432 19557 8466 19733
rect 8550 19557 8584 19733
rect 5517 18864 5551 19240
rect 5635 18864 5669 19240
rect 5753 18864 5787 19240
rect 5871 18864 5905 19240
rect 5989 18864 6023 19240
rect 6107 18864 6141 19240
rect 6225 18864 6259 19240
rect 11535 19553 11569 19729
rect 11653 19553 11687 19729
rect 11771 19553 11805 19729
rect 11889 19553 11923 19729
rect 12018 19553 12052 19929
rect 12136 19553 12170 19929
rect 12254 19553 12288 19929
rect 12372 19553 12406 19929
rect 12490 19553 12524 19929
rect 12608 19553 12642 19929
rect 12726 19553 12760 19929
rect 12856 19553 12890 19729
rect 12974 19553 13008 19729
rect 13092 19553 13126 19729
rect 13210 19553 13244 19729
rect 13433 19553 13467 19729
rect 13551 19553 13585 19729
rect 13669 19553 13703 19729
rect 13787 19553 13821 19729
rect 13916 19553 13950 19929
rect 14034 19553 14068 19929
rect 14152 19553 14186 19929
rect 14270 19553 14304 19929
rect 14388 19553 14422 19929
rect 14506 19553 14540 19929
rect 14624 19553 14658 19929
rect 14754 19553 14788 19729
rect 14872 19553 14906 19729
rect 14990 19553 15024 19729
rect 15108 19553 15142 19729
rect 7415 18864 7449 19240
rect 7533 18864 7567 19240
rect 7651 18864 7685 19240
rect 7769 18864 7803 19240
rect 7887 18864 7921 19240
rect 8005 18864 8039 19240
rect 8123 18864 8157 19240
rect 8957 18570 8991 18746
rect 9075 18570 9109 18746
rect 9193 18570 9227 18746
rect 9311 18570 9345 18746
rect 9429 18570 9463 18746
rect 9547 18570 9581 18746
rect 9665 18570 9699 18746
rect 9783 18570 9817 18746
rect 9901 18570 9935 18746
rect 10019 18570 10053 18746
rect 12075 18860 12109 19236
rect 12193 18860 12227 19236
rect 12311 18860 12345 19236
rect 12429 18860 12463 19236
rect 12547 18860 12581 19236
rect 12665 18860 12699 19236
rect 12783 18860 12817 19236
rect 18069 19558 18103 19734
rect 18187 19558 18221 19734
rect 18305 19558 18339 19734
rect 18423 19558 18457 19734
rect 18552 19558 18586 19934
rect 18670 19558 18704 19934
rect 18788 19558 18822 19934
rect 18906 19558 18940 19934
rect 19024 19558 19058 19934
rect 19142 19558 19176 19934
rect 19260 19558 19294 19934
rect 19390 19558 19424 19734
rect 19508 19558 19542 19734
rect 19626 19558 19660 19734
rect 19744 19558 19778 19734
rect 19967 19558 20001 19734
rect 20085 19558 20119 19734
rect 20203 19558 20237 19734
rect 20321 19558 20355 19734
rect 20450 19558 20484 19934
rect 20568 19558 20602 19934
rect 20686 19558 20720 19934
rect 20804 19558 20838 19934
rect 20922 19558 20956 19934
rect 21040 19558 21074 19934
rect 21158 19558 21192 19934
rect 21288 19558 21322 19734
rect 21406 19558 21440 19734
rect 21524 19558 21558 19734
rect 21642 19558 21676 19734
rect 13973 18860 14007 19236
rect 14091 18860 14125 19236
rect 14209 18860 14243 19236
rect 14327 18860 14361 19236
rect 14445 18860 14479 19236
rect 14563 18860 14597 19236
rect 14681 18860 14715 19236
rect 15515 18566 15549 18742
rect 15633 18566 15667 18742
rect 15751 18566 15785 18742
rect 15869 18566 15903 18742
rect 15987 18566 16021 18742
rect 16105 18566 16139 18742
rect 16223 18566 16257 18742
rect 16341 18566 16375 18742
rect 16459 18566 16493 18742
rect 16577 18566 16611 18742
rect 18609 18865 18643 19241
rect 18727 18865 18761 19241
rect 18845 18865 18879 19241
rect 18963 18865 18997 19241
rect 19081 18865 19115 19241
rect 19199 18865 19233 19241
rect 19317 18865 19351 19241
rect 24582 19561 24616 19737
rect 24700 19561 24734 19737
rect 24818 19561 24852 19737
rect 24936 19561 24970 19737
rect 25065 19561 25099 19937
rect 25183 19561 25217 19937
rect 25301 19561 25335 19937
rect 25419 19561 25453 19937
rect 25537 19561 25571 19937
rect 25655 19561 25689 19937
rect 25773 19561 25807 19937
rect 25903 19561 25937 19737
rect 26021 19561 26055 19737
rect 26139 19561 26173 19737
rect 26257 19561 26291 19737
rect 26480 19561 26514 19737
rect 26598 19561 26632 19737
rect 26716 19561 26750 19737
rect 26834 19561 26868 19737
rect 26963 19561 26997 19937
rect 27081 19561 27115 19937
rect 27199 19561 27233 19937
rect 27317 19561 27351 19937
rect 27435 19561 27469 19937
rect 27553 19561 27587 19937
rect 27671 19561 27705 19937
rect 36767 20117 37143 20151
rect 36767 19999 37143 20033
rect 27801 19561 27835 19737
rect 27919 19561 27953 19737
rect 28037 19561 28071 19737
rect 28155 19561 28189 19737
rect 20507 18865 20541 19241
rect 20625 18865 20659 19241
rect 20743 18865 20777 19241
rect 20861 18865 20895 19241
rect 20979 18865 21013 19241
rect 21097 18865 21131 19241
rect 21215 18865 21249 19241
rect 22049 18571 22083 18747
rect 22167 18571 22201 18747
rect 22285 18571 22319 18747
rect 22403 18571 22437 18747
rect 22521 18571 22555 18747
rect 22639 18571 22673 18747
rect 22757 18571 22791 18747
rect 22875 18571 22909 18747
rect 22993 18571 23027 18747
rect 23111 18571 23145 18747
rect 25122 18868 25156 19244
rect 25240 18868 25274 19244
rect 25358 18868 25392 19244
rect 25476 18868 25510 19244
rect 25594 18868 25628 19244
rect 25712 18868 25746 19244
rect 25830 18868 25864 19244
rect 36767 19881 37143 19915
rect 36967 19762 37143 19796
rect 36967 19644 37143 19678
rect 36967 19526 37143 19560
rect 36967 19408 37143 19442
rect 27020 18868 27054 19244
rect 27138 18868 27172 19244
rect 27256 18868 27290 19244
rect 27374 18868 27408 19244
rect 27492 18868 27526 19244
rect 27610 18868 27644 19244
rect 27728 18868 27762 19244
rect 36963 18838 37139 18872
rect 28562 18574 28596 18750
rect 28680 18574 28714 18750
rect 28798 18574 28832 18750
rect 28916 18574 28950 18750
rect 29034 18574 29068 18750
rect 29152 18574 29186 18750
rect 29270 18574 29304 18750
rect 29388 18574 29422 18750
rect 29506 18574 29540 18750
rect 29624 18574 29658 18750
rect 36963 18720 37139 18754
rect 36963 18602 37139 18636
rect 36963 18484 37139 18518
rect 36763 18397 37139 18431
rect 36763 18279 37139 18313
rect 36763 18161 37139 18195
rect 36763 18043 37139 18077
rect 36763 17930 37139 17964
rect 36763 17812 37139 17846
rect 36763 17694 37139 17728
rect 36763 17576 37139 17610
rect 36763 17458 37139 17492
rect 36763 17340 37139 17374
rect 36763 17222 37139 17256
rect 36763 17103 37139 17137
rect 36763 16985 37139 17019
rect 36763 16867 37139 16901
rect 36763 16749 37139 16783
rect 36963 16630 37139 16664
rect 36963 16512 37139 16546
rect 36963 16394 37139 16428
rect 36963 16276 37139 16310
rect -3592 16221 -3416 16255
rect -3592 16103 -3416 16137
rect -3592 15985 -3416 16019
rect -3592 15867 -3416 15901
rect -3792 15737 -3416 15771
rect -3099 15794 -2723 15828
rect -3792 15619 -3416 15653
rect -3099 15676 -2723 15710
rect 36963 15694 37139 15728
rect -3792 15501 -3416 15535
rect -3099 15558 -2723 15592
rect 36963 15576 37139 15610
rect -3099 15440 -2723 15474
rect -3792 15383 -3416 15417
rect -3792 15265 -3416 15299
rect -3792 15147 -3416 15181
rect -3099 15322 -2723 15356
rect 36963 15458 37139 15492
rect -3099 15204 -2723 15238
rect -3792 15029 -3416 15063
rect -3592 14900 -3416 14934
rect -3099 15086 -2723 15120
rect 7812 15048 7846 15224
rect 7930 15048 7964 15224
rect 8048 15048 8082 15224
rect 8166 15048 8200 15224
rect 8284 15048 8318 15224
rect 8402 15048 8436 15224
rect 8520 15048 8554 15224
rect 8638 15048 8672 15224
rect 8756 15048 8790 15224
rect 8874 15048 8908 15224
rect 14361 15047 14395 15223
rect -3592 14782 -3416 14816
rect 14479 15047 14513 15223
rect 14597 15047 14631 15223
rect 14715 15047 14749 15223
rect 14833 15047 14867 15223
rect 14951 15047 14985 15223
rect 15069 15047 15103 15223
rect 15187 15047 15221 15223
rect 15305 15047 15339 15223
rect 15423 15047 15457 15223
rect 21015 15068 21049 15244
rect 21133 15068 21167 15244
rect 21251 15068 21285 15244
rect 21369 15068 21403 15244
rect 21487 15068 21521 15244
rect 21605 15068 21639 15244
rect 21723 15068 21757 15244
rect 21841 15068 21875 15244
rect 21959 15068 21993 15244
rect 22077 15068 22111 15244
rect 36963 15340 37139 15374
rect 36763 15253 37139 15287
rect 36763 15135 37139 15169
rect -3592 14664 -3416 14698
rect -3592 14546 -3416 14580
rect 29668 14901 29702 15077
rect 29786 14901 29820 15077
rect 29904 14901 29938 15077
rect 30022 14901 30056 15077
rect 30140 14901 30174 15077
rect 30258 14901 30292 15077
rect 30376 14901 30410 15077
rect 30494 14901 30528 15077
rect 30612 14901 30646 15077
rect 30730 14901 30764 15077
rect 36763 15017 37139 15051
rect -3594 14153 -3418 14187
rect 31476 14496 31510 14672
rect 31594 14496 31628 14672
rect 31712 14496 31746 14672
rect 31830 14496 31864 14672
rect 31960 14496 31994 14872
rect 32078 14496 32112 14872
rect 32196 14496 32230 14872
rect 32314 14496 32348 14872
rect 32432 14496 32466 14872
rect 32550 14496 32584 14872
rect 32668 14496 32702 14872
rect 36763 14899 37139 14933
rect 36763 14786 37139 14820
rect 32797 14496 32831 14672
rect 32915 14496 32949 14672
rect 33033 14496 33067 14672
rect 33151 14496 33185 14672
rect 33269 14493 33303 14669
rect 33387 14493 33421 14669
rect 33505 14493 33539 14669
rect 33623 14493 33657 14669
rect 33741 14493 33775 14669
rect 33859 14493 33893 14669
rect 33977 14493 34011 14669
rect 34095 14493 34129 14669
rect 34213 14493 34247 14669
rect 34331 14493 34365 14669
rect 36763 14668 37139 14702
rect -3594 14035 -3418 14069
rect -3594 13917 -3418 13951
rect -3594 13799 -3418 13833
rect -3794 13669 -3418 13703
rect -3101 13726 -2725 13760
rect -3794 13551 -3418 13585
rect -3101 13608 -2725 13642
rect -3794 13433 -3418 13467
rect -3101 13490 -2725 13524
rect -3101 13372 -2725 13406
rect -3794 13315 -3418 13349
rect -3794 13197 -3418 13231
rect -3794 13079 -3418 13113
rect -3101 13254 -2725 13288
rect -3101 13136 -2725 13170
rect 1148 13148 1182 13324
rect 1266 13148 1300 13324
rect 1384 13148 1418 13324
rect 1502 13148 1536 13324
rect 1620 13148 1654 13324
rect 1738 13148 1772 13324
rect 1856 13148 1890 13324
rect 1974 13148 2008 13324
rect 2092 13148 2126 13324
rect 2210 13148 2244 13324
rect 31903 13803 31937 14179
rect 32021 13803 32055 14179
rect 32139 13803 32173 14179
rect 32257 13803 32291 14179
rect 32375 13803 32409 14179
rect 32493 13803 32527 14179
rect 32611 13803 32645 14179
rect 36763 14550 37139 14584
rect 36763 14432 37139 14466
rect 36763 14314 37139 14348
rect 36763 14196 37139 14230
rect 36763 14078 37139 14112
rect 36763 13959 37139 13993
rect 36763 13841 37139 13875
rect 36763 13723 37139 13757
rect 36763 13605 37139 13639
rect 36963 13486 37139 13520
rect -3794 12961 -3418 12995
rect -3594 12832 -3418 12866
rect -3101 13018 -2725 13052
rect -3594 12714 -3418 12748
rect -3594 12596 -3418 12630
rect -3594 12478 -3418 12512
rect 4038 12881 4072 13057
rect 4156 12881 4190 13057
rect 4274 12881 4308 13057
rect 4392 12881 4426 13057
rect 4510 12881 4544 13057
rect 4628 12881 4662 13057
rect 4746 12881 4780 13057
rect 4864 12881 4898 13057
rect 4982 12881 5016 13057
rect 5100 12881 5134 13057
rect 6363 12753 6397 13129
rect 6481 12753 6515 13129
rect 6599 12753 6633 13129
rect 6717 12753 6751 13129
rect 6835 12753 6869 13129
rect 6953 12753 6987 13129
rect 7071 12753 7105 13129
rect 7505 12757 7539 13133
rect 7623 12757 7657 13133
rect 7741 12757 7775 13133
rect 7859 12757 7893 13133
rect 7977 12757 8011 13133
rect 8095 12757 8129 13133
rect 8213 12757 8247 13133
rect 10587 12969 10621 13145
rect 10705 12969 10739 13145
rect 10823 12969 10857 13145
rect 10941 12969 10975 13145
rect 11059 12969 11093 13145
rect 11177 12969 11211 13145
rect 11295 12969 11329 13145
rect 11413 12969 11447 13145
rect 11531 12969 11565 13145
rect 11649 12969 11683 13145
rect 12912 12841 12946 13217
rect 13030 12841 13064 13217
rect 13148 12841 13182 13217
rect 13266 12841 13300 13217
rect 13384 12841 13418 13217
rect 13502 12841 13536 13217
rect 13620 12841 13654 13217
rect 14054 12845 14088 13221
rect 14172 12845 14206 13221
rect 14290 12845 14324 13221
rect 14408 12845 14442 13221
rect 14526 12845 14560 13221
rect 14644 12845 14678 13221
rect 14762 12845 14796 13221
rect 17241 12901 17275 13077
rect 17359 12901 17393 13077
rect 17477 12901 17511 13077
rect 17595 12901 17629 13077
rect 17713 12901 17747 13077
rect 17831 12901 17865 13077
rect 17949 12901 17983 13077
rect 18067 12901 18101 13077
rect 18185 12901 18219 13077
rect 18303 12901 18337 13077
rect 6792 12170 6826 12346
rect 6910 12170 6944 12346
rect 7028 12170 7062 12346
rect 7146 12170 7180 12346
rect 7934 12174 7968 12350
rect 8052 12174 8086 12350
rect 8170 12174 8204 12350
rect 8288 12174 8322 12350
rect 19566 12773 19600 13149
rect 19684 12773 19718 13149
rect 19802 12773 19836 13149
rect 19920 12773 19954 13149
rect 20038 12773 20072 13149
rect 20156 12773 20190 13149
rect 20274 12773 20308 13149
rect 20708 12777 20742 13153
rect 20826 12777 20860 13153
rect 20944 12777 20978 13153
rect 21062 12777 21096 13153
rect 21180 12777 21214 13153
rect 21298 12777 21332 13153
rect 21416 12777 21450 13153
rect 23866 12969 23900 13145
rect 23984 12969 24018 13145
rect 24102 12969 24136 13145
rect 24220 12969 24254 13145
rect 24338 12969 24372 13145
rect 24456 12969 24490 13145
rect 24574 12969 24608 13145
rect 24692 12969 24726 13145
rect 24810 12969 24844 13145
rect 24928 12969 24962 13145
rect 13341 12258 13375 12434
rect 13459 12258 13493 12434
rect 13577 12258 13611 12434
rect 13695 12258 13729 12434
rect 14483 12262 14517 12438
rect 14601 12262 14635 12438
rect 14719 12262 14753 12438
rect 14837 12262 14871 12438
rect 26191 12841 26225 13217
rect 26309 12841 26343 13217
rect 26427 12841 26461 13217
rect 26545 12841 26579 13217
rect 26663 12841 26697 13217
rect 26781 12841 26815 13217
rect 26899 12841 26933 13217
rect 27333 12845 27367 13221
rect 27451 12845 27485 13221
rect 27569 12845 27603 13221
rect 27687 12845 27721 13221
rect 27805 12845 27839 13221
rect 27923 12845 27957 13221
rect 28041 12845 28075 13221
rect 36963 13368 37139 13402
rect 36963 13250 37139 13284
rect 36963 13132 37139 13166
rect 19995 12190 20029 12366
rect 20113 12190 20147 12366
rect 20231 12190 20265 12366
rect 20349 12190 20383 12366
rect 21137 12194 21171 12370
rect 21255 12194 21289 12370
rect 21373 12194 21407 12370
rect 21491 12194 21525 12370
rect 26620 12258 26654 12434
rect 26738 12258 26772 12434
rect 26856 12258 26890 12434
rect 26974 12258 27008 12434
rect 27762 12262 27796 12438
rect 27880 12262 27914 12438
rect 27998 12262 28032 12438
rect 28116 12262 28150 12438
rect 29663 12330 29697 12506
rect 29781 12330 29815 12506
rect 29899 12330 29933 12506
rect 30017 12330 30051 12506
rect 30135 12330 30169 12506
rect 30253 12330 30287 12506
rect 30371 12330 30405 12506
rect 30489 12330 30523 12506
rect 30607 12330 30641 12506
rect 30725 12330 30759 12506
rect 36967 12492 37143 12526
rect 36967 12374 37143 12408
rect -3592 12084 -3416 12118
rect -3592 11966 -3416 12000
rect 36967 12256 37143 12290
rect 36967 12138 37143 12172
rect -3592 11848 -3416 11882
rect -3592 11730 -3416 11764
rect -3792 11600 -3416 11634
rect -3099 11657 -2723 11691
rect -3792 11482 -3416 11516
rect -3099 11539 -2723 11573
rect 36767 12051 37143 12085
rect 36767 11933 37143 11967
rect 36767 11815 37143 11849
rect 36767 11697 37143 11731
rect -3792 11364 -3416 11398
rect -3099 11421 -2723 11455
rect -3099 11303 -2723 11337
rect -3792 11246 -3416 11280
rect -3792 11128 -3416 11162
rect -3792 11010 -3416 11044
rect -3099 11185 -2723 11219
rect 4052 11231 4086 11407
rect 4170 11231 4204 11407
rect 4288 11231 4322 11407
rect 4406 11231 4440 11407
rect 4524 11231 4558 11407
rect 4642 11231 4676 11407
rect 4760 11231 4794 11407
rect 4878 11231 4912 11407
rect 4996 11231 5030 11407
rect 5114 11231 5148 11407
rect 10601 11319 10635 11495
rect 10719 11319 10753 11495
rect 10837 11319 10871 11495
rect 10955 11319 10989 11495
rect 11073 11319 11107 11495
rect 11191 11319 11225 11495
rect 11309 11319 11343 11495
rect 11427 11319 11461 11495
rect 11545 11319 11579 11495
rect 11663 11319 11697 11495
rect 36767 11584 37143 11618
rect -3099 11067 -2723 11101
rect -3792 10892 -3416 10926
rect -3592 10763 -3416 10797
rect -3099 10949 -2723 10983
rect 17255 11251 17289 11427
rect 17373 11251 17407 11427
rect 17491 11251 17525 11427
rect 17609 11251 17643 11427
rect 17727 11251 17761 11427
rect 17845 11251 17879 11427
rect 17963 11251 17997 11427
rect 18081 11251 18115 11427
rect 18199 11251 18233 11427
rect 18317 11251 18351 11427
rect 23880 11319 23914 11495
rect 23998 11319 24032 11495
rect 24116 11319 24150 11495
rect 24234 11319 24268 11495
rect 24352 11319 24386 11495
rect 24470 11319 24504 11495
rect 24588 11319 24622 11495
rect 24706 11319 24740 11495
rect 24824 11319 24858 11495
rect 24942 11319 24976 11495
rect 36767 11466 37143 11500
rect -3592 10645 -3416 10679
rect -3592 10527 -3416 10561
rect 1140 10563 1174 10739
rect 1258 10563 1292 10739
rect 1376 10563 1410 10739
rect 1494 10563 1528 10739
rect 1612 10563 1646 10739
rect 1730 10563 1764 10739
rect 1848 10563 1882 10739
rect 1966 10563 2000 10739
rect 2084 10563 2118 10739
rect 2202 10563 2236 10739
rect -3592 10409 -3416 10443
rect 5516 10614 5550 10790
rect 5634 10614 5668 10790
rect 5752 10614 5786 10790
rect 5870 10614 5904 10790
rect 6000 10614 6034 10990
rect 6118 10614 6152 10990
rect 6236 10614 6270 10990
rect 6354 10614 6388 10990
rect 6472 10614 6506 10990
rect 6590 10614 6624 10990
rect 6708 10614 6742 10990
rect 6837 10614 6871 10790
rect 6955 10614 6989 10790
rect 7073 10614 7107 10790
rect 7191 10614 7225 10790
rect 7414 10614 7448 10790
rect 7532 10614 7566 10790
rect 7650 10614 7684 10790
rect 7768 10614 7802 10790
rect 7898 10614 7932 10990
rect 8016 10614 8050 10990
rect 8134 10614 8168 10990
rect 8252 10614 8286 10990
rect 8370 10614 8404 10990
rect 8488 10614 8522 10990
rect 8606 10614 8640 10990
rect 8735 10614 8769 10790
rect 8853 10614 8887 10790
rect 8971 10614 9005 10790
rect 9089 10614 9123 10790
rect -3594 10016 -3418 10050
rect -3594 9898 -3418 9932
rect -3594 9780 -3418 9814
rect -3594 9662 -3418 9696
rect -3794 9532 -3418 9566
rect -3101 9589 -2725 9623
rect 4047 9627 4081 9803
rect 4165 9627 4199 9803
rect 4283 9627 4317 9803
rect 4401 9627 4435 9803
rect 4519 9627 4553 9803
rect 4637 9627 4671 9803
rect 4755 9627 4789 9803
rect 4873 9627 4907 9803
rect 4991 9627 5025 9803
rect 5109 9627 5143 9803
rect 5943 9921 5977 10297
rect 6061 9921 6095 10297
rect 6179 9921 6213 10297
rect 6297 9921 6331 10297
rect 6415 9921 6449 10297
rect 6533 9921 6567 10297
rect 6651 9921 6685 10297
rect -3794 9414 -3418 9448
rect -3101 9471 -2725 9505
rect -3794 9296 -3418 9330
rect -3101 9353 -2725 9387
rect 12065 10702 12099 10878
rect 12183 10702 12217 10878
rect 12301 10702 12335 10878
rect 12419 10702 12453 10878
rect 12549 10702 12583 11078
rect 12667 10702 12701 11078
rect 12785 10702 12819 11078
rect 12903 10702 12937 11078
rect 13021 10702 13055 11078
rect 13139 10702 13173 11078
rect 13257 10702 13291 11078
rect 13386 10702 13420 10878
rect 13504 10702 13538 10878
rect 13622 10702 13656 10878
rect 13740 10702 13774 10878
rect 13963 10702 13997 10878
rect 14081 10702 14115 10878
rect 14199 10702 14233 10878
rect 14317 10702 14351 10878
rect 14447 10702 14481 11078
rect 14565 10702 14599 11078
rect 14683 10702 14717 11078
rect 14801 10702 14835 11078
rect 14919 10702 14953 11078
rect 15037 10702 15071 11078
rect 15155 10702 15189 11078
rect 36767 11348 37143 11382
rect 36767 11230 37143 11264
rect 36767 11112 37143 11146
rect 15284 10702 15318 10878
rect 15402 10702 15436 10878
rect 15520 10702 15554 10878
rect 15638 10702 15672 10878
rect 7841 9921 7875 10297
rect 7959 9921 7993 10297
rect 8077 9921 8111 10297
rect 8195 9921 8229 10297
rect 8313 9921 8347 10297
rect 8431 9921 8465 10297
rect 8549 9921 8583 10297
rect 10596 9715 10630 9891
rect 10714 9715 10748 9891
rect 10832 9715 10866 9891
rect 10950 9715 10984 9891
rect 11068 9715 11102 9891
rect 11186 9715 11220 9891
rect 11304 9715 11338 9891
rect 11422 9715 11456 9891
rect 11540 9715 11574 9891
rect 11658 9715 11692 9891
rect 12492 10009 12526 10385
rect 12610 10009 12644 10385
rect 12728 10009 12762 10385
rect 12846 10009 12880 10385
rect 12964 10009 12998 10385
rect 13082 10009 13116 10385
rect 13200 10009 13234 10385
rect -3101 9235 -2725 9269
rect -3794 9178 -3418 9212
rect -3794 9060 -3418 9094
rect -3794 8942 -3418 8976
rect -3101 9117 -2725 9151
rect -3101 8999 -2725 9033
rect 18719 10634 18753 10810
rect 18837 10634 18871 10810
rect 18955 10634 18989 10810
rect 19073 10634 19107 10810
rect 19203 10634 19237 11010
rect 19321 10634 19355 11010
rect 19439 10634 19473 11010
rect 19557 10634 19591 11010
rect 19675 10634 19709 11010
rect 19793 10634 19827 11010
rect 19911 10634 19945 11010
rect 20040 10634 20074 10810
rect 20158 10634 20192 10810
rect 20276 10634 20310 10810
rect 20394 10634 20428 10810
rect 20617 10634 20651 10810
rect 20735 10634 20769 10810
rect 20853 10634 20887 10810
rect 20971 10634 21005 10810
rect 21101 10634 21135 11010
rect 21219 10634 21253 11010
rect 21337 10634 21371 11010
rect 21455 10634 21489 11010
rect 21573 10634 21607 11010
rect 21691 10634 21725 11010
rect 21809 10634 21843 11010
rect 21938 10634 21972 10810
rect 22056 10634 22090 10810
rect 22174 10634 22208 10810
rect 22292 10634 22326 10810
rect 14390 10009 14424 10385
rect 14508 10009 14542 10385
rect 14626 10009 14660 10385
rect 14744 10009 14778 10385
rect 14862 10009 14896 10385
rect 14980 10009 15014 10385
rect 15098 10009 15132 10385
rect 17250 9647 17284 9823
rect 17368 9647 17402 9823
rect 17486 9647 17520 9823
rect 17604 9647 17638 9823
rect 17722 9647 17756 9823
rect 17840 9647 17874 9823
rect 17958 9647 17992 9823
rect 18076 9647 18110 9823
rect 18194 9647 18228 9823
rect 18312 9647 18346 9823
rect 19146 9941 19180 10317
rect 19264 9941 19298 10317
rect 19382 9941 19416 10317
rect 19500 9941 19534 10317
rect 19618 9941 19652 10317
rect 19736 9941 19770 10317
rect 19854 9941 19888 10317
rect 25344 10702 25378 10878
rect 25462 10702 25496 10878
rect 25580 10702 25614 10878
rect 25698 10702 25732 10878
rect 25828 10702 25862 11078
rect 25946 10702 25980 11078
rect 26064 10702 26098 11078
rect 26182 10702 26216 11078
rect 26300 10702 26334 11078
rect 26418 10702 26452 11078
rect 26536 10702 26570 11078
rect 26665 10702 26699 10878
rect 26783 10702 26817 10878
rect 26901 10702 26935 10878
rect 27019 10702 27053 10878
rect 27242 10702 27276 10878
rect 27360 10702 27394 10878
rect 27478 10702 27512 10878
rect 27596 10702 27630 10878
rect 27726 10702 27760 11078
rect 27844 10702 27878 11078
rect 27962 10702 27996 11078
rect 28080 10702 28114 11078
rect 28198 10702 28232 11078
rect 28316 10702 28350 11078
rect 28434 10702 28468 11078
rect 36767 10994 37143 11028
rect 28563 10702 28597 10878
rect 28681 10702 28715 10878
rect 28799 10702 28833 10878
rect 28917 10702 28951 10878
rect 36767 10876 37143 10910
rect 21044 9941 21078 10317
rect 21162 9941 21196 10317
rect 21280 9941 21314 10317
rect 21398 9941 21432 10317
rect 21516 9941 21550 10317
rect 21634 9941 21668 10317
rect 21752 9941 21786 10317
rect 23875 9715 23909 9891
rect 23993 9715 24027 9891
rect 24111 9715 24145 9891
rect 24229 9715 24263 9891
rect 24347 9715 24381 9891
rect 24465 9715 24499 9891
rect 24583 9715 24617 9891
rect 24701 9715 24735 9891
rect 24819 9715 24853 9891
rect 24937 9715 24971 9891
rect 25771 10009 25805 10385
rect 25889 10009 25923 10385
rect 26007 10009 26041 10385
rect 26125 10009 26159 10385
rect 26243 10009 26277 10385
rect 26361 10009 26395 10385
rect 26479 10009 26513 10385
rect -3794 8824 -3418 8858
rect -3594 8695 -3418 8729
rect -3101 8881 -2725 8915
rect 27669 10009 27703 10385
rect 27787 10009 27821 10385
rect 27905 10009 27939 10385
rect 28023 10009 28057 10385
rect 28141 10009 28175 10385
rect 28259 10009 28293 10385
rect 28377 10009 28411 10385
rect 31478 10405 31512 10581
rect 31596 10405 31630 10581
rect 31714 10405 31748 10581
rect 31832 10405 31866 10581
rect 31962 10405 31996 10781
rect 32080 10405 32114 10781
rect 32198 10405 32232 10781
rect 32316 10405 32350 10781
rect 32434 10405 32468 10781
rect 32552 10405 32586 10781
rect 32670 10405 32704 10781
rect 36767 10757 37143 10791
rect 32799 10405 32833 10581
rect 32917 10405 32951 10581
rect 33035 10405 33069 10581
rect 36767 10639 37143 10673
rect 33153 10405 33187 10581
rect 33271 10402 33305 10578
rect 33389 10402 33423 10578
rect 33507 10402 33541 10578
rect 33625 10402 33659 10578
rect 33743 10402 33777 10578
rect 33861 10402 33895 10578
rect 33979 10402 34013 10578
rect 34097 10402 34131 10578
rect 34215 10402 34249 10578
rect 34333 10402 34367 10578
rect 36767 10521 37143 10555
rect 36767 10403 37143 10437
rect 29663 9297 29697 9473
rect 29781 9297 29815 9473
rect 29899 9297 29933 9473
rect 30017 9297 30051 9473
rect 30135 9297 30169 9473
rect 30253 9297 30287 9473
rect 30371 9297 30405 9473
rect 30489 9297 30523 9473
rect 30607 9297 30641 9473
rect 30725 9297 30759 9473
rect 31905 9712 31939 10088
rect 32023 9712 32057 10088
rect 32141 9712 32175 10088
rect 32259 9712 32293 10088
rect 32377 9712 32411 10088
rect 32495 9712 32529 10088
rect 32613 9712 32647 10088
rect 36967 10284 37143 10318
rect 36967 10166 37143 10200
rect 36967 10048 37143 10082
rect 36967 9930 37143 9964
rect -3594 8577 -3418 8611
rect 36967 9348 37143 9382
rect 36967 9230 37143 9264
rect 36967 9112 37143 9146
rect 36967 8994 37143 9028
rect 36767 8907 37143 8941
rect 36767 8789 37143 8823
rect 36767 8671 37143 8705
rect 36767 8553 37143 8587
rect -3594 8459 -3418 8493
rect 36767 8440 37143 8474
rect -3594 8341 -3418 8375
rect 36767 8322 37143 8356
rect 36767 8204 37143 8238
rect 36767 8086 37143 8120
rect -3594 7947 -3418 7981
rect -3594 7829 -3418 7863
rect 36767 7968 37143 8002
rect 36767 7850 37143 7884
rect -3594 7711 -3418 7745
rect -3594 7593 -3418 7627
rect -3794 7463 -3418 7497
rect -3101 7520 -2725 7554
rect -3794 7345 -3418 7379
rect -3101 7402 -2725 7436
rect -3794 7227 -3418 7261
rect -3101 7284 -2725 7318
rect 1121 7285 1155 7461
rect 1239 7285 1273 7461
rect 1357 7285 1391 7461
rect 1475 7285 1509 7461
rect 1593 7285 1627 7461
rect 1711 7285 1745 7461
rect 1829 7285 1863 7461
rect 1947 7285 1981 7461
rect 2065 7285 2099 7461
rect 2183 7285 2217 7461
rect -3101 7166 -2725 7200
rect -3794 7109 -3418 7143
rect -3794 6991 -3418 7025
rect -3794 6873 -3418 6907
rect -3101 7048 -2725 7082
rect 4030 7101 4064 7277
rect 4148 7101 4182 7277
rect 4266 7101 4300 7277
rect 4384 7101 4418 7277
rect 4502 7101 4536 7277
rect 4620 7101 4654 7277
rect 4738 7101 4772 7277
rect 4856 7101 4890 7277
rect 4974 7101 5008 7277
rect 5092 7101 5126 7277
rect -3101 6930 -2725 6964
rect -3794 6755 -3418 6789
rect -3594 6626 -3418 6660
rect -3101 6812 -2725 6846
rect 6355 6973 6389 7349
rect 6473 6973 6507 7349
rect 6591 6973 6625 7349
rect 6709 6973 6743 7349
rect 6827 6973 6861 7349
rect 6945 6973 6979 7349
rect 7063 6973 7097 7349
rect 7497 6977 7531 7353
rect 7615 6977 7649 7353
rect 7733 6977 7767 7353
rect 7851 6977 7885 7353
rect 7969 6977 8003 7353
rect 8087 6977 8121 7353
rect 36767 7732 37143 7766
rect 36767 7613 37143 7647
rect 8205 6977 8239 7353
rect 10581 7099 10615 7275
rect 10699 7099 10733 7275
rect 10817 7099 10851 7275
rect 10935 7099 10969 7275
rect 11053 7099 11087 7275
rect 11171 7099 11205 7275
rect 11289 7099 11323 7275
rect 11407 7099 11441 7275
rect 11525 7099 11559 7275
rect 11643 7099 11677 7275
rect -3594 6508 -3418 6542
rect -3594 6390 -3418 6424
rect 12906 6971 12940 7347
rect 13024 6971 13058 7347
rect 13142 6971 13176 7347
rect 13260 6971 13294 7347
rect 13378 6971 13412 7347
rect 13496 6971 13530 7347
rect 13614 6971 13648 7347
rect 14048 6975 14082 7351
rect 14166 6975 14200 7351
rect 14284 6975 14318 7351
rect 14402 6975 14436 7351
rect 14520 6975 14554 7351
rect 14638 6975 14672 7351
rect 14756 6975 14790 7351
rect 17236 7100 17270 7276
rect 17354 7100 17388 7276
rect 17472 7100 17506 7276
rect 17590 7100 17624 7276
rect 17708 7100 17742 7276
rect 17826 7100 17860 7276
rect 17944 7100 17978 7276
rect 18062 7100 18096 7276
rect 18180 7100 18214 7276
rect 18298 7100 18332 7276
rect 6784 6390 6818 6566
rect 6902 6390 6936 6566
rect 7020 6390 7054 6566
rect 7138 6390 7172 6566
rect 7926 6394 7960 6570
rect 8044 6394 8078 6570
rect 8162 6394 8196 6570
rect 8280 6394 8314 6570
rect 19561 6972 19595 7348
rect 19679 6972 19713 7348
rect 19797 6972 19831 7348
rect 19915 6972 19949 7348
rect 20033 6972 20067 7348
rect 20151 6972 20185 7348
rect 20269 6972 20303 7348
rect 20703 6976 20737 7352
rect 20821 6976 20855 7352
rect 20939 6976 20973 7352
rect 21057 6976 21091 7352
rect 21175 6976 21209 7352
rect 21293 6976 21327 7352
rect 29734 7377 29768 7553
rect 29852 7377 29886 7553
rect 29970 7377 30004 7553
rect 30088 7377 30122 7553
rect 30206 7377 30240 7553
rect 30324 7377 30358 7553
rect 30442 7377 30476 7553
rect 30560 7377 30594 7553
rect 30678 7377 30712 7553
rect 30796 7377 30830 7553
rect 36767 7495 37143 7529
rect 36767 7377 37143 7411
rect 21411 6976 21445 7352
rect 23858 7101 23892 7277
rect 23976 7101 24010 7277
rect 24094 7101 24128 7277
rect 24212 7101 24246 7277
rect 24330 7101 24364 7277
rect 24448 7101 24482 7277
rect 24566 7101 24600 7277
rect 24684 7101 24718 7277
rect 24802 7101 24836 7277
rect 24920 7101 24954 7277
rect -3594 6272 -3418 6306
rect 13335 6388 13369 6564
rect 13453 6388 13487 6564
rect 13571 6388 13605 6564
rect 13689 6388 13723 6564
rect 14477 6392 14511 6568
rect 14595 6392 14629 6568
rect 14713 6392 14747 6568
rect 14831 6392 14865 6568
rect 26183 6973 26217 7349
rect 26301 6973 26335 7349
rect 26419 6973 26453 7349
rect 26537 6973 26571 7349
rect 26655 6973 26689 7349
rect 26773 6973 26807 7349
rect 26891 6973 26925 7349
rect 27325 6977 27359 7353
rect 27443 6977 27477 7353
rect 27561 6977 27595 7353
rect 27679 6977 27713 7353
rect 27797 6977 27831 7353
rect 27915 6977 27949 7353
rect 28033 6977 28067 7353
rect 19990 6389 20024 6565
rect 20108 6389 20142 6565
rect 20226 6389 20260 6565
rect 20344 6389 20378 6565
rect 21132 6393 21166 6569
rect 21250 6393 21284 6569
rect 21368 6393 21402 6569
rect 21486 6393 21520 6569
rect 31478 6910 31512 7086
rect 31596 6910 31630 7086
rect 31714 6910 31748 7086
rect 31832 6910 31866 7086
rect 31962 6910 31996 7286
rect 32080 6910 32114 7286
rect 32198 6910 32232 7286
rect 32316 6910 32350 7286
rect 32434 6910 32468 7286
rect 32552 6910 32586 7286
rect 32670 6910 32704 7286
rect 36767 7259 37143 7293
rect 32799 6910 32833 7086
rect 32917 6910 32951 7086
rect 33035 6910 33069 7086
rect 36967 7140 37143 7174
rect 33153 6910 33187 7086
rect 33271 6907 33305 7083
rect 33389 6907 33423 7083
rect 33507 6907 33541 7083
rect 33625 6907 33659 7083
rect 33743 6907 33777 7083
rect 33861 6907 33895 7083
rect 33979 6907 34013 7083
rect 34097 6907 34131 7083
rect 34215 6907 34249 7083
rect 34333 6907 34367 7083
rect 36967 7022 37143 7056
rect 26612 6390 26646 6566
rect 26730 6390 26764 6566
rect 26848 6390 26882 6566
rect 26966 6390 27000 6566
rect 27754 6394 27788 6570
rect 27872 6394 27906 6570
rect 27990 6394 28024 6570
rect 28108 6394 28142 6570
rect -3596 5879 -3420 5913
rect -3596 5761 -3420 5795
rect 31905 6217 31939 6593
rect 32023 6217 32057 6593
rect 32141 6217 32175 6593
rect 32259 6217 32293 6593
rect 32377 6217 32411 6593
rect 32495 6217 32529 6593
rect 32613 6217 32647 6593
rect 36967 6904 37143 6938
rect 36967 6786 37143 6820
rect 36963 6216 37139 6250
rect 36963 6098 37139 6132
rect 36963 5980 37139 6014
rect -3596 5643 -3420 5677
rect -3596 5525 -3420 5559
rect -3796 5395 -3420 5429
rect -3103 5452 -2727 5486
rect 4044 5451 4078 5627
rect 4162 5451 4196 5627
rect 4280 5451 4314 5627
rect 4398 5451 4432 5627
rect 4516 5451 4550 5627
rect 4634 5451 4668 5627
rect 4752 5451 4786 5627
rect 4870 5451 4904 5627
rect 4988 5451 5022 5627
rect 5106 5451 5140 5627
rect 10595 5449 10629 5625
rect -3796 5277 -3420 5311
rect -3103 5334 -2727 5368
rect -3796 5159 -3420 5193
rect -3103 5216 -2727 5250
rect 10713 5449 10747 5625
rect 10831 5449 10865 5625
rect 10949 5449 10983 5625
rect 11067 5449 11101 5625
rect 11185 5449 11219 5625
rect 11303 5449 11337 5625
rect 11421 5449 11455 5625
rect 11539 5449 11573 5625
rect 11657 5449 11691 5625
rect 17250 5450 17284 5626
rect 17368 5450 17402 5626
rect 17486 5450 17520 5626
rect 17604 5450 17638 5626
rect 17722 5450 17756 5626
rect 17840 5450 17874 5626
rect 17958 5450 17992 5626
rect 18076 5450 18110 5626
rect 18194 5450 18228 5626
rect 18312 5450 18346 5626
rect 23872 5451 23906 5627
rect 23990 5451 24024 5627
rect 24108 5451 24142 5627
rect 24226 5451 24260 5627
rect 24344 5451 24378 5627
rect 24462 5451 24496 5627
rect 24580 5451 24614 5627
rect 24698 5451 24732 5627
rect 24816 5451 24850 5627
rect 24934 5451 24968 5627
rect 36963 5862 37139 5896
rect 36763 5775 37139 5809
rect 36763 5657 37139 5691
rect 36763 5539 37139 5573
rect -3103 5098 -2727 5132
rect -3796 5041 -3420 5075
rect -3796 4923 -3420 4957
rect -3796 4805 -3420 4839
rect -3103 4980 -2727 5014
rect -3103 4862 -2727 4896
rect -3796 4687 -3420 4721
rect -3596 4558 -3420 4592
rect -3103 4744 -2727 4778
rect 5508 4834 5542 5010
rect 5626 4834 5660 5010
rect 5744 4834 5778 5010
rect 5862 4834 5896 5010
rect 5992 4834 6026 5210
rect 6110 4834 6144 5210
rect 6228 4834 6262 5210
rect 6346 4834 6380 5210
rect 6464 4834 6498 5210
rect 6582 4834 6616 5210
rect 6700 4834 6734 5210
rect 6829 4834 6863 5010
rect 6947 4834 6981 5010
rect 7065 4834 7099 5010
rect 7183 4834 7217 5010
rect 7406 4834 7440 5010
rect 7524 4834 7558 5010
rect 7642 4834 7676 5010
rect 7760 4834 7794 5010
rect 7890 4834 7924 5210
rect 8008 4834 8042 5210
rect 8126 4834 8160 5210
rect 8244 4834 8278 5210
rect 8362 4834 8396 5210
rect 8480 4834 8514 5210
rect 8598 4834 8632 5210
rect 8727 4834 8761 5010
rect 8845 4834 8879 5010
rect 8963 4834 8997 5010
rect 9081 4834 9115 5010
rect -3596 4440 -3420 4474
rect 1137 4525 1171 4701
rect 1255 4525 1289 4701
rect 1373 4525 1407 4701
rect 1491 4525 1525 4701
rect 1609 4525 1643 4701
rect 1727 4525 1761 4701
rect 1845 4525 1879 4701
rect 1963 4525 1997 4701
rect 2081 4525 2115 4701
rect 2199 4525 2233 4701
rect -3596 4322 -3420 4356
rect -3596 4204 -3420 4238
rect -3594 3810 -3418 3844
rect -3594 3692 -3418 3726
rect 4039 3847 4073 4023
rect 4157 3847 4191 4023
rect 4275 3847 4309 4023
rect 4393 3847 4427 4023
rect 4511 3847 4545 4023
rect 4629 3847 4663 4023
rect 4747 3847 4781 4023
rect 4865 3847 4899 4023
rect 4983 3847 5017 4023
rect 5101 3847 5135 4023
rect 5935 4141 5969 4517
rect 6053 4141 6087 4517
rect 6171 4141 6205 4517
rect 6289 4141 6323 4517
rect 6407 4141 6441 4517
rect 6525 4141 6559 4517
rect 6643 4141 6677 4517
rect -3594 3574 -3418 3608
rect 12059 4832 12093 5008
rect 12177 4832 12211 5008
rect 12295 4832 12329 5008
rect 12413 4832 12447 5008
rect 12543 4832 12577 5208
rect 12661 4832 12695 5208
rect 12779 4832 12813 5208
rect 12897 4832 12931 5208
rect 13015 4832 13049 5208
rect 13133 4832 13167 5208
rect 13251 4832 13285 5208
rect 13380 4832 13414 5008
rect 13498 4832 13532 5008
rect 13616 4832 13650 5008
rect 13734 4832 13768 5008
rect 13957 4832 13991 5008
rect 14075 4832 14109 5008
rect 14193 4832 14227 5008
rect 14311 4832 14345 5008
rect 14441 4832 14475 5208
rect 14559 4832 14593 5208
rect 14677 4832 14711 5208
rect 14795 4832 14829 5208
rect 14913 4832 14947 5208
rect 15031 4832 15065 5208
rect 15149 4832 15183 5208
rect 15278 4832 15312 5008
rect 15396 4832 15430 5008
rect 15514 4832 15548 5008
rect 15632 4832 15666 5008
rect 7833 4141 7867 4517
rect 7951 4141 7985 4517
rect 8069 4141 8103 4517
rect 8187 4141 8221 4517
rect 8305 4141 8339 4517
rect 8423 4141 8457 4517
rect 8541 4141 8575 4517
rect 10590 3845 10624 4021
rect 10708 3845 10742 4021
rect 10826 3845 10860 4021
rect 10944 3845 10978 4021
rect 11062 3845 11096 4021
rect 11180 3845 11214 4021
rect 11298 3845 11332 4021
rect 11416 3845 11450 4021
rect 11534 3845 11568 4021
rect 11652 3845 11686 4021
rect 12486 4139 12520 4515
rect 12604 4139 12638 4515
rect 12722 4139 12756 4515
rect 12840 4139 12874 4515
rect 12958 4139 12992 4515
rect 13076 4139 13110 4515
rect 13194 4139 13228 4515
rect -3594 3456 -3418 3490
rect -3794 3326 -3418 3360
rect -3101 3383 -2725 3417
rect -3794 3208 -3418 3242
rect -3101 3265 -2725 3299
rect 18714 4833 18748 5009
rect 18832 4833 18866 5009
rect 18950 4833 18984 5009
rect 19068 4833 19102 5009
rect 19198 4833 19232 5209
rect 19316 4833 19350 5209
rect 19434 4833 19468 5209
rect 19552 4833 19586 5209
rect 19670 4833 19704 5209
rect 19788 4833 19822 5209
rect 19906 4833 19940 5209
rect 20035 4833 20069 5009
rect 20153 4833 20187 5009
rect 20271 4833 20305 5009
rect 20389 4833 20423 5009
rect 20612 4833 20646 5009
rect 20730 4833 20764 5009
rect 20848 4833 20882 5009
rect 20966 4833 21000 5009
rect 21096 4833 21130 5209
rect 21214 4833 21248 5209
rect 21332 4833 21366 5209
rect 21450 4833 21484 5209
rect 21568 4833 21602 5209
rect 21686 4833 21720 5209
rect 21804 4833 21838 5209
rect 36763 5421 37139 5455
rect 21933 4833 21967 5009
rect 22051 4833 22085 5009
rect 22169 4833 22203 5009
rect 22287 4833 22321 5009
rect 14384 4139 14418 4515
rect 14502 4139 14536 4515
rect 14620 4139 14654 4515
rect 14738 4139 14772 4515
rect 14856 4139 14890 4515
rect 14974 4139 15008 4515
rect 15092 4139 15126 4515
rect 17245 3846 17279 4022
rect 17363 3846 17397 4022
rect 17481 3846 17515 4022
rect 17599 3846 17633 4022
rect 17717 3846 17751 4022
rect 17835 3846 17869 4022
rect 17953 3846 17987 4022
rect 18071 3846 18105 4022
rect 18189 3846 18223 4022
rect 18307 3846 18341 4022
rect 19141 4140 19175 4516
rect 19259 4140 19293 4516
rect 19377 4140 19411 4516
rect 19495 4140 19529 4516
rect 19613 4140 19647 4516
rect 19731 4140 19765 4516
rect 19849 4140 19883 4516
rect -3794 3090 -3418 3124
rect -3101 3147 -2725 3181
rect 25336 4834 25370 5010
rect 25454 4834 25488 5010
rect 25572 4834 25606 5010
rect 25690 4834 25724 5010
rect 25820 4834 25854 5210
rect 25938 4834 25972 5210
rect 26056 4834 26090 5210
rect 26174 4834 26208 5210
rect 26292 4834 26326 5210
rect 26410 4834 26444 5210
rect 26528 4834 26562 5210
rect 26657 4834 26691 5010
rect 26775 4834 26809 5010
rect 26893 4834 26927 5010
rect 27011 4834 27045 5010
rect 27234 4834 27268 5010
rect 27352 4834 27386 5010
rect 27470 4834 27504 5010
rect 27588 4834 27622 5010
rect 27718 4834 27752 5210
rect 27836 4834 27870 5210
rect 27954 4834 27988 5210
rect 28072 4834 28106 5210
rect 28190 4834 28224 5210
rect 28308 4834 28342 5210
rect 28426 4834 28460 5210
rect 36763 5308 37139 5342
rect 36763 5190 37139 5224
rect 28555 4834 28589 5010
rect 28673 4834 28707 5010
rect 28791 4834 28825 5010
rect 28909 4834 28943 5010
rect 36763 5072 37139 5106
rect 36763 4954 37139 4988
rect 21039 4140 21073 4516
rect 21157 4140 21191 4516
rect 21275 4140 21309 4516
rect 21393 4140 21427 4516
rect 21511 4140 21545 4516
rect 21629 4140 21663 4516
rect 21747 4140 21781 4516
rect 23867 3847 23901 4023
rect 23985 3847 24019 4023
rect 24103 3847 24137 4023
rect 24221 3847 24255 4023
rect 24339 3847 24373 4023
rect 24457 3847 24491 4023
rect 24575 3847 24609 4023
rect 24693 3847 24727 4023
rect 24811 3847 24845 4023
rect 24929 3847 24963 4023
rect 25763 4141 25797 4517
rect 25881 4141 25915 4517
rect 25999 4141 26033 4517
rect 26117 4141 26151 4517
rect 26235 4141 26269 4517
rect 26353 4141 26387 4517
rect 26471 4141 26505 4517
rect -3101 3029 -2725 3063
rect -3794 2972 -3418 3006
rect -3794 2854 -3418 2888
rect -3794 2736 -3418 2770
rect -3101 2911 -2725 2945
rect 36763 4836 37139 4870
rect 36763 4718 37139 4752
rect 36763 4600 37139 4634
rect 27661 4141 27695 4517
rect 27779 4141 27813 4517
rect 27897 4141 27931 4517
rect 28015 4141 28049 4517
rect 28133 4141 28167 4517
rect 28251 4141 28285 4517
rect 28369 4141 28403 4517
rect 29731 4307 29765 4483
rect 29849 4307 29883 4483
rect 29967 4307 30001 4483
rect 30085 4307 30119 4483
rect 30203 4307 30237 4483
rect 30321 4307 30355 4483
rect 30439 4307 30473 4483
rect 30557 4307 30591 4483
rect 30675 4307 30709 4483
rect 30793 4307 30827 4483
rect 36763 4481 37139 4515
rect 36763 4363 37139 4397
rect 36763 4245 37139 4279
rect 36763 4127 37139 4161
rect 36963 4008 37139 4042
rect 36963 3890 37139 3924
rect 36963 3772 37139 3806
rect 36963 3654 37139 3688
rect 36963 3072 37139 3106
rect -3101 2793 -2725 2827
rect -3794 2618 -3418 2652
rect -3594 2489 -3418 2523
rect -3101 2675 -2725 2709
rect 31478 2562 31512 2738
rect 31596 2562 31630 2738
rect 31714 2562 31748 2738
rect 31832 2562 31866 2738
rect 31962 2562 31996 2938
rect 32080 2562 32114 2938
rect 32198 2562 32232 2938
rect 32316 2562 32350 2938
rect 32434 2562 32468 2938
rect 32552 2562 32586 2938
rect 32670 2562 32704 2938
rect 36963 2954 37139 2988
rect 36963 2836 37139 2870
rect 32799 2562 32833 2738
rect 32917 2562 32951 2738
rect 33035 2562 33069 2738
rect 33153 2562 33187 2738
rect 33271 2559 33305 2735
rect -3594 2371 -3418 2405
rect -3594 2253 -3418 2287
rect 33389 2559 33423 2735
rect 33507 2559 33541 2735
rect 33625 2559 33659 2735
rect 33743 2559 33777 2735
rect 33861 2559 33895 2735
rect 33979 2559 34013 2735
rect 34097 2559 34131 2735
rect 34215 2559 34249 2735
rect 34333 2559 34367 2735
rect 36963 2718 37139 2752
rect 36763 2631 37139 2665
rect -3594 2135 -3418 2169
rect -3596 1742 -3420 1776
rect -3596 1624 -3420 1658
rect -3596 1506 -3420 1540
rect -3596 1388 -3420 1422
rect -3796 1258 -3420 1292
rect -3103 1315 -2727 1349
rect 7847 1344 7881 1520
rect 7965 1344 7999 1520
rect 8083 1344 8117 1520
rect 8201 1344 8235 1520
rect 8319 1344 8353 1520
rect 8437 1344 8471 1520
rect 8555 1344 8589 1520
rect 8673 1344 8707 1520
rect 8791 1344 8825 1520
rect 8909 1344 8943 1520
rect 14401 1349 14435 1525
rect 14519 1349 14553 1525
rect 14637 1349 14671 1525
rect 14755 1349 14789 1525
rect 14873 1349 14907 1525
rect 14991 1349 15025 1525
rect 15109 1349 15143 1525
rect 15227 1349 15261 1525
rect 15345 1349 15379 1525
rect 15463 1349 15497 1525
rect 21050 1337 21084 1513
rect 21168 1337 21202 1513
rect 21286 1337 21320 1513
rect 21404 1337 21438 1513
rect 21522 1337 21556 1513
rect 21640 1337 21674 1513
rect 21758 1337 21792 1513
rect 21876 1337 21910 1513
rect 21994 1337 22028 1513
rect 22112 1337 22146 1513
rect 29738 1462 29772 1638
rect 29856 1462 29890 1638
rect 29974 1462 30008 1638
rect 30092 1462 30126 1638
rect 30210 1462 30244 1638
rect 30328 1462 30362 1638
rect 30446 1462 30480 1638
rect 30564 1462 30598 1638
rect 30682 1462 30716 1638
rect 30800 1462 30834 1638
rect 31905 1869 31939 2245
rect 32023 1869 32057 2245
rect 32141 1869 32175 2245
rect 32259 1869 32293 2245
rect 32377 1869 32411 2245
rect 32495 1869 32529 2245
rect 32613 1869 32647 2245
rect 36763 2513 37139 2547
rect 36763 2395 37139 2429
rect 36763 2277 37139 2311
rect 36763 2164 37139 2198
rect 36763 2046 37139 2080
rect 36763 1928 37139 1962
rect 36763 1810 37139 1844
rect 36763 1692 37139 1726
rect 36763 1574 37139 1608
rect -3796 1140 -3420 1174
rect -3103 1197 -2727 1231
rect -3796 1022 -3420 1056
rect -3103 1079 -2727 1113
rect -3103 961 -2727 995
rect -3796 904 -3420 938
rect -3796 786 -3420 820
rect -3796 668 -3420 702
rect -3103 843 -2727 877
rect 36763 1456 37139 1490
rect 36763 1337 37139 1371
rect 36763 1219 37139 1253
rect 36763 1101 37139 1135
rect 36763 983 37139 1017
rect 36963 864 37139 898
rect -3103 725 -2727 759
rect 36963 746 37139 780
rect -3796 550 -3420 584
rect -3596 421 -3420 455
rect -3103 607 -2727 641
rect 36963 628 37139 662
rect 36963 510 37139 544
rect -3596 303 -3420 337
rect -3596 185 -3420 219
rect -3596 67 -3420 101
<< psubdiff >>
rect 6603 26845 6837 26879
rect 6603 26755 6649 26845
rect 6812 26755 6837 26845
rect 6603 26724 6837 26755
rect 13116 26842 13350 26876
rect 13116 26752 13162 26842
rect 13325 26752 13350 26842
rect 13116 26721 13350 26752
rect 19650 26837 19884 26871
rect 19650 26747 19696 26837
rect 19859 26747 19884 26837
rect 19650 26716 19884 26747
rect 26208 26841 26442 26875
rect 26208 26751 26254 26841
rect 26417 26751 26442 26841
rect 26208 26720 26442 26751
rect 8100 26474 8255 26520
rect 8100 26311 8131 26474
rect 8221 26311 8255 26474
rect 8100 26286 8255 26311
rect 9242 26472 9397 26518
rect 9242 26309 9273 26472
rect 9363 26309 9397 26472
rect 14613 26471 14768 26517
rect 9242 26284 9397 26309
rect 14613 26308 14644 26471
rect 14734 26308 14768 26471
rect 14613 26283 14768 26308
rect 15755 26469 15910 26515
rect 15755 26306 15786 26469
rect 15876 26306 15910 26469
rect 21147 26466 21302 26512
rect 15755 26281 15910 26306
rect 21147 26303 21178 26466
rect 21268 26303 21302 26466
rect 21147 26278 21302 26303
rect 22289 26464 22444 26510
rect 22289 26301 22320 26464
rect 22410 26301 22444 26464
rect 27705 26470 27860 26516
rect 22289 26276 22444 26301
rect 27705 26307 27736 26470
rect 27826 26307 27860 26470
rect 27705 26282 27860 26307
rect 28847 26468 29002 26514
rect 28847 26305 28878 26468
rect 28968 26305 29002 26468
rect 28847 26280 29002 26305
rect 6617 25195 6851 25229
rect 6617 25105 6663 25195
rect 6826 25105 6851 25195
rect 6617 25074 6851 25105
rect 13130 25192 13364 25226
rect 13130 25102 13176 25192
rect 13339 25102 13364 25192
rect 13130 25071 13364 25102
rect 19664 25187 19898 25221
rect 19664 25097 19710 25187
rect 19873 25097 19898 25187
rect 19664 25066 19898 25097
rect 6612 23591 6846 23625
rect 6612 23501 6658 23591
rect 6821 23501 6846 23591
rect 26222 25191 26456 25225
rect 26222 25101 26268 25191
rect 26431 25101 26456 25191
rect 26222 25070 26456 25101
rect 13125 23588 13359 23622
rect 6612 23470 6846 23501
rect 8044 23431 8199 23477
rect 13125 23498 13171 23588
rect 13334 23498 13359 23588
rect 19659 23583 19893 23617
rect 13125 23467 13359 23498
rect 8044 23268 8075 23431
rect 8165 23268 8199 23431
rect 8044 23243 8199 23268
rect 14557 23428 14712 23474
rect 19659 23493 19705 23583
rect 19868 23493 19893 23583
rect 38719 23904 38825 23946
rect 26217 23587 26451 23621
rect 19659 23462 19893 23493
rect 14557 23265 14588 23428
rect 14678 23265 14712 23428
rect 14557 23240 14712 23265
rect 21091 23423 21246 23469
rect 26217 23497 26263 23587
rect 26426 23497 26451 23587
rect 26217 23466 26451 23497
rect 21091 23260 21122 23423
rect 21212 23260 21246 23423
rect 21091 23235 21246 23260
rect 27649 23427 27804 23473
rect 27649 23264 27680 23427
rect 27770 23264 27804 23427
rect 27649 23239 27804 23264
rect 38719 23800 38743 23904
rect 38789 23800 38825 23904
rect 38719 23760 38825 23800
rect 9067 21237 9301 21271
rect 9067 21147 9092 21237
rect 9255 21147 9301 21237
rect 9067 21116 9301 21147
rect 15625 21233 15859 21267
rect 15625 21143 15650 21233
rect 15813 21143 15859 21233
rect 15625 21112 15859 21143
rect 22159 21238 22393 21272
rect 22159 21148 22184 21238
rect 22347 21148 22393 21238
rect 22159 21117 22393 21148
rect 28672 21241 28906 21275
rect 28672 21151 28697 21241
rect 28860 21151 28906 21241
rect 28672 21120 28906 21151
rect 6507 20864 6662 20910
rect 6507 20701 6541 20864
rect 6631 20701 6662 20864
rect 6507 20676 6662 20701
rect 7649 20866 7804 20912
rect 7649 20703 7683 20866
rect 7773 20703 7804 20866
rect 13065 20860 13220 20906
rect 7649 20678 7804 20703
rect 13065 20697 13099 20860
rect 13189 20697 13220 20860
rect 13065 20672 13220 20697
rect 14207 20862 14362 20908
rect 14207 20699 14241 20862
rect 14331 20699 14362 20862
rect 19599 20865 19754 20911
rect 14207 20674 14362 20699
rect 19599 20702 19633 20865
rect 19723 20702 19754 20865
rect 19599 20677 19754 20702
rect 20741 20867 20896 20913
rect 20741 20704 20775 20867
rect 20865 20704 20896 20867
rect 26112 20868 26267 20914
rect 20741 20679 20896 20704
rect 26112 20705 26146 20868
rect 26236 20705 26267 20868
rect 26112 20680 26267 20705
rect 27254 20870 27409 20916
rect 27254 20707 27288 20870
rect 27378 20707 27409 20870
rect 27254 20682 27409 20707
rect 38719 20760 38825 20802
rect 9053 19587 9287 19621
rect 9053 19497 9078 19587
rect 9241 19497 9287 19587
rect 15611 19583 15845 19617
rect 9053 19466 9287 19497
rect 15611 19493 15636 19583
rect 15799 19493 15845 19583
rect 22145 19588 22379 19622
rect 15611 19462 15845 19493
rect 9058 17983 9292 18017
rect 9058 17893 9083 17983
rect 9246 17893 9292 17983
rect 22145 19498 22170 19588
rect 22333 19498 22379 19588
rect 38719 20656 38743 20760
rect 38789 20656 38825 20760
rect 38719 20616 38825 20656
rect 28658 19591 28892 19625
rect 22145 19467 22379 19498
rect 15616 17979 15850 18013
rect 7705 17823 7860 17869
rect 9058 17862 9292 17893
rect 15616 17889 15641 17979
rect 15804 17889 15850 17979
rect 28658 19501 28683 19591
rect 28846 19501 28892 19591
rect 28658 19470 28892 19501
rect 22150 17984 22384 18018
rect 7705 17660 7739 17823
rect 7829 17660 7860 17823
rect 7705 17635 7860 17660
rect 14263 17819 14418 17865
rect 15616 17858 15850 17889
rect 22150 17894 22175 17984
rect 22338 17894 22384 17984
rect 28663 17987 28897 18021
rect 14263 17656 14297 17819
rect 14387 17656 14418 17819
rect 14263 17631 14418 17656
rect 20797 17824 20952 17870
rect 22150 17863 22384 17894
rect 28663 17897 28688 17987
rect 28851 17897 28897 17987
rect 20797 17661 20831 17824
rect 20921 17661 20952 17824
rect 20797 17636 20952 17661
rect 27310 17827 27465 17873
rect 28663 17866 28897 17897
rect 27310 17664 27344 17827
rect 27434 17664 27465 17827
rect 27310 17639 27465 17664
rect 38715 17628 38821 17670
rect 38715 17524 38739 17628
rect 38785 17524 38821 17628
rect 38715 17484 38821 17524
rect -1823 15520 -1725 15578
rect -1823 15388 -1803 15520
rect -1747 15388 -1725 15520
rect -1823 15326 -1725 15388
rect 8301 14256 8513 14286
rect 8301 14200 8341 14256
rect 8475 14200 8513 14256
rect 8301 14178 8513 14200
rect 14850 14255 15062 14285
rect 14850 14199 14890 14255
rect 15024 14199 15062 14255
rect 14850 14177 15062 14199
rect 21504 14276 21716 14306
rect 21504 14220 21544 14276
rect 21678 14220 21716 14276
rect 21504 14198 21716 14220
rect 30157 14109 30369 14139
rect 30157 14053 30197 14109
rect 30331 14053 30369 14109
rect 30157 14031 30369 14053
rect -1825 13452 -1727 13510
rect -1825 13320 -1805 13452
rect -1749 13320 -1727 13452
rect -1825 13258 -1727 13320
rect 38715 14484 38821 14526
rect 38715 14380 38739 14484
rect 38785 14380 38821 14484
rect 38715 14340 38821 14380
rect 33758 13701 33970 13731
rect 33758 13645 33798 13701
rect 33932 13645 33970 13701
rect 33758 13623 33970 13645
rect 1637 12356 1849 12386
rect 1637 12300 1677 12356
rect 1811 12300 1849 12356
rect 1637 12278 1849 12300
rect 4799 12294 5033 12328
rect 4799 12204 4845 12294
rect 5008 12204 5033 12294
rect 4799 12173 5033 12204
rect 11348 12382 11582 12416
rect 11348 12292 11394 12382
rect 11557 12292 11582 12382
rect 11348 12261 11582 12292
rect 32168 12900 32410 12912
rect 18002 12314 18236 12348
rect 18002 12224 18048 12314
rect 18211 12224 18236 12314
rect 18002 12193 18236 12224
rect 32168 12798 32215 12900
rect 32350 12798 32410 12900
rect 32168 12781 32410 12798
rect 24627 12382 24861 12416
rect 24627 12292 24673 12382
rect 24836 12292 24861 12382
rect 24627 12261 24861 12292
rect 12845 12011 13000 12057
rect 6296 11923 6451 11969
rect 6296 11760 6327 11923
rect 6417 11760 6451 11923
rect 6296 11735 6451 11760
rect 7438 11921 7593 11967
rect 7438 11758 7469 11921
rect 7559 11758 7593 11921
rect 7438 11733 7593 11758
rect 12845 11848 12876 12011
rect 12966 11848 13000 12011
rect 12845 11823 13000 11848
rect 13987 12009 14142 12055
rect 13987 11846 14018 12009
rect 14108 11846 14142 12009
rect 26124 12011 26279 12057
rect 19499 11943 19654 11989
rect 13987 11821 14142 11846
rect 19499 11780 19530 11943
rect 19620 11780 19654 11943
rect 19499 11755 19654 11780
rect 20641 11941 20796 11987
rect 20641 11778 20672 11941
rect 20762 11778 20796 11941
rect 20641 11753 20796 11778
rect 26124 11848 26155 12011
rect 26245 11848 26279 12011
rect 26124 11823 26279 11848
rect 27266 12009 27421 12055
rect 27266 11846 27297 12009
rect 27387 11846 27421 12009
rect 27266 11821 27421 11846
rect -1823 11383 -1725 11441
rect -1823 11251 -1803 11383
rect -1747 11251 -1725 11383
rect -1823 11189 -1725 11251
rect 30152 11538 30364 11568
rect 30152 11482 30192 11538
rect 30326 11482 30364 11538
rect 30152 11460 30364 11482
rect 4813 10644 5047 10678
rect 4813 10554 4859 10644
rect 5022 10554 5047 10644
rect 11362 10732 11596 10766
rect 4813 10523 5047 10554
rect 1629 9771 1841 9801
rect 1629 9715 1669 9771
rect 1803 9715 1841 9771
rect 1629 9693 1841 9715
rect 11362 10642 11408 10732
rect 11571 10642 11596 10732
rect 38719 11282 38825 11324
rect 11362 10611 11596 10642
rect -1825 9315 -1727 9373
rect -1825 9183 -1805 9315
rect -1749 9183 -1727 9315
rect -1825 9121 -1727 9183
rect 18016 10664 18250 10698
rect 18016 10574 18062 10664
rect 18225 10574 18250 10664
rect 24641 10732 24875 10766
rect 18016 10543 18250 10574
rect 4808 9040 5042 9074
rect 24641 10642 24687 10732
rect 24850 10642 24875 10732
rect 24641 10611 24875 10642
rect 11357 9128 11591 9162
rect 4808 8950 4854 9040
rect 5017 8950 5042 9040
rect 11357 9038 11403 9128
rect 11566 9038 11591 9128
rect 11357 9007 11591 9038
rect 4808 8919 5042 8950
rect 12789 8968 12944 9014
rect 38719 11178 38743 11282
rect 38789 11178 38825 11282
rect 38719 11138 38825 11178
rect 18011 9060 18245 9094
rect 33760 9610 33972 9640
rect 33760 9554 33800 9610
rect 33934 9554 33972 9610
rect 33760 9532 33972 9554
rect 24636 9128 24870 9162
rect 6240 8880 6395 8926
rect 6240 8717 6271 8880
rect 6361 8717 6395 8880
rect 12789 8805 12820 8968
rect 12910 8805 12944 8968
rect 18011 8970 18057 9060
rect 18220 8970 18245 9060
rect 24636 9038 24682 9128
rect 24845 9038 24870 9128
rect 24636 9007 24870 9038
rect 18011 8939 18245 8970
rect 26068 8968 26223 9014
rect 12789 8780 12944 8805
rect 19443 8900 19598 8946
rect 6240 8692 6395 8717
rect 19443 8737 19474 8900
rect 19564 8737 19598 8900
rect 26068 8805 26099 8968
rect 26189 8805 26223 8968
rect 26068 8780 26223 8805
rect 19443 8712 19598 8737
rect 32170 8809 32412 8821
rect 32170 8707 32217 8809
rect 32352 8707 32412 8809
rect 32170 8690 32412 8707
rect 30152 8505 30364 8535
rect 30152 8449 30192 8505
rect 30326 8449 30364 8505
rect 30152 8427 30364 8449
rect 38719 8138 38825 8180
rect -1825 7246 -1727 7304
rect -1825 7114 -1805 7246
rect -1749 7114 -1727 7246
rect -1825 7052 -1727 7114
rect 1610 6493 1822 6523
rect 1610 6437 1650 6493
rect 1784 6437 1822 6493
rect 4791 6514 5025 6548
rect 1610 6415 1822 6437
rect 4791 6424 4837 6514
rect 5000 6424 5025 6514
rect 4791 6393 5025 6424
rect 38719 8034 38743 8138
rect 38789 8034 38825 8138
rect 38719 7994 38825 8034
rect 11342 6512 11576 6546
rect 11342 6422 11388 6512
rect 11551 6422 11576 6512
rect 11342 6391 11576 6422
rect 17997 6513 18231 6547
rect 17997 6423 18043 6513
rect 18206 6423 18231 6513
rect 17997 6392 18231 6423
rect 30223 6585 30435 6615
rect 24619 6514 24853 6548
rect 24619 6424 24665 6514
rect 24828 6424 24853 6514
rect 24619 6393 24853 6424
rect 30223 6529 30263 6585
rect 30397 6529 30435 6585
rect 30223 6507 30435 6529
rect 6288 6143 6443 6189
rect 6288 5980 6319 6143
rect 6409 5980 6443 6143
rect 6288 5955 6443 5980
rect 7430 6141 7585 6187
rect 7430 5978 7461 6141
rect 7551 5978 7585 6141
rect 12839 6141 12994 6187
rect 7430 5953 7585 5978
rect 12839 5978 12870 6141
rect 12960 5978 12994 6141
rect 12839 5953 12994 5978
rect 13981 6139 14136 6185
rect 13981 5976 14012 6139
rect 14102 5976 14136 6139
rect 19494 6142 19649 6188
rect 13981 5951 14136 5976
rect 19494 5979 19525 6142
rect 19615 5979 19649 6142
rect 19494 5954 19649 5979
rect 20636 6140 20791 6186
rect 20636 5977 20667 6140
rect 20757 5977 20791 6140
rect 26116 6143 26271 6189
rect 20636 5952 20791 5977
rect 26116 5980 26147 6143
rect 26237 5980 26271 6143
rect 26116 5955 26271 5980
rect 27258 6141 27413 6187
rect 27258 5978 27289 6141
rect 27379 5978 27413 6141
rect 27258 5953 27413 5978
rect 33760 6115 33972 6145
rect 33760 6059 33800 6115
rect 33934 6059 33972 6115
rect 33760 6037 33972 6059
rect -1827 5178 -1729 5236
rect -1827 5046 -1807 5178
rect -1751 5046 -1729 5178
rect -1827 4984 -1729 5046
rect 4805 4864 5039 4898
rect 4805 4774 4851 4864
rect 5014 4774 5039 4864
rect 4805 4743 5039 4774
rect 1626 3733 1838 3763
rect 1626 3677 1666 3733
rect 1800 3677 1838 3733
rect 1626 3655 1838 3677
rect 11356 4862 11590 4896
rect 11356 4772 11402 4862
rect 11565 4772 11590 4862
rect 11356 4741 11590 4772
rect 18011 4863 18245 4897
rect 18011 4773 18057 4863
rect 18220 4773 18245 4863
rect 32170 5314 32412 5326
rect 18011 4742 18245 4773
rect 4800 3260 5034 3294
rect -1825 3109 -1727 3167
rect 4800 3170 4846 3260
rect 5009 3170 5034 3260
rect 24633 4864 24867 4898
rect 24633 4774 24679 4864
rect 24842 4774 24867 4864
rect 32170 5212 32217 5314
rect 32352 5212 32412 5314
rect 32170 5195 32412 5212
rect 38715 5006 38821 5048
rect 24633 4743 24867 4774
rect 11351 3258 11585 3292
rect 4800 3139 5034 3170
rect -1825 2977 -1805 3109
rect -1749 2977 -1727 3109
rect -1825 2915 -1727 2977
rect 6232 3100 6387 3146
rect 11351 3168 11397 3258
rect 11560 3168 11585 3258
rect 38715 4902 38739 5006
rect 38785 4902 38821 5006
rect 38715 4862 38821 4902
rect 18006 3259 18240 3293
rect 11351 3137 11585 3168
rect 6232 2937 6263 3100
rect 6353 2937 6387 3100
rect 6232 2912 6387 2937
rect 12783 3098 12938 3144
rect 18006 3169 18052 3259
rect 18215 3169 18240 3259
rect 30220 3515 30432 3545
rect 30220 3459 30260 3515
rect 30394 3459 30432 3515
rect 30220 3437 30432 3459
rect 24628 3260 24862 3294
rect 18006 3138 18240 3169
rect 12783 2935 12814 3098
rect 12904 2935 12938 3098
rect 12783 2910 12938 2935
rect 19438 3099 19593 3145
rect 24628 3170 24674 3260
rect 24837 3170 24862 3260
rect 24628 3139 24862 3170
rect 19438 2936 19469 3099
rect 19559 2936 19593 3099
rect 19438 2911 19593 2936
rect 26060 3100 26215 3146
rect 26060 2937 26091 3100
rect 26181 2937 26215 3100
rect 26060 2912 26215 2937
rect 8336 2368 8548 2390
rect 8336 2312 8376 2368
rect 8510 2312 8548 2368
rect 8336 2282 8548 2312
rect 14890 2373 15102 2395
rect 14890 2317 14930 2373
rect 15064 2317 15102 2373
rect 14890 2287 15102 2317
rect 21539 2361 21751 2383
rect 21539 2305 21579 2361
rect 21713 2305 21751 2361
rect 21539 2275 21751 2305
rect 33760 1767 33972 1797
rect 33760 1711 33800 1767
rect 33934 1711 33972 1767
rect 33760 1689 33972 1711
rect 38715 1862 38821 1904
rect -1827 1041 -1729 1099
rect -1827 909 -1807 1041
rect -1751 909 -1729 1041
rect -1827 847 -1729 909
rect 38715 1758 38739 1862
rect 38785 1758 38821 1862
rect 38715 1718 38821 1758
rect 32170 966 32412 978
rect 32170 864 32217 966
rect 32352 864 32412 966
rect 32170 847 32412 864
rect 30227 670 30439 700
rect 30227 614 30267 670
rect 30401 614 30439 670
rect 30227 592 30439 614
<< nsubdiff >>
rect 8755 28076 8908 28116
rect 6273 28022 6426 28062
rect 6273 27873 6316 28022
rect 6383 27873 6426 28022
rect 6273 27804 6426 27873
rect 8755 27927 8798 28076
rect 8865 27927 8908 28076
rect 8755 27858 8908 27927
rect 9902 28076 10055 28116
rect 9902 27927 9945 28076
rect 10012 27927 10055 28076
rect 15268 28073 15421 28113
rect 9902 27858 10055 27927
rect 12786 28019 12939 28059
rect 12786 27870 12829 28019
rect 12896 27870 12939 28019
rect 12786 27801 12939 27870
rect 15268 27924 15311 28073
rect 15378 27924 15421 28073
rect 15268 27855 15421 27924
rect 16415 28073 16568 28113
rect 16415 27924 16458 28073
rect 16525 27924 16568 28073
rect 21802 28068 21955 28108
rect 16415 27855 16568 27924
rect 19320 28014 19473 28054
rect 19320 27865 19363 28014
rect 19430 27865 19473 28014
rect 19320 27796 19473 27865
rect 21802 27919 21845 28068
rect 21912 27919 21955 28068
rect 21802 27850 21955 27919
rect 22949 28068 23102 28108
rect 22949 27919 22992 28068
rect 23059 27919 23102 28068
rect 28360 28072 28513 28112
rect 22949 27850 23102 27919
rect 25878 28018 26031 28058
rect 25878 27869 25921 28018
rect 25988 27869 26031 28018
rect 25878 27800 26031 27869
rect 28360 27923 28403 28072
rect 28470 27923 28513 28072
rect 28360 27854 28513 27923
rect 29507 28072 29660 28112
rect 29507 27923 29550 28072
rect 29617 27923 29660 28072
rect 29507 27854 29660 27923
rect 6287 26372 6440 26412
rect 6287 26223 6330 26372
rect 6397 26223 6440 26372
rect 12800 26369 12953 26409
rect 6287 26154 6440 26223
rect 12800 26220 12843 26369
rect 12910 26220 12953 26369
rect 19334 26364 19487 26404
rect 12800 26151 12953 26220
rect 19334 26215 19377 26364
rect 19444 26215 19487 26364
rect 25892 26368 26045 26408
rect 19334 26146 19487 26215
rect 25892 26219 25935 26368
rect 26002 26219 26045 26368
rect 25892 26150 26045 26219
rect 9998 26029 10151 26069
rect 9998 25880 10041 26029
rect 10108 25880 10151 26029
rect 16511 26026 16664 26066
rect 9998 25811 10151 25880
rect 16511 25877 16554 26026
rect 16621 25877 16664 26026
rect 23045 26021 23198 26061
rect 29603 26025 29756 26065
rect 16511 25808 16664 25877
rect 23045 25872 23088 26021
rect 23155 25872 23198 26021
rect 23045 25803 23198 25872
rect 29603 25876 29646 26025
rect 29713 25876 29756 26025
rect 29603 25807 29756 25876
rect 6282 24768 6435 24808
rect 6282 24619 6325 24768
rect 6392 24619 6435 24768
rect 6282 24550 6435 24619
rect 12795 24765 12948 24805
rect 12795 24616 12838 24765
rect 12905 24616 12948 24765
rect 12795 24547 12948 24616
rect 19329 24760 19482 24800
rect 19329 24611 19372 24760
rect 19439 24611 19482 24760
rect 19329 24542 19482 24611
rect 25887 24764 26040 24804
rect 25887 24615 25930 24764
rect 25997 24615 26040 24764
rect 25887 24546 26040 24615
rect 36441 23962 36587 24016
rect 36441 23766 36497 23962
rect 36573 23766 36587 23962
rect 36441 23712 36587 23766
rect 5849 22468 6002 22508
rect 5849 22319 5892 22468
rect 5959 22319 6002 22468
rect 5849 22250 6002 22319
rect 6996 22468 7149 22508
rect 6996 22319 7039 22468
rect 7106 22319 7149 22468
rect 12407 22464 12560 22504
rect 6996 22250 7149 22319
rect 9478 22414 9631 22454
rect 9478 22265 9521 22414
rect 9588 22265 9631 22414
rect 9478 22196 9631 22265
rect 12407 22315 12450 22464
rect 12517 22315 12560 22464
rect 12407 22246 12560 22315
rect 13554 22464 13707 22504
rect 13554 22315 13597 22464
rect 13664 22315 13707 22464
rect 18941 22469 19094 22509
rect 13554 22246 13707 22315
rect 16036 22410 16189 22450
rect 16036 22261 16079 22410
rect 16146 22261 16189 22410
rect 16036 22192 16189 22261
rect 18941 22320 18984 22469
rect 19051 22320 19094 22469
rect 18941 22251 19094 22320
rect 20088 22469 20241 22509
rect 20088 22320 20131 22469
rect 20198 22320 20241 22469
rect 25454 22472 25607 22512
rect 20088 22251 20241 22320
rect 22570 22415 22723 22455
rect 22570 22266 22613 22415
rect 22680 22266 22723 22415
rect 22570 22197 22723 22266
rect 25454 22323 25497 22472
rect 25564 22323 25607 22472
rect 25454 22254 25607 22323
rect 26601 22472 26754 22512
rect 26601 22323 26644 22472
rect 26711 22323 26754 22472
rect 26601 22254 26754 22323
rect 29083 22418 29236 22458
rect 29083 22269 29126 22418
rect 29193 22269 29236 22418
rect 29083 22200 29236 22269
rect 9464 20764 9617 20804
rect 9464 20615 9507 20764
rect 9574 20615 9617 20764
rect 16022 20760 16175 20800
rect 9464 20546 9617 20615
rect 16022 20611 16065 20760
rect 16132 20611 16175 20760
rect 22556 20765 22709 20805
rect 16022 20542 16175 20611
rect 22556 20616 22599 20765
rect 22666 20616 22709 20765
rect 36441 20818 36587 20872
rect 29069 20768 29222 20808
rect 22556 20547 22709 20616
rect 29069 20619 29112 20768
rect 29179 20619 29222 20768
rect 29069 20550 29222 20619
rect 36441 20622 36497 20818
rect 36573 20622 36587 20818
rect 36441 20568 36587 20622
rect 5753 20421 5906 20461
rect 5753 20272 5796 20421
rect 5863 20272 5906 20421
rect 12311 20417 12464 20457
rect 5753 20203 5906 20272
rect 12311 20268 12354 20417
rect 12421 20268 12464 20417
rect 18845 20422 18998 20462
rect 12311 20199 12464 20268
rect 18845 20273 18888 20422
rect 18955 20273 18998 20422
rect 25358 20425 25511 20465
rect 18845 20204 18998 20273
rect 25358 20276 25401 20425
rect 25468 20276 25511 20425
rect 25358 20207 25511 20276
rect 9469 19160 9622 19200
rect 9469 19011 9512 19160
rect 9579 19011 9622 19160
rect 9469 18942 9622 19011
rect 16027 19156 16180 19196
rect 16027 19007 16070 19156
rect 16137 19007 16180 19156
rect 16027 18938 16180 19007
rect 22561 19161 22714 19201
rect 22561 19012 22604 19161
rect 22671 19012 22714 19161
rect 22561 18943 22714 19012
rect 29074 19164 29227 19204
rect 29074 19015 29117 19164
rect 29184 19015 29227 19164
rect 29074 18946 29227 19015
rect 36437 17686 36583 17740
rect 36437 17490 36493 17686
rect 36569 17490 36583 17686
rect 36437 17436 36583 17490
rect -4115 15470 -3971 15594
rect -4115 15348 -4063 15470
rect -4019 15348 -3971 15470
rect -4115 15194 -3971 15348
rect 8061 15464 8305 15502
rect 8061 15394 8117 15464
rect 8253 15394 8305 15464
rect 8061 15372 8305 15394
rect 14610 15463 14854 15501
rect 14610 15393 14666 15463
rect 14802 15393 14854 15463
rect 14610 15371 14854 15393
rect 21264 15484 21508 15522
rect 21264 15414 21320 15484
rect 21456 15414 21508 15484
rect 21264 15392 21508 15414
rect 32110 15376 32531 15410
rect 29917 15317 30161 15355
rect 29917 15247 29973 15317
rect 30109 15247 30161 15317
rect 29917 15225 30161 15247
rect 32110 15231 32173 15376
rect 32482 15231 32531 15376
rect 32110 15210 32531 15231
rect 33518 14909 33762 14947
rect 33518 14839 33574 14909
rect 33710 14839 33762 14909
rect 33518 14817 33762 14839
rect 36437 14542 36583 14596
rect 13500 13613 13653 13653
rect -4117 13402 -3973 13526
rect -4117 13280 -4065 13402
rect -4021 13280 -3973 13402
rect 1397 13564 1641 13602
rect 1397 13494 1453 13564
rect 1589 13494 1641 13564
rect 6951 13525 7104 13565
rect 1397 13472 1641 13494
rect -4117 13126 -3973 13280
rect 4469 13471 4622 13511
rect 4469 13322 4512 13471
rect 4579 13322 4622 13471
rect 4469 13253 4622 13322
rect 6951 13376 6994 13525
rect 7061 13376 7104 13525
rect 6951 13307 7104 13376
rect 8098 13525 8251 13565
rect 8098 13376 8141 13525
rect 8208 13376 8251 13525
rect 8098 13307 8251 13376
rect 11018 13559 11171 13599
rect 11018 13410 11061 13559
rect 11128 13410 11171 13559
rect 11018 13341 11171 13410
rect 13500 13464 13543 13613
rect 13610 13464 13653 13613
rect 13500 13395 13653 13464
rect 14647 13613 14800 13653
rect 14647 13464 14690 13613
rect 14757 13464 14800 13613
rect 26779 13613 26932 13653
rect 20154 13545 20307 13585
rect 14647 13395 14800 13464
rect 17672 13491 17825 13531
rect 17672 13342 17715 13491
rect 17782 13342 17825 13491
rect 17672 13273 17825 13342
rect 20154 13396 20197 13545
rect 20264 13396 20307 13545
rect 20154 13327 20307 13396
rect 21301 13545 21454 13585
rect 21301 13396 21344 13545
rect 21411 13396 21454 13545
rect 21301 13327 21454 13396
rect 24297 13559 24450 13599
rect 24297 13410 24340 13559
rect 24407 13410 24450 13559
rect 24297 13341 24450 13410
rect 26779 13464 26822 13613
rect 26889 13464 26932 13613
rect 26779 13395 26932 13464
rect 27926 13613 28079 13653
rect 27926 13464 27969 13613
rect 28036 13464 28079 13613
rect 27926 13395 28079 13464
rect 36437 14346 36493 14542
rect 36569 14346 36583 14542
rect 36437 14292 36583 14346
rect 29912 12746 30156 12784
rect 29912 12676 29968 12746
rect 30104 12676 30156 12746
rect 29912 12654 30156 12676
rect 4483 11821 4636 11861
rect 4483 11672 4526 11821
rect 4593 11672 4636 11821
rect 11032 11909 11185 11949
rect 11032 11760 11075 11909
rect 11142 11760 11185 11909
rect 17686 11841 17839 11881
rect 11032 11691 11185 11760
rect 17686 11692 17729 11841
rect 17796 11692 17839 11841
rect 24311 11909 24464 11949
rect 24311 11760 24354 11909
rect 24421 11760 24464 11909
rect 4483 11603 4636 11672
rect 17686 11623 17839 11692
rect 24311 11691 24464 11760
rect 14743 11566 14896 11606
rect -4115 11333 -3971 11457
rect -4115 11211 -4063 11333
rect -4019 11211 -3971 11333
rect 8194 11478 8347 11518
rect -4115 11057 -3971 11211
rect 8194 11329 8237 11478
rect 8304 11329 8347 11478
rect 8194 11260 8347 11329
rect 14743 11417 14786 11566
rect 14853 11417 14896 11566
rect 28022 11566 28175 11606
rect 21397 11498 21550 11538
rect 14743 11348 14896 11417
rect 1389 10979 1633 11017
rect 21397 11349 21440 11498
rect 21507 11349 21550 11498
rect 21397 11280 21550 11349
rect 28022 11417 28065 11566
rect 28132 11417 28175 11566
rect 28022 11348 28175 11417
rect 36441 11340 36587 11394
rect 1389 10909 1445 10979
rect 1581 10909 1633 10979
rect 1389 10887 1633 10909
rect 4478 10217 4631 10257
rect 4478 10068 4521 10217
rect 4588 10068 4631 10217
rect 4478 9999 4631 10068
rect -4117 9265 -3973 9389
rect -4117 9143 -4065 9265
rect -4021 9143 -3973 9265
rect 32112 11285 32533 11319
rect 32112 11140 32175 11285
rect 32484 11140 32533 11285
rect 32112 11119 32533 11140
rect 36441 11144 36497 11340
rect 36573 11144 36587 11340
rect 36441 11090 36587 11144
rect 11027 10305 11180 10345
rect 11027 10156 11070 10305
rect 11137 10156 11180 10305
rect 11027 10087 11180 10156
rect -4117 8989 -3973 9143
rect 17681 10237 17834 10277
rect 17681 10088 17724 10237
rect 17791 10088 17834 10237
rect 17681 10019 17834 10088
rect 33520 10818 33764 10856
rect 24306 10305 24459 10345
rect 24306 10156 24349 10305
rect 24416 10156 24459 10305
rect 24306 10087 24459 10156
rect 33520 10748 33576 10818
rect 33712 10748 33764 10818
rect 33520 10726 33764 10748
rect 29912 9713 30156 9751
rect 29912 9643 29968 9713
rect 30104 9643 30156 9713
rect 29912 9621 30156 9643
rect 36441 8196 36587 8250
rect 36441 8000 36497 8196
rect 36573 8000 36587 8196
rect 36441 7946 36587 8000
rect 29983 7793 30227 7831
rect 6943 7745 7096 7785
rect 1370 7701 1614 7739
rect 1370 7631 1426 7701
rect 1562 7631 1614 7701
rect 1370 7609 1614 7631
rect 4461 7691 4614 7731
rect 4461 7542 4504 7691
rect 4571 7542 4614 7691
rect 4461 7473 4614 7542
rect 6943 7596 6986 7745
rect 7053 7596 7096 7745
rect 6943 7527 7096 7596
rect 8090 7745 8243 7785
rect 8090 7596 8133 7745
rect 8200 7596 8243 7745
rect 13494 7743 13647 7783
rect 8090 7527 8243 7596
rect 11012 7689 11165 7729
rect 11012 7540 11055 7689
rect 11122 7540 11165 7689
rect -4117 7196 -3973 7320
rect -4117 7074 -4065 7196
rect -4021 7074 -3973 7196
rect 11012 7471 11165 7540
rect 13494 7594 13537 7743
rect 13604 7594 13647 7743
rect 13494 7525 13647 7594
rect 14641 7743 14794 7783
rect 14641 7594 14684 7743
rect 14751 7594 14794 7743
rect 20149 7744 20302 7784
rect 14641 7525 14794 7594
rect 17667 7690 17820 7730
rect 17667 7541 17710 7690
rect 17777 7541 17820 7690
rect 17667 7472 17820 7541
rect 20149 7595 20192 7744
rect 20259 7595 20302 7744
rect 20149 7526 20302 7595
rect 21296 7744 21449 7784
rect 21296 7595 21339 7744
rect 21406 7595 21449 7744
rect 26771 7745 26924 7785
rect 21296 7526 21449 7595
rect 24289 7691 24442 7731
rect 24289 7542 24332 7691
rect 24399 7542 24442 7691
rect -4117 6920 -3973 7074
rect 24289 7473 24442 7542
rect 26771 7596 26814 7745
rect 26881 7596 26924 7745
rect 26771 7527 26924 7596
rect 27918 7745 28071 7785
rect 27918 7596 27961 7745
rect 28028 7596 28071 7745
rect 29983 7723 30039 7793
rect 30175 7723 30227 7793
rect 29983 7701 30227 7723
rect 32112 7790 32533 7824
rect 32112 7645 32175 7790
rect 32484 7645 32533 7790
rect 32112 7624 32533 7645
rect 27918 7527 28071 7596
rect 33520 7323 33764 7361
rect 33520 7253 33576 7323
rect 33712 7253 33764 7323
rect 33520 7231 33764 7253
rect 4475 6041 4628 6081
rect 4475 5892 4518 6041
rect 4585 5892 4628 6041
rect 11026 6039 11179 6079
rect 4475 5823 4628 5892
rect 11026 5890 11069 6039
rect 11136 5890 11179 6039
rect 17681 6040 17834 6080
rect 11026 5821 11179 5890
rect 17681 5891 17724 6040
rect 17791 5891 17834 6040
rect 24303 6041 24456 6081
rect 17681 5822 17834 5891
rect 24303 5892 24346 6041
rect 24413 5892 24456 6041
rect 24303 5823 24456 5892
rect 8186 5698 8339 5738
rect 8186 5549 8229 5698
rect 8296 5549 8339 5698
rect 14737 5696 14890 5736
rect 8186 5480 8339 5549
rect -4119 5128 -3975 5252
rect -4119 5006 -4067 5128
rect -4023 5006 -3975 5128
rect 14737 5547 14780 5696
rect 14847 5547 14890 5696
rect 21392 5697 21545 5737
rect 14737 5478 14890 5547
rect 21392 5548 21435 5697
rect 21502 5548 21545 5697
rect 28014 5698 28167 5738
rect 21392 5479 21545 5548
rect 28014 5549 28057 5698
rect 28124 5549 28167 5698
rect 28014 5480 28167 5549
rect -4119 4852 -3975 5006
rect 1386 4941 1630 4979
rect 1386 4871 1442 4941
rect 1578 4871 1630 4941
rect 1386 4849 1630 4871
rect 4470 4437 4623 4477
rect 4470 4288 4513 4437
rect 4580 4288 4623 4437
rect 4470 4219 4623 4288
rect 11021 4435 11174 4475
rect 11021 4286 11064 4435
rect 11131 4286 11174 4435
rect 11021 4217 11174 4286
rect -4117 3059 -3973 3183
rect -4117 2937 -4065 3059
rect -4021 2937 -3973 3059
rect 17676 4436 17829 4476
rect 17676 4287 17719 4436
rect 17786 4287 17829 4436
rect 17676 4218 17829 4287
rect 36437 5064 36583 5118
rect 36437 4868 36493 5064
rect 36569 4868 36583 5064
rect 24298 4437 24451 4477
rect 24298 4288 24341 4437
rect 24408 4288 24451 4437
rect 24298 4219 24451 4288
rect -4117 2783 -3973 2937
rect 36437 4814 36583 4868
rect 29980 4723 30224 4761
rect 29980 4653 30036 4723
rect 30172 4653 30224 4723
rect 29980 4631 30224 4653
rect 32112 3442 32533 3476
rect 32112 3297 32175 3442
rect 32484 3297 32533 3442
rect 32112 3276 32533 3297
rect 33520 2975 33764 3013
rect 33520 2905 33576 2975
rect 33712 2905 33764 2975
rect 33520 2883 33764 2905
rect 29987 1878 30231 1916
rect 29987 1808 30043 1878
rect 30179 1808 30231 1878
rect 29987 1786 30231 1808
rect 36437 1920 36583 1974
rect 36437 1724 36493 1920
rect 36569 1724 36583 1920
rect 36437 1670 36583 1724
rect -4119 991 -3975 1115
rect -4119 869 -4067 991
rect -4023 869 -3975 991
rect 8096 1174 8340 1196
rect 8096 1104 8152 1174
rect 8288 1104 8340 1174
rect 8096 1066 8340 1104
rect 14650 1179 14894 1201
rect 14650 1109 14706 1179
rect 14842 1109 14894 1179
rect 14650 1071 14894 1109
rect 21299 1167 21543 1189
rect 21299 1097 21355 1167
rect 21491 1097 21543 1167
rect 21299 1059 21543 1097
rect -4119 715 -3975 869
<< psubdiffcont >>
rect 6649 26755 6812 26845
rect 13162 26752 13325 26842
rect 19696 26747 19859 26837
rect 26254 26751 26417 26841
rect 8131 26311 8221 26474
rect 9273 26309 9363 26472
rect 14644 26308 14734 26471
rect 15786 26306 15876 26469
rect 21178 26303 21268 26466
rect 22320 26301 22410 26464
rect 27736 26307 27826 26470
rect 28878 26305 28968 26468
rect 6663 25105 6826 25195
rect 13176 25102 13339 25192
rect 19710 25097 19873 25187
rect 6658 23501 6821 23591
rect 26268 25101 26431 25191
rect 13171 23498 13334 23588
rect 8075 23268 8165 23431
rect 19705 23493 19868 23583
rect 14588 23265 14678 23428
rect 26263 23497 26426 23587
rect 21122 23260 21212 23423
rect 27680 23264 27770 23427
rect 38743 23800 38789 23904
rect 9092 21147 9255 21237
rect 15650 21143 15813 21233
rect 22184 21148 22347 21238
rect 28697 21151 28860 21241
rect 6541 20701 6631 20864
rect 7683 20703 7773 20866
rect 13099 20697 13189 20860
rect 14241 20699 14331 20862
rect 19633 20702 19723 20865
rect 20775 20704 20865 20867
rect 26146 20705 26236 20868
rect 27288 20707 27378 20870
rect 9078 19497 9241 19587
rect 15636 19493 15799 19583
rect 9083 17893 9246 17983
rect 22170 19498 22333 19588
rect 38743 20656 38789 20760
rect 15641 17889 15804 17979
rect 28683 19501 28846 19591
rect 7739 17660 7829 17823
rect 22175 17894 22338 17984
rect 14297 17656 14387 17819
rect 28688 17897 28851 17987
rect 20831 17661 20921 17824
rect 27344 17664 27434 17827
rect 38739 17524 38785 17628
rect -1803 15388 -1747 15520
rect 8341 14200 8475 14256
rect 14890 14199 15024 14255
rect 21544 14220 21678 14276
rect 30197 14053 30331 14109
rect -1805 13320 -1749 13452
rect 38739 14380 38785 14484
rect 33798 13645 33932 13701
rect 1677 12300 1811 12356
rect 4845 12204 5008 12294
rect 11394 12292 11557 12382
rect 18048 12224 18211 12314
rect 32215 12798 32350 12900
rect 24673 12292 24836 12382
rect 6327 11760 6417 11923
rect 7469 11758 7559 11921
rect 12876 11848 12966 12011
rect 14018 11846 14108 12009
rect 19530 11780 19620 11943
rect 20672 11778 20762 11941
rect 26155 11848 26245 12011
rect 27297 11846 27387 12009
rect -1803 11251 -1747 11383
rect 30192 11482 30326 11538
rect 4859 10554 5022 10644
rect 1669 9715 1803 9771
rect 11408 10642 11571 10732
rect -1805 9183 -1749 9315
rect 18062 10574 18225 10664
rect 24687 10642 24850 10732
rect 4854 8950 5017 9040
rect 11403 9038 11566 9128
rect 38743 11178 38789 11282
rect 33800 9554 33934 9610
rect 6271 8717 6361 8880
rect 12820 8805 12910 8968
rect 18057 8970 18220 9060
rect 24682 9038 24845 9128
rect 19474 8737 19564 8900
rect 26099 8805 26189 8968
rect 32217 8707 32352 8809
rect 30192 8449 30326 8505
rect -1805 7114 -1749 7246
rect 1650 6437 1784 6493
rect 4837 6424 5000 6514
rect 38743 8034 38789 8138
rect 11388 6422 11551 6512
rect 18043 6423 18206 6513
rect 24665 6424 24828 6514
rect 30263 6529 30397 6585
rect 6319 5980 6409 6143
rect 7461 5978 7551 6141
rect 12870 5978 12960 6141
rect 14012 5976 14102 6139
rect 19525 5979 19615 6142
rect 20667 5977 20757 6140
rect 26147 5980 26237 6143
rect 27289 5978 27379 6141
rect 33800 6059 33934 6115
rect -1807 5046 -1751 5178
rect 4851 4774 5014 4864
rect 1666 3677 1800 3733
rect 11402 4772 11565 4862
rect 18057 4773 18220 4863
rect 4846 3170 5009 3260
rect 24679 4774 24842 4864
rect 32217 5212 32352 5314
rect -1805 2977 -1749 3109
rect 11397 3168 11560 3258
rect 38739 4902 38785 5006
rect 6263 2937 6353 3100
rect 18052 3169 18215 3259
rect 30260 3459 30394 3515
rect 12814 2935 12904 3098
rect 24674 3170 24837 3260
rect 19469 2936 19559 3099
rect 26091 2937 26181 3100
rect 8376 2312 8510 2368
rect 14930 2317 15064 2373
rect 21579 2305 21713 2361
rect 33800 1711 33934 1767
rect -1807 909 -1751 1041
rect 38739 1758 38785 1862
rect 32217 864 32352 966
rect 30267 614 30401 670
<< nsubdiffcont >>
rect 6316 27873 6383 28022
rect 8798 27927 8865 28076
rect 9945 27927 10012 28076
rect 12829 27870 12896 28019
rect 15311 27924 15378 28073
rect 16458 27924 16525 28073
rect 19363 27865 19430 28014
rect 21845 27919 21912 28068
rect 22992 27919 23059 28068
rect 25921 27869 25988 28018
rect 28403 27923 28470 28072
rect 29550 27923 29617 28072
rect 6330 26223 6397 26372
rect 12843 26220 12910 26369
rect 19377 26215 19444 26364
rect 25935 26219 26002 26368
rect 10041 25880 10108 26029
rect 16554 25877 16621 26026
rect 23088 25872 23155 26021
rect 29646 25876 29713 26025
rect 6325 24619 6392 24768
rect 12838 24616 12905 24765
rect 19372 24611 19439 24760
rect 25930 24615 25997 24764
rect 36497 23766 36573 23962
rect 5892 22319 5959 22468
rect 7039 22319 7106 22468
rect 9521 22265 9588 22414
rect 12450 22315 12517 22464
rect 13597 22315 13664 22464
rect 16079 22261 16146 22410
rect 18984 22320 19051 22469
rect 20131 22320 20198 22469
rect 22613 22266 22680 22415
rect 25497 22323 25564 22472
rect 26644 22323 26711 22472
rect 29126 22269 29193 22418
rect 9507 20615 9574 20764
rect 16065 20611 16132 20760
rect 22599 20616 22666 20765
rect 29112 20619 29179 20768
rect 36497 20622 36573 20818
rect 5796 20272 5863 20421
rect 12354 20268 12421 20417
rect 18888 20273 18955 20422
rect 25401 20276 25468 20425
rect 9512 19011 9579 19160
rect 16070 19007 16137 19156
rect 22604 19012 22671 19161
rect 29117 19015 29184 19164
rect 36493 17490 36569 17686
rect -4063 15348 -4019 15470
rect 8117 15394 8253 15464
rect 14666 15393 14802 15463
rect 21320 15414 21456 15484
rect 29973 15247 30109 15317
rect 32173 15231 32482 15376
rect 33574 14839 33710 14909
rect -4065 13280 -4021 13402
rect 1453 13494 1589 13564
rect 4512 13322 4579 13471
rect 6994 13376 7061 13525
rect 8141 13376 8208 13525
rect 11061 13410 11128 13559
rect 13543 13464 13610 13613
rect 14690 13464 14757 13613
rect 17715 13342 17782 13491
rect 20197 13396 20264 13545
rect 21344 13396 21411 13545
rect 24340 13410 24407 13559
rect 26822 13464 26889 13613
rect 27969 13464 28036 13613
rect 36493 14346 36569 14542
rect 29968 12676 30104 12746
rect 4526 11672 4593 11821
rect 11075 11760 11142 11909
rect 17729 11692 17796 11841
rect 24354 11760 24421 11909
rect -4063 11211 -4019 11333
rect 8237 11329 8304 11478
rect 14786 11417 14853 11566
rect 21440 11349 21507 11498
rect 28065 11417 28132 11566
rect 1445 10909 1581 10979
rect 4521 10068 4588 10217
rect -4065 9143 -4021 9265
rect 32175 11140 32484 11285
rect 36497 11144 36573 11340
rect 11070 10156 11137 10305
rect 17724 10088 17791 10237
rect 24349 10156 24416 10305
rect 33576 10748 33712 10818
rect 29968 9643 30104 9713
rect 36497 8000 36573 8196
rect 1426 7631 1562 7701
rect 4504 7542 4571 7691
rect 6986 7596 7053 7745
rect 8133 7596 8200 7745
rect 11055 7540 11122 7689
rect -4065 7074 -4021 7196
rect 13537 7594 13604 7743
rect 14684 7594 14751 7743
rect 17710 7541 17777 7690
rect 20192 7595 20259 7744
rect 21339 7595 21406 7744
rect 24332 7542 24399 7691
rect 26814 7596 26881 7745
rect 27961 7596 28028 7745
rect 30039 7723 30175 7793
rect 32175 7645 32484 7790
rect 33576 7253 33712 7323
rect 4518 5892 4585 6041
rect 11069 5890 11136 6039
rect 17724 5891 17791 6040
rect 24346 5892 24413 6041
rect 8229 5549 8296 5698
rect -4067 5006 -4023 5128
rect 14780 5547 14847 5696
rect 21435 5548 21502 5697
rect 28057 5549 28124 5698
rect 1442 4871 1578 4941
rect 4513 4288 4580 4437
rect 11064 4286 11131 4435
rect -4065 2937 -4021 3059
rect 17719 4287 17786 4436
rect 36493 4868 36569 5064
rect 24341 4288 24408 4437
rect 30036 4653 30172 4723
rect 32175 3297 32484 3442
rect 33576 2905 33712 2975
rect 30043 1808 30179 1878
rect 36493 1724 36569 1920
rect -4067 869 -4023 991
rect 8152 1104 8288 1174
rect 14706 1109 14842 1179
rect 21355 1097 21491 1167
<< poly >>
rect 8036 27856 8102 27872
rect 9166 27862 9232 27878
rect 8036 27822 8052 27856
rect 8086 27849 8102 27856
rect 8086 27822 8611 27849
rect 8036 27806 8611 27822
rect 9166 27828 9182 27862
rect 9216 27853 9232 27862
rect 9216 27828 9753 27853
rect 9166 27810 9753 27828
rect 8567 27754 8611 27806
rect 9709 27758 9753 27810
rect 14549 27853 14615 27869
rect 15679 27859 15745 27875
rect 14549 27819 14565 27853
rect 14599 27846 14615 27853
rect 14599 27819 15124 27846
rect 14549 27803 15124 27819
rect 15679 27825 15695 27859
rect 15729 27850 15745 27859
rect 15729 27825 16266 27850
rect 15679 27807 16266 27825
rect 8036 27738 8509 27754
rect 8036 27704 8052 27738
rect 8086 27713 8509 27738
rect 8086 27712 8273 27713
rect 8086 27704 8102 27712
rect 8036 27688 8102 27704
rect 8213 27692 8273 27712
rect 8331 27692 8391 27713
rect 8449 27692 8509 27713
rect 8567 27713 8863 27754
rect 8567 27692 8627 27713
rect 8685 27692 8745 27713
rect 8803 27692 8863 27713
rect 9166 27742 9651 27758
rect 9166 27708 9182 27742
rect 9216 27717 9651 27742
rect 9216 27716 9415 27717
rect 9216 27708 9232 27716
rect 9166 27692 9232 27708
rect 9355 27696 9415 27716
rect 9473 27696 9533 27717
rect 9591 27696 9651 27717
rect 9709 27717 10005 27758
rect 15080 27751 15124 27803
rect 16222 27755 16266 27807
rect 21083 27848 21149 27864
rect 22213 27854 22279 27870
rect 21083 27814 21099 27848
rect 21133 27841 21149 27848
rect 21133 27814 21658 27841
rect 21083 27798 21658 27814
rect 22213 27820 22229 27854
rect 22263 27845 22279 27854
rect 22263 27820 22800 27845
rect 22213 27802 22800 27820
rect 9709 27696 9769 27717
rect 9827 27696 9887 27717
rect 9945 27696 10005 27717
rect 14549 27735 15022 27751
rect 14549 27701 14565 27735
rect 14599 27710 15022 27735
rect 14599 27709 14786 27710
rect 14599 27701 14615 27709
rect 5888 27641 6184 27677
rect 5888 27620 5948 27641
rect 6006 27620 6066 27641
rect 6124 27620 6184 27641
rect 6242 27640 6538 27676
rect 6242 27620 6302 27640
rect 6360 27620 6420 27640
rect 6478 27620 6538 27640
rect 6596 27640 6892 27676
rect 6596 27620 6656 27640
rect 6714 27620 6774 27640
rect 6832 27620 6892 27640
rect 5888 27394 5948 27420
rect 6006 27394 6066 27420
rect 6124 27394 6184 27420
rect 6242 27400 6302 27420
rect 6242 27394 6303 27400
rect 6360 27394 6420 27420
rect 6478 27394 6538 27420
rect 6125 27209 6183 27394
rect 6125 27183 6185 27209
rect 6243 27183 6303 27394
rect 6596 27388 6656 27420
rect 6714 27394 6774 27420
rect 6832 27394 6892 27420
rect 6593 27372 6659 27388
rect 6593 27338 6609 27372
rect 6643 27338 6659 27372
rect 6593 27322 6659 27338
rect 14549 27685 14615 27701
rect 14726 27689 14786 27709
rect 14844 27689 14904 27710
rect 14962 27689 15022 27710
rect 15080 27710 15376 27751
rect 15080 27689 15140 27710
rect 15198 27689 15258 27710
rect 15316 27689 15376 27710
rect 15679 27739 16164 27755
rect 15679 27705 15695 27739
rect 15729 27714 16164 27739
rect 15729 27713 15928 27714
rect 15729 27705 15745 27713
rect 15679 27689 15745 27705
rect 15868 27693 15928 27713
rect 15986 27693 16046 27714
rect 16104 27693 16164 27714
rect 16222 27714 16518 27755
rect 21614 27746 21658 27798
rect 22756 27750 22800 27802
rect 27641 27852 27707 27868
rect 28771 27858 28837 27874
rect 27641 27818 27657 27852
rect 27691 27845 27707 27852
rect 27691 27818 28216 27845
rect 27641 27802 28216 27818
rect 28771 27824 28787 27858
rect 28821 27849 28837 27858
rect 28821 27824 29358 27849
rect 28771 27806 29358 27824
rect 28172 27750 28216 27802
rect 29314 27754 29358 27806
rect 16222 27693 16282 27714
rect 16340 27693 16400 27714
rect 16458 27693 16518 27714
rect 21083 27730 21556 27746
rect 21083 27696 21099 27730
rect 21133 27705 21556 27730
rect 21133 27704 21320 27705
rect 21133 27696 21149 27704
rect 12401 27638 12697 27674
rect 12401 27617 12461 27638
rect 12519 27617 12579 27638
rect 12637 27617 12697 27638
rect 12755 27637 13051 27673
rect 12755 27617 12815 27637
rect 12873 27617 12933 27637
rect 12991 27617 13051 27637
rect 13109 27637 13405 27673
rect 13109 27617 13169 27637
rect 13227 27617 13287 27637
rect 13345 27617 13405 27637
rect 12401 27391 12461 27417
rect 12519 27391 12579 27417
rect 12637 27391 12697 27417
rect 12755 27397 12815 27417
rect 12755 27391 12816 27397
rect 12873 27391 12933 27417
rect 12991 27391 13051 27417
rect 8213 27275 8273 27292
rect 6475 27255 6541 27271
rect 6475 27221 6491 27255
rect 6525 27221 6541 27255
rect 6475 27205 6541 27221
rect 6478 27183 6538 27205
rect 8213 27186 8274 27275
rect 8331 27266 8391 27292
rect 8449 27266 8509 27292
rect 8123 27133 8274 27186
rect 6478 26957 6538 26983
rect 8123 26909 8183 27133
rect 8567 27091 8627 27292
rect 8685 27266 8745 27292
rect 8803 27266 8863 27292
rect 9355 27279 9415 27296
rect 9355 27190 9416 27279
rect 9473 27270 9533 27296
rect 9591 27270 9651 27296
rect 8241 27040 8627 27091
rect 9265 27137 9416 27190
rect 8241 26909 8301 27040
rect 8356 26982 8422 26998
rect 8356 26948 8372 26982
rect 8406 26948 8422 26982
rect 8356 26932 8422 26948
rect 8359 26909 8419 26932
rect 8642 26909 8702 26935
rect 8760 26909 8820 26935
rect 8878 26909 8938 26935
rect 9265 26913 9325 27137
rect 9709 27095 9769 27296
rect 9827 27270 9887 27296
rect 9945 27270 10005 27296
rect 12638 27206 12696 27391
rect 12638 27180 12698 27206
rect 12756 27180 12816 27391
rect 13109 27385 13169 27417
rect 13227 27391 13287 27417
rect 13345 27391 13405 27417
rect 13106 27369 13172 27385
rect 13106 27335 13122 27369
rect 13156 27335 13172 27369
rect 13106 27319 13172 27335
rect 21083 27680 21149 27696
rect 21260 27684 21320 27704
rect 21378 27684 21438 27705
rect 21496 27684 21556 27705
rect 21614 27705 21910 27746
rect 21614 27684 21674 27705
rect 21732 27684 21792 27705
rect 21850 27684 21910 27705
rect 22213 27734 22698 27750
rect 22213 27700 22229 27734
rect 22263 27709 22698 27734
rect 22263 27708 22462 27709
rect 22263 27700 22279 27708
rect 22213 27684 22279 27700
rect 22402 27688 22462 27708
rect 22520 27688 22580 27709
rect 22638 27688 22698 27709
rect 22756 27709 23052 27750
rect 22756 27688 22816 27709
rect 22874 27688 22934 27709
rect 22992 27688 23052 27709
rect 27641 27734 28114 27750
rect 27641 27700 27657 27734
rect 27691 27709 28114 27734
rect 27691 27708 27878 27709
rect 27691 27700 27707 27708
rect 18935 27633 19231 27669
rect 18935 27612 18995 27633
rect 19053 27612 19113 27633
rect 19171 27612 19231 27633
rect 19289 27632 19585 27668
rect 19289 27612 19349 27632
rect 19407 27612 19467 27632
rect 19525 27612 19585 27632
rect 19643 27632 19939 27668
rect 19643 27612 19703 27632
rect 19761 27612 19821 27632
rect 19879 27612 19939 27632
rect 18935 27386 18995 27412
rect 19053 27386 19113 27412
rect 19171 27386 19231 27412
rect 19289 27392 19349 27412
rect 19289 27386 19350 27392
rect 19407 27386 19467 27412
rect 19525 27386 19585 27412
rect 14726 27272 14786 27289
rect 12988 27252 13054 27268
rect 12988 27218 13004 27252
rect 13038 27218 13054 27252
rect 12988 27202 13054 27218
rect 12991 27180 13051 27202
rect 14726 27183 14787 27272
rect 14844 27263 14904 27289
rect 14962 27263 15022 27289
rect 9383 27044 9769 27095
rect 9383 26913 9443 27044
rect 9498 26986 9564 27002
rect 9498 26952 9514 26986
rect 9548 26952 9564 26986
rect 9498 26936 9564 26952
rect 9501 26913 9561 26936
rect 9784 26913 9844 26939
rect 9902 26913 9962 26939
rect 10020 26913 10080 26939
rect 6125 26761 6185 26783
rect 6243 26761 6303 26783
rect 6122 26745 6188 26761
rect 6122 26711 6138 26745
rect 6172 26711 6188 26745
rect 6122 26695 6188 26711
rect 6240 26745 6306 26761
rect 6240 26711 6256 26745
rect 6290 26711 6306 26745
rect 6240 26695 6306 26711
rect 14636 27130 14787 27183
rect 12991 26954 13051 26980
rect 14636 26906 14696 27130
rect 15080 27088 15140 27289
rect 15198 27263 15258 27289
rect 15316 27263 15376 27289
rect 15868 27276 15928 27293
rect 15868 27187 15929 27276
rect 15986 27267 16046 27293
rect 16104 27267 16164 27293
rect 14754 27037 15140 27088
rect 15778 27134 15929 27187
rect 14754 26906 14814 27037
rect 14869 26979 14935 26995
rect 14869 26945 14885 26979
rect 14919 26945 14935 26979
rect 14869 26929 14935 26945
rect 14872 26906 14932 26929
rect 15155 26906 15215 26932
rect 15273 26906 15333 26932
rect 15391 26906 15451 26932
rect 15778 26910 15838 27134
rect 16222 27092 16282 27293
rect 16340 27267 16400 27293
rect 16458 27267 16518 27293
rect 19172 27201 19230 27386
rect 19172 27175 19232 27201
rect 19290 27175 19350 27386
rect 19643 27380 19703 27412
rect 19761 27386 19821 27412
rect 19879 27386 19939 27412
rect 19640 27364 19706 27380
rect 19640 27330 19656 27364
rect 19690 27330 19706 27364
rect 19640 27314 19706 27330
rect 27641 27684 27707 27700
rect 27818 27688 27878 27708
rect 27936 27688 27996 27709
rect 28054 27688 28114 27709
rect 28172 27709 28468 27750
rect 28172 27688 28232 27709
rect 28290 27688 28350 27709
rect 28408 27688 28468 27709
rect 28771 27738 29256 27754
rect 28771 27704 28787 27738
rect 28821 27713 29256 27738
rect 28821 27712 29020 27713
rect 28821 27704 28837 27712
rect 28771 27688 28837 27704
rect 28960 27692 29020 27712
rect 29078 27692 29138 27713
rect 29196 27692 29256 27713
rect 29314 27713 29610 27754
rect 29314 27692 29374 27713
rect 29432 27692 29492 27713
rect 29550 27692 29610 27713
rect 25493 27637 25789 27673
rect 25493 27616 25553 27637
rect 25611 27616 25671 27637
rect 25729 27616 25789 27637
rect 25847 27636 26143 27672
rect 25847 27616 25907 27636
rect 25965 27616 26025 27636
rect 26083 27616 26143 27636
rect 26201 27636 26497 27672
rect 26201 27616 26261 27636
rect 26319 27616 26379 27636
rect 26437 27616 26497 27636
rect 25493 27390 25553 27416
rect 25611 27390 25671 27416
rect 25729 27390 25789 27416
rect 25847 27396 25907 27416
rect 25847 27390 25908 27396
rect 25965 27390 26025 27416
rect 26083 27390 26143 27416
rect 21260 27267 21320 27284
rect 19522 27247 19588 27263
rect 19522 27213 19538 27247
rect 19572 27213 19588 27247
rect 19522 27197 19588 27213
rect 19525 27175 19585 27197
rect 21260 27178 21321 27267
rect 21378 27258 21438 27284
rect 21496 27258 21556 27284
rect 15896 27041 16282 27092
rect 15896 26910 15956 27041
rect 16011 26983 16077 26999
rect 16011 26949 16027 26983
rect 16061 26949 16077 26983
rect 16011 26933 16077 26949
rect 16014 26910 16074 26933
rect 16297 26910 16357 26936
rect 16415 26910 16475 26936
rect 16533 26910 16593 26936
rect 12638 26758 12698 26780
rect 12756 26758 12816 26780
rect 12635 26742 12701 26758
rect 8123 26683 8183 26709
rect 8241 26683 8301 26709
rect 8359 26677 8419 26709
rect 8642 26677 8702 26709
rect 8760 26677 8820 26709
rect 8878 26677 8938 26709
rect 9265 26687 9325 26713
rect 9383 26687 9443 26713
rect 8359 26636 8938 26677
rect 9501 26681 9561 26713
rect 9784 26681 9844 26713
rect 9902 26681 9962 26713
rect 10020 26681 10080 26713
rect 12635 26708 12651 26742
rect 12685 26708 12701 26742
rect 12635 26692 12701 26708
rect 12753 26742 12819 26758
rect 12753 26708 12769 26742
rect 12803 26708 12819 26742
rect 12753 26692 12819 26708
rect 21170 27125 21321 27178
rect 19525 26949 19585 26975
rect 21170 26901 21230 27125
rect 21614 27083 21674 27284
rect 21732 27258 21792 27284
rect 21850 27258 21910 27284
rect 22402 27271 22462 27288
rect 22402 27182 22463 27271
rect 22520 27262 22580 27288
rect 22638 27262 22698 27288
rect 21288 27032 21674 27083
rect 22312 27129 22463 27182
rect 21288 26901 21348 27032
rect 21403 26974 21469 26990
rect 21403 26940 21419 26974
rect 21453 26940 21469 26974
rect 21403 26924 21469 26940
rect 21406 26901 21466 26924
rect 21689 26901 21749 26927
rect 21807 26901 21867 26927
rect 21925 26901 21985 26927
rect 22312 26905 22372 27129
rect 22756 27087 22816 27288
rect 22874 27262 22934 27288
rect 22992 27262 23052 27288
rect 25730 27205 25788 27390
rect 25730 27179 25790 27205
rect 25848 27179 25908 27390
rect 26201 27384 26261 27416
rect 26319 27390 26379 27416
rect 26437 27390 26497 27416
rect 26198 27368 26264 27384
rect 26198 27334 26214 27368
rect 26248 27334 26264 27368
rect 26198 27318 26264 27334
rect 27818 27271 27878 27288
rect 26080 27251 26146 27267
rect 26080 27217 26096 27251
rect 26130 27217 26146 27251
rect 26080 27201 26146 27217
rect 26083 27179 26143 27201
rect 27818 27182 27879 27271
rect 27936 27262 27996 27288
rect 28054 27262 28114 27288
rect 22430 27036 22816 27087
rect 22430 26905 22490 27036
rect 22545 26978 22611 26994
rect 22545 26944 22561 26978
rect 22595 26944 22611 26978
rect 22545 26928 22611 26944
rect 22548 26905 22608 26928
rect 22831 26905 22891 26931
rect 22949 26905 23009 26931
rect 23067 26905 23127 26931
rect 19172 26753 19232 26775
rect 19290 26753 19350 26775
rect 19169 26737 19235 26753
rect 9501 26640 10080 26681
rect 14636 26680 14696 26706
rect 14754 26680 14814 26706
rect 14872 26674 14932 26706
rect 15155 26674 15215 26706
rect 15273 26674 15333 26706
rect 15391 26674 15451 26706
rect 15778 26684 15838 26710
rect 15896 26684 15956 26710
rect 14872 26633 15451 26674
rect 16014 26678 16074 26710
rect 16297 26678 16357 26710
rect 16415 26678 16475 26710
rect 16533 26678 16593 26710
rect 19169 26703 19185 26737
rect 19219 26703 19235 26737
rect 19169 26687 19235 26703
rect 19287 26737 19353 26753
rect 19287 26703 19303 26737
rect 19337 26703 19353 26737
rect 19287 26687 19353 26703
rect 27728 27129 27879 27182
rect 26083 26953 26143 26979
rect 27728 26905 27788 27129
rect 28172 27087 28232 27288
rect 28290 27262 28350 27288
rect 28408 27262 28468 27288
rect 28960 27275 29020 27292
rect 28960 27186 29021 27275
rect 29078 27266 29138 27292
rect 29196 27266 29256 27292
rect 27846 27036 28232 27087
rect 28870 27133 29021 27186
rect 27846 26905 27906 27036
rect 27961 26978 28027 26994
rect 27961 26944 27977 26978
rect 28011 26944 28027 26978
rect 27961 26928 28027 26944
rect 27964 26905 28024 26928
rect 28247 26905 28307 26931
rect 28365 26905 28425 26931
rect 28483 26905 28543 26931
rect 28870 26909 28930 27133
rect 29314 27091 29374 27292
rect 29432 27266 29492 27292
rect 29550 27266 29610 27292
rect 28988 27040 29374 27091
rect 28988 26909 29048 27040
rect 29103 26982 29169 26998
rect 29103 26948 29119 26982
rect 29153 26948 29169 26982
rect 29103 26932 29169 26948
rect 29106 26909 29166 26932
rect 29389 26909 29449 26935
rect 29507 26909 29567 26935
rect 29625 26909 29685 26935
rect 25730 26757 25790 26779
rect 25848 26757 25908 26779
rect 25727 26741 25793 26757
rect 25727 26707 25743 26741
rect 25777 26707 25793 26741
rect 16014 26637 16593 26678
rect 21170 26675 21230 26701
rect 21288 26675 21348 26701
rect 21406 26669 21466 26701
rect 21689 26669 21749 26701
rect 21807 26669 21867 26701
rect 21925 26669 21985 26701
rect 22312 26679 22372 26705
rect 22430 26679 22490 26705
rect 21406 26628 21985 26669
rect 22548 26673 22608 26705
rect 22831 26673 22891 26705
rect 22949 26673 23009 26705
rect 23067 26673 23127 26705
rect 25727 26691 25793 26707
rect 25845 26741 25911 26757
rect 25845 26707 25861 26741
rect 25895 26707 25911 26741
rect 25845 26691 25911 26707
rect 27728 26679 27788 26705
rect 27846 26679 27906 26705
rect 22548 26632 23127 26673
rect 27964 26673 28024 26705
rect 28247 26673 28307 26705
rect 28365 26673 28425 26705
rect 28483 26673 28543 26705
rect 28870 26683 28930 26709
rect 28988 26683 29048 26709
rect 27964 26632 28543 26673
rect 29106 26677 29166 26709
rect 29389 26677 29449 26709
rect 29507 26677 29567 26709
rect 29625 26677 29685 26709
rect 29106 26636 29685 26677
rect 5902 25991 6198 26027
rect 5902 25970 5962 25991
rect 6020 25970 6080 25991
rect 6138 25970 6198 25991
rect 6256 25990 6552 26026
rect 6256 25970 6316 25990
rect 6374 25970 6434 25990
rect 6492 25970 6552 25990
rect 6610 25990 6906 26026
rect 6610 25970 6670 25990
rect 6728 25970 6788 25990
rect 6846 25970 6906 25990
rect 12415 25988 12711 26024
rect 12415 25967 12475 25988
rect 12533 25967 12593 25988
rect 12651 25967 12711 25988
rect 12769 25987 13065 26023
rect 12769 25967 12829 25987
rect 12887 25967 12947 25987
rect 13005 25967 13065 25987
rect 13123 25987 13419 26023
rect 13123 25967 13183 25987
rect 13241 25967 13301 25987
rect 13359 25967 13419 25987
rect 5902 25744 5962 25770
rect 6020 25744 6080 25770
rect 6138 25744 6198 25770
rect 6256 25750 6316 25770
rect 6256 25744 6317 25750
rect 6374 25744 6434 25770
rect 6492 25744 6552 25770
rect 6139 25559 6197 25744
rect 6139 25533 6199 25559
rect 6257 25533 6317 25744
rect 6610 25738 6670 25770
rect 6728 25744 6788 25770
rect 6846 25744 6906 25770
rect 18949 25983 19245 26019
rect 18949 25962 19009 25983
rect 19067 25962 19127 25983
rect 19185 25962 19245 25983
rect 19303 25982 19599 26018
rect 19303 25962 19363 25982
rect 19421 25962 19481 25982
rect 19539 25962 19599 25982
rect 19657 25982 19953 26018
rect 19657 25962 19717 25982
rect 19775 25962 19835 25982
rect 19893 25962 19953 25982
rect 12415 25741 12475 25767
rect 12533 25741 12593 25767
rect 12651 25741 12711 25767
rect 12769 25747 12829 25767
rect 12769 25741 12830 25747
rect 12887 25741 12947 25767
rect 13005 25741 13065 25767
rect 6607 25722 6673 25738
rect 6607 25688 6623 25722
rect 6657 25688 6673 25722
rect 6607 25672 6673 25688
rect 6489 25605 6555 25621
rect 6489 25571 6505 25605
rect 6539 25571 6555 25605
rect 6489 25555 6555 25571
rect 7850 25568 8146 25619
rect 6492 25533 6552 25555
rect 7850 25553 7910 25568
rect 7968 25553 8028 25568
rect 8086 25553 8146 25568
rect 8204 25553 8264 25579
rect 8322 25553 8382 25579
rect 8440 25553 8500 25579
rect 9748 25568 10044 25619
rect 9748 25553 9808 25568
rect 9866 25553 9926 25568
rect 9984 25553 10044 25568
rect 10102 25553 10162 25579
rect 10220 25553 10280 25579
rect 10338 25553 10398 25579
rect 12652 25556 12710 25741
rect 7366 25353 7426 25379
rect 7484 25353 7544 25379
rect 7602 25353 7662 25379
rect 6492 25307 6552 25333
rect 6139 25111 6199 25133
rect 6257 25117 6317 25133
rect 6136 25095 6202 25111
rect 6136 25061 6152 25095
rect 6186 25061 6202 25095
rect 6136 25045 6202 25061
rect 6251 25095 6325 25117
rect 6251 25061 6270 25095
rect 6304 25061 6325 25095
rect 8687 25370 8983 25421
rect 8687 25353 8747 25370
rect 8805 25353 8865 25370
rect 8923 25353 8983 25370
rect 9264 25353 9324 25379
rect 9382 25353 9442 25379
rect 9500 25353 9560 25379
rect 12652 25530 12712 25556
rect 12770 25530 12830 25741
rect 13123 25735 13183 25767
rect 13241 25741 13301 25767
rect 13359 25741 13419 25767
rect 25507 25987 25803 26023
rect 25507 25966 25567 25987
rect 25625 25966 25685 25987
rect 25743 25966 25803 25987
rect 25861 25986 26157 26022
rect 25861 25966 25921 25986
rect 25979 25966 26039 25986
rect 26097 25966 26157 25986
rect 26215 25986 26511 26022
rect 26215 25966 26275 25986
rect 26333 25966 26393 25986
rect 26451 25966 26511 25986
rect 18949 25736 19009 25762
rect 19067 25736 19127 25762
rect 19185 25736 19245 25762
rect 19303 25742 19363 25762
rect 19303 25736 19364 25742
rect 19421 25736 19481 25762
rect 19539 25736 19599 25762
rect 13120 25719 13186 25735
rect 13120 25685 13136 25719
rect 13170 25685 13186 25719
rect 13120 25669 13186 25685
rect 13002 25602 13068 25618
rect 13002 25568 13018 25602
rect 13052 25568 13068 25602
rect 13002 25552 13068 25568
rect 14363 25565 14659 25616
rect 13005 25530 13065 25552
rect 14363 25550 14423 25565
rect 14481 25550 14541 25565
rect 14599 25550 14659 25565
rect 14717 25550 14777 25576
rect 14835 25550 14895 25576
rect 14953 25550 15013 25576
rect 16261 25565 16557 25616
rect 16261 25550 16321 25565
rect 16379 25550 16439 25565
rect 16497 25550 16557 25565
rect 16615 25550 16675 25576
rect 16733 25550 16793 25576
rect 16851 25550 16911 25576
rect 19186 25551 19244 25736
rect 10585 25370 10881 25421
rect 10585 25353 10645 25370
rect 10703 25353 10763 25370
rect 10821 25353 10881 25370
rect 7366 25136 7426 25153
rect 7484 25136 7544 25153
rect 7602 25136 7662 25153
rect 7850 25136 7910 25153
rect 7366 25085 7910 25136
rect 7968 25127 8028 25153
rect 8086 25127 8146 25153
rect 8204 25134 8264 25153
rect 8322 25134 8382 25153
rect 8440 25134 8500 25153
rect 8687 25134 8747 25153
rect 8805 25134 8865 25153
rect 6251 25004 6325 25061
rect 7491 25004 7551 25085
rect 8204 25083 8747 25134
rect 8789 25127 8865 25134
rect 8923 25127 8983 25153
rect 9264 25136 9324 25153
rect 9382 25136 9442 25153
rect 9500 25136 9560 25153
rect 9748 25136 9808 25153
rect 8789 25083 8864 25127
rect 9264 25085 9808 25136
rect 9866 25127 9926 25153
rect 9984 25127 10044 25153
rect 10102 25134 10162 25153
rect 10220 25134 10280 25153
rect 10338 25134 10398 25153
rect 10585 25134 10645 25153
rect 10703 25134 10763 25153
rect 6251 24979 7551 25004
rect 6250 24931 7551 24979
rect 8789 24963 8849 25083
rect 5897 24387 6193 24423
rect 5897 24366 5957 24387
rect 6015 24366 6075 24387
rect 6133 24366 6193 24387
rect 6251 24386 6547 24422
rect 6251 24366 6311 24386
rect 6369 24366 6429 24386
rect 6487 24366 6547 24386
rect 6605 24386 6901 24422
rect 6605 24366 6665 24386
rect 6723 24366 6783 24386
rect 6841 24366 6901 24386
rect 7491 24233 7551 24931
rect 7793 24883 8089 24943
rect 7793 24860 7853 24883
rect 7911 24860 7971 24883
rect 8029 24860 8089 24883
rect 8147 24884 8443 24944
rect 8788 24943 8849 24963
rect 8147 24860 8207 24884
rect 8265 24860 8325 24884
rect 8383 24860 8443 24884
rect 8769 24927 8849 24943
rect 8769 24893 8784 24927
rect 8818 24893 8849 24927
rect 8769 24877 8849 24893
rect 8788 24854 8849 24877
rect 8789 24708 8849 24854
rect 8788 24535 8849 24708
rect 7793 24434 7853 24460
rect 7761 24293 7828 24300
rect 7911 24293 7971 24460
rect 8029 24434 8089 24460
rect 8147 24434 8207 24460
rect 7761 24284 7971 24293
rect 7761 24250 7777 24284
rect 7811 24250 7971 24284
rect 7761 24234 7971 24250
rect 7491 24217 7642 24233
rect 7491 24183 7592 24217
rect 7626 24183 7642 24217
rect 7491 24167 7642 24183
rect 5897 24140 5957 24166
rect 6015 24140 6075 24166
rect 6133 24140 6193 24166
rect 6251 24146 6311 24166
rect 6251 24140 6312 24146
rect 6369 24140 6429 24166
rect 6487 24140 6547 24166
rect 6134 23955 6192 24140
rect 6134 23929 6194 23955
rect 6252 23929 6312 24140
rect 6605 24134 6665 24166
rect 6723 24140 6783 24166
rect 6841 24140 6901 24166
rect 6602 24118 6668 24134
rect 7491 24128 7551 24167
rect 7911 24128 7971 24234
rect 8265 24293 8325 24460
rect 8383 24434 8443 24460
rect 8408 24293 8475 24300
rect 8265 24284 8475 24293
rect 8265 24250 8425 24284
rect 8459 24250 8475 24284
rect 8265 24234 8475 24250
rect 8027 24200 8093 24216
rect 8027 24166 8043 24200
rect 8077 24166 8093 24200
rect 8027 24150 8093 24166
rect 8145 24201 8211 24216
rect 8145 24167 8161 24201
rect 8195 24167 8211 24201
rect 8145 24151 8211 24167
rect 8029 24128 8089 24150
rect 8147 24128 8207 24151
rect 8265 24128 8325 24234
rect 8789 24232 8849 24535
rect 8699 24216 8849 24232
rect 8699 24182 8715 24216
rect 8749 24182 8849 24216
rect 8699 24166 8849 24182
rect 8789 24128 8849 24166
rect 9389 24427 9449 25085
rect 10102 25083 10645 25134
rect 10687 25127 10763 25134
rect 10821 25127 10881 25153
rect 13879 25350 13939 25376
rect 13997 25350 14057 25376
rect 14115 25350 14175 25376
rect 13005 25304 13065 25330
rect 10687 25083 10762 25127
rect 12652 25108 12712 25130
rect 12770 25114 12830 25130
rect 12649 25092 12715 25108
rect 9691 24883 9987 24943
rect 9691 24860 9751 24883
rect 9809 24860 9869 24883
rect 9927 24860 9987 24883
rect 10045 24884 10341 24944
rect 10045 24860 10105 24884
rect 10163 24860 10223 24884
rect 10281 24860 10341 24884
rect 10687 24930 10747 25083
rect 12649 25058 12665 25092
rect 12699 25058 12715 25092
rect 12649 25042 12715 25058
rect 12764 25092 12838 25114
rect 12764 25058 12783 25092
rect 12817 25058 12838 25092
rect 15200 25367 15496 25418
rect 15200 25350 15260 25367
rect 15318 25350 15378 25367
rect 15436 25350 15496 25367
rect 15777 25350 15837 25376
rect 15895 25350 15955 25376
rect 16013 25350 16073 25376
rect 19186 25525 19246 25551
rect 19304 25525 19364 25736
rect 19657 25730 19717 25762
rect 19775 25736 19835 25762
rect 19893 25736 19953 25762
rect 25507 25740 25567 25766
rect 25625 25740 25685 25766
rect 25743 25740 25803 25766
rect 25861 25746 25921 25766
rect 25861 25740 25922 25746
rect 25979 25740 26039 25766
rect 26097 25740 26157 25766
rect 19654 25714 19720 25730
rect 19654 25680 19670 25714
rect 19704 25680 19720 25714
rect 19654 25664 19720 25680
rect 19536 25597 19602 25613
rect 19536 25563 19552 25597
rect 19586 25563 19602 25597
rect 19536 25547 19602 25563
rect 20897 25560 21193 25611
rect 19539 25525 19599 25547
rect 20897 25545 20957 25560
rect 21015 25545 21075 25560
rect 21133 25545 21193 25560
rect 21251 25545 21311 25571
rect 21369 25545 21429 25571
rect 21487 25545 21547 25571
rect 22795 25560 23091 25611
rect 22795 25545 22855 25560
rect 22913 25545 22973 25560
rect 23031 25545 23091 25560
rect 23149 25545 23209 25571
rect 23267 25545 23327 25571
rect 23385 25545 23445 25571
rect 25744 25555 25802 25740
rect 17098 25367 17394 25418
rect 17098 25350 17158 25367
rect 17216 25350 17276 25367
rect 17334 25350 17394 25367
rect 13879 25133 13939 25150
rect 13997 25133 14057 25150
rect 14115 25133 14175 25150
rect 14363 25133 14423 25150
rect 13879 25082 14423 25133
rect 14481 25124 14541 25150
rect 14599 25124 14659 25150
rect 14717 25131 14777 25150
rect 14835 25131 14895 25150
rect 14953 25131 15013 25150
rect 15200 25131 15260 25150
rect 15318 25131 15378 25150
rect 12764 25001 12838 25058
rect 14004 25001 14064 25082
rect 14717 25080 15260 25131
rect 15302 25124 15378 25131
rect 15436 25124 15496 25150
rect 15777 25133 15837 25150
rect 15895 25133 15955 25150
rect 16013 25133 16073 25150
rect 16261 25133 16321 25150
rect 15302 25080 15377 25124
rect 15777 25082 16321 25133
rect 16379 25124 16439 25150
rect 16497 25124 16557 25150
rect 16615 25131 16675 25150
rect 16733 25131 16793 25150
rect 16851 25131 16911 25150
rect 17098 25131 17158 25150
rect 17216 25131 17276 25150
rect 12764 24976 14064 25001
rect 10687 24906 10941 24930
rect 12763 24928 14064 24976
rect 15302 24960 15362 25080
rect 10687 24872 10891 24906
rect 10925 24872 10941 24906
rect 10687 24856 10941 24872
rect 9691 24434 9751 24460
rect 9389 24411 9456 24427
rect 9389 24377 9405 24411
rect 9439 24377 9456 24411
rect 9389 24361 9456 24377
rect 9389 24233 9449 24361
rect 9659 24293 9726 24300
rect 9809 24293 9869 24460
rect 9927 24434 9987 24460
rect 10045 24434 10105 24460
rect 9659 24284 9869 24293
rect 9659 24250 9675 24284
rect 9709 24250 9869 24284
rect 9659 24234 9869 24250
rect 9389 24217 9540 24233
rect 9389 24183 9490 24217
rect 9524 24183 9540 24217
rect 9389 24167 9540 24183
rect 9389 24128 9449 24167
rect 9809 24128 9869 24234
rect 10163 24293 10223 24460
rect 10281 24434 10341 24460
rect 10304 24294 10371 24301
rect 10298 24293 10371 24294
rect 10163 24285 10371 24293
rect 10163 24251 10321 24285
rect 10355 24251 10371 24285
rect 10163 24235 10371 24251
rect 10163 24234 10360 24235
rect 9925 24200 9991 24216
rect 9925 24166 9941 24200
rect 9975 24166 9991 24200
rect 9925 24150 9991 24166
rect 10043 24201 10109 24216
rect 10043 24167 10059 24201
rect 10093 24167 10109 24201
rect 10043 24151 10109 24167
rect 9927 24128 9987 24150
rect 10045 24128 10105 24151
rect 10163 24128 10223 24234
rect 10687 24232 10747 24856
rect 12410 24384 12706 24420
rect 12410 24363 12470 24384
rect 12528 24363 12588 24384
rect 12646 24363 12706 24384
rect 12764 24383 13060 24419
rect 12764 24363 12824 24383
rect 12882 24363 12942 24383
rect 13000 24363 13060 24383
rect 13118 24383 13414 24419
rect 13118 24363 13178 24383
rect 13236 24363 13296 24383
rect 13354 24363 13414 24383
rect 10597 24216 10747 24232
rect 10597 24182 10613 24216
rect 10647 24182 10747 24216
rect 10597 24166 10747 24182
rect 10687 24128 10747 24166
rect 14004 24230 14064 24928
rect 14306 24880 14602 24940
rect 14306 24857 14366 24880
rect 14424 24857 14484 24880
rect 14542 24857 14602 24880
rect 14660 24881 14956 24941
rect 15301 24940 15362 24960
rect 14660 24857 14720 24881
rect 14778 24857 14838 24881
rect 14896 24857 14956 24881
rect 15282 24924 15362 24940
rect 15282 24890 15297 24924
rect 15331 24890 15362 24924
rect 15282 24874 15362 24890
rect 15301 24851 15362 24874
rect 15302 24705 15362 24851
rect 15301 24532 15362 24705
rect 14306 24431 14366 24457
rect 14274 24290 14341 24297
rect 14424 24290 14484 24457
rect 14542 24431 14602 24457
rect 14660 24431 14720 24457
rect 14274 24281 14484 24290
rect 14274 24247 14290 24281
rect 14324 24247 14484 24281
rect 14274 24231 14484 24247
rect 14004 24214 14155 24230
rect 14004 24180 14105 24214
rect 14139 24180 14155 24214
rect 14004 24164 14155 24180
rect 12410 24137 12470 24163
rect 12528 24137 12588 24163
rect 12646 24137 12706 24163
rect 12764 24143 12824 24163
rect 12764 24137 12825 24143
rect 12882 24137 12942 24163
rect 13000 24137 13060 24163
rect 6602 24084 6618 24118
rect 6652 24084 6668 24118
rect 6602 24068 6668 24084
rect 6484 24001 6550 24017
rect 6484 23967 6500 24001
rect 6534 23967 6550 24001
rect 6484 23951 6550 23967
rect 6487 23929 6547 23951
rect 7491 23902 7551 23928
rect 6487 23703 6547 23729
rect 8789 23902 8849 23928
rect 9389 23902 9449 23928
rect 12647 23952 12705 24137
rect 10687 23902 10747 23928
rect 12647 23926 12707 23952
rect 12765 23926 12825 24137
rect 13118 24131 13178 24163
rect 13236 24137 13296 24163
rect 13354 24137 13414 24163
rect 13115 24115 13181 24131
rect 14004 24125 14064 24164
rect 14424 24125 14484 24231
rect 14778 24290 14838 24457
rect 14896 24431 14956 24457
rect 14921 24290 14988 24297
rect 14778 24281 14988 24290
rect 14778 24247 14938 24281
rect 14972 24247 14988 24281
rect 14778 24231 14988 24247
rect 14540 24197 14606 24213
rect 14540 24163 14556 24197
rect 14590 24163 14606 24197
rect 14540 24147 14606 24163
rect 14658 24198 14724 24213
rect 14658 24164 14674 24198
rect 14708 24164 14724 24198
rect 14658 24148 14724 24164
rect 14542 24125 14602 24147
rect 14660 24125 14720 24148
rect 14778 24125 14838 24231
rect 15302 24229 15362 24532
rect 15212 24213 15362 24229
rect 15212 24179 15228 24213
rect 15262 24179 15362 24213
rect 15212 24163 15362 24179
rect 15302 24125 15362 24163
rect 15902 24424 15962 25082
rect 16615 25080 17158 25131
rect 17200 25124 17276 25131
rect 17334 25124 17394 25150
rect 20413 25345 20473 25371
rect 20531 25345 20591 25371
rect 20649 25345 20709 25371
rect 19539 25299 19599 25325
rect 17200 25080 17275 25124
rect 19186 25103 19246 25125
rect 19304 25109 19364 25125
rect 19183 25087 19249 25103
rect 16204 24880 16500 24940
rect 16204 24857 16264 24880
rect 16322 24857 16382 24880
rect 16440 24857 16500 24880
rect 16558 24881 16854 24941
rect 16558 24857 16618 24881
rect 16676 24857 16736 24881
rect 16794 24857 16854 24881
rect 17200 24927 17260 25080
rect 19183 25053 19199 25087
rect 19233 25053 19249 25087
rect 19183 25037 19249 25053
rect 19298 25087 19372 25109
rect 19298 25053 19317 25087
rect 19351 25053 19372 25087
rect 21734 25362 22030 25413
rect 21734 25345 21794 25362
rect 21852 25345 21912 25362
rect 21970 25345 22030 25362
rect 22311 25345 22371 25371
rect 22429 25345 22489 25371
rect 22547 25345 22607 25371
rect 25744 25529 25804 25555
rect 25862 25529 25922 25740
rect 26215 25734 26275 25766
rect 26333 25740 26393 25766
rect 26451 25740 26511 25766
rect 26212 25718 26278 25734
rect 26212 25684 26228 25718
rect 26262 25684 26278 25718
rect 26212 25668 26278 25684
rect 26094 25601 26160 25617
rect 26094 25567 26110 25601
rect 26144 25567 26160 25601
rect 26094 25551 26160 25567
rect 27455 25564 27751 25615
rect 26097 25529 26157 25551
rect 27455 25549 27515 25564
rect 27573 25549 27633 25564
rect 27691 25549 27751 25564
rect 27809 25549 27869 25575
rect 27927 25549 27987 25575
rect 28045 25549 28105 25575
rect 29353 25564 29649 25615
rect 29353 25549 29413 25564
rect 29471 25549 29531 25564
rect 29589 25549 29649 25564
rect 29707 25549 29767 25575
rect 29825 25549 29885 25575
rect 29943 25549 30003 25575
rect 23632 25362 23928 25413
rect 23632 25345 23692 25362
rect 23750 25345 23810 25362
rect 23868 25345 23928 25362
rect 20413 25128 20473 25145
rect 20531 25128 20591 25145
rect 20649 25128 20709 25145
rect 20897 25128 20957 25145
rect 20413 25077 20957 25128
rect 21015 25119 21075 25145
rect 21133 25119 21193 25145
rect 21251 25126 21311 25145
rect 21369 25126 21429 25145
rect 21487 25126 21547 25145
rect 21734 25126 21794 25145
rect 21852 25126 21912 25145
rect 19298 24996 19372 25053
rect 20538 24996 20598 25077
rect 21251 25075 21794 25126
rect 21836 25119 21912 25126
rect 21970 25119 22030 25145
rect 22311 25128 22371 25145
rect 22429 25128 22489 25145
rect 22547 25128 22607 25145
rect 22795 25128 22855 25145
rect 21836 25075 21911 25119
rect 22311 25077 22855 25128
rect 22913 25119 22973 25145
rect 23031 25119 23091 25145
rect 23149 25126 23209 25145
rect 23267 25126 23327 25145
rect 23385 25126 23445 25145
rect 23632 25126 23692 25145
rect 23750 25126 23810 25145
rect 19298 24971 20598 24996
rect 17200 24903 17454 24927
rect 19297 24923 20598 24971
rect 21836 24955 21896 25075
rect 17200 24869 17404 24903
rect 17438 24869 17454 24903
rect 17200 24853 17454 24869
rect 16204 24431 16264 24457
rect 15902 24408 15969 24424
rect 15902 24374 15918 24408
rect 15952 24374 15969 24408
rect 15902 24358 15969 24374
rect 15902 24230 15962 24358
rect 16172 24290 16239 24297
rect 16322 24290 16382 24457
rect 16440 24431 16500 24457
rect 16558 24431 16618 24457
rect 16172 24281 16382 24290
rect 16172 24247 16188 24281
rect 16222 24247 16382 24281
rect 16172 24231 16382 24247
rect 15902 24214 16053 24230
rect 15902 24180 16003 24214
rect 16037 24180 16053 24214
rect 15902 24164 16053 24180
rect 15902 24125 15962 24164
rect 16322 24125 16382 24231
rect 16676 24290 16736 24457
rect 16794 24431 16854 24457
rect 16817 24291 16884 24298
rect 16811 24290 16884 24291
rect 16676 24282 16884 24290
rect 16676 24248 16834 24282
rect 16868 24248 16884 24282
rect 16676 24232 16884 24248
rect 16676 24231 16873 24232
rect 16438 24197 16504 24213
rect 16438 24163 16454 24197
rect 16488 24163 16504 24197
rect 16438 24147 16504 24163
rect 16556 24198 16622 24213
rect 16556 24164 16572 24198
rect 16606 24164 16622 24198
rect 16556 24148 16622 24164
rect 16440 24125 16500 24147
rect 16558 24125 16618 24148
rect 16676 24125 16736 24231
rect 17200 24229 17260 24853
rect 18944 24379 19240 24415
rect 18944 24358 19004 24379
rect 19062 24358 19122 24379
rect 19180 24358 19240 24379
rect 19298 24378 19594 24414
rect 19298 24358 19358 24378
rect 19416 24358 19476 24378
rect 19534 24358 19594 24378
rect 19652 24378 19948 24414
rect 19652 24358 19712 24378
rect 19770 24358 19830 24378
rect 19888 24358 19948 24378
rect 17110 24213 17260 24229
rect 17110 24179 17126 24213
rect 17160 24179 17260 24213
rect 17110 24163 17260 24179
rect 17200 24125 17260 24163
rect 20538 24225 20598 24923
rect 20840 24875 21136 24935
rect 20840 24852 20900 24875
rect 20958 24852 21018 24875
rect 21076 24852 21136 24875
rect 21194 24876 21490 24936
rect 21835 24935 21896 24955
rect 21194 24852 21254 24876
rect 21312 24852 21372 24876
rect 21430 24852 21490 24876
rect 21816 24919 21896 24935
rect 21816 24885 21831 24919
rect 21865 24885 21896 24919
rect 21816 24869 21896 24885
rect 21835 24846 21896 24869
rect 21836 24700 21896 24846
rect 21835 24527 21896 24700
rect 20840 24426 20900 24452
rect 20808 24285 20875 24292
rect 20958 24285 21018 24452
rect 21076 24426 21136 24452
rect 21194 24426 21254 24452
rect 20808 24276 21018 24285
rect 20808 24242 20824 24276
rect 20858 24242 21018 24276
rect 20808 24226 21018 24242
rect 20538 24209 20689 24225
rect 20538 24175 20639 24209
rect 20673 24175 20689 24209
rect 20538 24159 20689 24175
rect 18944 24132 19004 24158
rect 19062 24132 19122 24158
rect 19180 24132 19240 24158
rect 19298 24138 19358 24158
rect 19298 24132 19359 24138
rect 19416 24132 19476 24158
rect 19534 24132 19594 24158
rect 13115 24081 13131 24115
rect 13165 24081 13181 24115
rect 13115 24065 13181 24081
rect 12997 23998 13063 24014
rect 12997 23964 13013 23998
rect 13047 23964 13063 23998
rect 12997 23948 13063 23964
rect 13000 23926 13060 23948
rect 7911 23702 7971 23728
rect 8029 23702 8089 23728
rect 8147 23702 8207 23728
rect 8265 23702 8325 23728
rect 9809 23702 9869 23728
rect 9927 23702 9987 23728
rect 10045 23702 10105 23728
rect 10163 23702 10223 23728
rect 6134 23507 6194 23529
rect 6252 23507 6312 23529
rect 6131 23491 6197 23507
rect 6131 23457 6147 23491
rect 6181 23457 6197 23491
rect 6131 23441 6197 23457
rect 6249 23491 6315 23507
rect 6249 23457 6265 23491
rect 6299 23457 6315 23491
rect 14004 23899 14064 23925
rect 13000 23700 13060 23726
rect 15302 23899 15362 23925
rect 15902 23899 15962 23925
rect 19181 23947 19239 24132
rect 17200 23899 17260 23925
rect 19181 23921 19241 23947
rect 19299 23921 19359 24132
rect 19652 24126 19712 24158
rect 19770 24132 19830 24158
rect 19888 24132 19948 24158
rect 19649 24110 19715 24126
rect 20538 24120 20598 24159
rect 20958 24120 21018 24226
rect 21312 24285 21372 24452
rect 21430 24426 21490 24452
rect 21455 24285 21522 24292
rect 21312 24276 21522 24285
rect 21312 24242 21472 24276
rect 21506 24242 21522 24276
rect 21312 24226 21522 24242
rect 21074 24192 21140 24208
rect 21074 24158 21090 24192
rect 21124 24158 21140 24192
rect 21074 24142 21140 24158
rect 21192 24193 21258 24208
rect 21192 24159 21208 24193
rect 21242 24159 21258 24193
rect 21192 24143 21258 24159
rect 21076 24120 21136 24142
rect 21194 24120 21254 24143
rect 21312 24120 21372 24226
rect 21836 24224 21896 24527
rect 21746 24208 21896 24224
rect 21746 24174 21762 24208
rect 21796 24174 21896 24208
rect 21746 24158 21896 24174
rect 21836 24120 21896 24158
rect 22436 24419 22496 25077
rect 23149 25075 23692 25126
rect 23734 25119 23810 25126
rect 23868 25119 23928 25145
rect 26971 25349 27031 25375
rect 27089 25349 27149 25375
rect 27207 25349 27267 25375
rect 26097 25303 26157 25329
rect 23734 25075 23809 25119
rect 25744 25107 25804 25129
rect 25862 25113 25922 25129
rect 25741 25091 25807 25107
rect 22738 24875 23034 24935
rect 22738 24852 22798 24875
rect 22856 24852 22916 24875
rect 22974 24852 23034 24875
rect 23092 24876 23388 24936
rect 23092 24852 23152 24876
rect 23210 24852 23270 24876
rect 23328 24852 23388 24876
rect 23734 24922 23794 25075
rect 25741 25057 25757 25091
rect 25791 25057 25807 25091
rect 25741 25041 25807 25057
rect 25856 25091 25930 25113
rect 25856 25057 25875 25091
rect 25909 25057 25930 25091
rect 28292 25366 28588 25417
rect 28292 25349 28352 25366
rect 28410 25349 28470 25366
rect 28528 25349 28588 25366
rect 28869 25349 28929 25375
rect 28987 25349 29047 25375
rect 29105 25349 29165 25375
rect 30190 25366 30486 25417
rect 30190 25349 30250 25366
rect 30308 25349 30368 25366
rect 30426 25349 30486 25366
rect 26971 25132 27031 25149
rect 27089 25132 27149 25149
rect 27207 25132 27267 25149
rect 27455 25132 27515 25149
rect 26971 25081 27515 25132
rect 27573 25123 27633 25149
rect 27691 25123 27751 25149
rect 27809 25130 27869 25149
rect 27927 25130 27987 25149
rect 28045 25130 28105 25149
rect 28292 25130 28352 25149
rect 28410 25130 28470 25149
rect 25856 25000 25930 25057
rect 27096 25000 27156 25081
rect 27809 25079 28352 25130
rect 28394 25123 28470 25130
rect 28528 25123 28588 25149
rect 28869 25132 28929 25149
rect 28987 25132 29047 25149
rect 29105 25132 29165 25149
rect 29353 25132 29413 25149
rect 28394 25079 28469 25123
rect 28869 25081 29413 25132
rect 29471 25123 29531 25149
rect 29589 25123 29649 25149
rect 29707 25130 29767 25149
rect 29825 25130 29885 25149
rect 29943 25130 30003 25149
rect 30190 25130 30250 25149
rect 30308 25130 30368 25149
rect 25856 24975 27156 25000
rect 25855 24927 27156 24975
rect 28394 24959 28454 25079
rect 23734 24898 23988 24922
rect 23734 24864 23938 24898
rect 23972 24864 23988 24898
rect 23734 24848 23988 24864
rect 22738 24426 22798 24452
rect 22436 24403 22503 24419
rect 22436 24369 22452 24403
rect 22486 24369 22503 24403
rect 22436 24353 22503 24369
rect 22436 24225 22496 24353
rect 22706 24285 22773 24292
rect 22856 24285 22916 24452
rect 22974 24426 23034 24452
rect 23092 24426 23152 24452
rect 22706 24276 22916 24285
rect 22706 24242 22722 24276
rect 22756 24242 22916 24276
rect 22706 24226 22916 24242
rect 22436 24209 22587 24225
rect 22436 24175 22537 24209
rect 22571 24175 22587 24209
rect 22436 24159 22587 24175
rect 22436 24120 22496 24159
rect 22856 24120 22916 24226
rect 23210 24285 23270 24452
rect 23328 24426 23388 24452
rect 23351 24286 23418 24293
rect 23345 24285 23418 24286
rect 23210 24277 23418 24285
rect 23210 24243 23368 24277
rect 23402 24243 23418 24277
rect 23210 24227 23418 24243
rect 23210 24226 23407 24227
rect 22972 24192 23038 24208
rect 22972 24158 22988 24192
rect 23022 24158 23038 24192
rect 22972 24142 23038 24158
rect 23090 24193 23156 24208
rect 23090 24159 23106 24193
rect 23140 24159 23156 24193
rect 23090 24143 23156 24159
rect 22974 24120 23034 24142
rect 23092 24120 23152 24143
rect 23210 24120 23270 24226
rect 23734 24224 23794 24848
rect 25502 24383 25798 24419
rect 25502 24362 25562 24383
rect 25620 24362 25680 24383
rect 25738 24362 25798 24383
rect 25856 24382 26152 24418
rect 25856 24362 25916 24382
rect 25974 24362 26034 24382
rect 26092 24362 26152 24382
rect 26210 24382 26506 24418
rect 26210 24362 26270 24382
rect 26328 24362 26388 24382
rect 26446 24362 26506 24382
rect 23644 24208 23794 24224
rect 23644 24174 23660 24208
rect 23694 24174 23794 24208
rect 23644 24158 23794 24174
rect 27096 24229 27156 24927
rect 27398 24879 27694 24939
rect 27398 24856 27458 24879
rect 27516 24856 27576 24879
rect 27634 24856 27694 24879
rect 27752 24880 28048 24940
rect 28393 24939 28454 24959
rect 27752 24856 27812 24880
rect 27870 24856 27930 24880
rect 27988 24856 28048 24880
rect 28374 24923 28454 24939
rect 28374 24889 28389 24923
rect 28423 24889 28454 24923
rect 28374 24873 28454 24889
rect 28393 24850 28454 24873
rect 28394 24704 28454 24850
rect 28393 24531 28454 24704
rect 27398 24430 27458 24456
rect 27366 24289 27433 24296
rect 27516 24289 27576 24456
rect 27634 24430 27694 24456
rect 27752 24430 27812 24456
rect 27366 24280 27576 24289
rect 27366 24246 27382 24280
rect 27416 24246 27576 24280
rect 27366 24230 27576 24246
rect 27096 24213 27247 24229
rect 27096 24179 27197 24213
rect 27231 24179 27247 24213
rect 27096 24163 27247 24179
rect 23734 24120 23794 24158
rect 25502 24136 25562 24162
rect 25620 24136 25680 24162
rect 25738 24136 25798 24162
rect 25856 24142 25916 24162
rect 25856 24136 25917 24142
rect 25974 24136 26034 24162
rect 26092 24136 26152 24162
rect 19649 24076 19665 24110
rect 19699 24076 19715 24110
rect 19649 24060 19715 24076
rect 19531 23993 19597 24009
rect 19531 23959 19547 23993
rect 19581 23959 19597 23993
rect 19531 23943 19597 23959
rect 19534 23921 19594 23943
rect 14424 23699 14484 23725
rect 14542 23699 14602 23725
rect 14660 23699 14720 23725
rect 14778 23699 14838 23725
rect 16322 23699 16382 23725
rect 16440 23699 16500 23725
rect 16558 23699 16618 23725
rect 16676 23699 16736 23725
rect 12647 23504 12707 23526
rect 12765 23504 12825 23526
rect 12644 23488 12710 23504
rect 6249 23441 6315 23457
rect 12644 23454 12660 23488
rect 12694 23454 12710 23488
rect 12644 23438 12710 23454
rect 12762 23488 12828 23504
rect 12762 23454 12778 23488
rect 12812 23454 12828 23488
rect 20538 23894 20598 23920
rect 19534 23695 19594 23721
rect 21836 23894 21896 23920
rect 22436 23894 22496 23920
rect 25739 23951 25797 24136
rect 25739 23925 25799 23951
rect 25857 23925 25917 24136
rect 26210 24130 26270 24162
rect 26328 24136 26388 24162
rect 26446 24136 26506 24162
rect 26207 24114 26273 24130
rect 27096 24124 27156 24163
rect 27516 24124 27576 24230
rect 27870 24289 27930 24456
rect 27988 24430 28048 24456
rect 28013 24289 28080 24296
rect 27870 24280 28080 24289
rect 27870 24246 28030 24280
rect 28064 24246 28080 24280
rect 27870 24230 28080 24246
rect 27632 24196 27698 24212
rect 27632 24162 27648 24196
rect 27682 24162 27698 24196
rect 27632 24146 27698 24162
rect 27750 24197 27816 24212
rect 27750 24163 27766 24197
rect 27800 24163 27816 24197
rect 27750 24147 27816 24163
rect 27634 24124 27694 24146
rect 27752 24124 27812 24147
rect 27870 24124 27930 24230
rect 28394 24228 28454 24531
rect 28304 24212 28454 24228
rect 28304 24178 28320 24212
rect 28354 24178 28454 24212
rect 28304 24162 28454 24178
rect 28394 24124 28454 24162
rect 28994 24423 29054 25081
rect 29707 25079 30250 25130
rect 30292 25123 30368 25130
rect 30426 25123 30486 25149
rect 30292 25079 30367 25123
rect 29296 24879 29592 24939
rect 29296 24856 29356 24879
rect 29414 24856 29474 24879
rect 29532 24856 29592 24879
rect 29650 24880 29946 24940
rect 29650 24856 29710 24880
rect 29768 24856 29828 24880
rect 29886 24856 29946 24880
rect 30292 24926 30352 25079
rect 36900 25042 36955 25102
rect 37155 25043 37885 25102
rect 37155 25042 37458 25043
rect 36900 24984 36939 25042
rect 37441 24985 37458 25042
rect 37513 25042 37885 25043
rect 37513 24985 37528 25042
rect 30292 24902 30546 24926
rect 30292 24868 30496 24902
rect 30530 24868 30546 24902
rect 30292 24852 30546 24868
rect 36900 24924 36955 24984
rect 37155 24924 37181 24984
rect 37441 24966 37528 24985
rect 36900 24866 36939 24924
rect 29296 24430 29356 24456
rect 28994 24407 29061 24423
rect 28994 24373 29010 24407
rect 29044 24373 29061 24407
rect 28994 24357 29061 24373
rect 28994 24229 29054 24357
rect 29264 24289 29331 24296
rect 29414 24289 29474 24456
rect 29532 24430 29592 24456
rect 29650 24430 29710 24456
rect 29264 24280 29474 24289
rect 29264 24246 29280 24280
rect 29314 24246 29474 24280
rect 29264 24230 29474 24246
rect 28994 24213 29145 24229
rect 28994 24179 29095 24213
rect 29129 24179 29145 24213
rect 28994 24163 29145 24179
rect 28994 24124 29054 24163
rect 29414 24124 29474 24230
rect 29768 24289 29828 24456
rect 29886 24430 29946 24456
rect 29909 24290 29976 24297
rect 29903 24289 29976 24290
rect 29768 24281 29976 24289
rect 29768 24247 29926 24281
rect 29960 24247 29976 24281
rect 29768 24231 29976 24247
rect 29768 24230 29965 24231
rect 29530 24196 29596 24212
rect 29530 24162 29546 24196
rect 29580 24162 29596 24196
rect 29530 24146 29596 24162
rect 29648 24197 29714 24212
rect 29648 24163 29664 24197
rect 29698 24163 29714 24197
rect 29648 24147 29714 24163
rect 29532 24124 29592 24146
rect 29650 24124 29710 24147
rect 29768 24124 29828 24230
rect 30292 24228 30352 24852
rect 36900 24806 36955 24866
rect 37155 24806 37181 24866
rect 36701 24601 36755 24661
rect 37155 24601 37181 24661
rect 36701 24543 36740 24601
rect 36701 24483 36755 24543
rect 37155 24483 37630 24543
rect 36701 24425 36740 24483
rect 36701 24365 36755 24425
rect 37155 24365 37181 24425
rect 30202 24212 30352 24228
rect 30202 24178 30218 24212
rect 30252 24178 30352 24212
rect 30202 24162 30352 24178
rect 30292 24124 30352 24162
rect 36701 24134 36755 24194
rect 37155 24134 37181 24194
rect 26207 24080 26223 24114
rect 26257 24080 26273 24114
rect 26207 24064 26273 24080
rect 26089 23997 26155 24013
rect 26089 23963 26105 23997
rect 26139 23963 26155 23997
rect 26089 23947 26155 23963
rect 26092 23925 26152 23947
rect 23734 23894 23794 23920
rect 20958 23694 21018 23720
rect 21076 23694 21136 23720
rect 21194 23694 21254 23720
rect 21312 23694 21372 23720
rect 22856 23694 22916 23720
rect 22974 23694 23034 23720
rect 23092 23694 23152 23720
rect 23210 23694 23270 23720
rect 19181 23499 19241 23521
rect 19299 23499 19359 23521
rect 19178 23483 19244 23499
rect 12762 23438 12828 23454
rect 19178 23449 19194 23483
rect 19228 23449 19244 23483
rect 19178 23433 19244 23449
rect 19296 23483 19362 23499
rect 19296 23449 19312 23483
rect 19346 23449 19362 23483
rect 27096 23898 27156 23924
rect 26092 23699 26152 23725
rect 28394 23898 28454 23924
rect 28994 23898 29054 23924
rect 36701 24076 36740 24134
rect 36701 24016 36755 24076
rect 37155 24075 37181 24076
rect 37342 24075 37408 24078
rect 37155 24062 37408 24075
rect 37155 24028 37358 24062
rect 37392 24028 37408 24062
rect 37155 24016 37408 24028
rect 37573 24076 37630 24483
rect 37840 24268 37885 25042
rect 37840 24208 38088 24268
rect 38288 24208 38314 24268
rect 37729 24076 37808 24087
rect 37573 24074 38088 24076
rect 37573 24016 37742 24074
rect 37797 24016 38088 24074
rect 38488 24016 38514 24076
rect 30292 23898 30352 23924
rect 36701 23958 36740 24016
rect 37341 24012 37408 24016
rect 37729 24006 37808 24016
rect 37442 23958 37529 23975
rect 36701 23898 36755 23958
rect 37155 23898 37181 23958
rect 37442 23956 38088 23958
rect 37442 23898 37457 23956
rect 37512 23898 38088 23956
rect 38488 23898 38514 23958
rect 37442 23880 37529 23898
rect 27516 23698 27576 23724
rect 27634 23698 27694 23724
rect 27752 23698 27812 23724
rect 27870 23698 27930 23724
rect 29414 23698 29474 23724
rect 29532 23698 29592 23724
rect 29650 23698 29710 23724
rect 29768 23698 29828 23724
rect 36701 23780 36755 23840
rect 37155 23780 37181 23840
rect 36701 23722 36740 23780
rect 37480 23722 37529 23880
rect 37962 23840 38028 23843
rect 38561 23885 38627 23901
rect 38561 23851 38577 23885
rect 38611 23851 38627 23885
rect 37962 23827 38088 23840
rect 37962 23793 37978 23827
rect 38012 23793 38088 23827
rect 37962 23780 38088 23793
rect 38488 23780 38514 23840
rect 38561 23835 38627 23851
rect 37962 23777 38028 23780
rect 36701 23662 36755 23722
rect 37155 23662 37529 23722
rect 37571 23722 37640 23727
rect 37571 23708 38088 23722
rect 37571 23674 37588 23708
rect 37622 23674 38088 23708
rect 37571 23662 38088 23674
rect 38488 23662 38514 23722
rect 25739 23503 25799 23525
rect 25857 23503 25917 23525
rect 25736 23487 25802 23503
rect 19296 23433 19362 23449
rect 25736 23453 25752 23487
rect 25786 23453 25802 23487
rect 25736 23437 25802 23453
rect 25854 23487 25920 23503
rect 25854 23453 25870 23487
rect 25904 23453 25920 23487
rect 36701 23604 36740 23662
rect 37571 23658 37638 23662
rect 36701 23544 36755 23604
rect 37155 23544 37181 23604
rect 25854 23437 25920 23453
rect 36701 23307 36755 23367
rect 37155 23307 37181 23367
rect 36701 23249 36740 23307
rect 37571 23249 37628 23658
rect 38569 23526 38620 23835
rect 36701 23189 36755 23249
rect 37155 23189 37628 23249
rect 37840 23466 38088 23526
rect 38288 23466 38620 23526
rect 36701 23131 36740 23189
rect 36701 23071 36755 23131
rect 37155 23071 37181 23131
rect 36900 22834 36955 22894
rect 37155 22834 37181 22894
rect 36900 22776 36939 22834
rect 36900 22716 36955 22776
rect 37155 22716 37181 22776
rect 37301 22752 37367 22768
rect 37301 22718 37317 22752
rect 37351 22718 37367 22752
rect 36900 22658 36939 22716
rect 37301 22702 37367 22718
rect 37304 22658 37364 22702
rect 37840 22658 37885 23466
rect 36900 22598 36955 22658
rect 37155 22598 37885 22658
rect 6672 22254 6738 22270
rect 6672 22245 6688 22254
rect 6151 22220 6688 22245
rect 6722 22220 6738 22254
rect 7802 22248 7868 22264
rect 7802 22241 7818 22248
rect 6151 22202 6738 22220
rect 7293 22214 7818 22241
rect 7852 22214 7868 22248
rect 6151 22150 6195 22202
rect 7293 22198 7868 22214
rect 5899 22109 6195 22150
rect 5899 22088 5959 22109
rect 6017 22088 6077 22109
rect 6135 22088 6195 22109
rect 6253 22134 6738 22150
rect 7293 22146 7337 22198
rect 13230 22250 13296 22266
rect 13230 22241 13246 22250
rect 12709 22216 13246 22241
rect 13280 22216 13296 22250
rect 14360 22244 14426 22260
rect 14360 22237 14376 22244
rect 12709 22198 13296 22216
rect 13851 22210 14376 22237
rect 14410 22210 14426 22244
rect 12709 22146 12753 22198
rect 13851 22194 14426 22210
rect 6253 22109 6688 22134
rect 6253 22088 6313 22109
rect 6371 22088 6431 22109
rect 6489 22108 6688 22109
rect 6489 22088 6549 22108
rect 6672 22100 6688 22108
rect 6722 22100 6738 22134
rect 6672 22084 6738 22100
rect 7041 22105 7337 22146
rect 7041 22084 7101 22105
rect 7159 22084 7219 22105
rect 7277 22084 7337 22105
rect 7395 22130 7868 22146
rect 7395 22105 7818 22130
rect 7395 22084 7455 22105
rect 7513 22084 7573 22105
rect 7631 22104 7818 22105
rect 7631 22084 7691 22104
rect 7802 22096 7818 22104
rect 7852 22096 7868 22130
rect 5899 21662 5959 21688
rect 6017 21662 6077 21688
rect 6135 21487 6195 21688
rect 6253 21662 6313 21688
rect 6371 21662 6431 21688
rect 6489 21671 6549 21688
rect 7802 22080 7868 22096
rect 12457 22105 12753 22146
rect 12457 22084 12517 22105
rect 12575 22084 12635 22105
rect 12693 22084 12753 22105
rect 12811 22130 13296 22146
rect 13851 22142 13895 22194
rect 19764 22255 19830 22271
rect 19764 22246 19780 22255
rect 19243 22221 19780 22246
rect 19814 22221 19830 22255
rect 20894 22249 20960 22265
rect 20894 22242 20910 22249
rect 19243 22203 19830 22221
rect 20385 22215 20910 22242
rect 20944 22215 20960 22249
rect 19243 22151 19287 22203
rect 20385 22199 20960 22215
rect 12811 22105 13246 22130
rect 12811 22084 12871 22105
rect 12929 22084 12989 22105
rect 13047 22104 13246 22105
rect 13047 22084 13107 22104
rect 13230 22096 13246 22104
rect 13280 22096 13296 22130
rect 9012 22032 9308 22068
rect 9012 22012 9072 22032
rect 9130 22012 9190 22032
rect 9248 22012 9308 22032
rect 9366 22032 9662 22068
rect 9366 22012 9426 22032
rect 9484 22012 9544 22032
rect 9602 22012 9662 22032
rect 9720 22033 10016 22069
rect 9720 22012 9780 22033
rect 9838 22012 9898 22033
rect 9956 22012 10016 22033
rect 9012 21786 9072 21812
rect 9130 21786 9190 21812
rect 9248 21780 9308 21812
rect 9366 21786 9426 21812
rect 9484 21786 9544 21812
rect 9602 21792 9662 21812
rect 9601 21786 9662 21792
rect 9720 21786 9780 21812
rect 9838 21786 9898 21812
rect 9956 21786 10016 21812
rect 9245 21764 9311 21780
rect 9245 21730 9261 21764
rect 9295 21730 9311 21764
rect 9245 21714 9311 21730
rect 6488 21582 6549 21671
rect 7041 21658 7101 21684
rect 7159 21658 7219 21684
rect 6488 21529 6639 21582
rect 6135 21436 6521 21487
rect 6340 21378 6406 21394
rect 6340 21344 6356 21378
rect 6390 21344 6406 21378
rect 5824 21305 5884 21331
rect 5942 21305 6002 21331
rect 6060 21305 6120 21331
rect 6340 21328 6406 21344
rect 6343 21305 6403 21328
rect 6461 21305 6521 21436
rect 6579 21305 6639 21529
rect 7277 21483 7337 21684
rect 7395 21658 7455 21684
rect 7513 21658 7573 21684
rect 7631 21667 7691 21684
rect 7630 21578 7691 21667
rect 9363 21647 9429 21663
rect 9363 21613 9379 21647
rect 9413 21613 9429 21647
rect 9363 21597 9429 21613
rect 7630 21525 7781 21578
rect 9366 21575 9426 21597
rect 9601 21575 9661 21786
rect 9721 21601 9779 21786
rect 13230 22080 13296 22096
rect 13599 22101 13895 22142
rect 13599 22080 13659 22101
rect 13717 22080 13777 22101
rect 13835 22080 13895 22101
rect 13953 22126 14426 22142
rect 13953 22101 14376 22126
rect 13953 22080 14013 22101
rect 14071 22080 14131 22101
rect 14189 22100 14376 22101
rect 14189 22080 14249 22100
rect 14360 22092 14376 22100
rect 14410 22092 14426 22126
rect 12457 21658 12517 21684
rect 12575 21658 12635 21684
rect 9719 21575 9779 21601
rect 7277 21432 7663 21483
rect 7482 21374 7548 21390
rect 7482 21340 7498 21374
rect 7532 21340 7548 21374
rect 6966 21301 7026 21327
rect 7084 21301 7144 21327
rect 7202 21301 7262 21327
rect 7482 21324 7548 21340
rect 7485 21301 7545 21324
rect 7603 21301 7663 21432
rect 7721 21301 7781 21525
rect 9366 21349 9426 21375
rect 5824 21073 5884 21105
rect 5942 21073 6002 21105
rect 6060 21073 6120 21105
rect 6343 21073 6403 21105
rect 6461 21079 6521 21105
rect 6579 21079 6639 21105
rect 12693 21483 12753 21684
rect 12811 21658 12871 21684
rect 12929 21658 12989 21684
rect 13047 21667 13107 21684
rect 14360 22076 14426 22092
rect 18991 22110 19287 22151
rect 18991 22089 19051 22110
rect 19109 22089 19169 22110
rect 19227 22089 19287 22110
rect 19345 22135 19830 22151
rect 20385 22147 20429 22199
rect 26277 22258 26343 22274
rect 26277 22249 26293 22258
rect 25756 22224 26293 22249
rect 26327 22224 26343 22258
rect 27407 22252 27473 22268
rect 27407 22245 27423 22252
rect 25756 22206 26343 22224
rect 26898 22218 27423 22245
rect 27457 22218 27473 22252
rect 25756 22154 25800 22206
rect 26898 22202 27473 22218
rect 19345 22110 19780 22135
rect 19345 22089 19405 22110
rect 19463 22089 19523 22110
rect 19581 22109 19780 22110
rect 19581 22089 19641 22109
rect 19764 22101 19780 22109
rect 19814 22101 19830 22135
rect 15570 22028 15866 22064
rect 15570 22008 15630 22028
rect 15688 22008 15748 22028
rect 15806 22008 15866 22028
rect 15924 22028 16220 22064
rect 15924 22008 15984 22028
rect 16042 22008 16102 22028
rect 16160 22008 16220 22028
rect 16278 22029 16574 22065
rect 16278 22008 16338 22029
rect 16396 22008 16456 22029
rect 16514 22008 16574 22029
rect 15570 21782 15630 21808
rect 15688 21782 15748 21808
rect 15806 21776 15866 21808
rect 15924 21782 15984 21808
rect 16042 21782 16102 21808
rect 16160 21788 16220 21808
rect 16159 21782 16220 21788
rect 16278 21782 16338 21808
rect 16396 21782 16456 21808
rect 16514 21782 16574 21808
rect 15803 21760 15869 21776
rect 15803 21726 15819 21760
rect 15853 21726 15869 21760
rect 15803 21710 15869 21726
rect 13046 21578 13107 21667
rect 13599 21654 13659 21680
rect 13717 21654 13777 21680
rect 13046 21525 13197 21578
rect 12693 21432 13079 21483
rect 12898 21374 12964 21390
rect 12898 21340 12914 21374
rect 12948 21340 12964 21374
rect 12382 21301 12442 21327
rect 12500 21301 12560 21327
rect 12618 21301 12678 21327
rect 12898 21324 12964 21340
rect 12901 21301 12961 21324
rect 13019 21301 13079 21432
rect 13137 21301 13197 21525
rect 13835 21479 13895 21680
rect 13953 21654 14013 21680
rect 14071 21654 14131 21680
rect 14189 21663 14249 21680
rect 14188 21574 14249 21663
rect 15921 21643 15987 21659
rect 15921 21609 15937 21643
rect 15971 21609 15987 21643
rect 15921 21593 15987 21609
rect 14188 21521 14339 21574
rect 15924 21571 15984 21593
rect 16159 21571 16219 21782
rect 16279 21597 16337 21782
rect 19764 22085 19830 22101
rect 20133 22106 20429 22147
rect 20133 22085 20193 22106
rect 20251 22085 20311 22106
rect 20369 22085 20429 22106
rect 20487 22131 20960 22147
rect 20487 22106 20910 22131
rect 20487 22085 20547 22106
rect 20605 22085 20665 22106
rect 20723 22105 20910 22106
rect 20723 22085 20783 22105
rect 20894 22097 20910 22105
rect 20944 22097 20960 22131
rect 18991 21663 19051 21689
rect 19109 21663 19169 21689
rect 16277 21571 16337 21597
rect 13835 21428 14221 21479
rect 14040 21370 14106 21386
rect 14040 21336 14056 21370
rect 14090 21336 14106 21370
rect 9601 21153 9661 21175
rect 9719 21153 9779 21175
rect 9598 21137 9664 21153
rect 9598 21103 9614 21137
rect 9648 21103 9664 21137
rect 5824 21032 6403 21073
rect 6966 21069 7026 21101
rect 7084 21069 7144 21101
rect 7202 21069 7262 21101
rect 7485 21069 7545 21101
rect 7603 21075 7663 21101
rect 7721 21075 7781 21101
rect 9598 21087 9664 21103
rect 9716 21137 9782 21153
rect 9716 21103 9732 21137
rect 9766 21103 9782 21137
rect 9716 21087 9782 21103
rect 13524 21297 13584 21323
rect 13642 21297 13702 21323
rect 13760 21297 13820 21323
rect 14040 21320 14106 21336
rect 14043 21297 14103 21320
rect 14161 21297 14221 21428
rect 14279 21297 14339 21521
rect 15924 21345 15984 21371
rect 6966 21028 7545 21069
rect 12382 21069 12442 21101
rect 12500 21069 12560 21101
rect 12618 21069 12678 21101
rect 12901 21069 12961 21101
rect 13019 21075 13079 21101
rect 13137 21075 13197 21101
rect 19227 21488 19287 21689
rect 19345 21663 19405 21689
rect 19463 21663 19523 21689
rect 19581 21672 19641 21689
rect 20894 22081 20960 22097
rect 25504 22113 25800 22154
rect 25504 22092 25564 22113
rect 25622 22092 25682 22113
rect 25740 22092 25800 22113
rect 25858 22138 26343 22154
rect 26898 22150 26942 22202
rect 25858 22113 26293 22138
rect 25858 22092 25918 22113
rect 25976 22092 26036 22113
rect 26094 22112 26293 22113
rect 26094 22092 26154 22112
rect 26277 22104 26293 22112
rect 26327 22104 26343 22138
rect 22104 22033 22400 22069
rect 22104 22013 22164 22033
rect 22222 22013 22282 22033
rect 22340 22013 22400 22033
rect 22458 22033 22754 22069
rect 22458 22013 22518 22033
rect 22576 22013 22636 22033
rect 22694 22013 22754 22033
rect 22812 22034 23108 22070
rect 22812 22013 22872 22034
rect 22930 22013 22990 22034
rect 23048 22013 23108 22034
rect 22104 21787 22164 21813
rect 22222 21787 22282 21813
rect 22340 21781 22400 21813
rect 22458 21787 22518 21813
rect 22576 21787 22636 21813
rect 22694 21793 22754 21813
rect 22693 21787 22754 21793
rect 22812 21787 22872 21813
rect 22930 21787 22990 21813
rect 23048 21787 23108 21813
rect 22337 21765 22403 21781
rect 22337 21731 22353 21765
rect 22387 21731 22403 21765
rect 22337 21715 22403 21731
rect 19580 21583 19641 21672
rect 20133 21659 20193 21685
rect 20251 21659 20311 21685
rect 19580 21530 19731 21583
rect 19227 21437 19613 21488
rect 19432 21379 19498 21395
rect 19432 21345 19448 21379
rect 19482 21345 19498 21379
rect 18916 21306 18976 21332
rect 19034 21306 19094 21332
rect 19152 21306 19212 21332
rect 19432 21329 19498 21345
rect 19435 21306 19495 21329
rect 19553 21306 19613 21437
rect 19671 21306 19731 21530
rect 20369 21484 20429 21685
rect 20487 21659 20547 21685
rect 20605 21659 20665 21685
rect 20723 21668 20783 21685
rect 20722 21579 20783 21668
rect 22455 21648 22521 21664
rect 22455 21614 22471 21648
rect 22505 21614 22521 21648
rect 22455 21598 22521 21614
rect 20722 21526 20873 21579
rect 22458 21576 22518 21598
rect 22693 21576 22753 21787
rect 22813 21602 22871 21787
rect 26277 22088 26343 22104
rect 26646 22109 26942 22150
rect 26646 22088 26706 22109
rect 26764 22088 26824 22109
rect 26882 22088 26942 22109
rect 27000 22134 27473 22150
rect 27000 22109 27423 22134
rect 27000 22088 27060 22109
rect 27118 22088 27178 22109
rect 27236 22108 27423 22109
rect 27236 22088 27296 22108
rect 27407 22100 27423 22108
rect 27457 22100 27473 22134
rect 25504 21666 25564 21692
rect 25622 21666 25682 21692
rect 22811 21576 22871 21602
rect 20369 21433 20755 21484
rect 20574 21375 20640 21391
rect 20574 21341 20590 21375
rect 20624 21341 20640 21375
rect 16159 21149 16219 21171
rect 16277 21149 16337 21171
rect 16156 21133 16222 21149
rect 16156 21099 16172 21133
rect 16206 21099 16222 21133
rect 12382 21028 12961 21069
rect 13524 21065 13584 21097
rect 13642 21065 13702 21097
rect 13760 21065 13820 21097
rect 14043 21065 14103 21097
rect 14161 21071 14221 21097
rect 14279 21071 14339 21097
rect 16156 21083 16222 21099
rect 16274 21133 16340 21149
rect 16274 21099 16290 21133
rect 16324 21099 16340 21133
rect 20058 21302 20118 21328
rect 20176 21302 20236 21328
rect 20294 21302 20354 21328
rect 20574 21325 20640 21341
rect 20577 21302 20637 21325
rect 20695 21302 20755 21433
rect 20813 21302 20873 21526
rect 22458 21350 22518 21376
rect 16274 21083 16340 21099
rect 18916 21074 18976 21106
rect 19034 21074 19094 21106
rect 19152 21074 19212 21106
rect 19435 21074 19495 21106
rect 19553 21080 19613 21106
rect 19671 21080 19731 21106
rect 25740 21491 25800 21692
rect 25858 21666 25918 21692
rect 25976 21666 26036 21692
rect 26094 21675 26154 21692
rect 27407 22084 27473 22100
rect 28617 22036 28913 22072
rect 28617 22016 28677 22036
rect 28735 22016 28795 22036
rect 28853 22016 28913 22036
rect 28971 22036 29267 22072
rect 28971 22016 29031 22036
rect 29089 22016 29149 22036
rect 29207 22016 29267 22036
rect 29325 22037 29621 22073
rect 29325 22016 29385 22037
rect 29443 22016 29503 22037
rect 29561 22016 29621 22037
rect 36900 21898 36955 21958
rect 37155 21899 37885 21958
rect 37155 21898 37458 21899
rect 36900 21840 36939 21898
rect 37441 21841 37458 21898
rect 37513 21898 37885 21899
rect 37513 21841 37528 21898
rect 28617 21790 28677 21816
rect 28735 21790 28795 21816
rect 28853 21784 28913 21816
rect 28971 21790 29031 21816
rect 29089 21790 29149 21816
rect 29207 21796 29267 21816
rect 29206 21790 29267 21796
rect 29325 21790 29385 21816
rect 29443 21790 29503 21816
rect 29561 21790 29621 21816
rect 28850 21768 28916 21784
rect 28850 21734 28866 21768
rect 28900 21734 28916 21768
rect 28850 21718 28916 21734
rect 26093 21586 26154 21675
rect 26646 21662 26706 21688
rect 26764 21662 26824 21688
rect 26093 21533 26244 21586
rect 25740 21440 26126 21491
rect 25945 21382 26011 21398
rect 25945 21348 25961 21382
rect 25995 21348 26011 21382
rect 25429 21309 25489 21335
rect 25547 21309 25607 21335
rect 25665 21309 25725 21335
rect 25945 21332 26011 21348
rect 25948 21309 26008 21332
rect 26066 21309 26126 21440
rect 26184 21309 26244 21533
rect 26882 21487 26942 21688
rect 27000 21662 27060 21688
rect 27118 21662 27178 21688
rect 27236 21671 27296 21688
rect 27235 21582 27296 21671
rect 28968 21651 29034 21667
rect 28968 21617 28984 21651
rect 29018 21617 29034 21651
rect 28968 21601 29034 21617
rect 27235 21529 27386 21582
rect 28971 21579 29031 21601
rect 29206 21579 29266 21790
rect 29326 21605 29384 21790
rect 36900 21780 36955 21840
rect 37155 21780 37181 21840
rect 37441 21822 37528 21841
rect 36900 21722 36939 21780
rect 36900 21662 36955 21722
rect 37155 21662 37181 21722
rect 29324 21579 29384 21605
rect 26882 21436 27268 21487
rect 27087 21378 27153 21394
rect 27087 21344 27103 21378
rect 27137 21344 27153 21378
rect 22693 21154 22753 21176
rect 22811 21154 22871 21176
rect 22690 21138 22756 21154
rect 22690 21104 22706 21138
rect 22740 21104 22756 21138
rect 13524 21024 14103 21065
rect 18916 21033 19495 21074
rect 20058 21070 20118 21102
rect 20176 21070 20236 21102
rect 20294 21070 20354 21102
rect 20577 21070 20637 21102
rect 20695 21076 20755 21102
rect 20813 21076 20873 21102
rect 22690 21088 22756 21104
rect 22808 21138 22874 21154
rect 22808 21104 22824 21138
rect 22858 21104 22874 21138
rect 26571 21305 26631 21331
rect 26689 21305 26749 21331
rect 26807 21305 26867 21331
rect 27087 21328 27153 21344
rect 27090 21305 27150 21328
rect 27208 21305 27268 21436
rect 27326 21305 27386 21529
rect 28971 21353 29031 21379
rect 22808 21088 22874 21104
rect 25429 21077 25489 21109
rect 25547 21077 25607 21109
rect 25665 21077 25725 21109
rect 25948 21077 26008 21109
rect 26066 21083 26126 21109
rect 26184 21083 26244 21109
rect 36701 21457 36755 21517
rect 37155 21457 37181 21517
rect 36701 21399 36740 21457
rect 36701 21339 36755 21399
rect 37155 21339 37630 21399
rect 36701 21281 36740 21339
rect 36701 21221 36755 21281
rect 37155 21221 37181 21281
rect 29206 21157 29266 21179
rect 29324 21157 29384 21179
rect 29203 21141 29269 21157
rect 29203 21107 29219 21141
rect 29253 21107 29269 21141
rect 20058 21029 20637 21070
rect 25429 21036 26008 21077
rect 26571 21073 26631 21105
rect 26689 21073 26749 21105
rect 26807 21073 26867 21105
rect 27090 21073 27150 21105
rect 27208 21079 27268 21105
rect 27326 21079 27386 21105
rect 29203 21091 29269 21107
rect 29321 21141 29387 21157
rect 29321 21107 29337 21141
rect 29371 21107 29387 21141
rect 29321 21091 29387 21107
rect 26571 21032 27150 21073
rect 36701 20990 36755 21050
rect 37155 20990 37181 21050
rect 36701 20932 36740 20990
rect 36701 20872 36755 20932
rect 37155 20931 37181 20932
rect 37342 20931 37408 20934
rect 37155 20918 37408 20931
rect 37155 20884 37358 20918
rect 37392 20884 37408 20918
rect 37155 20872 37408 20884
rect 37573 20932 37630 21339
rect 37840 21124 37885 21898
rect 37840 21064 38088 21124
rect 38288 21064 38314 21124
rect 37729 20932 37808 20943
rect 37573 20930 38088 20932
rect 37573 20872 37742 20930
rect 37797 20872 38088 20930
rect 38488 20872 38514 20932
rect 36701 20814 36740 20872
rect 37341 20868 37408 20872
rect 37729 20862 37808 20872
rect 37442 20814 37529 20831
rect 36701 20754 36755 20814
rect 37155 20754 37181 20814
rect 37442 20812 38088 20814
rect 37442 20754 37457 20812
rect 37512 20754 38088 20812
rect 38488 20754 38514 20814
rect 37442 20736 37529 20754
rect 36701 20636 36755 20696
rect 37155 20636 37181 20696
rect 36701 20578 36740 20636
rect 37480 20578 37529 20736
rect 37962 20696 38028 20699
rect 38561 20741 38627 20757
rect 38561 20707 38577 20741
rect 38611 20707 38627 20741
rect 37962 20683 38088 20696
rect 37962 20649 37978 20683
rect 38012 20649 38088 20683
rect 37962 20636 38088 20649
rect 38488 20636 38514 20696
rect 38561 20691 38627 20707
rect 37962 20633 38028 20636
rect 36701 20518 36755 20578
rect 37155 20518 37529 20578
rect 37571 20578 37640 20583
rect 37571 20564 38088 20578
rect 37571 20530 37588 20564
rect 37622 20530 38088 20564
rect 37571 20518 38088 20530
rect 38488 20518 38514 20578
rect 8998 20382 9294 20418
rect 8998 20362 9058 20382
rect 9116 20362 9176 20382
rect 9234 20362 9294 20382
rect 9352 20382 9648 20418
rect 9352 20362 9412 20382
rect 9470 20362 9530 20382
rect 9588 20362 9648 20382
rect 9706 20383 10002 20419
rect 9706 20362 9766 20383
rect 9824 20362 9884 20383
rect 9942 20362 10002 20383
rect 15556 20378 15852 20414
rect 15556 20358 15616 20378
rect 15674 20358 15734 20378
rect 15792 20358 15852 20378
rect 15910 20378 16206 20414
rect 15910 20358 15970 20378
rect 16028 20358 16088 20378
rect 16146 20358 16206 20378
rect 16264 20379 16560 20415
rect 16264 20358 16324 20379
rect 16382 20358 16442 20379
rect 16500 20358 16560 20379
rect 8998 20136 9058 20162
rect 9116 20136 9176 20162
rect 9234 20130 9294 20162
rect 9352 20136 9412 20162
rect 9470 20136 9530 20162
rect 9588 20142 9648 20162
rect 9587 20136 9648 20142
rect 9706 20136 9766 20162
rect 9824 20136 9884 20162
rect 9942 20136 10002 20162
rect 22090 20383 22386 20419
rect 22090 20363 22150 20383
rect 22208 20363 22268 20383
rect 22326 20363 22386 20383
rect 22444 20383 22740 20419
rect 22444 20363 22504 20383
rect 22562 20363 22622 20383
rect 22680 20363 22740 20383
rect 22798 20384 23094 20420
rect 22798 20363 22858 20384
rect 22916 20363 22976 20384
rect 23034 20363 23094 20384
rect 36701 20460 36740 20518
rect 37571 20514 37638 20518
rect 28603 20386 28899 20422
rect 28603 20366 28663 20386
rect 28721 20366 28781 20386
rect 28839 20366 28899 20386
rect 28957 20386 29253 20422
rect 28957 20366 29017 20386
rect 29075 20366 29135 20386
rect 29193 20366 29253 20386
rect 29311 20387 29607 20423
rect 36701 20400 36755 20460
rect 37155 20400 37181 20460
rect 29311 20366 29371 20387
rect 29429 20366 29489 20387
rect 29547 20366 29607 20387
rect 9231 20114 9297 20130
rect 9231 20080 9247 20114
rect 9281 20080 9297 20114
rect 9231 20064 9297 20080
rect 5506 19945 5566 19971
rect 5624 19945 5684 19971
rect 5742 19945 5802 19971
rect 5860 19960 6156 20011
rect 5860 19945 5920 19960
rect 5978 19945 6038 19960
rect 6096 19945 6156 19960
rect 7404 19945 7464 19971
rect 7522 19945 7582 19971
rect 7640 19945 7700 19971
rect 7758 19960 8054 20011
rect 7758 19945 7818 19960
rect 7876 19945 7936 19960
rect 7994 19945 8054 19960
rect 9349 19997 9415 20013
rect 9349 19963 9365 19997
rect 9399 19963 9415 19997
rect 9349 19947 9415 19963
rect 5023 19762 5319 19813
rect 5023 19745 5083 19762
rect 5141 19745 5201 19762
rect 5259 19745 5319 19762
rect 6344 19745 6404 19771
rect 6462 19745 6522 19771
rect 6580 19745 6640 19771
rect 6921 19762 7217 19813
rect 6921 19745 6981 19762
rect 7039 19745 7099 19762
rect 7157 19745 7217 19762
rect 9352 19925 9412 19947
rect 9587 19925 9647 20136
rect 9707 19951 9765 20136
rect 15556 20132 15616 20158
rect 15674 20132 15734 20158
rect 15792 20126 15852 20158
rect 15910 20132 15970 20158
rect 16028 20132 16088 20158
rect 16146 20138 16206 20158
rect 16145 20132 16206 20138
rect 16264 20132 16324 20158
rect 16382 20132 16442 20158
rect 16500 20132 16560 20158
rect 22090 20137 22150 20163
rect 22208 20137 22268 20163
rect 15789 20110 15855 20126
rect 15789 20076 15805 20110
rect 15839 20076 15855 20110
rect 15789 20060 15855 20076
rect 9705 19925 9765 19951
rect 12064 19941 12124 19967
rect 12182 19941 12242 19967
rect 12300 19941 12360 19967
rect 12418 19956 12714 20007
rect 12418 19941 12478 19956
rect 12536 19941 12596 19956
rect 12654 19941 12714 19956
rect 13962 19941 14022 19967
rect 14080 19941 14140 19967
rect 14198 19941 14258 19967
rect 14316 19956 14612 20007
rect 14316 19941 14376 19956
rect 14434 19941 14494 19956
rect 14552 19941 14612 19956
rect 15907 19993 15973 20009
rect 15907 19959 15923 19993
rect 15957 19959 15973 19993
rect 15907 19943 15973 19959
rect 8242 19745 8302 19771
rect 8360 19745 8420 19771
rect 8478 19745 8538 19771
rect 9352 19699 9412 19725
rect 5023 19519 5083 19545
rect 5141 19526 5201 19545
rect 5259 19526 5319 19545
rect 5506 19526 5566 19545
rect 5624 19526 5684 19545
rect 5742 19526 5802 19545
rect 5141 19519 5217 19526
rect 5142 19475 5217 19519
rect 5259 19475 5802 19526
rect 5860 19519 5920 19545
rect 5978 19519 6038 19545
rect 6096 19528 6156 19545
rect 6344 19528 6404 19545
rect 6462 19528 6522 19545
rect 6580 19528 6640 19545
rect 6096 19477 6640 19528
rect 6921 19519 6981 19545
rect 7039 19526 7099 19545
rect 7157 19526 7217 19545
rect 7404 19526 7464 19545
rect 7522 19526 7582 19545
rect 7640 19526 7700 19545
rect 7039 19519 7115 19526
rect 5157 19322 5217 19475
rect 4963 19298 5217 19322
rect 4963 19264 4979 19298
rect 5013 19264 5217 19298
rect 4963 19248 5217 19264
rect 5563 19276 5859 19336
rect 5563 19252 5623 19276
rect 5681 19252 5741 19276
rect 5799 19252 5859 19276
rect 5917 19275 6213 19335
rect 5917 19252 5977 19275
rect 6035 19252 6095 19275
rect 6153 19252 6213 19275
rect 5157 18624 5217 19248
rect 5563 18826 5623 18852
rect 5533 18686 5600 18693
rect 5533 18685 5606 18686
rect 5681 18685 5741 18852
rect 5799 18826 5859 18852
rect 5917 18826 5977 18852
rect 5533 18677 5741 18685
rect 5533 18643 5549 18677
rect 5583 18643 5741 18677
rect 5533 18627 5741 18643
rect 5544 18626 5741 18627
rect 5157 18608 5307 18624
rect 5157 18574 5257 18608
rect 5291 18574 5307 18608
rect 5157 18558 5307 18574
rect 5157 18520 5217 18558
rect 5681 18520 5741 18626
rect 6035 18685 6095 18852
rect 6153 18826 6213 18852
rect 6455 18819 6515 19477
rect 7040 19475 7115 19519
rect 7157 19475 7700 19526
rect 7758 19519 7818 19545
rect 7876 19519 7936 19545
rect 7994 19528 8054 19545
rect 8242 19528 8302 19545
rect 8360 19528 8420 19545
rect 8478 19528 8538 19545
rect 7994 19477 8538 19528
rect 11581 19758 11877 19809
rect 11581 19741 11641 19758
rect 11699 19741 11759 19758
rect 11817 19741 11877 19758
rect 12902 19741 12962 19767
rect 13020 19741 13080 19767
rect 13138 19741 13198 19767
rect 13479 19758 13775 19809
rect 13479 19741 13539 19758
rect 13597 19741 13657 19758
rect 13715 19741 13775 19758
rect 15910 19921 15970 19943
rect 16145 19921 16205 20132
rect 16265 19947 16323 20132
rect 22326 20131 22386 20163
rect 22444 20137 22504 20163
rect 22562 20137 22622 20163
rect 22680 20143 22740 20163
rect 22679 20137 22740 20143
rect 22798 20137 22858 20163
rect 22916 20137 22976 20163
rect 23034 20137 23094 20163
rect 28603 20140 28663 20166
rect 28721 20140 28781 20166
rect 22323 20115 22389 20131
rect 22323 20081 22339 20115
rect 22373 20081 22389 20115
rect 22323 20065 22389 20081
rect 16263 19921 16323 19947
rect 18598 19946 18658 19972
rect 18716 19946 18776 19972
rect 18834 19946 18894 19972
rect 18952 19961 19248 20012
rect 18952 19946 19012 19961
rect 19070 19946 19130 19961
rect 19188 19946 19248 19961
rect 20496 19946 20556 19972
rect 20614 19946 20674 19972
rect 20732 19946 20792 19972
rect 20850 19961 21146 20012
rect 20850 19946 20910 19961
rect 20968 19946 21028 19961
rect 21086 19946 21146 19961
rect 22441 19998 22507 20014
rect 22441 19964 22457 19998
rect 22491 19964 22507 19998
rect 22441 19948 22507 19964
rect 14800 19741 14860 19767
rect 14918 19741 14978 19767
rect 15036 19741 15096 19767
rect 15910 19695 15970 19721
rect 9587 19509 9647 19525
rect 6448 18803 6515 18819
rect 6448 18769 6465 18803
rect 6499 18769 6515 18803
rect 6448 18753 6515 18769
rect 6178 18685 6245 18692
rect 6035 18676 6245 18685
rect 6035 18642 6195 18676
rect 6229 18642 6245 18676
rect 6035 18626 6245 18642
rect 5795 18593 5861 18608
rect 5795 18559 5811 18593
rect 5845 18559 5861 18593
rect 5795 18543 5861 18559
rect 5913 18592 5979 18608
rect 5913 18558 5929 18592
rect 5963 18558 5979 18592
rect 5799 18520 5859 18543
rect 5913 18542 5979 18558
rect 5917 18520 5977 18542
rect 6035 18520 6095 18626
rect 6455 18625 6515 18753
rect 6364 18609 6515 18625
rect 6364 18575 6380 18609
rect 6414 18575 6515 18609
rect 6364 18559 6515 18575
rect 6455 18520 6515 18559
rect 7055 19355 7115 19475
rect 8353 19396 8413 19477
rect 9579 19487 9653 19509
rect 9705 19503 9765 19525
rect 11581 19515 11641 19541
rect 11699 19522 11759 19541
rect 11817 19522 11877 19541
rect 12064 19522 12124 19541
rect 12182 19522 12242 19541
rect 12300 19522 12360 19541
rect 11699 19515 11775 19522
rect 9579 19453 9600 19487
rect 9634 19453 9653 19487
rect 9579 19396 9653 19453
rect 9702 19487 9768 19503
rect 9702 19453 9718 19487
rect 9752 19453 9768 19487
rect 11700 19471 11775 19515
rect 11817 19471 12360 19522
rect 12418 19515 12478 19541
rect 12536 19515 12596 19541
rect 12654 19524 12714 19541
rect 12902 19524 12962 19541
rect 13020 19524 13080 19541
rect 13138 19524 13198 19541
rect 12654 19473 13198 19524
rect 13479 19515 13539 19541
rect 13597 19522 13657 19541
rect 13715 19522 13775 19541
rect 13962 19522 14022 19541
rect 14080 19522 14140 19541
rect 14198 19522 14258 19541
rect 13597 19515 13673 19522
rect 9702 19437 9768 19453
rect 8353 19371 9653 19396
rect 7055 19335 7116 19355
rect 7055 19319 7135 19335
rect 7055 19285 7086 19319
rect 7120 19285 7135 19319
rect 7055 19269 7135 19285
rect 7461 19276 7757 19336
rect 7055 19246 7116 19269
rect 7461 19252 7521 19276
rect 7579 19252 7639 19276
rect 7697 19252 7757 19276
rect 7815 19275 8111 19335
rect 7815 19252 7875 19275
rect 7933 19252 7993 19275
rect 8051 19252 8111 19275
rect 8353 19323 9654 19371
rect 7055 19100 7115 19246
rect 7055 18927 7116 19100
rect 7055 18624 7115 18927
rect 7461 18826 7521 18852
rect 7429 18685 7496 18692
rect 7579 18685 7639 18852
rect 7697 18826 7757 18852
rect 7815 18826 7875 18852
rect 7429 18676 7639 18685
rect 7429 18642 7445 18676
rect 7479 18642 7639 18676
rect 7429 18626 7639 18642
rect 7055 18608 7205 18624
rect 7055 18574 7155 18608
rect 7189 18574 7205 18608
rect 7055 18558 7205 18574
rect 7055 18520 7115 18558
rect 7579 18520 7639 18626
rect 7933 18685 7993 18852
rect 8051 18826 8111 18852
rect 8076 18685 8143 18692
rect 7933 18676 8143 18685
rect 7933 18642 8093 18676
rect 8127 18642 8143 18676
rect 7933 18626 8143 18642
rect 7693 18593 7759 18608
rect 7693 18559 7709 18593
rect 7743 18559 7759 18593
rect 7693 18543 7759 18559
rect 7811 18592 7877 18608
rect 7811 18558 7827 18592
rect 7861 18558 7877 18592
rect 7697 18520 7757 18543
rect 7811 18542 7877 18558
rect 7815 18520 7875 18542
rect 7933 18520 7993 18626
rect 8353 18625 8413 19323
rect 11715 19318 11775 19471
rect 11521 19294 11775 19318
rect 11521 19260 11537 19294
rect 11571 19260 11775 19294
rect 11521 19244 11775 19260
rect 12121 19272 12417 19332
rect 12121 19248 12181 19272
rect 12239 19248 12299 19272
rect 12357 19248 12417 19272
rect 12475 19271 12771 19331
rect 12475 19248 12535 19271
rect 12593 19248 12653 19271
rect 12711 19248 12771 19271
rect 9003 18778 9299 18814
rect 9003 18758 9063 18778
rect 9121 18758 9181 18778
rect 9239 18758 9299 18778
rect 9357 18778 9653 18814
rect 9357 18758 9417 18778
rect 9475 18758 9535 18778
rect 9593 18758 9653 18778
rect 9711 18779 10007 18815
rect 9711 18758 9771 18779
rect 9829 18758 9889 18779
rect 9947 18758 10007 18779
rect 8262 18609 8413 18625
rect 8262 18575 8278 18609
rect 8312 18575 8413 18609
rect 8262 18559 8413 18575
rect 8353 18520 8413 18559
rect 11715 18620 11775 19244
rect 12121 18822 12181 18848
rect 12091 18682 12158 18689
rect 12091 18681 12164 18682
rect 12239 18681 12299 18848
rect 12357 18822 12417 18848
rect 12475 18822 12535 18848
rect 12091 18673 12299 18681
rect 12091 18639 12107 18673
rect 12141 18639 12299 18673
rect 12091 18623 12299 18639
rect 12102 18622 12299 18623
rect 11715 18604 11865 18620
rect 11715 18570 11815 18604
rect 11849 18570 11865 18604
rect 9003 18532 9063 18558
rect 9121 18532 9181 18558
rect 9239 18526 9299 18558
rect 9357 18532 9417 18558
rect 9475 18532 9535 18558
rect 9593 18538 9653 18558
rect 9592 18532 9653 18538
rect 9711 18532 9771 18558
rect 9829 18532 9889 18558
rect 9947 18532 10007 18558
rect 11715 18554 11865 18570
rect 5157 18294 5217 18320
rect 6455 18294 6515 18320
rect 7055 18294 7115 18320
rect 9236 18510 9302 18526
rect 9236 18476 9252 18510
rect 9286 18476 9302 18510
rect 9236 18460 9302 18476
rect 9354 18393 9420 18409
rect 9354 18359 9370 18393
rect 9404 18359 9420 18393
rect 9354 18343 9420 18359
rect 9357 18321 9417 18343
rect 9592 18321 9652 18532
rect 9712 18347 9770 18532
rect 11715 18516 11775 18554
rect 12239 18516 12299 18622
rect 12593 18681 12653 18848
rect 12711 18822 12771 18848
rect 13013 18815 13073 19473
rect 13598 19471 13673 19515
rect 13715 19471 14258 19522
rect 14316 19515 14376 19541
rect 14434 19515 14494 19541
rect 14552 19524 14612 19541
rect 14800 19524 14860 19541
rect 14918 19524 14978 19541
rect 15036 19524 15096 19541
rect 14552 19473 15096 19524
rect 18115 19763 18411 19814
rect 18115 19746 18175 19763
rect 18233 19746 18293 19763
rect 18351 19746 18411 19763
rect 19436 19746 19496 19772
rect 19554 19746 19614 19772
rect 19672 19746 19732 19772
rect 20013 19763 20309 19814
rect 20013 19746 20073 19763
rect 20131 19746 20191 19763
rect 20249 19746 20309 19763
rect 22444 19926 22504 19948
rect 22679 19926 22739 20137
rect 22799 19952 22857 20137
rect 28839 20134 28899 20166
rect 28957 20140 29017 20166
rect 29075 20140 29135 20166
rect 29193 20146 29253 20166
rect 29192 20140 29253 20146
rect 29311 20140 29371 20166
rect 29429 20140 29489 20166
rect 29547 20140 29607 20166
rect 36701 20163 36755 20223
rect 37155 20163 37181 20223
rect 28836 20118 28902 20134
rect 28836 20084 28852 20118
rect 28886 20084 28902 20118
rect 28836 20068 28902 20084
rect 22797 19926 22857 19952
rect 25111 19949 25171 19975
rect 25229 19949 25289 19975
rect 25347 19949 25407 19975
rect 25465 19964 25761 20015
rect 25465 19949 25525 19964
rect 25583 19949 25643 19964
rect 25701 19949 25761 19964
rect 27009 19949 27069 19975
rect 27127 19949 27187 19975
rect 27245 19949 27305 19975
rect 27363 19964 27659 20015
rect 27363 19949 27423 19964
rect 27481 19949 27541 19964
rect 27599 19949 27659 19964
rect 28954 20001 29020 20017
rect 28954 19967 28970 20001
rect 29004 19967 29020 20001
rect 28954 19951 29020 19967
rect 21334 19746 21394 19772
rect 21452 19746 21512 19772
rect 21570 19746 21630 19772
rect 22444 19700 22504 19726
rect 16145 19505 16205 19521
rect 13006 18799 13073 18815
rect 13006 18765 13023 18799
rect 13057 18765 13073 18799
rect 13006 18749 13073 18765
rect 12736 18681 12803 18688
rect 12593 18672 12803 18681
rect 12593 18638 12753 18672
rect 12787 18638 12803 18672
rect 12593 18622 12803 18638
rect 12353 18589 12419 18604
rect 12353 18555 12369 18589
rect 12403 18555 12419 18589
rect 12353 18539 12419 18555
rect 12471 18588 12537 18604
rect 12471 18554 12487 18588
rect 12521 18554 12537 18588
rect 12357 18516 12417 18539
rect 12471 18538 12537 18554
rect 12475 18516 12535 18538
rect 12593 18516 12653 18622
rect 13013 18621 13073 18749
rect 12922 18605 13073 18621
rect 12922 18571 12938 18605
rect 12972 18571 13073 18605
rect 12922 18555 13073 18571
rect 13013 18516 13073 18555
rect 13613 19351 13673 19471
rect 14911 19392 14971 19473
rect 16137 19483 16211 19505
rect 16263 19499 16323 19521
rect 18115 19520 18175 19546
rect 18233 19527 18293 19546
rect 18351 19527 18411 19546
rect 18598 19527 18658 19546
rect 18716 19527 18776 19546
rect 18834 19527 18894 19546
rect 18233 19520 18309 19527
rect 16137 19449 16158 19483
rect 16192 19449 16211 19483
rect 16137 19392 16211 19449
rect 16260 19483 16326 19499
rect 16260 19449 16276 19483
rect 16310 19449 16326 19483
rect 18234 19476 18309 19520
rect 18351 19476 18894 19527
rect 18952 19520 19012 19546
rect 19070 19520 19130 19546
rect 19188 19529 19248 19546
rect 19436 19529 19496 19546
rect 19554 19529 19614 19546
rect 19672 19529 19732 19546
rect 19188 19478 19732 19529
rect 20013 19520 20073 19546
rect 20131 19527 20191 19546
rect 20249 19527 20309 19546
rect 20496 19527 20556 19546
rect 20614 19527 20674 19546
rect 20732 19527 20792 19546
rect 20131 19520 20207 19527
rect 16260 19433 16326 19449
rect 14911 19367 16211 19392
rect 13613 19331 13674 19351
rect 13613 19315 13693 19331
rect 13613 19281 13644 19315
rect 13678 19281 13693 19315
rect 13613 19265 13693 19281
rect 14019 19272 14315 19332
rect 13613 19242 13674 19265
rect 14019 19248 14079 19272
rect 14137 19248 14197 19272
rect 14255 19248 14315 19272
rect 14373 19271 14669 19331
rect 14373 19248 14433 19271
rect 14491 19248 14551 19271
rect 14609 19248 14669 19271
rect 14911 19319 16212 19367
rect 18249 19323 18309 19476
rect 13613 19096 13673 19242
rect 13613 18923 13674 19096
rect 13613 18620 13673 18923
rect 14019 18822 14079 18848
rect 13987 18681 14054 18688
rect 14137 18681 14197 18848
rect 14255 18822 14315 18848
rect 14373 18822 14433 18848
rect 13987 18672 14197 18681
rect 13987 18638 14003 18672
rect 14037 18638 14197 18672
rect 13987 18622 14197 18638
rect 13613 18604 13763 18620
rect 13613 18570 13713 18604
rect 13747 18570 13763 18604
rect 13613 18554 13763 18570
rect 13613 18516 13673 18554
rect 14137 18516 14197 18622
rect 14491 18681 14551 18848
rect 14609 18822 14669 18848
rect 14634 18681 14701 18688
rect 14491 18672 14701 18681
rect 14491 18638 14651 18672
rect 14685 18638 14701 18672
rect 14491 18622 14701 18638
rect 14251 18589 14317 18604
rect 14251 18555 14267 18589
rect 14301 18555 14317 18589
rect 14251 18539 14317 18555
rect 14369 18588 14435 18604
rect 14369 18554 14385 18588
rect 14419 18554 14435 18588
rect 14255 18516 14315 18539
rect 14369 18538 14435 18554
rect 14373 18516 14433 18538
rect 14491 18516 14551 18622
rect 14911 18621 14971 19319
rect 18055 19299 18309 19323
rect 18055 19265 18071 19299
rect 18105 19265 18309 19299
rect 18055 19249 18309 19265
rect 18655 19277 18951 19337
rect 18655 19253 18715 19277
rect 18773 19253 18833 19277
rect 18891 19253 18951 19277
rect 19009 19276 19305 19336
rect 19009 19253 19069 19276
rect 19127 19253 19187 19276
rect 19245 19253 19305 19276
rect 15561 18774 15857 18810
rect 15561 18754 15621 18774
rect 15679 18754 15739 18774
rect 15797 18754 15857 18774
rect 15915 18774 16211 18810
rect 15915 18754 15975 18774
rect 16033 18754 16093 18774
rect 16151 18754 16211 18774
rect 16269 18775 16565 18811
rect 16269 18754 16329 18775
rect 16387 18754 16447 18775
rect 16505 18754 16565 18775
rect 14820 18605 14971 18621
rect 14820 18571 14836 18605
rect 14870 18571 14971 18605
rect 14820 18555 14971 18571
rect 14911 18516 14971 18555
rect 18249 18625 18309 19249
rect 18655 18827 18715 18853
rect 18625 18687 18692 18694
rect 18625 18686 18698 18687
rect 18773 18686 18833 18853
rect 18891 18827 18951 18853
rect 19009 18827 19069 18853
rect 18625 18678 18833 18686
rect 18625 18644 18641 18678
rect 18675 18644 18833 18678
rect 18625 18628 18833 18644
rect 18636 18627 18833 18628
rect 18249 18609 18399 18625
rect 18249 18575 18349 18609
rect 18383 18575 18399 18609
rect 18249 18559 18399 18575
rect 15561 18528 15621 18554
rect 15679 18528 15739 18554
rect 15797 18522 15857 18554
rect 15915 18528 15975 18554
rect 16033 18528 16093 18554
rect 16151 18534 16211 18554
rect 16150 18528 16211 18534
rect 16269 18528 16329 18554
rect 16387 18528 16447 18554
rect 16505 18528 16565 18554
rect 9710 18321 9770 18347
rect 8353 18294 8413 18320
rect 5681 18094 5741 18120
rect 5799 18094 5859 18120
rect 5917 18094 5977 18120
rect 6035 18094 6095 18120
rect 7579 18094 7639 18120
rect 7697 18094 7757 18120
rect 7815 18094 7875 18120
rect 7933 18094 7993 18120
rect 9357 18095 9417 18121
rect 11715 18290 11775 18316
rect 13013 18290 13073 18316
rect 13613 18290 13673 18316
rect 15794 18506 15860 18522
rect 15794 18472 15810 18506
rect 15844 18472 15860 18506
rect 15794 18456 15860 18472
rect 15912 18389 15978 18405
rect 15912 18355 15928 18389
rect 15962 18355 15978 18389
rect 15912 18339 15978 18355
rect 15915 18317 15975 18339
rect 16150 18317 16210 18528
rect 16270 18343 16328 18528
rect 18249 18521 18309 18559
rect 18773 18521 18833 18627
rect 19127 18686 19187 18853
rect 19245 18827 19305 18853
rect 19547 18820 19607 19478
rect 20132 19476 20207 19520
rect 20249 19476 20792 19527
rect 20850 19520 20910 19546
rect 20968 19520 21028 19546
rect 21086 19529 21146 19546
rect 21334 19529 21394 19546
rect 21452 19529 21512 19546
rect 21570 19529 21630 19546
rect 21086 19478 21630 19529
rect 24628 19766 24924 19817
rect 24628 19749 24688 19766
rect 24746 19749 24806 19766
rect 24864 19749 24924 19766
rect 25949 19749 26009 19775
rect 26067 19749 26127 19775
rect 26185 19749 26245 19775
rect 26526 19766 26822 19817
rect 26526 19749 26586 19766
rect 26644 19749 26704 19766
rect 26762 19749 26822 19766
rect 28957 19929 29017 19951
rect 29192 19929 29252 20140
rect 29312 19955 29370 20140
rect 29310 19929 29370 19955
rect 36701 20105 36740 20163
rect 37571 20105 37628 20514
rect 38569 20382 38620 20691
rect 36701 20045 36755 20105
rect 37155 20045 37628 20105
rect 37840 20322 38088 20382
rect 38288 20322 38620 20382
rect 36701 19987 36740 20045
rect 27847 19749 27907 19775
rect 27965 19749 28025 19775
rect 28083 19749 28143 19775
rect 28957 19703 29017 19729
rect 22679 19510 22739 19526
rect 19540 18804 19607 18820
rect 19540 18770 19557 18804
rect 19591 18770 19607 18804
rect 19540 18754 19607 18770
rect 19270 18686 19337 18693
rect 19127 18677 19337 18686
rect 19127 18643 19287 18677
rect 19321 18643 19337 18677
rect 19127 18627 19337 18643
rect 18887 18594 18953 18609
rect 18887 18560 18903 18594
rect 18937 18560 18953 18594
rect 18887 18544 18953 18560
rect 19005 18593 19071 18609
rect 19005 18559 19021 18593
rect 19055 18559 19071 18593
rect 18891 18521 18951 18544
rect 19005 18543 19071 18559
rect 19009 18521 19069 18543
rect 19127 18521 19187 18627
rect 19547 18626 19607 18754
rect 19456 18610 19607 18626
rect 19456 18576 19472 18610
rect 19506 18576 19607 18610
rect 19456 18560 19607 18576
rect 19547 18521 19607 18560
rect 20147 19356 20207 19476
rect 21445 19397 21505 19478
rect 22671 19488 22745 19510
rect 22797 19504 22857 19526
rect 24628 19523 24688 19549
rect 24746 19530 24806 19549
rect 24864 19530 24924 19549
rect 25111 19530 25171 19549
rect 25229 19530 25289 19549
rect 25347 19530 25407 19549
rect 24746 19523 24822 19530
rect 22671 19454 22692 19488
rect 22726 19454 22745 19488
rect 22671 19397 22745 19454
rect 22794 19488 22860 19504
rect 22794 19454 22810 19488
rect 22844 19454 22860 19488
rect 24747 19479 24822 19523
rect 24864 19479 25407 19530
rect 25465 19523 25525 19549
rect 25583 19523 25643 19549
rect 25701 19532 25761 19549
rect 25949 19532 26009 19549
rect 26067 19532 26127 19549
rect 26185 19532 26245 19549
rect 25701 19481 26245 19532
rect 26526 19523 26586 19549
rect 26644 19530 26704 19549
rect 26762 19530 26822 19549
rect 27009 19530 27069 19549
rect 27127 19530 27187 19549
rect 27245 19530 27305 19549
rect 26644 19523 26720 19530
rect 22794 19438 22860 19454
rect 21445 19372 22745 19397
rect 20147 19336 20208 19356
rect 20147 19320 20227 19336
rect 20147 19286 20178 19320
rect 20212 19286 20227 19320
rect 20147 19270 20227 19286
rect 20553 19277 20849 19337
rect 20147 19247 20208 19270
rect 20553 19253 20613 19277
rect 20671 19253 20731 19277
rect 20789 19253 20849 19277
rect 20907 19276 21203 19336
rect 20907 19253 20967 19276
rect 21025 19253 21085 19276
rect 21143 19253 21203 19276
rect 21445 19324 22746 19372
rect 24762 19326 24822 19479
rect 20147 19101 20207 19247
rect 20147 18928 20208 19101
rect 20147 18625 20207 18928
rect 20553 18827 20613 18853
rect 20521 18686 20588 18693
rect 20671 18686 20731 18853
rect 20789 18827 20849 18853
rect 20907 18827 20967 18853
rect 20521 18677 20731 18686
rect 20521 18643 20537 18677
rect 20571 18643 20731 18677
rect 20521 18627 20731 18643
rect 20147 18609 20297 18625
rect 20147 18575 20247 18609
rect 20281 18575 20297 18609
rect 20147 18559 20297 18575
rect 20147 18521 20207 18559
rect 20671 18521 20731 18627
rect 21025 18686 21085 18853
rect 21143 18827 21203 18853
rect 21168 18686 21235 18693
rect 21025 18677 21235 18686
rect 21025 18643 21185 18677
rect 21219 18643 21235 18677
rect 21025 18627 21235 18643
rect 20785 18594 20851 18609
rect 20785 18560 20801 18594
rect 20835 18560 20851 18594
rect 20785 18544 20851 18560
rect 20903 18593 20969 18609
rect 20903 18559 20919 18593
rect 20953 18559 20969 18593
rect 20789 18521 20849 18544
rect 20903 18543 20969 18559
rect 20907 18521 20967 18543
rect 21025 18521 21085 18627
rect 21445 18626 21505 19324
rect 24568 19302 24822 19326
rect 24568 19268 24584 19302
rect 24618 19268 24822 19302
rect 24568 19252 24822 19268
rect 25168 19280 25464 19340
rect 25168 19256 25228 19280
rect 25286 19256 25346 19280
rect 25404 19256 25464 19280
rect 25522 19279 25818 19339
rect 25522 19256 25582 19279
rect 25640 19256 25700 19279
rect 25758 19256 25818 19279
rect 22095 18779 22391 18815
rect 22095 18759 22155 18779
rect 22213 18759 22273 18779
rect 22331 18759 22391 18779
rect 22449 18779 22745 18815
rect 22449 18759 22509 18779
rect 22567 18759 22627 18779
rect 22685 18759 22745 18779
rect 22803 18780 23099 18816
rect 22803 18759 22863 18780
rect 22921 18759 22981 18780
rect 23039 18759 23099 18780
rect 21354 18610 21505 18626
rect 21354 18576 21370 18610
rect 21404 18576 21505 18610
rect 21354 18560 21505 18576
rect 21445 18521 21505 18560
rect 24762 18628 24822 19252
rect 25168 18830 25228 18856
rect 25138 18690 25205 18697
rect 25138 18689 25211 18690
rect 25286 18689 25346 18856
rect 25404 18830 25464 18856
rect 25522 18830 25582 18856
rect 25138 18681 25346 18689
rect 25138 18647 25154 18681
rect 25188 18647 25346 18681
rect 25138 18631 25346 18647
rect 25149 18630 25346 18631
rect 24762 18612 24912 18628
rect 24762 18578 24862 18612
rect 24896 18578 24912 18612
rect 24762 18562 24912 18578
rect 22095 18533 22155 18559
rect 22213 18533 22273 18559
rect 22331 18527 22391 18559
rect 22449 18533 22509 18559
rect 22567 18533 22627 18559
rect 22685 18539 22745 18559
rect 22684 18533 22745 18539
rect 22803 18533 22863 18559
rect 22921 18533 22981 18559
rect 23039 18533 23099 18559
rect 16268 18317 16328 18343
rect 14911 18290 14971 18316
rect 12239 18090 12299 18116
rect 12357 18090 12417 18116
rect 12475 18090 12535 18116
rect 12593 18090 12653 18116
rect 14137 18090 14197 18116
rect 14255 18090 14315 18116
rect 14373 18090 14433 18116
rect 14491 18090 14551 18116
rect 15915 18091 15975 18117
rect 9592 17899 9652 17921
rect 9710 17899 9770 17921
rect 9589 17883 9655 17899
rect 9589 17849 9605 17883
rect 9639 17849 9655 17883
rect 9589 17833 9655 17849
rect 9707 17883 9773 17899
rect 9707 17849 9723 17883
rect 9757 17849 9773 17883
rect 18249 18295 18309 18321
rect 19547 18295 19607 18321
rect 20147 18295 20207 18321
rect 22328 18511 22394 18527
rect 22328 18477 22344 18511
rect 22378 18477 22394 18511
rect 22328 18461 22394 18477
rect 22446 18394 22512 18410
rect 22446 18360 22462 18394
rect 22496 18360 22512 18394
rect 22446 18344 22512 18360
rect 22449 18322 22509 18344
rect 22684 18322 22744 18533
rect 22804 18348 22862 18533
rect 24762 18524 24822 18562
rect 25286 18524 25346 18630
rect 25640 18689 25700 18856
rect 25758 18830 25818 18856
rect 26060 18823 26120 19481
rect 26645 19479 26720 19523
rect 26762 19479 27305 19530
rect 27363 19523 27423 19549
rect 27481 19523 27541 19549
rect 27599 19532 27659 19549
rect 27847 19532 27907 19549
rect 27965 19532 28025 19549
rect 28083 19532 28143 19549
rect 27599 19481 28143 19532
rect 36701 19927 36755 19987
rect 37155 19927 37181 19987
rect 36900 19690 36955 19750
rect 37155 19690 37181 19750
rect 36900 19632 36939 19690
rect 36900 19572 36955 19632
rect 37155 19572 37181 19632
rect 37301 19608 37367 19624
rect 37301 19574 37317 19608
rect 37351 19574 37367 19608
rect 29192 19513 29252 19529
rect 26053 18807 26120 18823
rect 26053 18773 26070 18807
rect 26104 18773 26120 18807
rect 26053 18757 26120 18773
rect 25783 18689 25850 18696
rect 25640 18680 25850 18689
rect 25640 18646 25800 18680
rect 25834 18646 25850 18680
rect 25640 18630 25850 18646
rect 25400 18597 25466 18612
rect 25400 18563 25416 18597
rect 25450 18563 25466 18597
rect 25400 18547 25466 18563
rect 25518 18596 25584 18612
rect 25518 18562 25534 18596
rect 25568 18562 25584 18596
rect 25404 18524 25464 18547
rect 25518 18546 25584 18562
rect 25522 18524 25582 18546
rect 25640 18524 25700 18630
rect 26060 18629 26120 18757
rect 25969 18613 26120 18629
rect 25969 18579 25985 18613
rect 26019 18579 26120 18613
rect 25969 18563 26120 18579
rect 26060 18524 26120 18563
rect 26660 19359 26720 19479
rect 27958 19400 28018 19481
rect 29184 19491 29258 19513
rect 29310 19507 29370 19529
rect 36900 19514 36939 19572
rect 37301 19558 37367 19574
rect 37304 19514 37364 19558
rect 37840 19514 37885 20322
rect 29184 19457 29205 19491
rect 29239 19457 29258 19491
rect 29184 19400 29258 19457
rect 29307 19491 29373 19507
rect 29307 19457 29323 19491
rect 29357 19457 29373 19491
rect 29307 19441 29373 19457
rect 36900 19454 36955 19514
rect 37155 19454 37885 19514
rect 27958 19375 29258 19400
rect 26660 19339 26721 19359
rect 26660 19323 26740 19339
rect 26660 19289 26691 19323
rect 26725 19289 26740 19323
rect 26660 19273 26740 19289
rect 27066 19280 27362 19340
rect 26660 19250 26721 19273
rect 27066 19256 27126 19280
rect 27184 19256 27244 19280
rect 27302 19256 27362 19280
rect 27420 19279 27716 19339
rect 27420 19256 27480 19279
rect 27538 19256 27598 19279
rect 27656 19256 27716 19279
rect 27958 19327 29259 19375
rect 26660 19104 26720 19250
rect 26660 18931 26721 19104
rect 26660 18628 26720 18931
rect 27066 18830 27126 18856
rect 27034 18689 27101 18696
rect 27184 18689 27244 18856
rect 27302 18830 27362 18856
rect 27420 18830 27480 18856
rect 27034 18680 27244 18689
rect 27034 18646 27050 18680
rect 27084 18646 27244 18680
rect 27034 18630 27244 18646
rect 26660 18612 26810 18628
rect 26660 18578 26760 18612
rect 26794 18578 26810 18612
rect 26660 18562 26810 18578
rect 26660 18524 26720 18562
rect 27184 18524 27244 18630
rect 27538 18689 27598 18856
rect 27656 18830 27716 18856
rect 27681 18689 27748 18696
rect 27538 18680 27748 18689
rect 27538 18646 27698 18680
rect 27732 18646 27748 18680
rect 27538 18630 27748 18646
rect 27298 18597 27364 18612
rect 27298 18563 27314 18597
rect 27348 18563 27364 18597
rect 27298 18547 27364 18563
rect 27416 18596 27482 18612
rect 27416 18562 27432 18596
rect 27466 18562 27482 18596
rect 27302 18524 27362 18547
rect 27416 18546 27482 18562
rect 27420 18524 27480 18546
rect 27538 18524 27598 18630
rect 27958 18629 28018 19327
rect 28608 18782 28904 18818
rect 28608 18762 28668 18782
rect 28726 18762 28786 18782
rect 28844 18762 28904 18782
rect 28962 18782 29258 18818
rect 28962 18762 29022 18782
rect 29080 18762 29140 18782
rect 29198 18762 29258 18782
rect 29316 18783 29612 18819
rect 29316 18762 29376 18783
rect 29434 18762 29494 18783
rect 29552 18762 29612 18783
rect 36896 18766 36951 18826
rect 37151 18767 37881 18826
rect 37151 18766 37454 18767
rect 27867 18613 28018 18629
rect 27867 18579 27883 18613
rect 27917 18579 28018 18613
rect 27867 18563 28018 18579
rect 27958 18524 28018 18563
rect 36896 18708 36935 18766
rect 37437 18709 37454 18766
rect 37509 18766 37881 18767
rect 37509 18709 37524 18766
rect 36896 18648 36951 18708
rect 37151 18648 37177 18708
rect 37437 18690 37524 18709
rect 36896 18590 36935 18648
rect 28608 18536 28668 18562
rect 28726 18536 28786 18562
rect 28844 18530 28904 18562
rect 28962 18536 29022 18562
rect 29080 18536 29140 18562
rect 29198 18542 29258 18562
rect 29197 18536 29258 18542
rect 29316 18536 29376 18562
rect 29434 18536 29494 18562
rect 29552 18536 29612 18562
rect 22802 18322 22862 18348
rect 21445 18295 21505 18321
rect 18773 18095 18833 18121
rect 18891 18095 18951 18121
rect 19009 18095 19069 18121
rect 19127 18095 19187 18121
rect 20671 18095 20731 18121
rect 20789 18095 20849 18121
rect 20907 18095 20967 18121
rect 21025 18095 21085 18121
rect 22449 18096 22509 18122
rect 16150 17895 16210 17917
rect 16268 17895 16328 17917
rect 9707 17833 9773 17849
rect 16147 17879 16213 17895
rect 16147 17845 16163 17879
rect 16197 17845 16213 17879
rect 16147 17829 16213 17845
rect 16265 17879 16331 17895
rect 16265 17845 16281 17879
rect 16315 17845 16331 17879
rect 24762 18298 24822 18324
rect 26060 18298 26120 18324
rect 26660 18298 26720 18324
rect 28841 18514 28907 18530
rect 28841 18480 28857 18514
rect 28891 18480 28907 18514
rect 28841 18464 28907 18480
rect 28959 18397 29025 18413
rect 28959 18363 28975 18397
rect 29009 18363 29025 18397
rect 28959 18347 29025 18363
rect 28962 18325 29022 18347
rect 29197 18325 29257 18536
rect 29317 18351 29375 18536
rect 36896 18530 36951 18590
rect 37151 18530 37177 18590
rect 29315 18325 29375 18351
rect 36697 18325 36751 18385
rect 37151 18325 37177 18385
rect 27958 18298 28018 18324
rect 25286 18098 25346 18124
rect 25404 18098 25464 18124
rect 25522 18098 25582 18124
rect 25640 18098 25700 18124
rect 27184 18098 27244 18124
rect 27302 18098 27362 18124
rect 27420 18098 27480 18124
rect 27538 18098 27598 18124
rect 28962 18099 29022 18125
rect 22684 17900 22744 17922
rect 22802 17900 22862 17922
rect 16265 17829 16331 17845
rect 22681 17884 22747 17900
rect 22681 17850 22697 17884
rect 22731 17850 22747 17884
rect 22681 17834 22747 17850
rect 22799 17884 22865 17900
rect 22799 17850 22815 17884
rect 22849 17850 22865 17884
rect 36697 18267 36736 18325
rect 36697 18207 36751 18267
rect 37151 18207 37626 18267
rect 36697 18149 36736 18207
rect 36697 18089 36751 18149
rect 37151 18089 37177 18149
rect 29197 17903 29257 17925
rect 29315 17903 29375 17925
rect 22799 17834 22865 17850
rect 29194 17887 29260 17903
rect 29194 17853 29210 17887
rect 29244 17853 29260 17887
rect 29194 17837 29260 17853
rect 29312 17887 29378 17903
rect 29312 17853 29328 17887
rect 29362 17853 29378 17887
rect 29312 17837 29378 17853
rect 36697 17858 36751 17918
rect 37151 17858 37177 17918
rect 36697 17800 36736 17858
rect 36697 17740 36751 17800
rect 37151 17799 37177 17800
rect 37338 17799 37404 17802
rect 37151 17786 37404 17799
rect 37151 17752 37354 17786
rect 37388 17752 37404 17786
rect 37151 17740 37404 17752
rect 37569 17800 37626 18207
rect 37836 17992 37881 18766
rect 37836 17932 38084 17992
rect 38284 17932 38310 17992
rect 37725 17800 37804 17811
rect 37569 17798 38084 17800
rect 37569 17740 37738 17798
rect 37793 17740 38084 17798
rect 38484 17740 38510 17800
rect 36697 17682 36736 17740
rect 37337 17736 37404 17740
rect 37725 17730 37804 17740
rect 37438 17682 37525 17699
rect 36697 17622 36751 17682
rect 37151 17622 37177 17682
rect 37438 17680 38084 17682
rect 37438 17622 37453 17680
rect 37508 17622 38084 17680
rect 38484 17622 38510 17682
rect 37438 17604 37525 17622
rect 36697 17504 36751 17564
rect 37151 17504 37177 17564
rect 36697 17446 36736 17504
rect 37476 17446 37525 17604
rect 37958 17564 38024 17567
rect 38557 17609 38623 17625
rect 38557 17575 38573 17609
rect 38607 17575 38623 17609
rect 37958 17551 38084 17564
rect 37958 17517 37974 17551
rect 38008 17517 38084 17551
rect 37958 17504 38084 17517
rect 38484 17504 38510 17564
rect 38557 17559 38623 17575
rect 37958 17501 38024 17504
rect 36697 17386 36751 17446
rect 37151 17386 37525 17446
rect 37567 17446 37636 17451
rect 37567 17432 38084 17446
rect 37567 17398 37584 17432
rect 37618 17398 38084 17432
rect 37567 17386 38084 17398
rect 38484 17386 38510 17446
rect 36697 17328 36736 17386
rect 37567 17382 37634 17386
rect 36697 17268 36751 17328
rect 37151 17268 37177 17328
rect 36697 17031 36751 17091
rect 37151 17031 37177 17091
rect 36697 16973 36736 17031
rect 37567 16973 37624 17382
rect 38565 17250 38616 17559
rect 36697 16913 36751 16973
rect 37151 16913 37624 16973
rect 37836 17190 38084 17250
rect 38284 17190 38616 17250
rect 36697 16855 36736 16913
rect 36697 16795 36751 16855
rect 37151 16795 37177 16855
rect 36896 16558 36951 16618
rect 37151 16558 37177 16618
rect 36896 16500 36935 16558
rect 36896 16440 36951 16500
rect 37151 16440 37177 16500
rect 37297 16476 37363 16492
rect 37297 16442 37313 16476
rect 37347 16442 37363 16476
rect 36896 16382 36935 16440
rect 37297 16426 37363 16442
rect 37300 16382 37360 16426
rect 37836 16382 37881 17190
rect 36896 16322 36951 16382
rect 37151 16322 37881 16382
rect -3057 16232 -2997 16248
rect -3630 16149 -3604 16209
rect -3404 16149 -3336 16209
rect -3387 16091 -3336 16149
rect -3630 16031 -3604 16091
rect -3404 16084 -3336 16091
rect -3057 16198 -3043 16232
rect -3009 16198 -2997 16232
rect -3057 16084 -2997 16198
rect -3404 16031 -2379 16084
rect -3387 16024 -2379 16031
rect -2179 16024 -2153 16084
rect -3387 15973 -3336 16024
rect -3630 15913 -3604 15973
rect -3404 15913 -3336 15973
rect -2484 15983 -2418 16024
rect -2484 15949 -2468 15983
rect -2434 15949 -2418 15983
rect -2484 15933 -2418 15949
rect -3387 15725 -3336 15913
rect -2551 15798 -2485 15814
rect -3870 15665 -3804 15725
rect -3404 15665 -3336 15725
rect -3194 15722 -3111 15782
rect -2711 15722 -2685 15782
rect -2551 15764 -2535 15798
rect -2501 15764 -2485 15798
rect -2551 15747 -2485 15764
rect -3870 15607 -3819 15665
rect -3194 15664 -3134 15722
rect -2544 15664 -2485 15747
rect -3870 15547 -3804 15607
rect -3404 15547 -3378 15607
rect -3194 15604 -3111 15664
rect -2711 15604 -2379 15664
rect -1979 15604 -1953 15664
rect 36896 15622 36951 15682
rect 37151 15623 37881 15682
rect 37151 15622 37454 15623
rect -3870 15489 -3819 15547
rect -3194 15546 -3134 15604
rect -2467 15546 -2401 15548
rect -3870 15429 -3804 15489
rect -3404 15429 -3378 15489
rect -3194 15486 -3111 15546
rect -2711 15486 -2685 15546
rect -2467 15532 -2379 15546
rect -2467 15498 -2451 15532
rect -2417 15498 -2379 15532
rect -2467 15486 -2379 15498
rect -1979 15486 -1953 15546
rect 36896 15564 36935 15622
rect 37437 15565 37454 15622
rect 37509 15622 37881 15623
rect 37509 15565 37524 15622
rect -2467 15482 -2401 15486
rect -2467 15428 -2402 15430
rect -3830 15311 -3804 15371
rect -3404 15311 -3334 15371
rect -3385 15253 -3334 15311
rect -3830 15193 -3804 15253
rect -3404 15193 -3334 15253
rect -3385 15135 -3334 15193
rect -3830 15075 -3804 15135
rect -3404 15075 -3334 15135
rect -3195 15368 -3111 15428
rect -2711 15368 -2685 15428
rect -2467 15414 -2379 15428
rect -2467 15380 -2452 15414
rect -2418 15380 -2379 15414
rect -2467 15368 -2379 15380
rect -1979 15368 -1953 15428
rect -3195 15310 -3135 15368
rect -2467 15364 -2402 15368
rect 36896 15504 36951 15564
rect 37151 15504 37177 15564
rect 37437 15546 37524 15565
rect 36896 15446 36935 15504
rect 36896 15386 36951 15446
rect 37151 15386 37177 15446
rect -3195 15250 -3111 15310
rect -2711 15250 -2379 15310
rect -1979 15250 -1953 15310
rect 7858 15257 8154 15293
rect -3195 15192 -3135 15250
rect -3195 15132 -3111 15192
rect -2711 15132 -2685 15192
rect -2544 15167 -2485 15250
rect 7858 15236 7918 15257
rect 7976 15236 8036 15257
rect 8094 15236 8154 15257
rect 8212 15256 8508 15292
rect 8212 15236 8272 15256
rect 8330 15236 8390 15256
rect 8448 15236 8508 15256
rect 8566 15256 8862 15292
rect 8566 15236 8626 15256
rect 8684 15236 8744 15256
rect 8802 15236 8862 15256
rect 14407 15256 14703 15292
rect -2551 15150 -2485 15167
rect -3385 14888 -3334 15075
rect -2551 15116 -2535 15150
rect -2501 15116 -2485 15150
rect -2551 15100 -2485 15116
rect 14407 15235 14467 15256
rect 14525 15235 14585 15256
rect 14643 15235 14703 15256
rect 14761 15255 15057 15291
rect 14761 15235 14821 15255
rect 14879 15235 14939 15255
rect 14997 15235 15057 15255
rect 15115 15255 15411 15291
rect 21061 15277 21357 15313
rect 21061 15256 21121 15277
rect 21179 15256 21239 15277
rect 21297 15256 21357 15277
rect 21415 15276 21711 15312
rect 21415 15256 21475 15276
rect 21533 15256 21593 15276
rect 21651 15256 21711 15276
rect 21769 15276 22065 15312
rect 21769 15256 21829 15276
rect 21887 15256 21947 15276
rect 22005 15256 22065 15276
rect 15115 15235 15175 15255
rect 15233 15235 15293 15255
rect 15351 15235 15411 15255
rect 7858 15010 7918 15036
rect 7976 15010 8036 15036
rect 8094 15010 8154 15036
rect 8212 15016 8272 15036
rect 8212 15010 8273 15016
rect 8330 15010 8390 15036
rect 8448 15010 8508 15036
rect -3672 14828 -3604 14888
rect -3404 14828 -3334 14888
rect -2483 14860 -2417 14876
rect -3247 14838 -3193 14854
rect -3672 14770 -3621 14828
rect -3247 14804 -3237 14838
rect -3203 14804 -3193 14838
rect -3247 14786 -3193 14804
rect -2483 14826 -2467 14860
rect -2433 14826 -2417 14860
rect -2483 14786 -2417 14826
rect 8095 14825 8153 15010
rect 8095 14799 8155 14825
rect 8213 14799 8273 15010
rect 8566 15004 8626 15036
rect 8684 15010 8744 15036
rect 8802 15010 8862 15036
rect 36697 15181 36751 15241
rect 37151 15181 37177 15241
rect 29714 15110 30010 15146
rect 29714 15089 29774 15110
rect 29832 15089 29892 15110
rect 29950 15089 30010 15110
rect 30068 15109 30364 15145
rect 30068 15089 30128 15109
rect 30186 15089 30246 15109
rect 30304 15089 30364 15109
rect 30422 15109 30718 15145
rect 30422 15089 30482 15109
rect 30540 15089 30600 15109
rect 30658 15089 30718 15109
rect 36697 15123 36736 15181
rect 14407 15009 14467 15035
rect 14525 15009 14585 15035
rect 14643 15009 14703 15035
rect 14761 15015 14821 15035
rect 14761 15009 14822 15015
rect 14879 15009 14939 15035
rect 14997 15009 15057 15035
rect 8563 14988 8629 15004
rect 8563 14954 8579 14988
rect 8613 14954 8629 14988
rect 8563 14938 8629 14954
rect 8445 14871 8511 14887
rect 8445 14837 8461 14871
rect 8495 14837 8511 14871
rect 8445 14821 8511 14837
rect 14644 14824 14702 15009
rect 8448 14799 8508 14821
rect -3385 14770 -2379 14786
rect -3672 14710 -3604 14770
rect -3404 14726 -2379 14770
rect -2179 14726 -2153 14786
rect -3404 14711 -3334 14726
rect -3404 14710 -3378 14711
rect -3672 14652 -3621 14710
rect -3672 14592 -3604 14652
rect -3404 14592 -3378 14652
rect 14644 14798 14704 14824
rect 14762 14798 14822 15009
rect 15115 15003 15175 15035
rect 15233 15009 15293 15035
rect 15351 15009 15411 15035
rect 21061 15030 21121 15056
rect 21179 15030 21239 15056
rect 21297 15030 21357 15056
rect 21415 15036 21475 15056
rect 21415 15030 21476 15036
rect 21533 15030 21593 15056
rect 21651 15030 21711 15056
rect 15112 14987 15178 15003
rect 15112 14953 15128 14987
rect 15162 14953 15178 14987
rect 15112 14937 15178 14953
rect 14994 14870 15060 14886
rect 14994 14836 15010 14870
rect 15044 14836 15060 14870
rect 14994 14820 15060 14836
rect 21298 14845 21356 15030
rect 14997 14798 15057 14820
rect 21298 14819 21358 14845
rect 21416 14819 21476 15030
rect 21769 15024 21829 15056
rect 21887 15030 21947 15056
rect 22005 15030 22065 15056
rect 21766 15008 21832 15024
rect 21766 14974 21782 15008
rect 21816 14974 21832 15008
rect 21766 14958 21832 14974
rect 21648 14891 21714 14907
rect 21648 14857 21664 14891
rect 21698 14857 21714 14891
rect 36697 15063 36751 15123
rect 37151 15063 37626 15123
rect 36697 15005 36736 15063
rect 32006 14899 32302 14950
rect 29714 14863 29774 14889
rect 29832 14863 29892 14889
rect 29950 14863 30010 14889
rect 30068 14869 30128 14889
rect 30068 14863 30129 14869
rect 30186 14863 30246 14889
rect 30304 14863 30364 14889
rect 21648 14841 21714 14857
rect 21651 14819 21711 14841
rect 8448 14573 8508 14599
rect 8095 14377 8155 14399
rect 8213 14377 8273 14399
rect 14997 14572 15057 14598
rect 29951 14678 30009 14863
rect 29951 14652 30011 14678
rect 30069 14652 30129 14863
rect 30422 14857 30482 14889
rect 30540 14863 30600 14889
rect 30658 14863 30718 14889
rect 32006 14884 32066 14899
rect 32124 14884 32184 14899
rect 32242 14884 32302 14899
rect 32360 14884 32420 14910
rect 32478 14884 32538 14910
rect 32596 14884 32656 14910
rect 36697 14945 36751 15005
rect 37151 14945 37177 15005
rect 30419 14841 30485 14857
rect 30419 14807 30435 14841
rect 30469 14807 30485 14841
rect 30419 14791 30485 14807
rect 30301 14724 30367 14740
rect 30301 14690 30317 14724
rect 30351 14690 30367 14724
rect 30301 14674 30367 14690
rect 31522 14684 31582 14710
rect 31640 14684 31700 14710
rect 31758 14684 31818 14710
rect 30304 14652 30364 14674
rect 21651 14593 21711 14619
rect 8092 14361 8158 14377
rect 8092 14327 8108 14361
rect 8142 14327 8158 14361
rect 8092 14311 8158 14327
rect 8210 14361 8276 14377
rect 14644 14376 14704 14398
rect 14762 14376 14822 14398
rect 21298 14397 21358 14419
rect 21416 14397 21476 14419
rect 21295 14381 21361 14397
rect 8210 14327 8226 14361
rect 8260 14327 8276 14361
rect 8210 14311 8276 14327
rect 14641 14360 14707 14376
rect 14641 14326 14657 14360
rect 14691 14326 14707 14360
rect 14641 14310 14707 14326
rect 14759 14360 14825 14376
rect 14759 14326 14775 14360
rect 14809 14326 14825 14360
rect 21295 14347 21311 14381
rect 21345 14347 21361 14381
rect 21295 14331 21361 14347
rect 21413 14381 21479 14397
rect 21413 14347 21429 14381
rect 21463 14347 21479 14381
rect 21413 14331 21479 14347
rect 14759 14310 14825 14326
rect -3059 14164 -2999 14180
rect 32843 14701 33139 14752
rect 32843 14684 32903 14701
rect 32961 14684 33021 14701
rect 33079 14684 33139 14701
rect 33315 14702 33611 14738
rect 33315 14681 33375 14702
rect 33433 14681 33493 14702
rect 33551 14681 33611 14702
rect 33669 14701 33965 14737
rect 33669 14681 33729 14701
rect 33787 14681 33847 14701
rect 33905 14681 33965 14701
rect 34023 14701 34319 14737
rect 34023 14681 34083 14701
rect 34141 14681 34201 14701
rect 34259 14681 34319 14701
rect 36697 14714 36751 14774
rect 37151 14714 37177 14774
rect 31522 14467 31582 14484
rect 31640 14467 31700 14484
rect 31758 14467 31818 14484
rect 32006 14467 32066 14484
rect 30304 14426 30364 14452
rect 31522 14416 32066 14467
rect 32124 14458 32184 14484
rect 32242 14458 32302 14484
rect 32360 14465 32420 14484
rect 32478 14465 32538 14484
rect 32596 14465 32656 14484
rect 32843 14465 32903 14484
rect 32961 14465 33021 14484
rect 29951 14230 30011 14252
rect 30069 14230 30129 14252
rect 29948 14214 30014 14230
rect 29948 14180 29964 14214
rect 29998 14180 30014 14214
rect 29948 14164 30014 14180
rect 30066 14214 30132 14230
rect 30066 14180 30082 14214
rect 30116 14180 30132 14214
rect 30066 14164 30132 14180
rect 31647 14212 31707 14416
rect 32360 14414 32903 14465
rect 32945 14458 33021 14465
rect 33079 14458 33139 14484
rect 36697 14656 36736 14714
rect 36697 14596 36751 14656
rect 37151 14655 37177 14656
rect 37338 14655 37404 14658
rect 37151 14642 37404 14655
rect 37151 14608 37354 14642
rect 37388 14608 37404 14642
rect 37151 14596 37404 14608
rect 37569 14656 37626 15063
rect 37836 14848 37881 15622
rect 37836 14788 38084 14848
rect 38284 14788 38310 14848
rect 37725 14656 37804 14667
rect 37569 14654 38084 14656
rect 37569 14596 37738 14654
rect 37793 14596 38084 14654
rect 38484 14596 38510 14656
rect 32945 14414 33020 14458
rect 33315 14455 33375 14481
rect 33433 14455 33493 14481
rect 33551 14455 33611 14481
rect 33669 14461 33729 14481
rect 33669 14455 33730 14461
rect 33787 14455 33847 14481
rect 33905 14455 33965 14481
rect 32945 14332 33005 14414
rect 32945 14314 33179 14332
rect 32945 14280 33128 14314
rect 33162 14280 33179 14314
rect 31949 14214 32245 14274
rect 31647 14195 31778 14212
rect -3632 14081 -3606 14141
rect -3406 14081 -3338 14141
rect -3389 14023 -3338 14081
rect -3632 13963 -3606 14023
rect -3406 14016 -3338 14023
rect -3059 14130 -3045 14164
rect -3011 14130 -2999 14164
rect 31647 14161 31728 14195
rect 31762 14161 31778 14195
rect 31949 14191 32009 14214
rect 32067 14191 32127 14214
rect 32185 14191 32245 14214
rect 32303 14215 32599 14275
rect 32303 14191 32363 14215
rect 32421 14191 32481 14215
rect 32539 14191 32599 14215
rect 32945 14264 33179 14280
rect 33552 14270 33610 14455
rect 31647 14144 31778 14161
rect -3059 14016 -2999 14130
rect -3406 13963 -2381 14016
rect -3389 13956 -2381 13963
rect -2181 13956 -2155 14016
rect -3389 13905 -3338 13956
rect -3632 13845 -3606 13905
rect -3406 13845 -3338 13905
rect -2486 13915 -2420 13956
rect -2486 13881 -2470 13915
rect -2436 13881 -2420 13915
rect -2486 13865 -2420 13881
rect -3389 13657 -3338 13845
rect -2553 13730 -2487 13746
rect -3872 13597 -3806 13657
rect -3406 13597 -3338 13657
rect -3196 13654 -3113 13714
rect -2713 13654 -2687 13714
rect -2553 13696 -2537 13730
rect -2503 13696 -2487 13730
rect -2553 13679 -2487 13696
rect -3872 13539 -3821 13597
rect -3196 13596 -3136 13654
rect -2546 13596 -2487 13679
rect -3872 13479 -3806 13539
rect -3406 13479 -3380 13539
rect -3196 13536 -3113 13596
rect -2713 13536 -2381 13596
rect -1981 13536 -1955 13596
rect -3872 13421 -3821 13479
rect -3196 13478 -3136 13536
rect -2469 13478 -2403 13480
rect -3872 13361 -3806 13421
rect -3406 13361 -3380 13421
rect -3196 13418 -3113 13478
rect -2713 13418 -2687 13478
rect -2469 13464 -2381 13478
rect -2469 13430 -2453 13464
rect -2419 13430 -2381 13464
rect -2469 13418 -2381 13430
rect -1981 13418 -1955 13478
rect -2469 13414 -2403 13418
rect -2469 13360 -2404 13362
rect -3832 13243 -3806 13303
rect -3406 13243 -3336 13303
rect -3387 13185 -3336 13243
rect -3832 13125 -3806 13185
rect -3406 13125 -3336 13185
rect -3387 13067 -3336 13125
rect -3832 13007 -3806 13067
rect -3406 13007 -3336 13067
rect -3197 13300 -3113 13360
rect -2713 13300 -2687 13360
rect -2469 13346 -2381 13360
rect -2469 13312 -2454 13346
rect -2420 13312 -2381 13346
rect -2469 13300 -2381 13312
rect -1981 13300 -1955 13360
rect 1194 13357 1490 13393
rect 1194 13336 1254 13357
rect 1312 13336 1372 13357
rect 1430 13336 1490 13357
rect 1548 13356 1844 13392
rect 1548 13336 1608 13356
rect 1666 13336 1726 13356
rect 1784 13336 1844 13356
rect 1902 13356 2198 13392
rect 1902 13336 1962 13356
rect 2020 13336 2080 13356
rect 2138 13336 2198 13356
rect -3197 13242 -3137 13300
rect -2469 13296 -2404 13300
rect -3197 13182 -3113 13242
rect -2713 13182 -2381 13242
rect -1981 13182 -1955 13242
rect -3197 13124 -3137 13182
rect -3197 13064 -3113 13124
rect -2713 13064 -2687 13124
rect -2546 13099 -2487 13182
rect 6232 13305 6298 13321
rect 7362 13311 7428 13327
rect 6232 13271 6248 13305
rect 6282 13298 6298 13305
rect 6282 13271 6807 13298
rect 6232 13255 6807 13271
rect 7362 13277 7378 13311
rect 7412 13302 7428 13311
rect 12781 13393 12847 13409
rect 13911 13399 13977 13415
rect 12781 13359 12797 13393
rect 12831 13386 12847 13393
rect 12831 13359 13356 13386
rect 12781 13343 13356 13359
rect 13911 13365 13927 13399
rect 13961 13390 13977 13399
rect 13961 13365 14498 13390
rect 13911 13347 14498 13365
rect 7412 13277 7949 13302
rect 13312 13291 13356 13343
rect 14454 13295 14498 13347
rect 7362 13259 7949 13277
rect 6763 13203 6807 13255
rect 7905 13207 7949 13259
rect 12781 13275 13254 13291
rect 12781 13241 12797 13275
rect 12831 13250 13254 13275
rect 12831 13249 13018 13250
rect 12831 13241 12847 13249
rect 12781 13225 12847 13241
rect 12958 13229 13018 13249
rect 13076 13229 13136 13250
rect 13194 13229 13254 13250
rect 13312 13250 13608 13291
rect 13312 13229 13372 13250
rect 13430 13229 13490 13250
rect 13548 13229 13608 13250
rect 13911 13279 14396 13295
rect 13911 13245 13927 13279
rect 13961 13254 14396 13279
rect 13961 13253 14160 13254
rect 13961 13245 13977 13253
rect 13911 13229 13977 13245
rect 14100 13233 14160 13253
rect 14218 13233 14278 13254
rect 14336 13233 14396 13254
rect 14454 13254 14750 13295
rect 19435 13325 19501 13341
rect 20565 13331 20631 13347
rect 19435 13291 19451 13325
rect 19485 13318 19501 13325
rect 19485 13291 20010 13318
rect 19435 13275 20010 13291
rect 20565 13297 20581 13331
rect 20615 13322 20631 13331
rect 26060 13393 26126 13409
rect 27190 13399 27256 13415
rect 26060 13359 26076 13393
rect 26110 13386 26126 13393
rect 26110 13359 26635 13386
rect 26060 13343 26635 13359
rect 27190 13365 27206 13399
rect 27240 13390 27256 13399
rect 31647 13564 31707 14144
rect 31949 13765 32009 13791
rect 31917 13624 31984 13631
rect 32067 13624 32127 13791
rect 32185 13765 32245 13791
rect 32303 13765 32363 13791
rect 31917 13615 32127 13624
rect 31917 13581 31933 13615
rect 31967 13581 32127 13615
rect 31917 13565 32127 13581
rect 31647 13548 31798 13564
rect 31647 13514 31748 13548
rect 31782 13514 31798 13548
rect 31647 13498 31798 13514
rect 31647 13459 31707 13498
rect 32067 13459 32127 13565
rect 32421 13624 32481 13791
rect 32539 13765 32599 13791
rect 32564 13624 32631 13631
rect 32421 13615 32631 13624
rect 32421 13581 32581 13615
rect 32615 13581 32631 13615
rect 32421 13565 32631 13581
rect 32183 13531 32249 13547
rect 32183 13497 32199 13531
rect 32233 13497 32249 13531
rect 32183 13481 32249 13497
rect 32301 13532 32367 13547
rect 32301 13498 32317 13532
rect 32351 13498 32367 13532
rect 32301 13482 32367 13498
rect 32185 13459 32245 13481
rect 32303 13459 32363 13482
rect 32421 13459 32481 13565
rect 32945 13563 33005 14264
rect 33552 14244 33612 14270
rect 33670 14244 33730 14455
rect 34023 14449 34083 14481
rect 34141 14455 34201 14481
rect 34259 14455 34319 14481
rect 34020 14433 34086 14449
rect 34020 14399 34036 14433
rect 34070 14399 34086 14433
rect 34020 14383 34086 14399
rect 36697 14538 36736 14596
rect 37337 14592 37404 14596
rect 37725 14586 37804 14596
rect 37438 14538 37525 14555
rect 36697 14478 36751 14538
rect 37151 14478 37177 14538
rect 37438 14536 38084 14538
rect 37438 14478 37453 14536
rect 37508 14478 38084 14536
rect 38484 14478 38510 14538
rect 37438 14460 37525 14478
rect 33902 14316 33968 14332
rect 33902 14282 33918 14316
rect 33952 14282 33968 14316
rect 36697 14360 36751 14420
rect 37151 14360 37177 14420
rect 36697 14302 36736 14360
rect 37476 14302 37525 14460
rect 37958 14420 38024 14423
rect 38557 14465 38623 14481
rect 38557 14431 38573 14465
rect 38607 14431 38623 14465
rect 37958 14407 38084 14420
rect 37958 14373 37974 14407
rect 38008 14373 38084 14407
rect 37958 14360 38084 14373
rect 38484 14360 38510 14420
rect 38557 14415 38623 14431
rect 37958 14357 38024 14360
rect 33902 14266 33968 14282
rect 33905 14244 33965 14266
rect 36697 14242 36751 14302
rect 37151 14242 37525 14302
rect 37567 14302 37636 14307
rect 37567 14288 38084 14302
rect 37567 14254 37584 14288
rect 37618 14254 38084 14288
rect 37567 14242 38084 14254
rect 38484 14242 38510 14302
rect 36697 14184 36736 14242
rect 37567 14238 37634 14242
rect 36697 14124 36751 14184
rect 37151 14124 37177 14184
rect 33905 14018 33965 14044
rect 36697 13887 36751 13947
rect 37151 13887 37177 13947
rect 33552 13822 33612 13844
rect 33670 13822 33730 13844
rect 36697 13829 36736 13887
rect 37567 13829 37624 14238
rect 38565 14106 38616 14415
rect 33549 13806 33615 13822
rect 33549 13772 33565 13806
rect 33599 13772 33615 13806
rect 33549 13756 33615 13772
rect 33667 13806 33733 13822
rect 33667 13772 33683 13806
rect 33717 13772 33733 13806
rect 33667 13756 33733 13772
rect 36697 13769 36751 13829
rect 37151 13769 37624 13829
rect 37836 14046 38084 14106
rect 38284 14046 38616 14106
rect 36697 13711 36736 13769
rect 36697 13651 36751 13711
rect 37151 13651 37177 13711
rect 32855 13547 33005 13563
rect 32855 13513 32871 13547
rect 32905 13513 33005 13547
rect 32855 13497 33005 13513
rect 32945 13459 33005 13497
rect 27240 13365 27777 13390
rect 27190 13347 27777 13365
rect 20615 13297 21152 13322
rect 20565 13279 21152 13297
rect 26591 13291 26635 13343
rect 27733 13295 27777 13347
rect 14454 13233 14514 13254
rect 14572 13233 14632 13254
rect 14690 13233 14750 13254
rect 6232 13187 6705 13203
rect 6232 13153 6248 13187
rect 6282 13162 6705 13187
rect 6282 13161 6469 13162
rect 6282 13153 6298 13161
rect 6232 13137 6298 13153
rect 6409 13141 6469 13161
rect 6527 13141 6587 13162
rect 6645 13141 6705 13162
rect 6763 13162 7059 13203
rect 6763 13141 6823 13162
rect 6881 13141 6941 13162
rect 6999 13141 7059 13162
rect 7362 13191 7847 13207
rect 7362 13157 7378 13191
rect 7412 13166 7847 13191
rect 7412 13165 7611 13166
rect 7412 13157 7428 13165
rect 7362 13141 7428 13157
rect 7551 13145 7611 13165
rect 7669 13145 7729 13166
rect 7787 13145 7847 13166
rect 7905 13166 8201 13207
rect 7905 13145 7965 13166
rect 8023 13145 8083 13166
rect 8141 13145 8201 13166
rect 10633 13178 10929 13214
rect 10633 13157 10693 13178
rect 10751 13157 10811 13178
rect 10869 13157 10929 13178
rect 10987 13177 11283 13213
rect 10987 13157 11047 13177
rect 11105 13157 11165 13177
rect 11223 13157 11283 13177
rect 11341 13177 11637 13213
rect 11341 13157 11401 13177
rect 11459 13157 11519 13177
rect 11577 13157 11637 13177
rect 1194 13110 1254 13136
rect 1312 13110 1372 13136
rect 1430 13110 1490 13136
rect 1548 13116 1608 13136
rect 1548 13110 1609 13116
rect 1666 13110 1726 13136
rect 1784 13110 1844 13136
rect -2553 13082 -2487 13099
rect -3387 12820 -3336 13007
rect -2553 13048 -2537 13082
rect -2503 13048 -2487 13082
rect -2553 13032 -2487 13048
rect 1431 12925 1489 13110
rect 1431 12899 1491 12925
rect 1549 12899 1609 13110
rect 1902 13104 1962 13136
rect 2020 13110 2080 13136
rect 2138 13110 2198 13136
rect 1899 13088 1965 13104
rect 1899 13054 1915 13088
rect 1949 13054 1965 13088
rect 4084 13090 4380 13126
rect 4084 13069 4144 13090
rect 4202 13069 4262 13090
rect 4320 13069 4380 13090
rect 4438 13089 4734 13125
rect 4438 13069 4498 13089
rect 4556 13069 4616 13089
rect 4674 13069 4734 13089
rect 4792 13089 5088 13125
rect 4792 13069 4852 13089
rect 4910 13069 4970 13089
rect 5028 13069 5088 13089
rect 1899 13038 1965 13054
rect 1781 12971 1847 12987
rect 1781 12937 1797 12971
rect 1831 12937 1847 12971
rect 1781 12921 1847 12937
rect 1784 12899 1844 12921
rect -3674 12760 -3606 12820
rect -3406 12760 -3336 12820
rect -2485 12792 -2419 12808
rect -3249 12770 -3195 12786
rect -3674 12702 -3623 12760
rect -3249 12736 -3239 12770
rect -3205 12736 -3195 12770
rect -3249 12718 -3195 12736
rect -2485 12758 -2469 12792
rect -2435 12758 -2419 12792
rect -2485 12718 -2419 12758
rect -3387 12702 -2381 12718
rect -3674 12642 -3606 12702
rect -3406 12658 -2381 12702
rect -2181 12658 -2155 12718
rect -3406 12643 -3336 12658
rect -3406 12642 -3380 12643
rect -3674 12584 -3623 12642
rect -3674 12524 -3606 12584
rect -3406 12524 -3380 12584
rect 4084 12843 4144 12869
rect 4202 12843 4262 12869
rect 4320 12843 4380 12869
rect 4438 12849 4498 12869
rect 4438 12843 4499 12849
rect 4556 12843 4616 12869
rect 4674 12843 4734 12869
rect 1784 12673 1844 12699
rect 4321 12658 4379 12843
rect 4321 12632 4381 12658
rect 4439 12632 4499 12843
rect 4792 12837 4852 12869
rect 4910 12843 4970 12869
rect 5028 12843 5088 12869
rect 4789 12821 4855 12837
rect 4789 12787 4805 12821
rect 4839 12787 4855 12821
rect 4789 12771 4855 12787
rect 10633 12931 10693 12957
rect 10751 12931 10811 12957
rect 10869 12931 10929 12957
rect 10987 12937 11047 12957
rect 10987 12931 11048 12937
rect 11105 12931 11165 12957
rect 11223 12931 11283 12957
rect 10870 12746 10928 12931
rect 6409 12724 6469 12741
rect 4671 12704 4737 12720
rect 4671 12670 4687 12704
rect 4721 12670 4737 12704
rect 4671 12654 4737 12670
rect 4674 12632 4734 12654
rect 6409 12635 6470 12724
rect 6527 12715 6587 12741
rect 6645 12715 6705 12741
rect 1431 12477 1491 12499
rect 1549 12477 1609 12499
rect 1428 12461 1494 12477
rect 1428 12427 1444 12461
rect 1478 12427 1494 12461
rect 1428 12411 1494 12427
rect 1546 12461 1612 12477
rect 1546 12427 1562 12461
rect 1596 12427 1612 12461
rect 1546 12411 1612 12427
rect 6319 12582 6470 12635
rect 4674 12406 4734 12432
rect 6319 12358 6379 12582
rect 6763 12540 6823 12741
rect 6881 12715 6941 12741
rect 6999 12715 7059 12741
rect 7551 12728 7611 12745
rect 7551 12639 7612 12728
rect 7669 12719 7729 12745
rect 7787 12719 7847 12745
rect 6437 12489 6823 12540
rect 7461 12586 7612 12639
rect 6437 12358 6497 12489
rect 6552 12431 6618 12447
rect 6552 12397 6568 12431
rect 6602 12397 6618 12431
rect 6552 12381 6618 12397
rect 6555 12358 6615 12381
rect 6838 12358 6898 12384
rect 6956 12358 7016 12384
rect 7074 12358 7134 12384
rect 7461 12362 7521 12586
rect 7905 12544 7965 12745
rect 8023 12719 8083 12745
rect 8141 12719 8201 12745
rect 10870 12720 10930 12746
rect 10988 12720 11048 12931
rect 11341 12925 11401 12957
rect 11459 12931 11519 12957
rect 11577 12931 11637 12957
rect 11338 12909 11404 12925
rect 11338 12875 11354 12909
rect 11388 12875 11404 12909
rect 11338 12859 11404 12875
rect 19966 13223 20010 13275
rect 21108 13227 21152 13279
rect 26060 13275 26533 13291
rect 26060 13241 26076 13275
rect 26110 13250 26533 13275
rect 26110 13249 26297 13250
rect 26110 13241 26126 13249
rect 19435 13207 19908 13223
rect 19435 13173 19451 13207
rect 19485 13182 19908 13207
rect 19485 13181 19672 13182
rect 19485 13173 19501 13181
rect 19435 13157 19501 13173
rect 19612 13161 19672 13181
rect 19730 13161 19790 13182
rect 19848 13161 19908 13182
rect 19966 13182 20262 13223
rect 19966 13161 20026 13182
rect 20084 13161 20144 13182
rect 20202 13161 20262 13182
rect 20565 13211 21050 13227
rect 20565 13177 20581 13211
rect 20615 13186 21050 13211
rect 20615 13185 20814 13186
rect 20615 13177 20631 13185
rect 20565 13161 20631 13177
rect 20754 13165 20814 13185
rect 20872 13165 20932 13186
rect 20990 13165 21050 13186
rect 21108 13186 21404 13227
rect 26060 13225 26126 13241
rect 26237 13229 26297 13249
rect 26355 13229 26415 13250
rect 26473 13229 26533 13250
rect 26591 13250 26887 13291
rect 26591 13229 26651 13250
rect 26709 13229 26769 13250
rect 26827 13229 26887 13250
rect 27190 13279 27675 13295
rect 27190 13245 27206 13279
rect 27240 13254 27675 13279
rect 27240 13253 27439 13254
rect 27240 13245 27256 13253
rect 27190 13229 27256 13245
rect 27379 13233 27439 13253
rect 27497 13233 27557 13254
rect 27615 13233 27675 13254
rect 27733 13254 28029 13295
rect 27733 13233 27793 13254
rect 27851 13233 27911 13254
rect 27969 13233 28029 13254
rect 31647 13233 31707 13259
rect 21108 13165 21168 13186
rect 21226 13165 21286 13186
rect 21344 13165 21404 13186
rect 23912 13178 24208 13214
rect 17287 13110 17583 13146
rect 17287 13089 17347 13110
rect 17405 13089 17465 13110
rect 17523 13089 17583 13110
rect 17641 13109 17937 13145
rect 17641 13089 17701 13109
rect 17759 13089 17819 13109
rect 17877 13089 17937 13109
rect 17995 13109 18291 13145
rect 17995 13089 18055 13109
rect 18113 13089 18173 13109
rect 18231 13089 18291 13109
rect 17287 12863 17347 12889
rect 17405 12863 17465 12889
rect 17523 12863 17583 12889
rect 17641 12869 17701 12889
rect 17641 12863 17702 12869
rect 17759 12863 17819 12889
rect 17877 12863 17937 12889
rect 12958 12812 13018 12829
rect 11220 12792 11286 12808
rect 11220 12758 11236 12792
rect 11270 12758 11286 12792
rect 11220 12742 11286 12758
rect 11223 12720 11283 12742
rect 12958 12723 13019 12812
rect 13076 12803 13136 12829
rect 13194 12803 13254 12829
rect 7579 12493 7965 12544
rect 7579 12362 7639 12493
rect 7694 12435 7760 12451
rect 7694 12401 7710 12435
rect 7744 12401 7760 12435
rect 7694 12385 7760 12401
rect 7697 12362 7757 12385
rect 7980 12362 8040 12388
rect 8098 12362 8158 12388
rect 8216 12362 8276 12388
rect 4321 12210 4381 12232
rect 4439 12210 4499 12232
rect 4318 12194 4384 12210
rect 4318 12160 4334 12194
rect 4368 12160 4384 12194
rect 4318 12144 4384 12160
rect 4436 12194 4502 12210
rect 4436 12160 4452 12194
rect 4486 12160 4502 12194
rect 4436 12144 4502 12160
rect 12868 12670 13019 12723
rect 11223 12494 11283 12520
rect 12868 12446 12928 12670
rect 13312 12628 13372 12829
rect 13430 12803 13490 12829
rect 13548 12803 13608 12829
rect 14100 12816 14160 12833
rect 14100 12727 14161 12816
rect 14218 12807 14278 12833
rect 14336 12807 14396 12833
rect 12986 12577 13372 12628
rect 14010 12674 14161 12727
rect 12986 12446 13046 12577
rect 13101 12519 13167 12535
rect 13101 12485 13117 12519
rect 13151 12485 13167 12519
rect 13101 12469 13167 12485
rect 13104 12446 13164 12469
rect 13387 12446 13447 12472
rect 13505 12446 13565 12472
rect 13623 12446 13683 12472
rect 14010 12450 14070 12674
rect 14454 12632 14514 12833
rect 14572 12807 14632 12833
rect 14690 12807 14750 12833
rect 17524 12678 17582 12863
rect 17524 12652 17584 12678
rect 17642 12652 17702 12863
rect 17995 12857 18055 12889
rect 18113 12863 18173 12889
rect 18231 12863 18291 12889
rect 17992 12841 18058 12857
rect 17992 12807 18008 12841
rect 18042 12807 18058 12841
rect 17992 12791 18058 12807
rect 23912 13157 23972 13178
rect 24030 13157 24090 13178
rect 24148 13157 24208 13178
rect 24266 13177 24562 13213
rect 24266 13157 24326 13177
rect 24384 13157 24444 13177
rect 24502 13157 24562 13177
rect 24620 13177 24916 13213
rect 24620 13157 24680 13177
rect 24738 13157 24798 13177
rect 24856 13157 24916 13177
rect 23912 12931 23972 12957
rect 24030 12931 24090 12957
rect 24148 12931 24208 12957
rect 24266 12937 24326 12957
rect 24266 12931 24327 12937
rect 24384 12931 24444 12957
rect 24502 12931 24562 12957
rect 19612 12744 19672 12761
rect 17874 12724 17940 12740
rect 17874 12690 17890 12724
rect 17924 12690 17940 12724
rect 17874 12674 17940 12690
rect 17877 12652 17937 12674
rect 19612 12655 19673 12744
rect 19730 12735 19790 12761
rect 19848 12735 19908 12761
rect 14128 12581 14514 12632
rect 14128 12450 14188 12581
rect 14243 12523 14309 12539
rect 14243 12489 14259 12523
rect 14293 12489 14309 12523
rect 14243 12473 14309 12489
rect 14246 12450 14306 12473
rect 14529 12450 14589 12476
rect 14647 12450 14707 12476
rect 14765 12450 14825 12476
rect 10870 12298 10930 12320
rect 10988 12298 11048 12320
rect 10867 12282 10933 12298
rect 10867 12248 10883 12282
rect 10917 12248 10933 12282
rect 10867 12232 10933 12248
rect 10985 12282 11051 12298
rect 10985 12248 11001 12282
rect 11035 12248 11051 12282
rect 10985 12232 11051 12248
rect 19522 12602 19673 12655
rect 17877 12426 17937 12452
rect 19522 12378 19582 12602
rect 19966 12560 20026 12761
rect 20084 12735 20144 12761
rect 20202 12735 20262 12761
rect 20754 12748 20814 12765
rect 20754 12659 20815 12748
rect 20872 12739 20932 12765
rect 20990 12739 21050 12765
rect 19640 12509 20026 12560
rect 20664 12606 20815 12659
rect 19640 12378 19700 12509
rect 19755 12451 19821 12467
rect 19755 12417 19771 12451
rect 19805 12417 19821 12451
rect 19755 12401 19821 12417
rect 19758 12378 19818 12401
rect 20041 12378 20101 12404
rect 20159 12378 20219 12404
rect 20277 12378 20337 12404
rect 20664 12382 20724 12606
rect 21108 12564 21168 12765
rect 21226 12739 21286 12765
rect 21344 12739 21404 12765
rect 24149 12746 24207 12931
rect 24149 12720 24209 12746
rect 24267 12720 24327 12931
rect 24620 12925 24680 12957
rect 24738 12931 24798 12957
rect 24856 12931 24916 12957
rect 24617 12909 24683 12925
rect 24617 12875 24633 12909
rect 24667 12875 24683 12909
rect 24617 12859 24683 12875
rect 36896 13414 36951 13474
rect 37151 13414 37177 13474
rect 36896 13356 36935 13414
rect 36896 13296 36951 13356
rect 37151 13296 37177 13356
rect 37297 13332 37363 13348
rect 37297 13298 37313 13332
rect 37347 13298 37363 13332
rect 32945 13233 33005 13259
rect 36896 13238 36935 13296
rect 37297 13282 37363 13298
rect 37300 13238 37360 13282
rect 37836 13238 37881 14046
rect 36896 13178 36951 13238
rect 37151 13178 37881 13238
rect 32067 13033 32127 13059
rect 32185 13033 32245 13059
rect 32303 13033 32363 13059
rect 32421 13033 32481 13059
rect 26237 12812 26297 12829
rect 24499 12792 24565 12808
rect 24499 12758 24515 12792
rect 24549 12758 24565 12792
rect 24499 12742 24565 12758
rect 24502 12720 24562 12742
rect 26237 12723 26298 12812
rect 26355 12803 26415 12829
rect 26473 12803 26533 12829
rect 20782 12513 21168 12564
rect 20782 12382 20842 12513
rect 20897 12455 20963 12471
rect 20897 12421 20913 12455
rect 20947 12421 20963 12455
rect 20897 12405 20963 12421
rect 20900 12382 20960 12405
rect 21183 12382 21243 12408
rect 21301 12382 21361 12408
rect 21419 12382 21479 12408
rect 12868 12220 12928 12246
rect 12986 12220 13046 12246
rect 13104 12214 13164 12246
rect 13387 12214 13447 12246
rect 13505 12214 13565 12246
rect 13623 12214 13683 12246
rect 14010 12224 14070 12250
rect 14128 12224 14188 12250
rect 13104 12173 13683 12214
rect 14246 12218 14306 12250
rect 14529 12218 14589 12250
rect 14647 12218 14707 12250
rect 14765 12218 14825 12250
rect 17524 12230 17584 12252
rect 17642 12230 17702 12252
rect 14246 12177 14825 12218
rect 17521 12214 17587 12230
rect 17521 12180 17537 12214
rect 17571 12180 17587 12214
rect 17521 12164 17587 12180
rect 17639 12214 17705 12230
rect 17639 12180 17655 12214
rect 17689 12180 17705 12214
rect 17639 12164 17705 12180
rect 26147 12670 26298 12723
rect 24502 12494 24562 12520
rect 26147 12446 26207 12670
rect 26591 12628 26651 12829
rect 26709 12803 26769 12829
rect 26827 12803 26887 12829
rect 27379 12816 27439 12833
rect 27379 12727 27440 12816
rect 27497 12807 27557 12833
rect 27615 12807 27675 12833
rect 26265 12577 26651 12628
rect 27289 12674 27440 12727
rect 26265 12446 26325 12577
rect 26380 12519 26446 12535
rect 26380 12485 26396 12519
rect 26430 12485 26446 12519
rect 26380 12469 26446 12485
rect 26383 12446 26443 12469
rect 26666 12446 26726 12472
rect 26784 12446 26844 12472
rect 26902 12446 26962 12472
rect 27289 12450 27349 12674
rect 27733 12632 27793 12833
rect 27851 12807 27911 12833
rect 27969 12807 28029 12833
rect 27407 12581 27793 12632
rect 27407 12450 27467 12581
rect 29709 12539 30005 12575
rect 27522 12523 27588 12539
rect 27522 12489 27538 12523
rect 27572 12489 27588 12523
rect 29709 12518 29769 12539
rect 29827 12518 29887 12539
rect 29945 12518 30005 12539
rect 30063 12538 30359 12574
rect 30063 12518 30123 12538
rect 30181 12518 30241 12538
rect 30299 12518 30359 12538
rect 30417 12538 30713 12574
rect 30417 12518 30477 12538
rect 30535 12518 30595 12538
rect 30653 12518 30713 12538
rect 27522 12473 27588 12489
rect 27525 12450 27585 12473
rect 27808 12450 27868 12476
rect 27926 12450 27986 12476
rect 28044 12450 28104 12476
rect 24149 12298 24209 12320
rect 24267 12298 24327 12320
rect 24146 12282 24212 12298
rect 24146 12248 24162 12282
rect 24196 12248 24212 12282
rect 24146 12232 24212 12248
rect 24264 12282 24330 12298
rect 24264 12248 24280 12282
rect 24314 12248 24330 12282
rect 24264 12232 24330 12248
rect 36900 12420 36955 12480
rect 37155 12421 37885 12480
rect 37155 12420 37458 12421
rect 36900 12362 36939 12420
rect 37441 12363 37458 12420
rect 37513 12420 37885 12421
rect 37513 12363 37528 12420
rect 29709 12292 29769 12318
rect 29827 12292 29887 12318
rect 29945 12292 30005 12318
rect 30063 12298 30123 12318
rect 30063 12292 30124 12298
rect 30181 12292 30241 12318
rect 30299 12292 30359 12318
rect 26147 12220 26207 12246
rect 26265 12220 26325 12246
rect 26383 12214 26443 12246
rect 26666 12214 26726 12246
rect 26784 12214 26844 12246
rect 26902 12214 26962 12246
rect 27289 12224 27349 12250
rect 27407 12224 27467 12250
rect 6319 12132 6379 12158
rect 6437 12132 6497 12158
rect 6555 12126 6615 12158
rect 6838 12126 6898 12158
rect 6956 12126 7016 12158
rect 7074 12126 7134 12158
rect 7461 12136 7521 12162
rect 7579 12136 7639 12162
rect -3057 12095 -2997 12111
rect -3630 12012 -3604 12072
rect -3404 12012 -3336 12072
rect -3387 11954 -3336 12012
rect -3630 11894 -3604 11954
rect -3404 11947 -3336 11954
rect -3057 12061 -3043 12095
rect -3009 12061 -2997 12095
rect 6555 12085 7134 12126
rect 7697 12130 7757 12162
rect 7980 12130 8040 12162
rect 8098 12130 8158 12162
rect 8216 12130 8276 12162
rect 19522 12152 19582 12178
rect 19640 12152 19700 12178
rect 7697 12089 8276 12130
rect 19758 12146 19818 12178
rect 20041 12146 20101 12178
rect 20159 12146 20219 12178
rect 20277 12146 20337 12178
rect 20664 12156 20724 12182
rect 20782 12156 20842 12182
rect 19758 12105 20337 12146
rect 20900 12150 20960 12182
rect 21183 12150 21243 12182
rect 21301 12150 21361 12182
rect 21419 12150 21479 12182
rect 26383 12173 26962 12214
rect 27525 12218 27585 12250
rect 27808 12218 27868 12250
rect 27926 12218 27986 12250
rect 28044 12218 28104 12250
rect 27525 12177 28104 12218
rect 20900 12109 21479 12150
rect 29946 12107 30004 12292
rect 29946 12081 30006 12107
rect 30064 12081 30124 12292
rect 30417 12286 30477 12318
rect 30535 12292 30595 12318
rect 30653 12292 30713 12318
rect 36900 12302 36955 12362
rect 37155 12302 37181 12362
rect 37441 12344 37528 12363
rect 30414 12270 30480 12286
rect 30414 12236 30430 12270
rect 30464 12236 30480 12270
rect 30414 12220 30480 12236
rect 36900 12244 36939 12302
rect 36900 12184 36955 12244
rect 37155 12184 37181 12244
rect 30296 12153 30362 12169
rect 30296 12119 30312 12153
rect 30346 12119 30362 12153
rect 30296 12103 30362 12119
rect 30299 12081 30359 12103
rect -3057 11947 -2997 12061
rect -3404 11894 -2379 11947
rect -3387 11887 -2379 11894
rect -2179 11887 -2153 11947
rect -3387 11836 -3336 11887
rect -3630 11776 -3604 11836
rect -3404 11776 -3336 11836
rect -2484 11846 -2418 11887
rect -2484 11812 -2468 11846
rect -2434 11812 -2418 11846
rect -2484 11796 -2418 11812
rect -3387 11588 -3336 11776
rect -2551 11661 -2485 11677
rect -3870 11528 -3804 11588
rect -3404 11528 -3336 11588
rect -3194 11585 -3111 11645
rect -2711 11585 -2685 11645
rect -2551 11627 -2535 11661
rect -2501 11627 -2485 11661
rect -2551 11610 -2485 11627
rect -3870 11470 -3819 11528
rect -3194 11527 -3134 11585
rect -2544 11527 -2485 11610
rect 36701 11979 36755 12039
rect 37155 11979 37181 12039
rect 36701 11921 36740 11979
rect 30299 11855 30359 11881
rect 36701 11861 36755 11921
rect 37155 11861 37630 11921
rect 36701 11803 36740 11861
rect 36701 11743 36755 11803
rect 37155 11743 37181 11803
rect 29946 11659 30006 11681
rect 30064 11659 30124 11681
rect 29943 11643 30009 11659
rect 29943 11609 29959 11643
rect 29993 11609 30009 11643
rect 10647 11528 10943 11564
rect -3870 11410 -3804 11470
rect -3404 11410 -3378 11470
rect -3194 11467 -3111 11527
rect -2711 11467 -2379 11527
rect -1979 11467 -1953 11527
rect 10647 11507 10707 11528
rect 10765 11507 10825 11528
rect 10883 11507 10943 11528
rect 11001 11527 11297 11563
rect 11001 11507 11061 11527
rect 11119 11507 11179 11527
rect 11237 11507 11297 11527
rect 11355 11527 11651 11563
rect 11355 11507 11415 11527
rect 11473 11507 11533 11527
rect 11591 11507 11651 11527
rect -3870 11352 -3819 11410
rect -3194 11409 -3134 11467
rect -2467 11409 -2401 11411
rect -3870 11292 -3804 11352
rect -3404 11292 -3378 11352
rect -3194 11349 -3111 11409
rect -2711 11349 -2685 11409
rect -2467 11395 -2379 11409
rect -2467 11361 -2451 11395
rect -2417 11361 -2379 11395
rect -2467 11349 -2379 11361
rect -1979 11349 -1953 11409
rect 4098 11440 4394 11476
rect 4098 11419 4158 11440
rect 4216 11419 4276 11440
rect 4334 11419 4394 11440
rect 4452 11439 4748 11475
rect 4452 11419 4512 11439
rect 4570 11419 4630 11439
rect 4688 11419 4748 11439
rect 4806 11439 5102 11475
rect 4806 11419 4866 11439
rect 4924 11419 4984 11439
rect 5042 11419 5102 11439
rect -2467 11345 -2401 11349
rect -2467 11291 -2402 11293
rect -3830 11174 -3804 11234
rect -3404 11174 -3334 11234
rect -3385 11116 -3334 11174
rect -3830 11056 -3804 11116
rect -3404 11056 -3334 11116
rect -3385 10998 -3334 11056
rect -3830 10938 -3804 10998
rect -3404 10938 -3334 10998
rect -3195 11231 -3111 11291
rect -2711 11231 -2685 11291
rect -2467 11277 -2379 11291
rect -2467 11243 -2452 11277
rect -2418 11243 -2379 11277
rect -2467 11231 -2379 11243
rect -1979 11231 -1953 11291
rect -3195 11173 -3135 11231
rect -2467 11227 -2402 11231
rect 29943 11593 30009 11609
rect 30061 11643 30127 11659
rect 30061 11609 30077 11643
rect 30111 11609 30127 11643
rect 30061 11593 30127 11609
rect 23926 11528 24222 11564
rect 23926 11507 23986 11528
rect 24044 11507 24104 11528
rect 24162 11507 24222 11528
rect 24280 11527 24576 11563
rect 24280 11507 24340 11527
rect 24398 11507 24458 11527
rect 24516 11507 24576 11527
rect 24634 11527 24930 11563
rect 24634 11507 24694 11527
rect 24752 11507 24812 11527
rect 24870 11507 24930 11527
rect 17301 11460 17597 11496
rect 17301 11439 17361 11460
rect 17419 11439 17479 11460
rect 17537 11439 17597 11460
rect 17655 11459 17951 11495
rect 17655 11439 17715 11459
rect 17773 11439 17833 11459
rect 17891 11439 17951 11459
rect 18009 11459 18305 11495
rect 18009 11439 18069 11459
rect 18127 11439 18187 11459
rect 18245 11439 18305 11459
rect 10647 11281 10707 11307
rect 10765 11281 10825 11307
rect 10883 11281 10943 11307
rect 11001 11287 11061 11307
rect 11001 11281 11062 11287
rect 11119 11281 11179 11307
rect 11237 11281 11297 11307
rect 4098 11193 4158 11219
rect 4216 11193 4276 11219
rect 4334 11193 4394 11219
rect 4452 11199 4512 11219
rect 4452 11193 4513 11199
rect 4570 11193 4630 11219
rect 4688 11193 4748 11219
rect -3195 11113 -3111 11173
rect -2711 11113 -2379 11173
rect -1979 11113 -1953 11173
rect -3195 11055 -3135 11113
rect -3195 10995 -3111 11055
rect -2711 10995 -2685 11055
rect -2544 11030 -2485 11113
rect -2551 11013 -2485 11030
rect -3385 10751 -3334 10938
rect -2551 10979 -2535 11013
rect -2501 10979 -2485 11013
rect -2551 10963 -2485 10979
rect 4335 11008 4393 11193
rect 4335 10982 4395 11008
rect 4453 10982 4513 11193
rect 4806 11187 4866 11219
rect 4924 11193 4984 11219
rect 5042 11193 5102 11219
rect 4803 11171 4869 11187
rect 4803 11137 4819 11171
rect 4853 11137 4869 11171
rect 4803 11121 4869 11137
rect 10884 11096 10942 11281
rect 10884 11070 10944 11096
rect 11002 11070 11062 11281
rect 11355 11275 11415 11307
rect 11473 11281 11533 11307
rect 11591 11281 11651 11307
rect 11352 11259 11418 11275
rect 11352 11225 11368 11259
rect 11402 11225 11418 11259
rect 36701 11512 36755 11572
rect 37155 11512 37181 11572
rect 36701 11454 36740 11512
rect 36701 11394 36755 11454
rect 37155 11453 37181 11454
rect 37342 11453 37408 11456
rect 37155 11440 37408 11453
rect 37155 11406 37358 11440
rect 37392 11406 37408 11440
rect 37155 11394 37408 11406
rect 37573 11454 37630 11861
rect 37840 11646 37885 12420
rect 37840 11586 38088 11646
rect 38288 11586 38314 11646
rect 37729 11454 37808 11465
rect 37573 11452 38088 11454
rect 37573 11394 37742 11452
rect 37797 11394 38088 11452
rect 38488 11394 38514 11454
rect 23926 11281 23986 11307
rect 24044 11281 24104 11307
rect 24162 11281 24222 11307
rect 24280 11287 24340 11307
rect 24280 11281 24341 11287
rect 24398 11281 24458 11307
rect 24516 11281 24576 11307
rect 11352 11209 11418 11225
rect 17301 11213 17361 11239
rect 17419 11213 17479 11239
rect 17537 11213 17597 11239
rect 17655 11219 17715 11239
rect 17655 11213 17716 11219
rect 17773 11213 17833 11239
rect 17891 11213 17951 11239
rect 11234 11142 11300 11158
rect 11234 11108 11250 11142
rect 11284 11108 11300 11142
rect 11234 11092 11300 11108
rect 12595 11105 12891 11156
rect 11237 11070 11297 11092
rect 12595 11090 12655 11105
rect 12713 11090 12773 11105
rect 12831 11090 12891 11105
rect 12949 11090 13009 11116
rect 13067 11090 13127 11116
rect 13185 11090 13245 11116
rect 14493 11105 14789 11156
rect 14493 11090 14553 11105
rect 14611 11090 14671 11105
rect 14729 11090 14789 11105
rect 14847 11090 14907 11116
rect 14965 11090 15025 11116
rect 15083 11090 15143 11116
rect 4685 11054 4751 11070
rect 4685 11020 4701 11054
rect 4735 11020 4751 11054
rect 4685 11004 4751 11020
rect 6046 11017 6342 11068
rect 4688 10982 4748 11004
rect 6046 11002 6106 11017
rect 6164 11002 6224 11017
rect 6282 11002 6342 11017
rect 6400 11002 6460 11028
rect 6518 11002 6578 11028
rect 6636 11002 6696 11028
rect 7944 11017 8240 11068
rect 7944 11002 8004 11017
rect 8062 11002 8122 11017
rect 8180 11002 8240 11017
rect 8298 11002 8358 11028
rect 8416 11002 8476 11028
rect 8534 11002 8594 11028
rect 1186 10772 1482 10808
rect 1186 10751 1246 10772
rect 1304 10751 1364 10772
rect 1422 10751 1482 10772
rect 1540 10771 1836 10807
rect 1540 10751 1600 10771
rect 1658 10751 1718 10771
rect 1776 10751 1836 10771
rect 1894 10771 2190 10807
rect 1894 10751 1954 10771
rect 2012 10751 2072 10771
rect 2130 10751 2190 10771
rect -3672 10691 -3604 10751
rect -3404 10691 -3334 10751
rect -2483 10723 -2417 10739
rect -3247 10701 -3193 10717
rect -3672 10633 -3621 10691
rect -3247 10667 -3237 10701
rect -3203 10667 -3193 10701
rect -3247 10649 -3193 10667
rect -2483 10689 -2467 10723
rect -2433 10689 -2417 10723
rect -2483 10649 -2417 10689
rect -3385 10633 -2379 10649
rect -3672 10573 -3604 10633
rect -3404 10589 -2379 10633
rect -2179 10589 -2153 10649
rect -3404 10574 -3334 10589
rect -3404 10573 -3378 10574
rect -3672 10515 -3621 10573
rect 5562 10802 5622 10828
rect 5680 10802 5740 10828
rect 5798 10802 5858 10828
rect 4688 10756 4748 10782
rect 4335 10560 4395 10582
rect 4453 10566 4513 10582
rect 1186 10525 1246 10551
rect 1304 10525 1364 10551
rect 1422 10525 1482 10551
rect 1540 10531 1600 10551
rect 1540 10525 1601 10531
rect 1658 10525 1718 10551
rect 1776 10525 1836 10551
rect -3672 10455 -3604 10515
rect -3404 10455 -3378 10515
rect 1423 10340 1481 10525
rect 1423 10314 1483 10340
rect 1541 10314 1601 10525
rect 1894 10519 1954 10551
rect 2012 10525 2072 10551
rect 2130 10525 2190 10551
rect 4332 10544 4398 10560
rect 1891 10503 1957 10519
rect 1891 10469 1907 10503
rect 1941 10469 1957 10503
rect 4332 10510 4348 10544
rect 4382 10510 4398 10544
rect 4332 10494 4398 10510
rect 4447 10544 4521 10566
rect 4447 10510 4466 10544
rect 4500 10510 4521 10544
rect 6883 10819 7179 10870
rect 6883 10802 6943 10819
rect 7001 10802 7061 10819
rect 7119 10802 7179 10819
rect 7460 10802 7520 10828
rect 7578 10802 7638 10828
rect 7696 10802 7756 10828
rect 8781 10819 9077 10870
rect 8781 10802 8841 10819
rect 8899 10802 8959 10819
rect 9017 10802 9077 10819
rect 12111 10890 12171 10916
rect 12229 10890 12289 10916
rect 12347 10890 12407 10916
rect 11237 10844 11297 10870
rect 10884 10648 10944 10670
rect 11002 10654 11062 10670
rect 10881 10632 10947 10648
rect 5562 10585 5622 10602
rect 5680 10585 5740 10602
rect 5798 10585 5858 10602
rect 6046 10585 6106 10602
rect 5562 10534 6106 10585
rect 6164 10576 6224 10602
rect 6282 10576 6342 10602
rect 6400 10583 6460 10602
rect 6518 10583 6578 10602
rect 6636 10583 6696 10602
rect 6883 10583 6943 10602
rect 7001 10583 7061 10602
rect 1891 10453 1957 10469
rect 4447 10453 4521 10510
rect 5687 10453 5747 10534
rect 6400 10532 6943 10583
rect 6985 10576 7061 10583
rect 7119 10576 7179 10602
rect 7460 10585 7520 10602
rect 7578 10585 7638 10602
rect 7696 10585 7756 10602
rect 7944 10585 8004 10602
rect 6985 10532 7060 10576
rect 7460 10534 8004 10585
rect 8062 10576 8122 10602
rect 8180 10576 8240 10602
rect 8298 10583 8358 10602
rect 8416 10583 8476 10602
rect 8534 10583 8594 10602
rect 8781 10583 8841 10602
rect 8899 10583 8959 10602
rect 4447 10428 5747 10453
rect 1773 10386 1839 10402
rect 1773 10352 1789 10386
rect 1823 10352 1839 10386
rect 4446 10380 5747 10428
rect 6985 10412 7045 10532
rect 1773 10336 1839 10352
rect 1776 10314 1836 10336
rect -3059 10027 -2999 10043
rect -3632 9944 -3606 10004
rect -3406 9944 -3338 10004
rect -3389 9886 -3338 9944
rect -3632 9826 -3606 9886
rect -3406 9879 -3338 9886
rect -3059 9993 -3045 10027
rect -3011 9993 -2999 10027
rect -3059 9879 -2999 9993
rect 1776 10088 1836 10114
rect 1423 9892 1483 9914
rect 1541 9892 1601 9914
rect -3406 9826 -2381 9879
rect -3389 9819 -2381 9826
rect -2181 9819 -2155 9879
rect 1420 9876 1486 9892
rect 1420 9842 1436 9876
rect 1470 9842 1486 9876
rect 1420 9826 1486 9842
rect 1538 9876 1604 9892
rect 1538 9842 1554 9876
rect 1588 9842 1604 9876
rect 1538 9826 1604 9842
rect 4093 9836 4389 9872
rect -3389 9768 -3338 9819
rect -3632 9708 -3606 9768
rect -3406 9708 -3338 9768
rect -2486 9778 -2420 9819
rect -2486 9744 -2470 9778
rect -2436 9744 -2420 9778
rect 4093 9815 4153 9836
rect 4211 9815 4271 9836
rect 4329 9815 4389 9836
rect 4447 9835 4743 9871
rect 4447 9815 4507 9835
rect 4565 9815 4625 9835
rect 4683 9815 4743 9835
rect 4801 9835 5097 9871
rect 4801 9815 4861 9835
rect 4919 9815 4979 9835
rect 5037 9815 5097 9835
rect -2486 9728 -2420 9744
rect -3389 9520 -3338 9708
rect 5687 9682 5747 10380
rect 5989 10332 6285 10392
rect 5989 10309 6049 10332
rect 6107 10309 6167 10332
rect 6225 10309 6285 10332
rect 6343 10333 6639 10393
rect 6984 10392 7045 10412
rect 6343 10309 6403 10333
rect 6461 10309 6521 10333
rect 6579 10309 6639 10333
rect 6965 10376 7045 10392
rect 6965 10342 6980 10376
rect 7014 10342 7045 10376
rect 6965 10326 7045 10342
rect 6984 10303 7045 10326
rect 6985 10157 7045 10303
rect 6984 9984 7045 10157
rect 5989 9883 6049 9909
rect 5957 9742 6024 9749
rect 6107 9742 6167 9909
rect 6225 9883 6285 9909
rect 6343 9883 6403 9909
rect 5957 9733 6167 9742
rect 5957 9699 5973 9733
rect 6007 9699 6167 9733
rect 5957 9683 6167 9699
rect 5687 9666 5838 9682
rect 5687 9632 5788 9666
rect 5822 9632 5838 9666
rect 5687 9616 5838 9632
rect -2553 9593 -2487 9609
rect -3872 9460 -3806 9520
rect -3406 9460 -3338 9520
rect -3196 9517 -3113 9577
rect -2713 9517 -2687 9577
rect -2553 9559 -2537 9593
rect -2503 9559 -2487 9593
rect 4093 9589 4153 9615
rect 4211 9589 4271 9615
rect 4329 9589 4389 9615
rect 4447 9595 4507 9615
rect 4447 9589 4508 9595
rect 4565 9589 4625 9615
rect 4683 9589 4743 9615
rect -2553 9542 -2487 9559
rect -3872 9402 -3821 9460
rect -3196 9459 -3136 9517
rect -2546 9459 -2487 9542
rect -3872 9342 -3806 9402
rect -3406 9342 -3380 9402
rect -3196 9399 -3113 9459
rect -2713 9399 -2381 9459
rect -1981 9399 -1955 9459
rect 4330 9404 4388 9589
rect -3872 9284 -3821 9342
rect -3196 9341 -3136 9399
rect 4330 9378 4390 9404
rect 4448 9378 4508 9589
rect 4801 9583 4861 9615
rect 4919 9589 4979 9615
rect 5037 9589 5097 9615
rect 4798 9567 4864 9583
rect 5687 9577 5747 9616
rect 6107 9577 6167 9683
rect 6461 9742 6521 9909
rect 6579 9883 6639 9909
rect 6604 9742 6671 9749
rect 6461 9733 6671 9742
rect 6461 9699 6621 9733
rect 6655 9699 6671 9733
rect 6461 9683 6671 9699
rect 6223 9649 6289 9665
rect 6223 9615 6239 9649
rect 6273 9615 6289 9649
rect 6223 9599 6289 9615
rect 6341 9650 6407 9665
rect 6341 9616 6357 9650
rect 6391 9616 6407 9650
rect 6341 9600 6407 9616
rect 6225 9577 6285 9599
rect 6343 9577 6403 9600
rect 6461 9577 6521 9683
rect 6985 9681 7045 9984
rect 6895 9665 7045 9681
rect 6895 9631 6911 9665
rect 6945 9631 7045 9665
rect 6895 9615 7045 9631
rect 6985 9577 7045 9615
rect 7585 9876 7645 10534
rect 8298 10532 8841 10583
rect 8883 10576 8959 10583
rect 9017 10576 9077 10602
rect 10881 10598 10897 10632
rect 10931 10598 10947 10632
rect 10881 10582 10947 10598
rect 10996 10632 11070 10654
rect 10996 10598 11015 10632
rect 11049 10598 11070 10632
rect 13432 10907 13728 10958
rect 13432 10890 13492 10907
rect 13550 10890 13610 10907
rect 13668 10890 13728 10907
rect 14009 10890 14069 10916
rect 14127 10890 14187 10916
rect 14245 10890 14305 10916
rect 17538 11028 17596 11213
rect 17538 11002 17598 11028
rect 17656 11002 17716 11213
rect 18009 11207 18069 11239
rect 18127 11213 18187 11239
rect 18245 11213 18305 11239
rect 18006 11191 18072 11207
rect 18006 11157 18022 11191
rect 18056 11157 18072 11191
rect 18006 11141 18072 11157
rect 24163 11096 24221 11281
rect 17888 11074 17954 11090
rect 17888 11040 17904 11074
rect 17938 11040 17954 11074
rect 17888 11024 17954 11040
rect 19249 11037 19545 11088
rect 17891 11002 17951 11024
rect 19249 11022 19309 11037
rect 19367 11022 19427 11037
rect 19485 11022 19545 11037
rect 19603 11022 19663 11048
rect 19721 11022 19781 11048
rect 19839 11022 19899 11048
rect 21147 11037 21443 11088
rect 24163 11070 24223 11096
rect 24281 11070 24341 11281
rect 24634 11275 24694 11307
rect 24752 11281 24812 11307
rect 24870 11281 24930 11307
rect 24631 11259 24697 11275
rect 24631 11225 24647 11259
rect 24681 11225 24697 11259
rect 24631 11209 24697 11225
rect 24513 11142 24579 11158
rect 24513 11108 24529 11142
rect 24563 11108 24579 11142
rect 24513 11092 24579 11108
rect 25874 11105 26170 11156
rect 24516 11070 24576 11092
rect 25874 11090 25934 11105
rect 25992 11090 26052 11105
rect 26110 11090 26170 11105
rect 26228 11090 26288 11116
rect 26346 11090 26406 11116
rect 26464 11090 26524 11116
rect 27772 11105 28068 11156
rect 36701 11336 36740 11394
rect 37341 11390 37408 11394
rect 37729 11384 37808 11394
rect 37442 11336 37529 11353
rect 36701 11276 36755 11336
rect 37155 11276 37181 11336
rect 37442 11334 38088 11336
rect 37442 11276 37457 11334
rect 37512 11276 38088 11334
rect 38488 11276 38514 11336
rect 37442 11258 37529 11276
rect 27772 11090 27832 11105
rect 27890 11090 27950 11105
rect 28008 11090 28068 11105
rect 28126 11090 28186 11116
rect 28244 11090 28304 11116
rect 28362 11090 28422 11116
rect 36701 11158 36755 11218
rect 37155 11158 37181 11218
rect 36701 11100 36740 11158
rect 37480 11100 37529 11258
rect 37962 11218 38028 11221
rect 38561 11263 38627 11279
rect 38561 11229 38577 11263
rect 38611 11229 38627 11263
rect 37962 11205 38088 11218
rect 37962 11171 37978 11205
rect 38012 11171 38088 11205
rect 37962 11158 38088 11171
rect 38488 11158 38514 11218
rect 38561 11213 38627 11229
rect 37962 11155 38028 11158
rect 21147 11022 21207 11037
rect 21265 11022 21325 11037
rect 21383 11022 21443 11037
rect 21501 11022 21561 11048
rect 21619 11022 21679 11048
rect 21737 11022 21797 11048
rect 15330 10907 15626 10958
rect 15330 10890 15390 10907
rect 15448 10890 15508 10907
rect 15566 10890 15626 10907
rect 12111 10673 12171 10690
rect 12229 10673 12289 10690
rect 12347 10673 12407 10690
rect 12595 10673 12655 10690
rect 12111 10622 12655 10673
rect 12713 10664 12773 10690
rect 12831 10664 12891 10690
rect 12949 10671 13009 10690
rect 13067 10671 13127 10690
rect 13185 10671 13245 10690
rect 13432 10671 13492 10690
rect 13550 10671 13610 10690
rect 8883 10532 8958 10576
rect 10996 10541 11070 10598
rect 12236 10541 12296 10622
rect 12949 10620 13492 10671
rect 13534 10664 13610 10671
rect 13668 10664 13728 10690
rect 14009 10673 14069 10690
rect 14127 10673 14187 10690
rect 14245 10673 14305 10690
rect 14493 10673 14553 10690
rect 13534 10620 13609 10664
rect 14009 10622 14553 10673
rect 14611 10664 14671 10690
rect 14729 10664 14789 10690
rect 14847 10671 14907 10690
rect 14965 10671 15025 10690
rect 15083 10671 15143 10690
rect 15330 10671 15390 10690
rect 15448 10671 15508 10690
rect 7887 10332 8183 10392
rect 7887 10309 7947 10332
rect 8005 10309 8065 10332
rect 8123 10309 8183 10332
rect 8241 10333 8537 10393
rect 8241 10309 8301 10333
rect 8359 10309 8419 10333
rect 8477 10309 8537 10333
rect 8883 10379 8943 10532
rect 10996 10516 12296 10541
rect 10995 10468 12296 10516
rect 13534 10500 13594 10620
rect 8883 10355 9137 10379
rect 8883 10321 9087 10355
rect 9121 10321 9137 10355
rect 8883 10305 9137 10321
rect 7887 9883 7947 9909
rect 7585 9860 7652 9876
rect 7585 9826 7601 9860
rect 7635 9826 7652 9860
rect 7585 9810 7652 9826
rect 7585 9682 7645 9810
rect 7855 9742 7922 9749
rect 8005 9742 8065 9909
rect 8123 9883 8183 9909
rect 8241 9883 8301 9909
rect 7855 9733 8065 9742
rect 7855 9699 7871 9733
rect 7905 9699 8065 9733
rect 7855 9683 8065 9699
rect 7585 9666 7736 9682
rect 7585 9632 7686 9666
rect 7720 9632 7736 9666
rect 7585 9616 7736 9632
rect 7585 9577 7645 9616
rect 8005 9577 8065 9683
rect 8359 9742 8419 9909
rect 8477 9883 8537 9909
rect 8500 9743 8567 9750
rect 8494 9742 8567 9743
rect 8359 9734 8567 9742
rect 8359 9700 8517 9734
rect 8551 9700 8567 9734
rect 8359 9684 8567 9700
rect 8359 9683 8556 9684
rect 8121 9649 8187 9665
rect 8121 9615 8137 9649
rect 8171 9615 8187 9649
rect 8121 9599 8187 9615
rect 8239 9650 8305 9665
rect 8239 9616 8255 9650
rect 8289 9616 8305 9650
rect 8239 9600 8305 9616
rect 8123 9577 8183 9599
rect 8241 9577 8301 9600
rect 8359 9577 8419 9683
rect 8883 9681 8943 10305
rect 10642 9924 10938 9960
rect 10642 9903 10702 9924
rect 10760 9903 10820 9924
rect 10878 9903 10938 9924
rect 10996 9923 11292 9959
rect 10996 9903 11056 9923
rect 11114 9903 11174 9923
rect 11232 9903 11292 9923
rect 11350 9923 11646 9959
rect 11350 9903 11410 9923
rect 11468 9903 11528 9923
rect 11586 9903 11646 9923
rect 12236 9770 12296 10468
rect 12538 10420 12834 10480
rect 12538 10397 12598 10420
rect 12656 10397 12716 10420
rect 12774 10397 12834 10420
rect 12892 10421 13188 10481
rect 13533 10480 13594 10500
rect 12892 10397 12952 10421
rect 13010 10397 13070 10421
rect 13128 10397 13188 10421
rect 13514 10464 13594 10480
rect 13514 10430 13529 10464
rect 13563 10430 13594 10464
rect 13514 10414 13594 10430
rect 13533 10391 13594 10414
rect 13534 10245 13594 10391
rect 13533 10072 13594 10245
rect 12538 9971 12598 9997
rect 12506 9830 12573 9837
rect 12656 9830 12716 9997
rect 12774 9971 12834 9997
rect 12892 9971 12952 9997
rect 12506 9821 12716 9830
rect 12506 9787 12522 9821
rect 12556 9787 12716 9821
rect 12506 9771 12716 9787
rect 12236 9754 12387 9770
rect 12236 9720 12337 9754
rect 12371 9720 12387 9754
rect 12236 9704 12387 9720
rect 8793 9665 8943 9681
rect 10642 9677 10702 9703
rect 10760 9677 10820 9703
rect 10878 9677 10938 9703
rect 10996 9683 11056 9703
rect 10996 9677 11057 9683
rect 11114 9677 11174 9703
rect 11232 9677 11292 9703
rect 8793 9631 8809 9665
rect 8843 9631 8943 9665
rect 8793 9615 8943 9631
rect 8883 9577 8943 9615
rect 4798 9533 4814 9567
rect 4848 9533 4864 9567
rect 4798 9517 4864 9533
rect 4680 9450 4746 9466
rect 4680 9416 4696 9450
rect 4730 9416 4746 9450
rect 4680 9400 4746 9416
rect 4683 9378 4743 9400
rect -2469 9341 -2403 9343
rect -3872 9224 -3806 9284
rect -3406 9224 -3380 9284
rect -3196 9281 -3113 9341
rect -2713 9281 -2687 9341
rect -2469 9327 -2381 9341
rect -2469 9293 -2453 9327
rect -2419 9293 -2381 9327
rect -2469 9281 -2381 9293
rect -1981 9281 -1955 9341
rect -2469 9277 -2403 9281
rect -2469 9223 -2404 9225
rect -3832 9106 -3806 9166
rect -3406 9106 -3336 9166
rect -3387 9048 -3336 9106
rect -3832 8988 -3806 9048
rect -3406 8988 -3336 9048
rect -3387 8930 -3336 8988
rect -3832 8870 -3806 8930
rect -3406 8870 -3336 8930
rect -3197 9163 -3113 9223
rect -2713 9163 -2687 9223
rect -2469 9209 -2381 9223
rect -2469 9175 -2454 9209
rect -2420 9175 -2381 9209
rect -2469 9163 -2381 9175
rect -1981 9163 -1955 9223
rect -3197 9105 -3137 9163
rect -2469 9159 -2404 9163
rect -3197 9045 -3113 9105
rect -2713 9045 -2381 9105
rect -1981 9045 -1955 9105
rect -3197 8987 -3137 9045
rect -3197 8927 -3113 8987
rect -2713 8927 -2687 8987
rect -2546 8962 -2487 9045
rect 5687 9351 5747 9377
rect 4683 9152 4743 9178
rect 6985 9351 7045 9377
rect 7585 9351 7645 9377
rect 10879 9492 10937 9677
rect 10879 9466 10939 9492
rect 10997 9466 11057 9677
rect 11350 9671 11410 9703
rect 11468 9677 11528 9703
rect 11586 9677 11646 9703
rect 11347 9655 11413 9671
rect 12236 9665 12296 9704
rect 12656 9665 12716 9771
rect 13010 9830 13070 9997
rect 13128 9971 13188 9997
rect 13153 9830 13220 9837
rect 13010 9821 13220 9830
rect 13010 9787 13170 9821
rect 13204 9787 13220 9821
rect 13010 9771 13220 9787
rect 12772 9737 12838 9753
rect 12772 9703 12788 9737
rect 12822 9703 12838 9737
rect 12772 9687 12838 9703
rect 12890 9738 12956 9753
rect 12890 9704 12906 9738
rect 12940 9704 12956 9738
rect 12890 9688 12956 9704
rect 12774 9665 12834 9687
rect 12892 9665 12952 9688
rect 13010 9665 13070 9771
rect 13534 9769 13594 10072
rect 13444 9753 13594 9769
rect 13444 9719 13460 9753
rect 13494 9719 13594 9753
rect 13444 9703 13594 9719
rect 13534 9665 13594 9703
rect 14134 9964 14194 10622
rect 14847 10620 15390 10671
rect 15432 10664 15508 10671
rect 15566 10664 15626 10690
rect 15432 10620 15507 10664
rect 14436 10420 14732 10480
rect 14436 10397 14496 10420
rect 14554 10397 14614 10420
rect 14672 10397 14732 10420
rect 14790 10421 15086 10481
rect 14790 10397 14850 10421
rect 14908 10397 14968 10421
rect 15026 10397 15086 10421
rect 15432 10467 15492 10620
rect 18765 10822 18825 10848
rect 18883 10822 18943 10848
rect 19001 10822 19061 10848
rect 17891 10776 17951 10802
rect 17538 10580 17598 10602
rect 17656 10586 17716 10602
rect 17535 10564 17601 10580
rect 17535 10530 17551 10564
rect 17585 10530 17601 10564
rect 17535 10514 17601 10530
rect 17650 10564 17724 10586
rect 17650 10530 17669 10564
rect 17703 10530 17724 10564
rect 20086 10839 20382 10890
rect 20086 10822 20146 10839
rect 20204 10822 20264 10839
rect 20322 10822 20382 10839
rect 20663 10822 20723 10848
rect 20781 10822 20841 10848
rect 20899 10822 20959 10848
rect 21984 10839 22280 10890
rect 21984 10822 22044 10839
rect 22102 10822 22162 10839
rect 22220 10822 22280 10839
rect 25390 10890 25450 10916
rect 25508 10890 25568 10916
rect 25626 10890 25686 10916
rect 24516 10844 24576 10870
rect 24163 10648 24223 10670
rect 24281 10654 24341 10670
rect 24160 10632 24226 10648
rect 18765 10605 18825 10622
rect 18883 10605 18943 10622
rect 19001 10605 19061 10622
rect 19249 10605 19309 10622
rect 18765 10554 19309 10605
rect 19367 10596 19427 10622
rect 19485 10596 19545 10622
rect 19603 10603 19663 10622
rect 19721 10603 19781 10622
rect 19839 10603 19899 10622
rect 20086 10603 20146 10622
rect 20204 10603 20264 10622
rect 17650 10473 17724 10530
rect 18890 10473 18950 10554
rect 19603 10552 20146 10603
rect 20188 10596 20264 10603
rect 20322 10596 20382 10622
rect 20663 10605 20723 10622
rect 20781 10605 20841 10622
rect 20899 10605 20959 10622
rect 21147 10605 21207 10622
rect 20188 10552 20263 10596
rect 20663 10554 21207 10605
rect 21265 10596 21325 10622
rect 21383 10596 21443 10622
rect 21501 10603 21561 10622
rect 21619 10603 21679 10622
rect 21737 10603 21797 10622
rect 21984 10603 22044 10622
rect 22102 10603 22162 10622
rect 15432 10443 15686 10467
rect 17650 10448 18950 10473
rect 15432 10409 15636 10443
rect 15670 10409 15686 10443
rect 15432 10393 15686 10409
rect 17649 10400 18950 10448
rect 20188 10432 20248 10552
rect 14436 9971 14496 9997
rect 14134 9948 14201 9964
rect 14134 9914 14150 9948
rect 14184 9914 14201 9948
rect 14134 9898 14201 9914
rect 14134 9770 14194 9898
rect 14404 9830 14471 9837
rect 14554 9830 14614 9997
rect 14672 9971 14732 9997
rect 14790 9971 14850 9997
rect 14404 9821 14614 9830
rect 14404 9787 14420 9821
rect 14454 9787 14614 9821
rect 14404 9771 14614 9787
rect 14134 9754 14285 9770
rect 14134 9720 14235 9754
rect 14269 9720 14285 9754
rect 14134 9704 14285 9720
rect 14134 9665 14194 9704
rect 14554 9665 14614 9771
rect 14908 9830 14968 9997
rect 15026 9971 15086 9997
rect 15049 9831 15116 9838
rect 15043 9830 15116 9831
rect 14908 9822 15116 9830
rect 14908 9788 15066 9822
rect 15100 9788 15116 9822
rect 14908 9772 15116 9788
rect 14908 9771 15105 9772
rect 14670 9737 14736 9753
rect 14670 9703 14686 9737
rect 14720 9703 14736 9737
rect 14670 9687 14736 9703
rect 14788 9738 14854 9753
rect 14788 9704 14804 9738
rect 14838 9704 14854 9738
rect 14788 9688 14854 9704
rect 14672 9665 14732 9687
rect 14790 9665 14850 9688
rect 14908 9665 14968 9771
rect 15432 9769 15492 10393
rect 17296 9856 17592 9892
rect 17296 9835 17356 9856
rect 17414 9835 17474 9856
rect 17532 9835 17592 9856
rect 17650 9855 17946 9891
rect 17650 9835 17710 9855
rect 17768 9835 17828 9855
rect 17886 9835 17946 9855
rect 18004 9855 18300 9891
rect 18004 9835 18064 9855
rect 18122 9835 18182 9855
rect 18240 9835 18300 9855
rect 15342 9753 15492 9769
rect 15342 9719 15358 9753
rect 15392 9719 15492 9753
rect 15342 9703 15492 9719
rect 15432 9665 15492 9703
rect 11347 9621 11363 9655
rect 11397 9621 11413 9655
rect 11347 9605 11413 9621
rect 11229 9538 11295 9554
rect 11229 9504 11245 9538
rect 11279 9504 11295 9538
rect 11229 9488 11295 9504
rect 11232 9466 11292 9488
rect 8883 9351 8943 9377
rect 6107 9151 6167 9177
rect 6225 9151 6285 9177
rect 6343 9151 6403 9177
rect 6461 9151 6521 9177
rect 8005 9151 8065 9177
rect 8123 9151 8183 9177
rect 8241 9151 8301 9177
rect 8359 9151 8419 9177
rect 12236 9439 12296 9465
rect 11232 9240 11292 9266
rect 13534 9439 13594 9465
rect 14134 9439 14194 9465
rect 18890 9702 18950 10400
rect 19192 10352 19488 10412
rect 19192 10329 19252 10352
rect 19310 10329 19370 10352
rect 19428 10329 19488 10352
rect 19546 10353 19842 10413
rect 20187 10412 20248 10432
rect 19546 10329 19606 10353
rect 19664 10329 19724 10353
rect 19782 10329 19842 10353
rect 20168 10396 20248 10412
rect 20168 10362 20183 10396
rect 20217 10362 20248 10396
rect 20168 10346 20248 10362
rect 20187 10323 20248 10346
rect 20188 10177 20248 10323
rect 20187 10004 20248 10177
rect 19192 9903 19252 9929
rect 19160 9762 19227 9769
rect 19310 9762 19370 9929
rect 19428 9903 19488 9929
rect 19546 9903 19606 9929
rect 19160 9753 19370 9762
rect 19160 9719 19176 9753
rect 19210 9719 19370 9753
rect 19160 9703 19370 9719
rect 18890 9686 19041 9702
rect 18890 9652 18991 9686
rect 19025 9652 19041 9686
rect 18890 9636 19041 9652
rect 17296 9609 17356 9635
rect 17414 9609 17474 9635
rect 17532 9609 17592 9635
rect 17650 9615 17710 9635
rect 17650 9609 17711 9615
rect 17768 9609 17828 9635
rect 17886 9609 17946 9635
rect 15432 9439 15492 9465
rect 17533 9424 17591 9609
rect 17533 9398 17593 9424
rect 17651 9398 17711 9609
rect 18004 9603 18064 9635
rect 18122 9609 18182 9635
rect 18240 9609 18300 9635
rect 18001 9587 18067 9603
rect 18890 9597 18950 9636
rect 19310 9597 19370 9703
rect 19664 9762 19724 9929
rect 19782 9903 19842 9929
rect 19807 9762 19874 9769
rect 19664 9753 19874 9762
rect 19664 9719 19824 9753
rect 19858 9719 19874 9753
rect 19664 9703 19874 9719
rect 19426 9669 19492 9685
rect 19426 9635 19442 9669
rect 19476 9635 19492 9669
rect 19426 9619 19492 9635
rect 19544 9670 19610 9685
rect 19544 9636 19560 9670
rect 19594 9636 19610 9670
rect 19544 9620 19610 9636
rect 19428 9597 19488 9619
rect 19546 9597 19606 9620
rect 19664 9597 19724 9703
rect 20188 9701 20248 10004
rect 20098 9685 20248 9701
rect 20098 9651 20114 9685
rect 20148 9651 20248 9685
rect 20098 9635 20248 9651
rect 20188 9597 20248 9635
rect 20788 9896 20848 10554
rect 21501 10552 22044 10603
rect 22086 10596 22162 10603
rect 22220 10596 22280 10622
rect 24160 10598 24176 10632
rect 24210 10598 24226 10632
rect 22086 10552 22161 10596
rect 24160 10582 24226 10598
rect 24275 10632 24349 10654
rect 24275 10598 24294 10632
rect 24328 10598 24349 10632
rect 26711 10907 27007 10958
rect 26711 10890 26771 10907
rect 26829 10890 26889 10907
rect 26947 10890 27007 10907
rect 27288 10890 27348 10916
rect 27406 10890 27466 10916
rect 27524 10890 27584 10916
rect 36701 11040 36755 11100
rect 37155 11040 37529 11100
rect 37571 11100 37640 11105
rect 37571 11086 38088 11100
rect 37571 11052 37588 11086
rect 37622 11052 38088 11086
rect 37571 11040 38088 11052
rect 38488 11040 38514 11100
rect 36701 10982 36740 11040
rect 37571 11036 37638 11040
rect 28609 10907 28905 10958
rect 36701 10922 36755 10982
rect 37155 10922 37181 10982
rect 28609 10890 28669 10907
rect 28727 10890 28787 10907
rect 28845 10890 28905 10907
rect 32008 10808 32304 10859
rect 32008 10793 32068 10808
rect 32126 10793 32186 10808
rect 32244 10793 32304 10808
rect 32362 10793 32422 10819
rect 32480 10793 32540 10819
rect 32598 10793 32658 10819
rect 25390 10673 25450 10690
rect 25508 10673 25568 10690
rect 25626 10673 25686 10690
rect 25874 10673 25934 10690
rect 25390 10622 25934 10673
rect 25992 10664 26052 10690
rect 26110 10664 26170 10690
rect 26228 10671 26288 10690
rect 26346 10671 26406 10690
rect 26464 10671 26524 10690
rect 26711 10671 26771 10690
rect 26829 10671 26889 10690
rect 21090 10352 21386 10412
rect 21090 10329 21150 10352
rect 21208 10329 21268 10352
rect 21326 10329 21386 10352
rect 21444 10353 21740 10413
rect 21444 10329 21504 10353
rect 21562 10329 21622 10353
rect 21680 10329 21740 10353
rect 22086 10399 22146 10552
rect 24275 10541 24349 10598
rect 25515 10541 25575 10622
rect 26228 10620 26771 10671
rect 26813 10664 26889 10671
rect 26947 10664 27007 10690
rect 27288 10673 27348 10690
rect 27406 10673 27466 10690
rect 27524 10673 27584 10690
rect 27772 10673 27832 10690
rect 26813 10620 26888 10664
rect 27288 10622 27832 10673
rect 27890 10664 27950 10690
rect 28008 10664 28068 10690
rect 28126 10671 28186 10690
rect 28244 10671 28304 10690
rect 28362 10671 28422 10690
rect 28609 10671 28669 10690
rect 28727 10671 28787 10690
rect 24275 10516 25575 10541
rect 24274 10468 25575 10516
rect 26813 10500 26873 10620
rect 22086 10375 22340 10399
rect 22086 10341 22290 10375
rect 22324 10341 22340 10375
rect 22086 10325 22340 10341
rect 21090 9903 21150 9929
rect 20788 9880 20855 9896
rect 20788 9846 20804 9880
rect 20838 9846 20855 9880
rect 20788 9830 20855 9846
rect 20788 9702 20848 9830
rect 21058 9762 21125 9769
rect 21208 9762 21268 9929
rect 21326 9903 21386 9929
rect 21444 9903 21504 9929
rect 21058 9753 21268 9762
rect 21058 9719 21074 9753
rect 21108 9719 21268 9753
rect 21058 9703 21268 9719
rect 20788 9686 20939 9702
rect 20788 9652 20889 9686
rect 20923 9652 20939 9686
rect 20788 9636 20939 9652
rect 20788 9597 20848 9636
rect 21208 9597 21268 9703
rect 21562 9762 21622 9929
rect 21680 9903 21740 9929
rect 21703 9763 21770 9770
rect 21697 9762 21770 9763
rect 21562 9754 21770 9762
rect 21562 9720 21720 9754
rect 21754 9720 21770 9754
rect 21562 9704 21770 9720
rect 21562 9703 21759 9704
rect 21324 9669 21390 9685
rect 21324 9635 21340 9669
rect 21374 9635 21390 9669
rect 21324 9619 21390 9635
rect 21442 9670 21508 9685
rect 21442 9636 21458 9670
rect 21492 9636 21508 9670
rect 21442 9620 21508 9636
rect 21326 9597 21386 9619
rect 21444 9597 21504 9620
rect 21562 9597 21622 9703
rect 22086 9701 22146 10325
rect 23921 9924 24217 9960
rect 23921 9903 23981 9924
rect 24039 9903 24099 9924
rect 24157 9903 24217 9924
rect 24275 9923 24571 9959
rect 24275 9903 24335 9923
rect 24393 9903 24453 9923
rect 24511 9903 24571 9923
rect 24629 9923 24925 9959
rect 24629 9903 24689 9923
rect 24747 9903 24807 9923
rect 24865 9903 24925 9923
rect 25515 9770 25575 10468
rect 25817 10420 26113 10480
rect 25817 10397 25877 10420
rect 25935 10397 25995 10420
rect 26053 10397 26113 10420
rect 26171 10421 26467 10481
rect 26812 10480 26873 10500
rect 26171 10397 26231 10421
rect 26289 10397 26349 10421
rect 26407 10397 26467 10421
rect 26793 10464 26873 10480
rect 26793 10430 26808 10464
rect 26842 10430 26873 10464
rect 26793 10414 26873 10430
rect 26812 10391 26873 10414
rect 26813 10245 26873 10391
rect 26812 10072 26873 10245
rect 25817 9971 25877 9997
rect 25785 9830 25852 9837
rect 25935 9830 25995 9997
rect 26053 9971 26113 9997
rect 26171 9971 26231 9997
rect 25785 9821 25995 9830
rect 25785 9787 25801 9821
rect 25835 9787 25995 9821
rect 25785 9771 25995 9787
rect 25515 9754 25666 9770
rect 25515 9720 25616 9754
rect 25650 9720 25666 9754
rect 25515 9704 25666 9720
rect 21996 9685 22146 9701
rect 21996 9651 22012 9685
rect 22046 9651 22146 9685
rect 23921 9677 23981 9703
rect 24039 9677 24099 9703
rect 24157 9677 24217 9703
rect 24275 9683 24335 9703
rect 24275 9677 24336 9683
rect 24393 9677 24453 9703
rect 24511 9677 24571 9703
rect 21996 9635 22146 9651
rect 22086 9597 22146 9635
rect 18001 9553 18017 9587
rect 18051 9553 18067 9587
rect 18001 9537 18067 9553
rect 17883 9470 17949 9486
rect 17883 9436 17899 9470
rect 17933 9436 17949 9470
rect 17883 9420 17949 9436
rect 17886 9398 17946 9420
rect 12656 9239 12716 9265
rect 12774 9239 12834 9265
rect 12892 9239 12952 9265
rect 13010 9239 13070 9265
rect 14554 9239 14614 9265
rect 14672 9239 14732 9265
rect 14790 9239 14850 9265
rect 14908 9239 14968 9265
rect 10879 9044 10939 9066
rect 10997 9044 11057 9066
rect -2553 8945 -2487 8962
rect 4330 8956 4390 8978
rect 4448 8956 4508 8978
rect -3387 8683 -3336 8870
rect -2553 8911 -2537 8945
rect -2503 8911 -2487 8945
rect -2553 8895 -2487 8911
rect 4327 8940 4393 8956
rect 4327 8906 4343 8940
rect 4377 8906 4393 8940
rect 4327 8890 4393 8906
rect 4445 8940 4511 8956
rect 4445 8906 4461 8940
rect 4495 8906 4511 8940
rect 10876 9028 10942 9044
rect 10876 8994 10892 9028
rect 10926 8994 10942 9028
rect 10876 8978 10942 8994
rect 10994 9028 11060 9044
rect 10994 8994 11010 9028
rect 11044 8994 11060 9028
rect 10994 8978 11060 8994
rect 18890 9371 18950 9397
rect 17886 9172 17946 9198
rect 20188 9371 20248 9397
rect 20788 9371 20848 9397
rect 24158 9492 24216 9677
rect 24158 9466 24218 9492
rect 24276 9466 24336 9677
rect 24629 9671 24689 9703
rect 24747 9677 24807 9703
rect 24865 9677 24925 9703
rect 24626 9655 24692 9671
rect 25515 9665 25575 9704
rect 25935 9665 25995 9771
rect 26289 9830 26349 9997
rect 26407 9971 26467 9997
rect 26432 9830 26499 9837
rect 26289 9821 26499 9830
rect 26289 9787 26449 9821
rect 26483 9787 26499 9821
rect 26289 9771 26499 9787
rect 26051 9737 26117 9753
rect 26051 9703 26067 9737
rect 26101 9703 26117 9737
rect 26051 9687 26117 9703
rect 26169 9738 26235 9753
rect 26169 9704 26185 9738
rect 26219 9704 26235 9738
rect 26169 9688 26235 9704
rect 26053 9665 26113 9687
rect 26171 9665 26231 9688
rect 26289 9665 26349 9771
rect 26813 9769 26873 10072
rect 26723 9753 26873 9769
rect 26723 9719 26739 9753
rect 26773 9719 26873 9753
rect 26723 9703 26873 9719
rect 26813 9665 26873 9703
rect 27413 9964 27473 10622
rect 28126 10620 28669 10671
rect 28711 10664 28787 10671
rect 28845 10664 28905 10690
rect 28711 10620 28786 10664
rect 27715 10420 28011 10480
rect 27715 10397 27775 10420
rect 27833 10397 27893 10420
rect 27951 10397 28011 10420
rect 28069 10421 28365 10481
rect 28069 10397 28129 10421
rect 28187 10397 28247 10421
rect 28305 10397 28365 10421
rect 28711 10467 28771 10620
rect 31524 10593 31584 10619
rect 31642 10593 31702 10619
rect 31760 10593 31820 10619
rect 28711 10443 28965 10467
rect 28711 10409 28915 10443
rect 28949 10409 28965 10443
rect 28711 10393 28965 10409
rect 36701 10685 36755 10745
rect 37155 10685 37181 10745
rect 32845 10610 33141 10661
rect 32845 10593 32905 10610
rect 32963 10593 33023 10610
rect 33081 10593 33141 10610
rect 33317 10611 33613 10647
rect 33317 10590 33377 10611
rect 33435 10590 33495 10611
rect 33553 10590 33613 10611
rect 33671 10610 33967 10646
rect 33671 10590 33731 10610
rect 33789 10590 33849 10610
rect 33907 10590 33967 10610
rect 34025 10610 34321 10646
rect 34025 10590 34085 10610
rect 34143 10590 34203 10610
rect 34261 10590 34321 10610
rect 36701 10627 36740 10685
rect 37571 10627 37628 11036
rect 38569 10904 38620 11213
rect 27715 9971 27775 9997
rect 27413 9948 27480 9964
rect 27413 9914 27429 9948
rect 27463 9914 27480 9948
rect 27413 9898 27480 9914
rect 27413 9770 27473 9898
rect 27683 9830 27750 9837
rect 27833 9830 27893 9997
rect 27951 9971 28011 9997
rect 28069 9971 28129 9997
rect 27683 9821 27893 9830
rect 27683 9787 27699 9821
rect 27733 9787 27893 9821
rect 27683 9771 27893 9787
rect 27413 9754 27564 9770
rect 27413 9720 27514 9754
rect 27548 9720 27564 9754
rect 27413 9704 27564 9720
rect 27413 9665 27473 9704
rect 27833 9665 27893 9771
rect 28187 9830 28247 9997
rect 28305 9971 28365 9997
rect 28328 9831 28395 9838
rect 28322 9830 28395 9831
rect 28187 9822 28395 9830
rect 28187 9788 28345 9822
rect 28379 9788 28395 9822
rect 28187 9772 28395 9788
rect 28187 9771 28384 9772
rect 27949 9737 28015 9753
rect 27949 9703 27965 9737
rect 27999 9703 28015 9737
rect 27949 9687 28015 9703
rect 28067 9738 28133 9753
rect 28067 9704 28083 9738
rect 28117 9704 28133 9738
rect 28067 9688 28133 9704
rect 27951 9665 28011 9687
rect 28069 9665 28129 9688
rect 28187 9665 28247 9771
rect 28711 9769 28771 10393
rect 31524 10376 31584 10393
rect 31642 10376 31702 10393
rect 31760 10376 31820 10393
rect 32008 10376 32068 10393
rect 31524 10325 32068 10376
rect 32126 10367 32186 10393
rect 32244 10367 32304 10393
rect 32362 10374 32422 10393
rect 32480 10374 32540 10393
rect 32598 10374 32658 10393
rect 32845 10374 32905 10393
rect 32963 10374 33023 10393
rect 28621 9753 28771 9769
rect 28621 9719 28637 9753
rect 28671 9719 28771 9753
rect 31649 10121 31709 10325
rect 32362 10323 32905 10374
rect 32947 10367 33023 10374
rect 33081 10367 33141 10393
rect 36701 10567 36755 10627
rect 37155 10567 37628 10627
rect 37840 10844 38088 10904
rect 38288 10844 38620 10904
rect 36701 10509 36740 10567
rect 36701 10449 36755 10509
rect 37155 10449 37181 10509
rect 32947 10323 33022 10367
rect 33317 10364 33377 10390
rect 33435 10364 33495 10390
rect 33553 10364 33613 10390
rect 33671 10370 33731 10390
rect 33671 10364 33732 10370
rect 33789 10364 33849 10390
rect 33907 10364 33967 10390
rect 32947 10241 33007 10323
rect 32947 10223 33181 10241
rect 32947 10189 33130 10223
rect 33164 10189 33181 10223
rect 31951 10123 32247 10183
rect 31649 10104 31780 10121
rect 31649 10070 31730 10104
rect 31764 10070 31780 10104
rect 31951 10100 32011 10123
rect 32069 10100 32129 10123
rect 32187 10100 32247 10123
rect 32305 10124 32601 10184
rect 32305 10100 32365 10124
rect 32423 10100 32483 10124
rect 32541 10100 32601 10124
rect 32947 10173 33181 10189
rect 33554 10179 33612 10364
rect 31649 10053 31780 10070
rect 28621 9703 28771 9719
rect 28711 9665 28771 9703
rect 24626 9621 24642 9655
rect 24676 9621 24692 9655
rect 24626 9605 24692 9621
rect 24508 9538 24574 9554
rect 24508 9504 24524 9538
rect 24558 9504 24574 9538
rect 24508 9488 24574 9504
rect 24511 9466 24571 9488
rect 22086 9371 22146 9397
rect 19310 9171 19370 9197
rect 19428 9171 19488 9197
rect 19546 9171 19606 9197
rect 19664 9171 19724 9197
rect 21208 9171 21268 9197
rect 21326 9171 21386 9197
rect 21444 9171 21504 9197
rect 21562 9171 21622 9197
rect 25515 9439 25575 9465
rect 24511 9240 24571 9266
rect 26813 9439 26873 9465
rect 27413 9439 27473 9465
rect 29709 9506 30005 9542
rect 29709 9485 29769 9506
rect 29827 9485 29887 9506
rect 29945 9485 30005 9506
rect 30063 9505 30359 9541
rect 30063 9485 30123 9505
rect 30181 9485 30241 9505
rect 30299 9485 30359 9505
rect 30417 9505 30713 9541
rect 30417 9485 30477 9505
rect 30535 9485 30595 9505
rect 30653 9485 30713 9505
rect 28711 9439 28771 9465
rect 31649 9473 31709 10053
rect 31951 9674 32011 9700
rect 31919 9533 31986 9540
rect 32069 9533 32129 9700
rect 32187 9674 32247 9700
rect 32305 9674 32365 9700
rect 31919 9524 32129 9533
rect 31919 9490 31935 9524
rect 31969 9490 32129 9524
rect 31919 9474 32129 9490
rect 31649 9457 31800 9473
rect 31649 9423 31750 9457
rect 31784 9423 31800 9457
rect 31649 9407 31800 9423
rect 31649 9368 31709 9407
rect 32069 9368 32129 9474
rect 32423 9533 32483 9700
rect 32541 9674 32601 9700
rect 32566 9533 32633 9540
rect 32423 9524 32633 9533
rect 32423 9490 32583 9524
rect 32617 9490 32633 9524
rect 32423 9474 32633 9490
rect 32185 9440 32251 9456
rect 32185 9406 32201 9440
rect 32235 9406 32251 9440
rect 32185 9390 32251 9406
rect 32303 9441 32369 9456
rect 32303 9407 32319 9441
rect 32353 9407 32369 9441
rect 32303 9391 32369 9407
rect 32187 9368 32247 9390
rect 32305 9368 32365 9391
rect 32423 9368 32483 9474
rect 32947 9472 33007 10173
rect 33554 10153 33614 10179
rect 33672 10153 33732 10364
rect 34025 10358 34085 10390
rect 34143 10364 34203 10390
rect 34261 10364 34321 10390
rect 34022 10342 34088 10358
rect 34022 10308 34038 10342
rect 34072 10308 34088 10342
rect 34022 10292 34088 10308
rect 33904 10225 33970 10241
rect 33904 10191 33920 10225
rect 33954 10191 33970 10225
rect 33904 10175 33970 10191
rect 36900 10212 36955 10272
rect 37155 10212 37181 10272
rect 33907 10153 33967 10175
rect 36900 10154 36939 10212
rect 36900 10094 36955 10154
rect 37155 10094 37181 10154
rect 37301 10130 37367 10146
rect 37301 10096 37317 10130
rect 37351 10096 37367 10130
rect 36900 10036 36939 10094
rect 37301 10080 37367 10096
rect 37304 10036 37364 10080
rect 37840 10036 37885 10844
rect 36900 9976 36955 10036
rect 37155 9976 37885 10036
rect 33907 9927 33967 9953
rect 33554 9731 33614 9753
rect 33672 9731 33732 9753
rect 33551 9715 33617 9731
rect 33551 9681 33567 9715
rect 33601 9681 33617 9715
rect 33551 9665 33617 9681
rect 33669 9715 33735 9731
rect 33669 9681 33685 9715
rect 33719 9681 33735 9715
rect 33669 9665 33735 9681
rect 32857 9456 33007 9472
rect 32857 9422 32873 9456
rect 32907 9422 33007 9456
rect 32857 9406 33007 9422
rect 32947 9368 33007 9406
rect 25935 9239 25995 9265
rect 26053 9239 26113 9265
rect 26171 9239 26231 9265
rect 26289 9239 26349 9265
rect 27833 9239 27893 9265
rect 27951 9239 28011 9265
rect 28069 9239 28129 9265
rect 28187 9239 28247 9265
rect 29709 9259 29769 9285
rect 29827 9259 29887 9285
rect 29945 9259 30005 9285
rect 30063 9265 30123 9285
rect 30063 9259 30124 9265
rect 30181 9259 30241 9285
rect 30299 9259 30359 9285
rect 17533 8976 17593 8998
rect 17651 8976 17711 8998
rect 4445 8890 4511 8906
rect 17530 8960 17596 8976
rect 17530 8926 17546 8960
rect 17580 8926 17596 8960
rect 17530 8910 17596 8926
rect 17648 8960 17714 8976
rect 17648 8926 17664 8960
rect 17698 8926 17714 8960
rect 24158 9044 24218 9066
rect 24276 9044 24336 9066
rect 24155 9028 24221 9044
rect 24155 8994 24171 9028
rect 24205 8994 24221 9028
rect 24155 8978 24221 8994
rect 24273 9028 24339 9044
rect 24273 8994 24289 9028
rect 24323 8994 24339 9028
rect 29946 9074 30004 9259
rect 29946 9048 30006 9074
rect 30064 9048 30124 9259
rect 30417 9253 30477 9285
rect 30535 9259 30595 9285
rect 30653 9259 30713 9285
rect 30414 9237 30480 9253
rect 30414 9203 30430 9237
rect 30464 9203 30480 9237
rect 30414 9187 30480 9203
rect 31649 9142 31709 9168
rect 30296 9120 30362 9136
rect 30296 9086 30312 9120
rect 30346 9086 30362 9120
rect 30296 9070 30362 9086
rect 30299 9048 30359 9070
rect 24273 8978 24339 8994
rect 17648 8910 17714 8926
rect -3674 8623 -3606 8683
rect -3406 8623 -3336 8683
rect -2485 8655 -2419 8671
rect -3249 8633 -3195 8649
rect -3674 8565 -3623 8623
rect -3249 8599 -3239 8633
rect -3205 8599 -3195 8633
rect -3249 8581 -3195 8599
rect -2485 8621 -2469 8655
rect -2435 8621 -2419 8655
rect 36900 9276 36955 9336
rect 37155 9277 37885 9336
rect 37155 9276 37458 9277
rect 36900 9218 36939 9276
rect 37441 9219 37458 9276
rect 37513 9276 37885 9277
rect 37513 9219 37528 9276
rect 32947 9142 33007 9168
rect 36900 9158 36955 9218
rect 37155 9158 37181 9218
rect 37441 9200 37528 9219
rect 36900 9100 36939 9158
rect 36900 9040 36955 9100
rect 37155 9040 37181 9100
rect 32069 8942 32129 8968
rect 32187 8942 32247 8968
rect 32305 8942 32365 8968
rect 32423 8942 32483 8968
rect 30299 8822 30359 8848
rect 36701 8835 36755 8895
rect 37155 8835 37181 8895
rect 36701 8777 36740 8835
rect 36701 8717 36755 8777
rect 37155 8717 37630 8777
rect 36701 8659 36740 8717
rect -2485 8581 -2419 8621
rect 29946 8626 30006 8648
rect 30064 8626 30124 8648
rect 29943 8610 30009 8626
rect -3387 8565 -2381 8581
rect -3674 8505 -3606 8565
rect -3406 8521 -2381 8565
rect -2181 8521 -2155 8581
rect 29943 8576 29959 8610
rect 29993 8576 30009 8610
rect 29943 8560 30009 8576
rect 30061 8610 30127 8626
rect 30061 8576 30077 8610
rect 30111 8576 30127 8610
rect 36701 8599 36755 8659
rect 37155 8599 37181 8659
rect 30061 8560 30127 8576
rect -3406 8506 -3336 8521
rect -3406 8505 -3380 8506
rect -3674 8447 -3623 8505
rect -3674 8387 -3606 8447
rect -3406 8387 -3380 8447
rect 36701 8368 36755 8428
rect 37155 8368 37181 8428
rect 36701 8310 36740 8368
rect 36701 8250 36755 8310
rect 37155 8309 37181 8310
rect 37342 8309 37408 8312
rect 37155 8296 37408 8309
rect 37155 8262 37358 8296
rect 37392 8262 37408 8296
rect 37155 8250 37408 8262
rect 37573 8310 37630 8717
rect 37840 8502 37885 9276
rect 37840 8442 38088 8502
rect 38288 8442 38314 8502
rect 37729 8310 37808 8321
rect 37573 8308 38088 8310
rect 37573 8250 37742 8308
rect 37797 8250 38088 8308
rect 38488 8250 38514 8310
rect 36701 8192 36740 8250
rect 37341 8246 37408 8250
rect 37729 8240 37808 8250
rect 37442 8192 37529 8209
rect 36701 8132 36755 8192
rect 37155 8132 37181 8192
rect 37442 8190 38088 8192
rect 37442 8132 37457 8190
rect 37512 8132 38088 8190
rect 38488 8132 38514 8192
rect 37442 8114 37529 8132
rect -3059 7958 -2999 7974
rect -3632 7875 -3606 7935
rect -3406 7875 -3338 7935
rect -3389 7817 -3338 7875
rect -3632 7757 -3606 7817
rect -3406 7810 -3338 7817
rect -3059 7924 -3045 7958
rect -3011 7924 -2999 7958
rect 36701 8014 36755 8074
rect 37155 8014 37181 8074
rect 36701 7956 36740 8014
rect 37480 7956 37529 8114
rect 37962 8074 38028 8077
rect 38561 8119 38627 8135
rect 38561 8085 38577 8119
rect 38611 8085 38627 8119
rect 37962 8061 38088 8074
rect 37962 8027 37978 8061
rect 38012 8027 38088 8061
rect 37962 8014 38088 8027
rect 38488 8014 38514 8074
rect 38561 8069 38627 8085
rect 37962 8011 38028 8014
rect -3059 7810 -2999 7924
rect 36701 7896 36755 7956
rect 37155 7896 37529 7956
rect 37571 7956 37640 7961
rect 37571 7942 38088 7956
rect 37571 7908 37588 7942
rect 37622 7908 38088 7942
rect 37571 7896 38088 7908
rect 38488 7896 38514 7956
rect 36701 7838 36740 7896
rect 37571 7892 37638 7896
rect -3406 7757 -2381 7810
rect -3389 7750 -2381 7757
rect -2181 7750 -2155 7810
rect -3389 7699 -3338 7750
rect -3632 7639 -3606 7699
rect -3406 7639 -3338 7699
rect -2486 7709 -2420 7750
rect -2486 7675 -2470 7709
rect -2436 7675 -2420 7709
rect -2486 7659 -2420 7675
rect -3389 7451 -3338 7639
rect -2553 7524 -2487 7540
rect -3872 7391 -3806 7451
rect -3406 7391 -3338 7451
rect -3196 7448 -3113 7508
rect -2713 7448 -2687 7508
rect -2553 7490 -2537 7524
rect -2503 7490 -2487 7524
rect -2553 7473 -2487 7490
rect 1167 7494 1463 7530
rect 1167 7473 1227 7494
rect 1285 7473 1345 7494
rect 1403 7473 1463 7494
rect 1521 7493 1817 7529
rect 1521 7473 1581 7493
rect 1639 7473 1699 7493
rect 1757 7473 1817 7493
rect 1875 7493 2171 7529
rect 1875 7473 1935 7493
rect 1993 7473 2053 7493
rect 2111 7473 2171 7493
rect 6224 7525 6290 7541
rect 7354 7531 7420 7547
rect 6224 7491 6240 7525
rect 6274 7518 6290 7525
rect 6274 7491 6799 7518
rect 6224 7475 6799 7491
rect 7354 7497 7370 7531
rect 7404 7522 7420 7531
rect 7404 7497 7941 7522
rect 7354 7479 7941 7497
rect -3872 7333 -3821 7391
rect -3196 7390 -3136 7448
rect -2546 7390 -2487 7473
rect -3872 7273 -3806 7333
rect -3406 7273 -3380 7333
rect -3196 7330 -3113 7390
rect -2713 7330 -2381 7390
rect -1981 7330 -1955 7390
rect -3872 7215 -3821 7273
rect -3196 7272 -3136 7330
rect -2469 7272 -2403 7274
rect -3872 7155 -3806 7215
rect -3406 7155 -3380 7215
rect -3196 7212 -3113 7272
rect -2713 7212 -2687 7272
rect -2469 7258 -2381 7272
rect -2469 7224 -2453 7258
rect -2419 7224 -2381 7258
rect -2469 7212 -2381 7224
rect -1981 7212 -1955 7272
rect 6755 7423 6799 7475
rect 7897 7427 7941 7479
rect 12775 7523 12841 7539
rect 13905 7529 13971 7545
rect 12775 7489 12791 7523
rect 12825 7516 12841 7523
rect 12825 7489 13350 7516
rect 12775 7473 13350 7489
rect 13905 7495 13921 7529
rect 13955 7520 13971 7529
rect 13955 7495 14492 7520
rect 13905 7477 14492 7495
rect 6224 7407 6697 7423
rect 6224 7373 6240 7407
rect 6274 7382 6697 7407
rect 6274 7381 6461 7382
rect 6274 7373 6290 7381
rect 6224 7357 6290 7373
rect 6401 7361 6461 7381
rect 6519 7361 6579 7382
rect 6637 7361 6697 7382
rect 6755 7382 7051 7423
rect 6755 7361 6815 7382
rect 6873 7361 6933 7382
rect 6991 7361 7051 7382
rect 7354 7411 7839 7427
rect 7354 7377 7370 7411
rect 7404 7386 7839 7411
rect 7404 7385 7603 7386
rect 7404 7377 7420 7385
rect 7354 7361 7420 7377
rect 7543 7365 7603 7385
rect 7661 7365 7721 7386
rect 7779 7365 7839 7386
rect 7897 7386 8193 7427
rect 13306 7421 13350 7473
rect 14448 7425 14492 7477
rect 19430 7524 19496 7540
rect 20560 7530 20626 7546
rect 19430 7490 19446 7524
rect 19480 7517 19496 7524
rect 19480 7490 20005 7517
rect 19430 7474 20005 7490
rect 20560 7496 20576 7530
rect 20610 7521 20626 7530
rect 20610 7496 21147 7521
rect 20560 7478 21147 7496
rect 7897 7365 7957 7386
rect 8015 7365 8075 7386
rect 8133 7365 8193 7386
rect 12775 7405 13248 7421
rect 12775 7371 12791 7405
rect 12825 7380 13248 7405
rect 12825 7379 13012 7380
rect 12825 7371 12841 7379
rect 4076 7310 4372 7346
rect 4076 7289 4136 7310
rect 4194 7289 4254 7310
rect 4312 7289 4372 7310
rect 4430 7309 4726 7345
rect 4430 7289 4490 7309
rect 4548 7289 4608 7309
rect 4666 7289 4726 7309
rect 4784 7309 5080 7345
rect 4784 7289 4844 7309
rect 4902 7289 4962 7309
rect 5020 7289 5080 7309
rect 1167 7247 1227 7273
rect 1285 7247 1345 7273
rect 1403 7247 1463 7273
rect 1521 7253 1581 7273
rect 1521 7247 1582 7253
rect 1639 7247 1699 7273
rect 1757 7247 1817 7273
rect -2469 7208 -2403 7212
rect -2469 7154 -2404 7156
rect -3832 7037 -3806 7097
rect -3406 7037 -3336 7097
rect -3387 6979 -3336 7037
rect -3832 6919 -3806 6979
rect -3406 6919 -3336 6979
rect -3387 6861 -3336 6919
rect -3832 6801 -3806 6861
rect -3406 6801 -3336 6861
rect -3197 7094 -3113 7154
rect -2713 7094 -2687 7154
rect -2469 7140 -2381 7154
rect -2469 7106 -2454 7140
rect -2420 7106 -2381 7140
rect -2469 7094 -2381 7106
rect -1981 7094 -1955 7154
rect -3197 7036 -3137 7094
rect -2469 7090 -2404 7094
rect 1404 7062 1462 7247
rect 1404 7036 1464 7062
rect 1522 7036 1582 7247
rect 1875 7241 1935 7273
rect 1993 7247 2053 7273
rect 2111 7247 2171 7273
rect 1872 7225 1938 7241
rect 1872 7191 1888 7225
rect 1922 7191 1938 7225
rect 1872 7175 1938 7191
rect 1754 7108 1820 7124
rect 1754 7074 1770 7108
rect 1804 7074 1820 7108
rect 1754 7058 1820 7074
rect 4076 7063 4136 7089
rect 4194 7063 4254 7089
rect 4312 7063 4372 7089
rect 4430 7069 4490 7089
rect 4430 7063 4491 7069
rect 4548 7063 4608 7089
rect 4666 7063 4726 7089
rect 1757 7036 1817 7058
rect -3197 6976 -3113 7036
rect -2713 6976 -2381 7036
rect -1981 6976 -1955 7036
rect -3197 6918 -3137 6976
rect -3197 6858 -3113 6918
rect -2713 6858 -2687 6918
rect -2546 6893 -2487 6976
rect -2553 6876 -2487 6893
rect -3387 6614 -3336 6801
rect -2553 6842 -2537 6876
rect -2503 6842 -2487 6876
rect -2553 6826 -2487 6842
rect 4313 6878 4371 7063
rect 4313 6852 4373 6878
rect 4431 6852 4491 7063
rect 4784 7057 4844 7089
rect 4902 7063 4962 7089
rect 5020 7063 5080 7089
rect 4781 7041 4847 7057
rect 4781 7007 4797 7041
rect 4831 7007 4847 7041
rect 4781 6991 4847 7007
rect 12775 7355 12841 7371
rect 12952 7359 13012 7379
rect 13070 7359 13130 7380
rect 13188 7359 13248 7380
rect 13306 7380 13602 7421
rect 13306 7359 13366 7380
rect 13424 7359 13484 7380
rect 13542 7359 13602 7380
rect 13905 7409 14390 7425
rect 13905 7375 13921 7409
rect 13955 7384 14390 7409
rect 13955 7383 14154 7384
rect 13955 7375 13971 7383
rect 13905 7359 13971 7375
rect 14094 7363 14154 7383
rect 14212 7363 14272 7384
rect 14330 7363 14390 7384
rect 14448 7384 14744 7425
rect 19961 7422 20005 7474
rect 21103 7426 21147 7478
rect 26052 7525 26118 7541
rect 36701 7778 36755 7838
rect 37155 7778 37181 7838
rect 27182 7531 27248 7547
rect 26052 7491 26068 7525
rect 26102 7518 26118 7525
rect 26102 7491 26627 7518
rect 26052 7475 26627 7491
rect 27182 7497 27198 7531
rect 27232 7522 27248 7531
rect 29780 7586 30076 7622
rect 29780 7565 29840 7586
rect 29898 7565 29958 7586
rect 30016 7565 30076 7586
rect 30134 7585 30430 7621
rect 30134 7565 30194 7585
rect 30252 7565 30312 7585
rect 30370 7565 30430 7585
rect 30488 7585 30784 7621
rect 30488 7565 30548 7585
rect 30606 7565 30666 7585
rect 30724 7565 30784 7585
rect 27232 7497 27769 7522
rect 27182 7479 27769 7497
rect 14448 7363 14508 7384
rect 14566 7363 14626 7384
rect 14684 7363 14744 7384
rect 19430 7406 19903 7422
rect 19430 7372 19446 7406
rect 19480 7381 19903 7406
rect 19480 7380 19667 7381
rect 19480 7372 19496 7380
rect 10627 7308 10923 7344
rect 10627 7287 10687 7308
rect 10745 7287 10805 7308
rect 10863 7287 10923 7308
rect 10981 7307 11277 7343
rect 10981 7287 11041 7307
rect 11099 7287 11159 7307
rect 11217 7287 11277 7307
rect 11335 7307 11631 7343
rect 11335 7287 11395 7307
rect 11453 7287 11513 7307
rect 11571 7287 11631 7307
rect 10627 7061 10687 7087
rect 10745 7061 10805 7087
rect 10863 7061 10923 7087
rect 10981 7067 11041 7087
rect 10981 7061 11042 7067
rect 11099 7061 11159 7087
rect 11217 7061 11277 7087
rect 6401 6944 6461 6961
rect 4663 6924 4729 6940
rect 4663 6890 4679 6924
rect 4713 6890 4729 6924
rect 4663 6874 4729 6890
rect 4666 6852 4726 6874
rect 6401 6855 6462 6944
rect 6519 6935 6579 6961
rect 6637 6935 6697 6961
rect 1757 6810 1817 6836
rect 1404 6614 1464 6636
rect 1522 6614 1582 6636
rect -3674 6554 -3606 6614
rect -3406 6554 -3336 6614
rect -2485 6586 -2419 6602
rect -3249 6564 -3195 6580
rect -3674 6496 -3623 6554
rect -3249 6530 -3239 6564
rect -3205 6530 -3195 6564
rect -3249 6512 -3195 6530
rect -2485 6552 -2469 6586
rect -2435 6552 -2419 6586
rect 1401 6598 1467 6614
rect -2485 6512 -2419 6552
rect 1401 6564 1417 6598
rect 1451 6564 1467 6598
rect 1401 6548 1467 6564
rect 1519 6598 1585 6614
rect 1519 6564 1535 6598
rect 1569 6564 1585 6598
rect 1519 6548 1585 6564
rect -3387 6496 -2381 6512
rect -3674 6436 -3606 6496
rect -3406 6452 -2381 6496
rect -2181 6452 -2155 6512
rect -3406 6437 -3336 6452
rect -3406 6436 -3380 6437
rect -3674 6378 -3623 6436
rect 6311 6802 6462 6855
rect 4666 6626 4726 6652
rect 6311 6578 6371 6802
rect 6755 6760 6815 6961
rect 6873 6935 6933 6961
rect 6991 6935 7051 6961
rect 7543 6948 7603 6965
rect 7543 6859 7604 6948
rect 7661 6939 7721 6965
rect 7779 6939 7839 6965
rect 6429 6709 6815 6760
rect 7453 6806 7604 6859
rect 6429 6578 6489 6709
rect 6544 6651 6610 6667
rect 6544 6617 6560 6651
rect 6594 6617 6610 6651
rect 6544 6601 6610 6617
rect 6547 6578 6607 6601
rect 6830 6578 6890 6604
rect 6948 6578 7008 6604
rect 7066 6578 7126 6604
rect 7453 6582 7513 6806
rect 7897 6764 7957 6965
rect 8015 6939 8075 6965
rect 8133 6939 8193 6965
rect 10864 6876 10922 7061
rect 10864 6850 10924 6876
rect 10982 6850 11042 7061
rect 11335 7055 11395 7087
rect 11453 7061 11513 7087
rect 11571 7061 11631 7087
rect 11332 7039 11398 7055
rect 11332 7005 11348 7039
rect 11382 7005 11398 7039
rect 11332 6989 11398 7005
rect 19430 7356 19496 7372
rect 19607 7360 19667 7380
rect 19725 7360 19785 7381
rect 19843 7360 19903 7381
rect 19961 7381 20257 7422
rect 19961 7360 20021 7381
rect 20079 7360 20139 7381
rect 20197 7360 20257 7381
rect 20560 7410 21045 7426
rect 20560 7376 20576 7410
rect 20610 7385 21045 7410
rect 20610 7384 20809 7385
rect 20610 7376 20626 7384
rect 20560 7360 20626 7376
rect 20749 7364 20809 7384
rect 20867 7364 20927 7385
rect 20985 7364 21045 7385
rect 21103 7385 21399 7426
rect 26583 7423 26627 7475
rect 27725 7427 27769 7479
rect 21103 7364 21163 7385
rect 21221 7364 21281 7385
rect 21339 7364 21399 7385
rect 26052 7407 26525 7423
rect 26052 7373 26068 7407
rect 26102 7382 26525 7407
rect 26102 7381 26289 7382
rect 26102 7373 26118 7381
rect 17282 7309 17578 7345
rect 17282 7288 17342 7309
rect 17400 7288 17460 7309
rect 17518 7288 17578 7309
rect 17636 7308 17932 7344
rect 17636 7288 17696 7308
rect 17754 7288 17814 7308
rect 17872 7288 17932 7308
rect 17990 7308 18286 7344
rect 17990 7288 18050 7308
rect 18108 7288 18168 7308
rect 18226 7288 18286 7308
rect 17282 7062 17342 7088
rect 17400 7062 17460 7088
rect 17518 7062 17578 7088
rect 17636 7068 17696 7088
rect 17636 7062 17697 7068
rect 17754 7062 17814 7088
rect 17872 7062 17932 7088
rect 12952 6942 13012 6959
rect 11214 6922 11280 6938
rect 11214 6888 11230 6922
rect 11264 6888 11280 6922
rect 11214 6872 11280 6888
rect 11217 6850 11277 6872
rect 12952 6853 13013 6942
rect 13070 6933 13130 6959
rect 13188 6933 13248 6959
rect 7571 6713 7957 6764
rect 7571 6582 7631 6713
rect 7686 6655 7752 6671
rect 7686 6621 7702 6655
rect 7736 6621 7752 6655
rect 7686 6605 7752 6621
rect 7689 6582 7749 6605
rect 7972 6582 8032 6608
rect 8090 6582 8150 6608
rect 8208 6582 8268 6608
rect 4313 6430 4373 6452
rect 4431 6430 4491 6452
rect 4310 6414 4376 6430
rect 4310 6380 4326 6414
rect 4360 6380 4376 6414
rect -3674 6318 -3606 6378
rect -3406 6318 -3380 6378
rect 4310 6364 4376 6380
rect 4428 6414 4494 6430
rect 4428 6380 4444 6414
rect 4478 6380 4494 6414
rect 4428 6364 4494 6380
rect 12862 6800 13013 6853
rect 11217 6624 11277 6650
rect 12862 6576 12922 6800
rect 13306 6758 13366 6959
rect 13424 6933 13484 6959
rect 13542 6933 13602 6959
rect 14094 6946 14154 6963
rect 14094 6857 14155 6946
rect 14212 6937 14272 6963
rect 14330 6937 14390 6963
rect 12980 6707 13366 6758
rect 14004 6804 14155 6857
rect 12980 6576 13040 6707
rect 13095 6649 13161 6665
rect 13095 6615 13111 6649
rect 13145 6615 13161 6649
rect 13095 6599 13161 6615
rect 13098 6576 13158 6599
rect 13381 6576 13441 6602
rect 13499 6576 13559 6602
rect 13617 6576 13677 6602
rect 14004 6580 14064 6804
rect 14448 6762 14508 6963
rect 14566 6937 14626 6963
rect 14684 6937 14744 6963
rect 17519 6877 17577 7062
rect 17519 6851 17579 6877
rect 17637 6851 17697 7062
rect 17990 7056 18050 7088
rect 18108 7062 18168 7088
rect 18226 7062 18286 7088
rect 17987 7040 18053 7056
rect 17987 7006 18003 7040
rect 18037 7006 18053 7040
rect 17987 6990 18053 7006
rect 26052 7357 26118 7373
rect 26229 7361 26289 7381
rect 26347 7361 26407 7382
rect 26465 7361 26525 7382
rect 26583 7382 26879 7423
rect 26583 7361 26643 7382
rect 26701 7361 26761 7382
rect 26819 7361 26879 7382
rect 27182 7411 27667 7427
rect 27182 7377 27198 7411
rect 27232 7386 27667 7411
rect 27232 7385 27431 7386
rect 27232 7377 27248 7385
rect 27182 7361 27248 7377
rect 27371 7365 27431 7385
rect 27489 7365 27549 7386
rect 27607 7365 27667 7386
rect 27725 7386 28021 7427
rect 27725 7365 27785 7386
rect 27843 7365 27903 7386
rect 27961 7365 28021 7386
rect 36701 7541 36755 7601
rect 37155 7541 37181 7601
rect 36701 7483 36740 7541
rect 37571 7483 37628 7892
rect 38569 7760 38620 8069
rect 36701 7423 36755 7483
rect 37155 7423 37628 7483
rect 37840 7700 38088 7760
rect 38288 7700 38620 7760
rect 36701 7365 36740 7423
rect 23904 7310 24200 7346
rect 23904 7289 23964 7310
rect 24022 7289 24082 7310
rect 24140 7289 24200 7310
rect 24258 7309 24554 7345
rect 24258 7289 24318 7309
rect 24376 7289 24436 7309
rect 24494 7289 24554 7309
rect 24612 7309 24908 7345
rect 24612 7289 24672 7309
rect 24730 7289 24790 7309
rect 24848 7289 24908 7309
rect 23904 7063 23964 7089
rect 24022 7063 24082 7089
rect 24140 7063 24200 7089
rect 24258 7069 24318 7089
rect 24258 7063 24319 7069
rect 24376 7063 24436 7089
rect 24494 7063 24554 7089
rect 19607 6943 19667 6960
rect 17869 6923 17935 6939
rect 17869 6889 17885 6923
rect 17919 6889 17935 6923
rect 17869 6873 17935 6889
rect 17872 6851 17932 6873
rect 19607 6854 19668 6943
rect 19725 6934 19785 6960
rect 19843 6934 19903 6960
rect 14122 6711 14508 6762
rect 14122 6580 14182 6711
rect 14237 6653 14303 6669
rect 14237 6619 14253 6653
rect 14287 6619 14303 6653
rect 14237 6603 14303 6619
rect 14240 6580 14300 6603
rect 14523 6580 14583 6606
rect 14641 6580 14701 6606
rect 14759 6580 14819 6606
rect 10864 6428 10924 6450
rect 10982 6428 11042 6450
rect 10861 6412 10927 6428
rect 6311 6352 6371 6378
rect 6429 6352 6489 6378
rect 6547 6346 6607 6378
rect 6830 6346 6890 6378
rect 6948 6346 7008 6378
rect 7066 6346 7126 6378
rect 7453 6356 7513 6382
rect 7571 6356 7631 6382
rect 6547 6305 7126 6346
rect 7689 6350 7749 6382
rect 7972 6350 8032 6382
rect 8090 6350 8150 6382
rect 8208 6350 8268 6382
rect 10861 6378 10877 6412
rect 10911 6378 10927 6412
rect 10861 6362 10927 6378
rect 10979 6412 11045 6428
rect 10979 6378 10995 6412
rect 11029 6378 11045 6412
rect 10979 6362 11045 6378
rect 19517 6801 19668 6854
rect 17872 6625 17932 6651
rect 19517 6577 19577 6801
rect 19961 6759 20021 6960
rect 20079 6934 20139 6960
rect 20197 6934 20257 6960
rect 20749 6947 20809 6964
rect 20749 6858 20810 6947
rect 20867 6938 20927 6964
rect 20985 6938 21045 6964
rect 19635 6708 20021 6759
rect 20659 6805 20810 6858
rect 19635 6577 19695 6708
rect 19750 6650 19816 6666
rect 19750 6616 19766 6650
rect 19800 6616 19816 6650
rect 19750 6600 19816 6616
rect 19753 6577 19813 6600
rect 20036 6577 20096 6603
rect 20154 6577 20214 6603
rect 20272 6577 20332 6603
rect 20659 6581 20719 6805
rect 21103 6763 21163 6964
rect 21221 6938 21281 6964
rect 21339 6938 21399 6964
rect 24141 6878 24199 7063
rect 24141 6852 24201 6878
rect 24259 6852 24319 7063
rect 24612 7057 24672 7089
rect 24730 7063 24790 7089
rect 24848 7063 24908 7089
rect 24609 7041 24675 7057
rect 24609 7007 24625 7041
rect 24659 7007 24675 7041
rect 24609 6991 24675 7007
rect 29780 7339 29840 7365
rect 29898 7339 29958 7365
rect 30016 7339 30076 7365
rect 30134 7345 30194 7365
rect 30134 7339 30195 7345
rect 30252 7339 30312 7365
rect 30370 7339 30430 7365
rect 30017 7154 30075 7339
rect 30017 7128 30077 7154
rect 30135 7128 30195 7339
rect 30488 7333 30548 7365
rect 30606 7339 30666 7365
rect 30724 7339 30784 7365
rect 30485 7317 30551 7333
rect 30485 7283 30501 7317
rect 30535 7283 30551 7317
rect 32008 7313 32304 7364
rect 32008 7298 32068 7313
rect 32126 7298 32186 7313
rect 32244 7298 32304 7313
rect 32362 7298 32422 7324
rect 32480 7298 32540 7324
rect 32598 7298 32658 7324
rect 30485 7267 30551 7283
rect 30367 7200 30433 7216
rect 30367 7166 30383 7200
rect 30417 7166 30433 7200
rect 30367 7150 30433 7166
rect 30370 7128 30430 7150
rect 26229 6944 26289 6961
rect 24491 6924 24557 6940
rect 24491 6890 24507 6924
rect 24541 6890 24557 6924
rect 24491 6874 24557 6890
rect 24494 6852 24554 6874
rect 26229 6855 26290 6944
rect 26347 6935 26407 6961
rect 26465 6935 26525 6961
rect 20777 6712 21163 6763
rect 20777 6581 20837 6712
rect 20892 6654 20958 6670
rect 20892 6620 20908 6654
rect 20942 6620 20958 6654
rect 20892 6604 20958 6620
rect 20895 6581 20955 6604
rect 21178 6581 21238 6607
rect 21296 6581 21356 6607
rect 21414 6581 21474 6607
rect 17519 6429 17579 6451
rect 17637 6429 17697 6451
rect 17516 6413 17582 6429
rect 12862 6350 12922 6376
rect 12980 6350 13040 6376
rect 7689 6309 8268 6350
rect 13098 6344 13158 6376
rect 13381 6344 13441 6376
rect 13499 6344 13559 6376
rect 13617 6344 13677 6376
rect 14004 6354 14064 6380
rect 14122 6354 14182 6380
rect 13098 6303 13677 6344
rect 14240 6348 14300 6380
rect 14523 6348 14583 6380
rect 14641 6348 14701 6380
rect 14759 6348 14819 6380
rect 17516 6379 17532 6413
rect 17566 6379 17582 6413
rect 17516 6363 17582 6379
rect 17634 6413 17700 6429
rect 17634 6379 17650 6413
rect 17684 6379 17700 6413
rect 17634 6363 17700 6379
rect 26139 6802 26290 6855
rect 24494 6626 24554 6652
rect 26139 6578 26199 6802
rect 26583 6760 26643 6961
rect 26701 6935 26761 6961
rect 26819 6935 26879 6961
rect 27371 6948 27431 6965
rect 27371 6859 27432 6948
rect 27489 6939 27549 6965
rect 27607 6939 27667 6965
rect 26257 6709 26643 6760
rect 27281 6806 27432 6859
rect 26257 6578 26317 6709
rect 26372 6651 26438 6667
rect 26372 6617 26388 6651
rect 26422 6617 26438 6651
rect 26372 6601 26438 6617
rect 26375 6578 26435 6601
rect 26658 6578 26718 6604
rect 26776 6578 26836 6604
rect 26894 6578 26954 6604
rect 27281 6582 27341 6806
rect 27725 6764 27785 6965
rect 27843 6939 27903 6965
rect 27961 6939 28021 6965
rect 27399 6713 27785 6764
rect 31524 7098 31584 7124
rect 31642 7098 31702 7124
rect 31760 7098 31820 7124
rect 30370 6902 30430 6928
rect 36701 7305 36755 7365
rect 37155 7305 37181 7365
rect 32845 7115 33141 7166
rect 32845 7098 32905 7115
rect 32963 7098 33023 7115
rect 33081 7098 33141 7115
rect 33317 7116 33613 7152
rect 33317 7095 33377 7116
rect 33435 7095 33495 7116
rect 33553 7095 33613 7116
rect 33671 7115 33967 7151
rect 33671 7095 33731 7115
rect 33789 7095 33849 7115
rect 33907 7095 33967 7115
rect 34025 7115 34321 7151
rect 34025 7095 34085 7115
rect 34143 7095 34203 7115
rect 34261 7095 34321 7115
rect 31524 6881 31584 6898
rect 31642 6881 31702 6898
rect 31760 6881 31820 6898
rect 32008 6881 32068 6898
rect 31524 6830 32068 6881
rect 32126 6872 32186 6898
rect 32244 6872 32304 6898
rect 32362 6879 32422 6898
rect 32480 6879 32540 6898
rect 32598 6879 32658 6898
rect 32845 6879 32905 6898
rect 32963 6879 33023 6898
rect 27399 6582 27459 6713
rect 30017 6706 30077 6728
rect 30135 6706 30195 6728
rect 30014 6690 30080 6706
rect 27514 6655 27580 6671
rect 27514 6621 27530 6655
rect 27564 6621 27580 6655
rect 30014 6656 30030 6690
rect 30064 6656 30080 6690
rect 30014 6640 30080 6656
rect 30132 6690 30198 6706
rect 30132 6656 30148 6690
rect 30182 6656 30198 6690
rect 30132 6640 30198 6656
rect 27514 6605 27580 6621
rect 31649 6626 31709 6830
rect 32362 6828 32905 6879
rect 32947 6872 33023 6879
rect 33081 6872 33141 6898
rect 36900 7068 36955 7128
rect 37155 7068 37181 7128
rect 36900 7010 36939 7068
rect 36900 6950 36955 7010
rect 37155 6950 37181 7010
rect 37301 6986 37367 7002
rect 37301 6952 37317 6986
rect 37351 6952 37367 6986
rect 32947 6828 33022 6872
rect 33317 6869 33377 6895
rect 33435 6869 33495 6895
rect 33553 6869 33613 6895
rect 33671 6875 33731 6895
rect 33671 6869 33732 6875
rect 33789 6869 33849 6895
rect 33907 6869 33967 6895
rect 32947 6746 33007 6828
rect 32947 6728 33181 6746
rect 32947 6694 33130 6728
rect 33164 6694 33181 6728
rect 31951 6628 32247 6688
rect 27517 6582 27577 6605
rect 27800 6582 27860 6608
rect 27918 6582 27978 6608
rect 28036 6582 28096 6608
rect 24141 6430 24201 6452
rect 24259 6430 24319 6452
rect 24138 6414 24204 6430
rect 19517 6351 19577 6377
rect 19635 6351 19695 6377
rect 14240 6307 14819 6348
rect 19753 6345 19813 6377
rect 20036 6345 20096 6377
rect 20154 6345 20214 6377
rect 20272 6345 20332 6377
rect 20659 6355 20719 6381
rect 20777 6355 20837 6381
rect 19753 6304 20332 6345
rect 20895 6349 20955 6381
rect 21178 6349 21238 6381
rect 21296 6349 21356 6381
rect 21414 6349 21474 6381
rect 24138 6380 24154 6414
rect 24188 6380 24204 6414
rect 24138 6364 24204 6380
rect 24256 6414 24322 6430
rect 24256 6380 24272 6414
rect 24306 6380 24322 6414
rect 24256 6364 24322 6380
rect 31649 6609 31780 6626
rect 31649 6575 31730 6609
rect 31764 6575 31780 6609
rect 31951 6605 32011 6628
rect 32069 6605 32129 6628
rect 32187 6605 32247 6628
rect 32305 6629 32601 6689
rect 32305 6605 32365 6629
rect 32423 6605 32483 6629
rect 32541 6605 32601 6629
rect 32947 6678 33181 6694
rect 33554 6684 33612 6869
rect 31649 6558 31780 6575
rect 26139 6352 26199 6378
rect 26257 6352 26317 6378
rect 20895 6308 21474 6349
rect 26375 6346 26435 6378
rect 26658 6346 26718 6378
rect 26776 6346 26836 6378
rect 26894 6346 26954 6378
rect 27281 6356 27341 6382
rect 27399 6356 27459 6382
rect 26375 6305 26954 6346
rect 27517 6350 27577 6382
rect 27800 6350 27860 6382
rect 27918 6350 27978 6382
rect 28036 6350 28096 6382
rect 27517 6309 28096 6350
rect -3061 5890 -3001 5906
rect -3634 5807 -3608 5867
rect -3408 5807 -3340 5867
rect -3391 5749 -3340 5807
rect -3634 5689 -3608 5749
rect -3408 5742 -3340 5749
rect -3061 5856 -3047 5890
rect -3013 5856 -3001 5890
rect -3061 5742 -3001 5856
rect 31649 5978 31709 6558
rect 31951 6179 32011 6205
rect 31919 6038 31986 6045
rect 32069 6038 32129 6205
rect 32187 6179 32247 6205
rect 32305 6179 32365 6205
rect 31919 6029 32129 6038
rect 31919 5995 31935 6029
rect 31969 5995 32129 6029
rect 31919 5979 32129 5995
rect 31649 5962 31800 5978
rect 31649 5928 31750 5962
rect 31784 5928 31800 5962
rect 31649 5912 31800 5928
rect 31649 5873 31709 5912
rect 32069 5873 32129 5979
rect 32423 6038 32483 6205
rect 32541 6179 32601 6205
rect 32566 6038 32633 6045
rect 32423 6029 32633 6038
rect 32423 5995 32583 6029
rect 32617 5995 32633 6029
rect 32423 5979 32633 5995
rect 32185 5945 32251 5961
rect 32185 5911 32201 5945
rect 32235 5911 32251 5945
rect 32185 5895 32251 5911
rect 32303 5946 32369 5961
rect 32303 5912 32319 5946
rect 32353 5912 32369 5946
rect 32303 5896 32369 5912
rect 32187 5873 32247 5895
rect 32305 5873 32365 5896
rect 32423 5873 32483 5979
rect 32947 5977 33007 6678
rect 33554 6658 33614 6684
rect 33672 6658 33732 6869
rect 34025 6863 34085 6895
rect 34143 6869 34203 6895
rect 34261 6869 34321 6895
rect 36900 6892 36939 6950
rect 37301 6936 37367 6952
rect 37304 6892 37364 6936
rect 37840 6892 37885 7700
rect 34022 6847 34088 6863
rect 34022 6813 34038 6847
rect 34072 6813 34088 6847
rect 36900 6832 36955 6892
rect 37155 6832 37885 6892
rect 34022 6797 34088 6813
rect 33904 6730 33970 6746
rect 33904 6696 33920 6730
rect 33954 6696 33970 6730
rect 33904 6680 33970 6696
rect 33907 6658 33967 6680
rect 33907 6432 33967 6458
rect 33554 6236 33614 6258
rect 33672 6236 33732 6258
rect 33551 6220 33617 6236
rect 33551 6186 33567 6220
rect 33601 6186 33617 6220
rect 33551 6170 33617 6186
rect 33669 6220 33735 6236
rect 33669 6186 33685 6220
rect 33719 6186 33735 6220
rect 33669 6170 33735 6186
rect 36896 6144 36951 6204
rect 37151 6145 37881 6204
rect 37151 6144 37454 6145
rect 36896 6086 36935 6144
rect 37437 6087 37454 6144
rect 37509 6144 37881 6145
rect 37509 6087 37524 6144
rect 32857 5961 33007 5977
rect 32857 5927 32873 5961
rect 32907 5927 33007 5961
rect 32857 5911 33007 5927
rect 32947 5873 33007 5911
rect 36896 6026 36951 6086
rect 37151 6026 37177 6086
rect 37437 6068 37524 6087
rect 36896 5968 36935 6026
rect 36896 5908 36951 5968
rect 37151 5908 37177 5968
rect -3408 5689 -2383 5742
rect -3391 5682 -2383 5689
rect -2183 5682 -2157 5742
rect -3391 5631 -3340 5682
rect -3634 5571 -3608 5631
rect -3408 5571 -3340 5631
rect -2488 5641 -2422 5682
rect -2488 5607 -2472 5641
rect -2438 5607 -2422 5641
rect 4090 5660 4386 5696
rect 4090 5639 4150 5660
rect 4208 5639 4268 5660
rect 4326 5639 4386 5660
rect 4444 5659 4740 5695
rect 4444 5639 4504 5659
rect 4562 5639 4622 5659
rect 4680 5639 4740 5659
rect 4798 5659 5094 5695
rect 4798 5639 4858 5659
rect 4916 5639 4976 5659
rect 5034 5639 5094 5659
rect -2488 5591 -2422 5607
rect -3391 5383 -3340 5571
rect -2555 5456 -2489 5472
rect -3874 5323 -3808 5383
rect -3408 5323 -3340 5383
rect -3198 5380 -3115 5440
rect -2715 5380 -2689 5440
rect -2555 5422 -2539 5456
rect -2505 5422 -2489 5456
rect 10641 5658 10937 5694
rect 10641 5637 10701 5658
rect 10759 5637 10819 5658
rect 10877 5637 10937 5658
rect 10995 5657 11291 5693
rect 10995 5637 11055 5657
rect 11113 5637 11173 5657
rect 11231 5637 11291 5657
rect 11349 5657 11645 5693
rect 11349 5637 11409 5657
rect 11467 5637 11527 5657
rect 11585 5637 11645 5657
rect -2555 5405 -2489 5422
rect 4090 5413 4150 5439
rect 4208 5413 4268 5439
rect 4326 5413 4386 5439
rect 4444 5419 4504 5439
rect 4444 5413 4505 5419
rect 4562 5413 4622 5439
rect 4680 5413 4740 5439
rect -3874 5265 -3823 5323
rect -3198 5322 -3138 5380
rect -2548 5322 -2489 5405
rect -3874 5205 -3808 5265
rect -3408 5205 -3382 5265
rect -3198 5262 -3115 5322
rect -2715 5262 -2383 5322
rect -1983 5262 -1957 5322
rect -3874 5147 -3823 5205
rect -3198 5204 -3138 5262
rect -2471 5204 -2405 5206
rect -3874 5087 -3808 5147
rect -3408 5087 -3382 5147
rect -3198 5144 -3115 5204
rect -2715 5144 -2689 5204
rect -2471 5190 -2383 5204
rect -2471 5156 -2455 5190
rect -2421 5156 -2383 5190
rect -2471 5144 -2383 5156
rect -1983 5144 -1957 5204
rect 4327 5228 4385 5413
rect 4327 5202 4387 5228
rect 4445 5202 4505 5413
rect 4798 5407 4858 5439
rect 4916 5413 4976 5439
rect 5034 5413 5094 5439
rect 17296 5659 17592 5695
rect 17296 5638 17356 5659
rect 17414 5638 17474 5659
rect 17532 5638 17592 5659
rect 17650 5658 17946 5694
rect 17650 5638 17710 5658
rect 17768 5638 17828 5658
rect 17886 5638 17946 5658
rect 18004 5658 18300 5694
rect 18004 5638 18064 5658
rect 18122 5638 18182 5658
rect 18240 5638 18300 5658
rect 23918 5660 24214 5696
rect 23918 5639 23978 5660
rect 24036 5639 24096 5660
rect 24154 5639 24214 5660
rect 24272 5659 24568 5695
rect 24272 5639 24332 5659
rect 24390 5639 24450 5659
rect 24508 5639 24568 5659
rect 24626 5659 24922 5695
rect 24626 5639 24686 5659
rect 24744 5639 24804 5659
rect 24862 5639 24922 5659
rect 31649 5647 31709 5673
rect 36697 5703 36751 5763
rect 37151 5703 37177 5763
rect 32947 5647 33007 5673
rect 36697 5645 36736 5703
rect 36697 5585 36751 5645
rect 37151 5585 37626 5645
rect 36697 5527 36736 5585
rect 32069 5447 32129 5473
rect 32187 5447 32247 5473
rect 32305 5447 32365 5473
rect 32423 5447 32483 5473
rect 36697 5467 36751 5527
rect 37151 5467 37177 5527
rect 10641 5411 10701 5437
rect 10759 5411 10819 5437
rect 10877 5411 10937 5437
rect 10995 5417 11055 5437
rect 10995 5411 11056 5417
rect 11113 5411 11173 5437
rect 11231 5411 11291 5437
rect 4795 5391 4861 5407
rect 4795 5357 4811 5391
rect 4845 5357 4861 5391
rect 4795 5341 4861 5357
rect 4677 5274 4743 5290
rect 4677 5240 4693 5274
rect 4727 5240 4743 5274
rect 4677 5224 4743 5240
rect 6038 5237 6334 5288
rect 4680 5202 4740 5224
rect 6038 5222 6098 5237
rect 6156 5222 6216 5237
rect 6274 5222 6334 5237
rect 6392 5222 6452 5248
rect 6510 5222 6570 5248
rect 6628 5222 6688 5248
rect 7936 5237 8232 5288
rect 7936 5222 7996 5237
rect 8054 5222 8114 5237
rect 8172 5222 8232 5237
rect 8290 5222 8350 5248
rect 8408 5222 8468 5248
rect 8526 5222 8586 5248
rect 10878 5226 10936 5411
rect -2471 5140 -2405 5144
rect -2471 5086 -2406 5088
rect -3834 4969 -3808 5029
rect -3408 4969 -3338 5029
rect -3389 4911 -3338 4969
rect -3834 4851 -3808 4911
rect -3408 4851 -3338 4911
rect -3389 4793 -3338 4851
rect -3834 4733 -3808 4793
rect -3408 4733 -3338 4793
rect -3199 5026 -3115 5086
rect -2715 5026 -2689 5086
rect -2471 5072 -2383 5086
rect -2471 5038 -2456 5072
rect -2422 5038 -2383 5072
rect -2471 5026 -2383 5038
rect -1983 5026 -1957 5086
rect -3199 4968 -3139 5026
rect -2471 5022 -2406 5026
rect -3199 4908 -3115 4968
rect -2715 4908 -2383 4968
rect -1983 4908 -1957 4968
rect -3199 4850 -3139 4908
rect -3199 4790 -3115 4850
rect -2715 4790 -2689 4850
rect -2548 4825 -2489 4908
rect -2555 4808 -2489 4825
rect -3389 4546 -3338 4733
rect -2555 4774 -2539 4808
rect -2505 4774 -2489 4808
rect 5554 5022 5614 5048
rect 5672 5022 5732 5048
rect 5790 5022 5850 5048
rect 4680 4976 4740 5002
rect 4327 4780 4387 4802
rect 4445 4786 4505 4802
rect -2555 4758 -2489 4774
rect 1183 4734 1479 4770
rect 1183 4713 1243 4734
rect 1301 4713 1361 4734
rect 1419 4713 1479 4734
rect 1537 4733 1833 4769
rect 1537 4713 1597 4733
rect 1655 4713 1715 4733
rect 1773 4713 1833 4733
rect 1891 4733 2187 4769
rect 1891 4713 1951 4733
rect 2009 4713 2069 4733
rect 2127 4713 2187 4733
rect 4324 4764 4390 4780
rect 4324 4730 4340 4764
rect 4374 4730 4390 4764
rect 4324 4714 4390 4730
rect 4439 4764 4513 4786
rect 4439 4730 4458 4764
rect 4492 4730 4513 4764
rect 6875 5039 7171 5090
rect 6875 5022 6935 5039
rect 6993 5022 7053 5039
rect 7111 5022 7171 5039
rect 7452 5022 7512 5048
rect 7570 5022 7630 5048
rect 7688 5022 7748 5048
rect 10878 5200 10938 5226
rect 10996 5200 11056 5411
rect 11349 5405 11409 5437
rect 11467 5411 11527 5437
rect 11585 5411 11645 5437
rect 17296 5412 17356 5438
rect 17414 5412 17474 5438
rect 17532 5412 17592 5438
rect 17650 5418 17710 5438
rect 17650 5412 17711 5418
rect 17768 5412 17828 5438
rect 17886 5412 17946 5438
rect 11346 5389 11412 5405
rect 11346 5355 11362 5389
rect 11396 5355 11412 5389
rect 11346 5339 11412 5355
rect 11228 5272 11294 5288
rect 11228 5238 11244 5272
rect 11278 5238 11294 5272
rect 11228 5222 11294 5238
rect 12589 5235 12885 5286
rect 11231 5200 11291 5222
rect 12589 5220 12649 5235
rect 12707 5220 12767 5235
rect 12825 5220 12885 5235
rect 12943 5220 13003 5246
rect 13061 5220 13121 5246
rect 13179 5220 13239 5246
rect 14487 5235 14783 5286
rect 14487 5220 14547 5235
rect 14605 5220 14665 5235
rect 14723 5220 14783 5235
rect 14841 5220 14901 5246
rect 14959 5220 15019 5246
rect 15077 5220 15137 5246
rect 17533 5227 17591 5412
rect 8773 5039 9069 5090
rect 8773 5022 8833 5039
rect 8891 5022 8951 5039
rect 9009 5022 9069 5039
rect 5554 4805 5614 4822
rect 5672 4805 5732 4822
rect 5790 4805 5850 4822
rect 6038 4805 6098 4822
rect 5554 4754 6098 4805
rect 6156 4796 6216 4822
rect 6274 4796 6334 4822
rect 6392 4803 6452 4822
rect 6510 4803 6570 4822
rect 6628 4803 6688 4822
rect 6875 4803 6935 4822
rect 6993 4803 7053 4822
rect -3676 4486 -3608 4546
rect -3408 4486 -3338 4546
rect -2487 4518 -2421 4534
rect -3251 4496 -3197 4512
rect -3676 4428 -3625 4486
rect -3251 4462 -3241 4496
rect -3207 4462 -3197 4496
rect -3251 4444 -3197 4462
rect -2487 4484 -2471 4518
rect -2437 4484 -2421 4518
rect 4439 4673 4513 4730
rect 5679 4673 5739 4754
rect 6392 4752 6935 4803
rect 6977 4796 7053 4803
rect 7111 4796 7171 4822
rect 7452 4805 7512 4822
rect 7570 4805 7630 4822
rect 7688 4805 7748 4822
rect 7936 4805 7996 4822
rect 6977 4752 7052 4796
rect 7452 4754 7996 4805
rect 8054 4796 8114 4822
rect 8172 4796 8232 4822
rect 8290 4803 8350 4822
rect 8408 4803 8468 4822
rect 8526 4803 8586 4822
rect 8773 4803 8833 4822
rect 8891 4803 8951 4822
rect 4439 4648 5739 4673
rect 4438 4600 5739 4648
rect 6977 4632 7037 4752
rect -2487 4444 -2421 4484
rect 1183 4487 1243 4513
rect 1301 4487 1361 4513
rect 1419 4487 1479 4513
rect 1537 4493 1597 4513
rect 1537 4487 1598 4493
rect 1655 4487 1715 4513
rect 1773 4487 1833 4513
rect -3389 4428 -2383 4444
rect -3676 4368 -3608 4428
rect -3408 4384 -2383 4428
rect -2183 4384 -2157 4444
rect -3408 4369 -3338 4384
rect -3408 4368 -3382 4369
rect -3676 4310 -3625 4368
rect -3676 4250 -3608 4310
rect -3408 4250 -3382 4310
rect 1420 4302 1478 4487
rect 1420 4276 1480 4302
rect 1538 4276 1598 4487
rect 1891 4481 1951 4513
rect 2009 4487 2069 4513
rect 2127 4487 2187 4513
rect 1888 4465 1954 4481
rect 1888 4431 1904 4465
rect 1938 4431 1954 4465
rect 1888 4415 1954 4431
rect 1770 4348 1836 4364
rect 1770 4314 1786 4348
rect 1820 4314 1836 4348
rect 1770 4298 1836 4314
rect 1773 4276 1833 4298
rect 1773 4050 1833 4076
rect 4085 4056 4381 4092
rect 4085 4035 4145 4056
rect 4203 4035 4263 4056
rect 4321 4035 4381 4056
rect 4439 4055 4735 4091
rect 4439 4035 4499 4055
rect 4557 4035 4617 4055
rect 4675 4035 4735 4055
rect 4793 4055 5089 4091
rect 4793 4035 4853 4055
rect 4911 4035 4971 4055
rect 5029 4035 5089 4055
rect 1420 3854 1480 3876
rect 1538 3854 1598 3876
rect 1417 3838 1483 3854
rect -3059 3821 -2999 3837
rect -3632 3738 -3606 3798
rect -3406 3738 -3338 3798
rect -3389 3680 -3338 3738
rect -3632 3620 -3606 3680
rect -3406 3673 -3338 3680
rect -3059 3787 -3045 3821
rect -3011 3787 -2999 3821
rect 1417 3804 1433 3838
rect 1467 3804 1483 3838
rect 1417 3788 1483 3804
rect 1535 3838 1601 3854
rect 1535 3804 1551 3838
rect 1585 3804 1601 3838
rect 5679 3902 5739 4600
rect 5981 4552 6277 4612
rect 5981 4529 6041 4552
rect 6099 4529 6159 4552
rect 6217 4529 6277 4552
rect 6335 4553 6631 4613
rect 6976 4612 7037 4632
rect 6335 4529 6395 4553
rect 6453 4529 6513 4553
rect 6571 4529 6631 4553
rect 6957 4596 7037 4612
rect 6957 4562 6972 4596
rect 7006 4562 7037 4596
rect 6957 4546 7037 4562
rect 6976 4523 7037 4546
rect 6977 4377 7037 4523
rect 6976 4204 7037 4377
rect 5981 4103 6041 4129
rect 5949 3962 6016 3969
rect 6099 3962 6159 4129
rect 6217 4103 6277 4129
rect 6335 4103 6395 4129
rect 5949 3953 6159 3962
rect 5949 3919 5965 3953
rect 5999 3919 6159 3953
rect 5949 3903 6159 3919
rect 5679 3886 5830 3902
rect 5679 3852 5780 3886
rect 5814 3852 5830 3886
rect 5679 3836 5830 3852
rect 4085 3809 4145 3835
rect 4203 3809 4263 3835
rect 4321 3809 4381 3835
rect 4439 3815 4499 3835
rect 4439 3809 4500 3815
rect 4557 3809 4617 3835
rect 4675 3809 4735 3835
rect 1535 3788 1601 3804
rect -3059 3673 -2999 3787
rect -3406 3620 -2381 3673
rect -3389 3613 -2381 3620
rect -2181 3613 -2155 3673
rect 4322 3624 4380 3809
rect -3389 3562 -3338 3613
rect -3632 3502 -3606 3562
rect -3406 3502 -3338 3562
rect -2486 3572 -2420 3613
rect -2486 3538 -2470 3572
rect -2436 3538 -2420 3572
rect 4322 3598 4382 3624
rect 4440 3598 4500 3809
rect 4793 3803 4853 3835
rect 4911 3809 4971 3835
rect 5029 3809 5089 3835
rect 4790 3787 4856 3803
rect 5679 3797 5739 3836
rect 6099 3797 6159 3903
rect 6453 3962 6513 4129
rect 6571 4103 6631 4129
rect 6596 3962 6663 3969
rect 6453 3953 6663 3962
rect 6453 3919 6613 3953
rect 6647 3919 6663 3953
rect 6453 3903 6663 3919
rect 6215 3869 6281 3885
rect 6215 3835 6231 3869
rect 6265 3835 6281 3869
rect 6215 3819 6281 3835
rect 6333 3870 6399 3885
rect 6333 3836 6349 3870
rect 6383 3836 6399 3870
rect 6333 3820 6399 3836
rect 6217 3797 6277 3819
rect 6335 3797 6395 3820
rect 6453 3797 6513 3903
rect 6977 3901 7037 4204
rect 6887 3885 7037 3901
rect 6887 3851 6903 3885
rect 6937 3851 7037 3885
rect 6887 3835 7037 3851
rect 6977 3797 7037 3835
rect 7577 4096 7637 4754
rect 8290 4752 8833 4803
rect 8875 4796 8951 4803
rect 9009 4796 9069 4822
rect 12105 5020 12165 5046
rect 12223 5020 12283 5046
rect 12341 5020 12401 5046
rect 11231 4974 11291 5000
rect 8875 4752 8950 4796
rect 10878 4778 10938 4800
rect 10996 4784 11056 4800
rect 10875 4762 10941 4778
rect 7879 4552 8175 4612
rect 7879 4529 7939 4552
rect 7997 4529 8057 4552
rect 8115 4529 8175 4552
rect 8233 4553 8529 4613
rect 8233 4529 8293 4553
rect 8351 4529 8411 4553
rect 8469 4529 8529 4553
rect 8875 4599 8935 4752
rect 10875 4728 10891 4762
rect 10925 4728 10941 4762
rect 10875 4712 10941 4728
rect 10990 4762 11064 4784
rect 10990 4728 11009 4762
rect 11043 4728 11064 4762
rect 13426 5037 13722 5088
rect 13426 5020 13486 5037
rect 13544 5020 13604 5037
rect 13662 5020 13722 5037
rect 14003 5020 14063 5046
rect 14121 5020 14181 5046
rect 14239 5020 14299 5046
rect 17533 5201 17593 5227
rect 17651 5201 17711 5412
rect 18004 5406 18064 5438
rect 18122 5412 18182 5438
rect 18240 5412 18300 5438
rect 23918 5413 23978 5439
rect 24036 5413 24096 5439
rect 24154 5413 24214 5439
rect 24272 5419 24332 5439
rect 24272 5413 24333 5419
rect 24390 5413 24450 5439
rect 24508 5413 24568 5439
rect 18001 5390 18067 5406
rect 18001 5356 18017 5390
rect 18051 5356 18067 5390
rect 18001 5340 18067 5356
rect 17883 5273 17949 5289
rect 17883 5239 17899 5273
rect 17933 5239 17949 5273
rect 17883 5223 17949 5239
rect 19244 5236 19540 5287
rect 17886 5201 17946 5223
rect 19244 5221 19304 5236
rect 19362 5221 19422 5236
rect 19480 5221 19540 5236
rect 19598 5221 19658 5247
rect 19716 5221 19776 5247
rect 19834 5221 19894 5247
rect 21142 5236 21438 5287
rect 21142 5221 21202 5236
rect 21260 5221 21320 5236
rect 21378 5221 21438 5236
rect 21496 5221 21556 5247
rect 21614 5221 21674 5247
rect 21732 5221 21792 5247
rect 24155 5228 24213 5413
rect 15324 5037 15620 5088
rect 15324 5020 15384 5037
rect 15442 5020 15502 5037
rect 15560 5020 15620 5037
rect 12105 4803 12165 4820
rect 12223 4803 12283 4820
rect 12341 4803 12401 4820
rect 12589 4803 12649 4820
rect 12105 4752 12649 4803
rect 12707 4794 12767 4820
rect 12825 4794 12885 4820
rect 12943 4801 13003 4820
rect 13061 4801 13121 4820
rect 13179 4801 13239 4820
rect 13426 4801 13486 4820
rect 13544 4801 13604 4820
rect 10990 4671 11064 4728
rect 12230 4671 12290 4752
rect 12943 4750 13486 4801
rect 13528 4794 13604 4801
rect 13662 4794 13722 4820
rect 14003 4803 14063 4820
rect 14121 4803 14181 4820
rect 14239 4803 14299 4820
rect 14487 4803 14547 4820
rect 13528 4750 13603 4794
rect 14003 4752 14547 4803
rect 14605 4794 14665 4820
rect 14723 4794 14783 4820
rect 14841 4801 14901 4820
rect 14959 4801 15019 4820
rect 15077 4801 15137 4820
rect 15324 4801 15384 4820
rect 15442 4801 15502 4820
rect 10990 4646 12290 4671
rect 8875 4575 9129 4599
rect 10989 4598 12290 4646
rect 13528 4630 13588 4750
rect 8875 4541 9079 4575
rect 9113 4541 9129 4575
rect 8875 4525 9129 4541
rect 7879 4103 7939 4129
rect 7577 4080 7644 4096
rect 7577 4046 7593 4080
rect 7627 4046 7644 4080
rect 7577 4030 7644 4046
rect 7577 3902 7637 4030
rect 7847 3962 7914 3969
rect 7997 3962 8057 4129
rect 8115 4103 8175 4129
rect 8233 4103 8293 4129
rect 7847 3953 8057 3962
rect 7847 3919 7863 3953
rect 7897 3919 8057 3953
rect 7847 3903 8057 3919
rect 7577 3886 7728 3902
rect 7577 3852 7678 3886
rect 7712 3852 7728 3886
rect 7577 3836 7728 3852
rect 7577 3797 7637 3836
rect 7997 3797 8057 3903
rect 8351 3962 8411 4129
rect 8469 4103 8529 4129
rect 8492 3963 8559 3970
rect 8486 3962 8559 3963
rect 8351 3954 8559 3962
rect 8351 3920 8509 3954
rect 8543 3920 8559 3954
rect 8351 3904 8559 3920
rect 8351 3903 8548 3904
rect 8113 3869 8179 3885
rect 8113 3835 8129 3869
rect 8163 3835 8179 3869
rect 8113 3819 8179 3835
rect 8231 3870 8297 3885
rect 8231 3836 8247 3870
rect 8281 3836 8297 3870
rect 8231 3820 8297 3836
rect 8115 3797 8175 3819
rect 8233 3797 8293 3820
rect 8351 3797 8411 3903
rect 8875 3901 8935 4525
rect 10636 4054 10932 4090
rect 10636 4033 10696 4054
rect 10754 4033 10814 4054
rect 10872 4033 10932 4054
rect 10990 4053 11286 4089
rect 10990 4033 11050 4053
rect 11108 4033 11168 4053
rect 11226 4033 11286 4053
rect 11344 4053 11640 4089
rect 11344 4033 11404 4053
rect 11462 4033 11522 4053
rect 11580 4033 11640 4053
rect 8785 3885 8935 3901
rect 8785 3851 8801 3885
rect 8835 3851 8935 3885
rect 8785 3835 8935 3851
rect 8875 3797 8935 3835
rect 12230 3900 12290 4598
rect 12532 4550 12828 4610
rect 12532 4527 12592 4550
rect 12650 4527 12710 4550
rect 12768 4527 12828 4550
rect 12886 4551 13182 4611
rect 13527 4610 13588 4630
rect 12886 4527 12946 4551
rect 13004 4527 13064 4551
rect 13122 4527 13182 4551
rect 13508 4594 13588 4610
rect 13508 4560 13523 4594
rect 13557 4560 13588 4594
rect 13508 4544 13588 4560
rect 13527 4521 13588 4544
rect 13528 4375 13588 4521
rect 13527 4202 13588 4375
rect 12532 4101 12592 4127
rect 12500 3960 12567 3967
rect 12650 3960 12710 4127
rect 12768 4101 12828 4127
rect 12886 4101 12946 4127
rect 12500 3951 12710 3960
rect 12500 3917 12516 3951
rect 12550 3917 12710 3951
rect 12500 3901 12710 3917
rect 12230 3884 12381 3900
rect 12230 3850 12331 3884
rect 12365 3850 12381 3884
rect 12230 3834 12381 3850
rect 10636 3807 10696 3833
rect 10754 3807 10814 3833
rect 10872 3807 10932 3833
rect 10990 3813 11050 3833
rect 10990 3807 11051 3813
rect 11108 3807 11168 3833
rect 11226 3807 11286 3833
rect 4790 3753 4806 3787
rect 4840 3753 4856 3787
rect 4790 3737 4856 3753
rect 4672 3670 4738 3686
rect 4672 3636 4688 3670
rect 4722 3636 4738 3670
rect 4672 3620 4738 3636
rect 4675 3598 4735 3620
rect -2486 3522 -2420 3538
rect -3389 3314 -3338 3502
rect -2553 3387 -2487 3403
rect -3872 3254 -3806 3314
rect -3406 3254 -3338 3314
rect -3196 3311 -3113 3371
rect -2713 3311 -2687 3371
rect -2553 3353 -2537 3387
rect -2503 3353 -2487 3387
rect -2553 3336 -2487 3353
rect -3872 3196 -3821 3254
rect -3196 3253 -3136 3311
rect -2546 3253 -2487 3336
rect -3872 3136 -3806 3196
rect -3406 3136 -3380 3196
rect -3196 3193 -3113 3253
rect -2713 3193 -2381 3253
rect -1981 3193 -1955 3253
rect 5679 3571 5739 3597
rect 4675 3372 4735 3398
rect 6977 3571 7037 3597
rect 7577 3571 7637 3597
rect 10873 3622 10931 3807
rect 8875 3571 8935 3597
rect 10873 3596 10933 3622
rect 10991 3596 11051 3807
rect 11344 3801 11404 3833
rect 11462 3807 11522 3833
rect 11580 3807 11640 3833
rect 11341 3785 11407 3801
rect 12230 3795 12290 3834
rect 12650 3795 12710 3901
rect 13004 3960 13064 4127
rect 13122 4101 13182 4127
rect 13147 3960 13214 3967
rect 13004 3951 13214 3960
rect 13004 3917 13164 3951
rect 13198 3917 13214 3951
rect 13004 3901 13214 3917
rect 12766 3867 12832 3883
rect 12766 3833 12782 3867
rect 12816 3833 12832 3867
rect 12766 3817 12832 3833
rect 12884 3868 12950 3883
rect 12884 3834 12900 3868
rect 12934 3834 12950 3868
rect 12884 3818 12950 3834
rect 12768 3795 12828 3817
rect 12886 3795 12946 3818
rect 13004 3795 13064 3901
rect 13528 3899 13588 4202
rect 13438 3883 13588 3899
rect 13438 3849 13454 3883
rect 13488 3849 13588 3883
rect 13438 3833 13588 3849
rect 13528 3795 13588 3833
rect 14128 4094 14188 4752
rect 14841 4750 15384 4801
rect 15426 4794 15502 4801
rect 15560 4794 15620 4820
rect 18760 5021 18820 5047
rect 18878 5021 18938 5047
rect 18996 5021 19056 5047
rect 17886 4975 17946 5001
rect 15426 4750 15501 4794
rect 17533 4779 17593 4801
rect 17651 4785 17711 4801
rect 17530 4763 17596 4779
rect 14430 4550 14726 4610
rect 14430 4527 14490 4550
rect 14548 4527 14608 4550
rect 14666 4527 14726 4550
rect 14784 4551 15080 4611
rect 14784 4527 14844 4551
rect 14902 4527 14962 4551
rect 15020 4527 15080 4551
rect 15426 4597 15486 4750
rect 17530 4729 17546 4763
rect 17580 4729 17596 4763
rect 17530 4713 17596 4729
rect 17645 4763 17719 4785
rect 17645 4729 17664 4763
rect 17698 4729 17719 4763
rect 20081 5038 20377 5089
rect 20081 5021 20141 5038
rect 20199 5021 20259 5038
rect 20317 5021 20377 5038
rect 20658 5021 20718 5047
rect 20776 5021 20836 5047
rect 20894 5021 20954 5047
rect 24155 5202 24215 5228
rect 24273 5202 24333 5413
rect 24626 5407 24686 5439
rect 24744 5413 24804 5439
rect 24862 5413 24922 5439
rect 24623 5391 24689 5407
rect 24623 5357 24639 5391
rect 24673 5357 24689 5391
rect 24623 5341 24689 5357
rect 24505 5274 24571 5290
rect 24505 5240 24521 5274
rect 24555 5240 24571 5274
rect 24505 5224 24571 5240
rect 25866 5237 26162 5288
rect 24508 5202 24568 5224
rect 25866 5222 25926 5237
rect 25984 5222 26044 5237
rect 26102 5222 26162 5237
rect 26220 5222 26280 5248
rect 26338 5222 26398 5248
rect 26456 5222 26516 5248
rect 27764 5237 28060 5288
rect 27764 5222 27824 5237
rect 27882 5222 27942 5237
rect 28000 5222 28060 5237
rect 28118 5222 28178 5248
rect 28236 5222 28296 5248
rect 28354 5222 28414 5248
rect 21979 5038 22275 5089
rect 21979 5021 22039 5038
rect 22097 5021 22157 5038
rect 22215 5021 22275 5038
rect 18760 4804 18820 4821
rect 18878 4804 18938 4821
rect 18996 4804 19056 4821
rect 19244 4804 19304 4821
rect 18760 4753 19304 4804
rect 19362 4795 19422 4821
rect 19480 4795 19540 4821
rect 19598 4802 19658 4821
rect 19716 4802 19776 4821
rect 19834 4802 19894 4821
rect 20081 4802 20141 4821
rect 20199 4802 20259 4821
rect 17645 4672 17719 4729
rect 18885 4672 18945 4753
rect 19598 4751 20141 4802
rect 20183 4795 20259 4802
rect 20317 4795 20377 4821
rect 20658 4804 20718 4821
rect 20776 4804 20836 4821
rect 20894 4804 20954 4821
rect 21142 4804 21202 4821
rect 20183 4751 20258 4795
rect 20658 4753 21202 4804
rect 21260 4795 21320 4821
rect 21378 4795 21438 4821
rect 21496 4802 21556 4821
rect 21614 4802 21674 4821
rect 21732 4802 21792 4821
rect 21979 4802 22039 4821
rect 22097 4802 22157 4821
rect 17645 4647 18945 4672
rect 17644 4599 18945 4647
rect 20183 4631 20243 4751
rect 15426 4573 15680 4597
rect 15426 4539 15630 4573
rect 15664 4539 15680 4573
rect 15426 4523 15680 4539
rect 14430 4101 14490 4127
rect 14128 4078 14195 4094
rect 14128 4044 14144 4078
rect 14178 4044 14195 4078
rect 14128 4028 14195 4044
rect 14128 3900 14188 4028
rect 14398 3960 14465 3967
rect 14548 3960 14608 4127
rect 14666 4101 14726 4127
rect 14784 4101 14844 4127
rect 14398 3951 14608 3960
rect 14398 3917 14414 3951
rect 14448 3917 14608 3951
rect 14398 3901 14608 3917
rect 14128 3884 14279 3900
rect 14128 3850 14229 3884
rect 14263 3850 14279 3884
rect 14128 3834 14279 3850
rect 14128 3795 14188 3834
rect 14548 3795 14608 3901
rect 14902 3960 14962 4127
rect 15020 4101 15080 4127
rect 15043 3961 15110 3968
rect 15037 3960 15110 3961
rect 14902 3952 15110 3960
rect 14902 3918 15060 3952
rect 15094 3918 15110 3952
rect 14902 3902 15110 3918
rect 14902 3901 15099 3902
rect 14664 3867 14730 3883
rect 14664 3833 14680 3867
rect 14714 3833 14730 3867
rect 14664 3817 14730 3833
rect 14782 3868 14848 3883
rect 14782 3834 14798 3868
rect 14832 3834 14848 3868
rect 14782 3818 14848 3834
rect 14666 3795 14726 3817
rect 14784 3795 14844 3818
rect 14902 3795 14962 3901
rect 15426 3899 15486 4523
rect 17291 4055 17587 4091
rect 17291 4034 17351 4055
rect 17409 4034 17469 4055
rect 17527 4034 17587 4055
rect 17645 4054 17941 4090
rect 17645 4034 17705 4054
rect 17763 4034 17823 4054
rect 17881 4034 17941 4054
rect 17999 4054 18295 4090
rect 17999 4034 18059 4054
rect 18117 4034 18177 4054
rect 18235 4034 18295 4054
rect 15336 3883 15486 3899
rect 15336 3849 15352 3883
rect 15386 3849 15486 3883
rect 15336 3833 15486 3849
rect 18885 3901 18945 4599
rect 19187 4551 19483 4611
rect 19187 4528 19247 4551
rect 19305 4528 19365 4551
rect 19423 4528 19483 4551
rect 19541 4552 19837 4612
rect 20182 4611 20243 4631
rect 19541 4528 19601 4552
rect 19659 4528 19719 4552
rect 19777 4528 19837 4552
rect 20163 4595 20243 4611
rect 20163 4561 20178 4595
rect 20212 4561 20243 4595
rect 20163 4545 20243 4561
rect 20182 4522 20243 4545
rect 20183 4376 20243 4522
rect 20182 4203 20243 4376
rect 19187 4102 19247 4128
rect 19155 3961 19222 3968
rect 19305 3961 19365 4128
rect 19423 4102 19483 4128
rect 19541 4102 19601 4128
rect 19155 3952 19365 3961
rect 19155 3918 19171 3952
rect 19205 3918 19365 3952
rect 19155 3902 19365 3918
rect 18885 3885 19036 3901
rect 18885 3851 18986 3885
rect 19020 3851 19036 3885
rect 18885 3835 19036 3851
rect 15426 3795 15486 3833
rect 17291 3808 17351 3834
rect 17409 3808 17469 3834
rect 17527 3808 17587 3834
rect 17645 3814 17705 3834
rect 17645 3808 17706 3814
rect 17763 3808 17823 3834
rect 17881 3808 17941 3834
rect 11341 3751 11357 3785
rect 11391 3751 11407 3785
rect 11341 3735 11407 3751
rect 11223 3668 11289 3684
rect 11223 3634 11239 3668
rect 11273 3634 11289 3668
rect 11223 3618 11289 3634
rect 11226 3596 11286 3618
rect 6099 3371 6159 3397
rect 6217 3371 6277 3397
rect 6335 3371 6395 3397
rect 6453 3371 6513 3397
rect 7997 3371 8057 3397
rect 8115 3371 8175 3397
rect 8233 3371 8293 3397
rect 8351 3371 8411 3397
rect -3872 3078 -3821 3136
rect -3196 3135 -3136 3193
rect 4322 3176 4382 3198
rect 4440 3176 4500 3198
rect -2469 3135 -2403 3137
rect -3872 3018 -3806 3078
rect -3406 3018 -3380 3078
rect -3196 3075 -3113 3135
rect -2713 3075 -2687 3135
rect -2469 3121 -2381 3135
rect -2469 3087 -2453 3121
rect -2419 3087 -2381 3121
rect -2469 3075 -2381 3087
rect -1981 3075 -1955 3135
rect 4319 3160 4385 3176
rect 4319 3126 4335 3160
rect 4369 3126 4385 3160
rect 4319 3110 4385 3126
rect 4437 3160 4503 3176
rect 4437 3126 4453 3160
rect 4487 3126 4503 3160
rect 12230 3569 12290 3595
rect 11226 3370 11286 3396
rect 13528 3569 13588 3595
rect 14128 3569 14188 3595
rect 17528 3623 17586 3808
rect 17528 3597 17588 3623
rect 17646 3597 17706 3808
rect 17999 3802 18059 3834
rect 18117 3808 18177 3834
rect 18235 3808 18295 3834
rect 17996 3786 18062 3802
rect 18885 3796 18945 3835
rect 19305 3796 19365 3902
rect 19659 3961 19719 4128
rect 19777 4102 19837 4128
rect 19802 3961 19869 3968
rect 19659 3952 19869 3961
rect 19659 3918 19819 3952
rect 19853 3918 19869 3952
rect 19659 3902 19869 3918
rect 19421 3868 19487 3884
rect 19421 3834 19437 3868
rect 19471 3834 19487 3868
rect 19421 3818 19487 3834
rect 19539 3869 19605 3884
rect 19539 3835 19555 3869
rect 19589 3835 19605 3869
rect 19539 3819 19605 3835
rect 19423 3796 19483 3818
rect 19541 3796 19601 3819
rect 19659 3796 19719 3902
rect 20183 3900 20243 4203
rect 20093 3884 20243 3900
rect 20093 3850 20109 3884
rect 20143 3850 20243 3884
rect 20093 3834 20243 3850
rect 20183 3796 20243 3834
rect 20783 4095 20843 4753
rect 21496 4751 22039 4802
rect 22081 4795 22157 4802
rect 22215 4795 22275 4821
rect 25382 5022 25442 5048
rect 25500 5022 25560 5048
rect 25618 5022 25678 5048
rect 24508 4976 24568 5002
rect 22081 4751 22156 4795
rect 24155 4780 24215 4802
rect 24273 4786 24333 4802
rect 24152 4764 24218 4780
rect 21085 4551 21381 4611
rect 21085 4528 21145 4551
rect 21203 4528 21263 4551
rect 21321 4528 21381 4551
rect 21439 4552 21735 4612
rect 21439 4528 21499 4552
rect 21557 4528 21617 4552
rect 21675 4528 21735 4552
rect 22081 4598 22141 4751
rect 24152 4730 24168 4764
rect 24202 4730 24218 4764
rect 24152 4714 24218 4730
rect 24267 4764 24341 4786
rect 24267 4730 24286 4764
rect 24320 4730 24341 4764
rect 26703 5039 26999 5090
rect 26703 5022 26763 5039
rect 26821 5022 26881 5039
rect 26939 5022 26999 5039
rect 27280 5022 27340 5048
rect 27398 5022 27458 5048
rect 27516 5022 27576 5048
rect 36697 5236 36751 5296
rect 37151 5236 37177 5296
rect 36697 5178 36736 5236
rect 36697 5118 36751 5178
rect 37151 5177 37177 5178
rect 37338 5177 37404 5180
rect 37151 5164 37404 5177
rect 37151 5130 37354 5164
rect 37388 5130 37404 5164
rect 37151 5118 37404 5130
rect 37569 5178 37626 5585
rect 37836 5370 37881 6144
rect 37836 5310 38084 5370
rect 38284 5310 38310 5370
rect 37725 5178 37804 5189
rect 37569 5176 38084 5178
rect 37569 5118 37738 5176
rect 37793 5118 38084 5176
rect 38484 5118 38510 5178
rect 28601 5039 28897 5090
rect 28601 5022 28661 5039
rect 28719 5022 28779 5039
rect 28837 5022 28897 5039
rect 36697 5060 36736 5118
rect 37337 5114 37404 5118
rect 37725 5108 37804 5118
rect 37438 5060 37525 5077
rect 36697 5000 36751 5060
rect 37151 5000 37177 5060
rect 37438 5058 38084 5060
rect 37438 5000 37453 5058
rect 37508 5000 38084 5058
rect 38484 5000 38510 5060
rect 37438 4982 37525 5000
rect 25382 4805 25442 4822
rect 25500 4805 25560 4822
rect 25618 4805 25678 4822
rect 25866 4805 25926 4822
rect 25382 4754 25926 4805
rect 25984 4796 26044 4822
rect 26102 4796 26162 4822
rect 26220 4803 26280 4822
rect 26338 4803 26398 4822
rect 26456 4803 26516 4822
rect 26703 4803 26763 4822
rect 26821 4803 26881 4822
rect 24267 4673 24341 4730
rect 25507 4673 25567 4754
rect 26220 4752 26763 4803
rect 26805 4796 26881 4803
rect 26939 4796 26999 4822
rect 27280 4805 27340 4822
rect 27398 4805 27458 4822
rect 27516 4805 27576 4822
rect 27764 4805 27824 4822
rect 26805 4752 26880 4796
rect 27280 4754 27824 4805
rect 27882 4796 27942 4822
rect 28000 4796 28060 4822
rect 28118 4803 28178 4822
rect 28236 4803 28296 4822
rect 28354 4803 28414 4822
rect 28601 4803 28661 4822
rect 28719 4803 28779 4822
rect 24267 4648 25567 4673
rect 24266 4600 25567 4648
rect 26805 4632 26865 4752
rect 22081 4574 22335 4598
rect 22081 4540 22285 4574
rect 22319 4540 22335 4574
rect 22081 4524 22335 4540
rect 21085 4102 21145 4128
rect 20783 4079 20850 4095
rect 20783 4045 20799 4079
rect 20833 4045 20850 4079
rect 20783 4029 20850 4045
rect 20783 3901 20843 4029
rect 21053 3961 21120 3968
rect 21203 3961 21263 4128
rect 21321 4102 21381 4128
rect 21439 4102 21499 4128
rect 21053 3952 21263 3961
rect 21053 3918 21069 3952
rect 21103 3918 21263 3952
rect 21053 3902 21263 3918
rect 20783 3885 20934 3901
rect 20783 3851 20884 3885
rect 20918 3851 20934 3885
rect 20783 3835 20934 3851
rect 20783 3796 20843 3835
rect 21203 3796 21263 3902
rect 21557 3961 21617 4128
rect 21675 4102 21735 4128
rect 21698 3962 21765 3969
rect 21692 3961 21765 3962
rect 21557 3953 21765 3961
rect 21557 3919 21715 3953
rect 21749 3919 21765 3953
rect 21557 3903 21765 3919
rect 21557 3902 21754 3903
rect 21319 3868 21385 3884
rect 21319 3834 21335 3868
rect 21369 3834 21385 3868
rect 21319 3818 21385 3834
rect 21437 3869 21503 3884
rect 21437 3835 21453 3869
rect 21487 3835 21503 3869
rect 21437 3819 21503 3835
rect 21321 3796 21381 3818
rect 21439 3796 21499 3819
rect 21557 3796 21617 3902
rect 22081 3900 22141 4524
rect 23913 4056 24209 4092
rect 23913 4035 23973 4056
rect 24031 4035 24091 4056
rect 24149 4035 24209 4056
rect 24267 4055 24563 4091
rect 24267 4035 24327 4055
rect 24385 4035 24445 4055
rect 24503 4035 24563 4055
rect 24621 4055 24917 4091
rect 24621 4035 24681 4055
rect 24739 4035 24799 4055
rect 24857 4035 24917 4055
rect 21991 3884 22141 3900
rect 21991 3850 22007 3884
rect 22041 3850 22141 3884
rect 21991 3834 22141 3850
rect 25507 3902 25567 4600
rect 25809 4552 26105 4612
rect 25809 4529 25869 4552
rect 25927 4529 25987 4552
rect 26045 4529 26105 4552
rect 26163 4553 26459 4613
rect 26804 4612 26865 4632
rect 26163 4529 26223 4553
rect 26281 4529 26341 4553
rect 26399 4529 26459 4553
rect 26785 4596 26865 4612
rect 26785 4562 26800 4596
rect 26834 4562 26865 4596
rect 26785 4546 26865 4562
rect 26804 4523 26865 4546
rect 26805 4377 26865 4523
rect 26804 4204 26865 4377
rect 25809 4103 25869 4129
rect 25777 3962 25844 3969
rect 25927 3962 25987 4129
rect 26045 4103 26105 4129
rect 26163 4103 26223 4129
rect 25777 3953 25987 3962
rect 25777 3919 25793 3953
rect 25827 3919 25987 3953
rect 25777 3903 25987 3919
rect 25507 3886 25658 3902
rect 25507 3852 25608 3886
rect 25642 3852 25658 3886
rect 25507 3836 25658 3852
rect 22081 3796 22141 3834
rect 23913 3809 23973 3835
rect 24031 3809 24091 3835
rect 24149 3809 24209 3835
rect 24267 3815 24327 3835
rect 24267 3809 24328 3815
rect 24385 3809 24445 3835
rect 24503 3809 24563 3835
rect 17996 3752 18012 3786
rect 18046 3752 18062 3786
rect 17996 3736 18062 3752
rect 17878 3669 17944 3685
rect 17878 3635 17894 3669
rect 17928 3635 17944 3669
rect 17878 3619 17944 3635
rect 17881 3597 17941 3619
rect 15426 3569 15486 3595
rect 12650 3369 12710 3395
rect 12768 3369 12828 3395
rect 12886 3369 12946 3395
rect 13004 3369 13064 3395
rect 14548 3369 14608 3395
rect 14666 3369 14726 3395
rect 14784 3369 14844 3395
rect 14902 3369 14962 3395
rect 10873 3174 10933 3196
rect 10991 3174 11051 3196
rect 10870 3158 10936 3174
rect 4437 3110 4503 3126
rect -2469 3071 -2403 3075
rect -2469 3017 -2404 3019
rect -3832 2900 -3806 2960
rect -3406 2900 -3336 2960
rect -3387 2842 -3336 2900
rect -3832 2782 -3806 2842
rect -3406 2782 -3336 2842
rect -3387 2724 -3336 2782
rect -3832 2664 -3806 2724
rect -3406 2664 -3336 2724
rect -3197 2957 -3113 3017
rect -2713 2957 -2687 3017
rect -2469 3003 -2381 3017
rect -2469 2969 -2454 3003
rect -2420 2969 -2381 3003
rect -2469 2957 -2381 2969
rect -1981 2957 -1955 3017
rect -3197 2899 -3137 2957
rect -2469 2953 -2404 2957
rect 10870 3124 10886 3158
rect 10920 3124 10936 3158
rect 10870 3108 10936 3124
rect 10988 3158 11054 3174
rect 10988 3124 11004 3158
rect 11038 3124 11054 3158
rect 18885 3570 18945 3596
rect 17881 3371 17941 3397
rect 20183 3570 20243 3596
rect 20783 3570 20843 3596
rect 24150 3624 24208 3809
rect 24150 3598 24210 3624
rect 24268 3598 24328 3809
rect 24621 3803 24681 3835
rect 24739 3809 24799 3835
rect 24857 3809 24917 3835
rect 24618 3787 24684 3803
rect 25507 3797 25567 3836
rect 25927 3797 25987 3903
rect 26281 3962 26341 4129
rect 26399 4103 26459 4129
rect 26424 3962 26491 3969
rect 26281 3953 26491 3962
rect 26281 3919 26441 3953
rect 26475 3919 26491 3953
rect 26281 3903 26491 3919
rect 26043 3869 26109 3885
rect 26043 3835 26059 3869
rect 26093 3835 26109 3869
rect 26043 3819 26109 3835
rect 26161 3870 26227 3885
rect 26161 3836 26177 3870
rect 26211 3836 26227 3870
rect 26161 3820 26227 3836
rect 26045 3797 26105 3819
rect 26163 3797 26223 3820
rect 26281 3797 26341 3903
rect 26805 3901 26865 4204
rect 26715 3885 26865 3901
rect 26715 3851 26731 3885
rect 26765 3851 26865 3885
rect 26715 3835 26865 3851
rect 26805 3797 26865 3835
rect 27405 4096 27465 4754
rect 28118 4752 28661 4803
rect 28703 4796 28779 4803
rect 28837 4796 28897 4822
rect 36697 4882 36751 4942
rect 37151 4882 37177 4942
rect 36697 4824 36736 4882
rect 37476 4824 37525 4982
rect 37958 4942 38024 4945
rect 38557 4987 38623 5003
rect 38557 4953 38573 4987
rect 38607 4953 38623 4987
rect 37958 4929 38084 4942
rect 37958 4895 37974 4929
rect 38008 4895 38084 4929
rect 37958 4882 38084 4895
rect 38484 4882 38510 4942
rect 38557 4937 38623 4953
rect 37958 4879 38024 4882
rect 28703 4752 28778 4796
rect 36697 4764 36751 4824
rect 37151 4764 37525 4824
rect 37567 4824 37636 4829
rect 37567 4810 38084 4824
rect 37567 4776 37584 4810
rect 37618 4776 38084 4810
rect 37567 4764 38084 4776
rect 38484 4764 38510 4824
rect 27707 4552 28003 4612
rect 27707 4529 27767 4552
rect 27825 4529 27885 4552
rect 27943 4529 28003 4552
rect 28061 4553 28357 4613
rect 28061 4529 28121 4553
rect 28179 4529 28239 4553
rect 28297 4529 28357 4553
rect 28703 4599 28763 4752
rect 36697 4706 36736 4764
rect 37567 4760 37634 4764
rect 36697 4646 36751 4706
rect 37151 4646 37177 4706
rect 28703 4575 28957 4599
rect 28703 4541 28907 4575
rect 28941 4541 28957 4575
rect 28703 4525 28957 4541
rect 27707 4103 27767 4129
rect 27405 4080 27472 4096
rect 27405 4046 27421 4080
rect 27455 4046 27472 4080
rect 27405 4030 27472 4046
rect 27405 3902 27465 4030
rect 27675 3962 27742 3969
rect 27825 3962 27885 4129
rect 27943 4103 28003 4129
rect 28061 4103 28121 4129
rect 27675 3953 27885 3962
rect 27675 3919 27691 3953
rect 27725 3919 27885 3953
rect 27675 3903 27885 3919
rect 27405 3886 27556 3902
rect 27405 3852 27506 3886
rect 27540 3852 27556 3886
rect 27405 3836 27556 3852
rect 27405 3797 27465 3836
rect 27825 3797 27885 3903
rect 28179 3962 28239 4129
rect 28297 4103 28357 4129
rect 28320 3963 28387 3970
rect 28314 3962 28387 3963
rect 28179 3954 28387 3962
rect 28179 3920 28337 3954
rect 28371 3920 28387 3954
rect 28179 3904 28387 3920
rect 28179 3903 28376 3904
rect 27941 3869 28007 3885
rect 27941 3835 27957 3869
rect 27991 3835 28007 3869
rect 27941 3819 28007 3835
rect 28059 3870 28125 3885
rect 28059 3836 28075 3870
rect 28109 3836 28125 3870
rect 28059 3820 28125 3836
rect 27943 3797 28003 3819
rect 28061 3797 28121 3820
rect 28179 3797 28239 3903
rect 28703 3901 28763 4525
rect 29777 4516 30073 4552
rect 29777 4495 29837 4516
rect 29895 4495 29955 4516
rect 30013 4495 30073 4516
rect 30131 4515 30427 4551
rect 30131 4495 30191 4515
rect 30249 4495 30309 4515
rect 30367 4495 30427 4515
rect 30485 4515 30781 4551
rect 30485 4495 30545 4515
rect 30603 4495 30663 4515
rect 30721 4495 30781 4515
rect 36697 4409 36751 4469
rect 37151 4409 37177 4469
rect 36697 4351 36736 4409
rect 37567 4351 37624 4760
rect 38565 4628 38616 4937
rect 29777 4269 29837 4295
rect 29895 4269 29955 4295
rect 30013 4269 30073 4295
rect 30131 4275 30191 4295
rect 30131 4269 30192 4275
rect 30249 4269 30309 4295
rect 30367 4269 30427 4295
rect 30014 4084 30072 4269
rect 30014 4058 30074 4084
rect 30132 4058 30192 4269
rect 30485 4263 30545 4295
rect 30603 4269 30663 4295
rect 30721 4269 30781 4295
rect 36697 4291 36751 4351
rect 37151 4291 37624 4351
rect 37836 4568 38084 4628
rect 38284 4568 38616 4628
rect 30482 4247 30548 4263
rect 30482 4213 30498 4247
rect 30532 4213 30548 4247
rect 30482 4197 30548 4213
rect 36697 4233 36736 4291
rect 36697 4173 36751 4233
rect 37151 4173 37177 4233
rect 30364 4130 30430 4146
rect 30364 4096 30380 4130
rect 30414 4096 30430 4130
rect 30364 4080 30430 4096
rect 30367 4058 30427 4080
rect 28613 3885 28763 3901
rect 28613 3851 28629 3885
rect 28663 3851 28763 3885
rect 28613 3835 28763 3851
rect 28703 3797 28763 3835
rect 24618 3753 24634 3787
rect 24668 3753 24684 3787
rect 24618 3737 24684 3753
rect 24500 3670 24566 3686
rect 24500 3636 24516 3670
rect 24550 3636 24566 3670
rect 24500 3620 24566 3636
rect 24503 3598 24563 3620
rect 22081 3570 22141 3596
rect 19305 3370 19365 3396
rect 19423 3370 19483 3396
rect 19541 3370 19601 3396
rect 19659 3370 19719 3396
rect 21203 3370 21263 3396
rect 21321 3370 21381 3396
rect 21439 3370 21499 3396
rect 21557 3370 21617 3396
rect 17528 3175 17588 3197
rect 17646 3175 17706 3197
rect 17525 3159 17591 3175
rect 10988 3108 11054 3124
rect 17525 3125 17541 3159
rect 17575 3125 17591 3159
rect 17525 3109 17591 3125
rect 17643 3159 17709 3175
rect 17643 3125 17659 3159
rect 17693 3125 17709 3159
rect 25507 3571 25567 3597
rect 24503 3372 24563 3398
rect 26805 3571 26865 3597
rect 27405 3571 27465 3597
rect 36896 3936 36951 3996
rect 37151 3936 37177 3996
rect 36896 3878 36935 3936
rect 30367 3832 30427 3858
rect 36896 3818 36951 3878
rect 37151 3818 37177 3878
rect 37297 3854 37363 3870
rect 37297 3820 37313 3854
rect 37347 3820 37363 3854
rect 36896 3760 36935 3818
rect 37297 3804 37363 3820
rect 37300 3760 37360 3804
rect 37836 3760 37881 4568
rect 36896 3700 36951 3760
rect 37151 3700 37881 3760
rect 30014 3636 30074 3658
rect 30132 3636 30192 3658
rect 30011 3620 30077 3636
rect 28703 3571 28763 3597
rect 30011 3586 30027 3620
rect 30061 3586 30077 3620
rect 30011 3570 30077 3586
rect 30129 3620 30195 3636
rect 30129 3586 30145 3620
rect 30179 3586 30195 3620
rect 30129 3570 30195 3586
rect 25927 3371 25987 3397
rect 26045 3371 26105 3397
rect 26163 3371 26223 3397
rect 26281 3371 26341 3397
rect 27825 3371 27885 3397
rect 27943 3371 28003 3397
rect 28061 3371 28121 3397
rect 28179 3371 28239 3397
rect 24150 3176 24210 3198
rect 24268 3176 24328 3198
rect 24147 3160 24213 3176
rect 17643 3109 17709 3125
rect 24147 3126 24163 3160
rect 24197 3126 24213 3160
rect 24147 3110 24213 3126
rect 24265 3160 24331 3176
rect 24265 3126 24281 3160
rect 24315 3126 24331 3160
rect 24265 3110 24331 3126
rect 32008 2965 32304 3016
rect 32008 2950 32068 2965
rect 32126 2950 32186 2965
rect 32244 2950 32304 2965
rect 32362 2950 32422 2976
rect 32480 2950 32540 2976
rect 32598 2950 32658 2976
rect -3197 2839 -3113 2899
rect -2713 2839 -2381 2899
rect -1981 2839 -1955 2899
rect -3197 2781 -3137 2839
rect -3197 2721 -3113 2781
rect -2713 2721 -2687 2781
rect -2546 2756 -2487 2839
rect -2553 2739 -2487 2756
rect 31524 2750 31584 2776
rect 31642 2750 31702 2776
rect 31760 2750 31820 2776
rect -3387 2477 -3336 2664
rect -2553 2705 -2537 2739
rect -2503 2705 -2487 2739
rect -2553 2689 -2487 2705
rect 36896 3000 36951 3060
rect 37151 3001 37881 3060
rect 37151 3000 37454 3001
rect 36896 2942 36935 3000
rect 37437 2943 37454 3000
rect 37509 3000 37881 3001
rect 37509 2943 37524 3000
rect 36896 2882 36951 2942
rect 37151 2882 37177 2942
rect 37437 2924 37524 2943
rect 36896 2824 36935 2882
rect 32845 2767 33141 2818
rect 32845 2750 32905 2767
rect 32963 2750 33023 2767
rect 33081 2750 33141 2767
rect 33317 2768 33613 2804
rect 33317 2747 33377 2768
rect 33435 2747 33495 2768
rect 33553 2747 33613 2768
rect 33671 2767 33967 2803
rect 33671 2747 33731 2767
rect 33789 2747 33849 2767
rect 33907 2747 33967 2767
rect 34025 2767 34321 2803
rect 34025 2747 34085 2767
rect 34143 2747 34203 2767
rect 34261 2747 34321 2767
rect 36896 2764 36951 2824
rect 37151 2764 37177 2824
rect 31524 2533 31584 2550
rect 31642 2533 31702 2550
rect 31760 2533 31820 2550
rect 32008 2533 32068 2550
rect 31524 2482 32068 2533
rect 32126 2524 32186 2550
rect 32244 2524 32304 2550
rect 32362 2531 32422 2550
rect 32480 2531 32540 2550
rect 32598 2531 32658 2550
rect 32845 2531 32905 2550
rect 32963 2531 33023 2550
rect -3674 2417 -3606 2477
rect -3406 2417 -3336 2477
rect -2485 2449 -2419 2465
rect -3249 2427 -3195 2443
rect -3674 2359 -3623 2417
rect -3249 2393 -3239 2427
rect -3205 2393 -3195 2427
rect -3249 2375 -3195 2393
rect -2485 2415 -2469 2449
rect -2435 2415 -2419 2449
rect -2485 2375 -2419 2415
rect -3387 2359 -2381 2375
rect -3674 2299 -3606 2359
rect -3406 2315 -2381 2359
rect -2181 2315 -2155 2375
rect -3406 2300 -3336 2315
rect -3406 2299 -3380 2300
rect -3674 2241 -3623 2299
rect 31649 2278 31709 2482
rect 32362 2480 32905 2531
rect 32947 2524 33023 2531
rect 33081 2524 33141 2550
rect 36697 2559 36751 2619
rect 37151 2559 37177 2619
rect 32947 2480 33022 2524
rect 33317 2521 33377 2547
rect 33435 2521 33495 2547
rect 33553 2521 33613 2547
rect 33671 2527 33731 2547
rect 33671 2521 33732 2527
rect 33789 2521 33849 2547
rect 33907 2521 33967 2547
rect 32947 2398 33007 2480
rect 32947 2380 33181 2398
rect 32947 2346 33130 2380
rect 33164 2346 33181 2380
rect 31951 2280 32247 2340
rect 8127 2241 8193 2257
rect -3674 2181 -3606 2241
rect -3406 2181 -3380 2241
rect 8127 2207 8143 2241
rect 8177 2207 8193 2241
rect 8127 2191 8193 2207
rect 8245 2241 8311 2257
rect 8245 2207 8261 2241
rect 8295 2207 8311 2241
rect 8245 2191 8311 2207
rect 14681 2246 14747 2262
rect 14681 2212 14697 2246
rect 14731 2212 14747 2246
rect 14681 2196 14747 2212
rect 14799 2246 14865 2262
rect 31649 2261 31780 2278
rect 14799 2212 14815 2246
rect 14849 2212 14865 2246
rect 14799 2196 14865 2212
rect 21330 2234 21396 2250
rect 21330 2200 21346 2234
rect 21380 2200 21396 2234
rect 8130 2169 8190 2191
rect 8248 2169 8308 2191
rect 14684 2174 14744 2196
rect 14802 2174 14862 2196
rect 21330 2184 21396 2200
rect 21448 2234 21514 2250
rect 21448 2200 21464 2234
rect 21498 2200 21514 2234
rect 21448 2184 21514 2200
rect 31649 2227 31730 2261
rect 31764 2227 31780 2261
rect 31951 2257 32011 2280
rect 32069 2257 32129 2280
rect 32187 2257 32247 2280
rect 32305 2281 32601 2341
rect 32305 2257 32365 2281
rect 32423 2257 32483 2281
rect 32541 2257 32601 2281
rect 32947 2330 33181 2346
rect 33554 2336 33612 2521
rect 31649 2210 31780 2227
rect 8483 1969 8543 1995
rect 21333 2162 21393 2184
rect 21451 2162 21511 2184
rect 15037 1974 15097 2000
rect -3061 1753 -3001 1769
rect -3634 1670 -3608 1730
rect -3408 1670 -3340 1730
rect -3391 1612 -3340 1670
rect -3634 1552 -3608 1612
rect -3408 1605 -3340 1612
rect -3061 1719 -3047 1753
rect -3013 1719 -3001 1753
rect -3061 1605 -3001 1719
rect 8130 1743 8190 1769
rect -3408 1552 -2383 1605
rect -3391 1545 -2383 1552
rect -2183 1545 -2157 1605
rect 8130 1558 8188 1743
rect 8248 1558 8308 1769
rect 8483 1747 8543 1769
rect 14684 1748 14744 1774
rect 8480 1731 8546 1747
rect 8480 1697 8496 1731
rect 8530 1697 8546 1731
rect 8480 1681 8546 1697
rect 8598 1614 8664 1630
rect 8598 1580 8614 1614
rect 8648 1580 8664 1614
rect 8598 1564 8664 1580
rect -3391 1494 -3340 1545
rect -3634 1434 -3608 1494
rect -3408 1434 -3340 1494
rect -2488 1504 -2422 1545
rect -2488 1470 -2472 1504
rect -2438 1470 -2422 1504
rect 7893 1532 7953 1558
rect 8011 1532 8071 1558
rect 8129 1532 8189 1558
rect 8247 1552 8308 1558
rect 8247 1532 8307 1552
rect 8365 1532 8425 1558
rect 8483 1532 8543 1558
rect 8601 1532 8661 1564
rect 14684 1563 14742 1748
rect 14802 1563 14862 1774
rect 15037 1752 15097 1774
rect 21686 1962 21746 1988
rect 15034 1736 15100 1752
rect 15034 1702 15050 1736
rect 15084 1702 15100 1736
rect 15034 1686 15100 1702
rect 21333 1736 21393 1762
rect 15152 1619 15218 1635
rect 15152 1585 15168 1619
rect 15202 1585 15218 1619
rect 15152 1569 15218 1585
rect 8719 1532 8779 1558
rect 8837 1532 8897 1558
rect 14447 1537 14507 1563
rect 14565 1537 14625 1563
rect 14683 1537 14743 1563
rect 14801 1557 14862 1563
rect 14801 1537 14861 1557
rect 14919 1537 14979 1563
rect 15037 1537 15097 1563
rect 15155 1537 15215 1569
rect 15273 1537 15333 1563
rect 15391 1537 15451 1563
rect 21333 1551 21391 1736
rect 21451 1551 21511 1762
rect 21686 1740 21746 1762
rect 21683 1724 21749 1740
rect 21683 1690 21699 1724
rect 21733 1690 21749 1724
rect 21683 1674 21749 1690
rect 29784 1671 30080 1707
rect 29784 1650 29844 1671
rect 29902 1650 29962 1671
rect 30020 1650 30080 1671
rect 30138 1670 30434 1706
rect 30138 1650 30198 1670
rect 30256 1650 30316 1670
rect 30374 1650 30434 1670
rect 30492 1670 30788 1706
rect 30492 1650 30552 1670
rect 30610 1650 30670 1670
rect 30728 1650 30788 1670
rect 21801 1607 21867 1623
rect 21801 1573 21817 1607
rect 21851 1573 21867 1607
rect 21801 1557 21867 1573
rect -2488 1454 -2422 1470
rect -3391 1246 -3340 1434
rect -2555 1319 -2489 1335
rect 21096 1525 21156 1551
rect 21214 1525 21274 1551
rect 21332 1525 21392 1551
rect 21450 1545 21511 1551
rect 21450 1525 21510 1545
rect 21568 1525 21628 1551
rect 21686 1525 21746 1551
rect 21804 1525 21864 1557
rect 21922 1525 21982 1551
rect 22040 1525 22100 1551
rect -3874 1186 -3808 1246
rect -3408 1186 -3340 1246
rect -3198 1243 -3115 1303
rect -2715 1243 -2689 1303
rect -2555 1285 -2539 1319
rect -2505 1285 -2489 1319
rect -2555 1268 -2489 1285
rect 7893 1311 7953 1332
rect 8011 1311 8071 1332
rect 8129 1311 8189 1332
rect 7893 1275 8189 1311
rect 8247 1312 8307 1332
rect 8365 1312 8425 1332
rect 8483 1312 8543 1332
rect 8247 1276 8543 1312
rect 8601 1312 8661 1332
rect 8719 1312 8779 1332
rect 8837 1312 8897 1332
rect 8601 1276 8897 1312
rect 14447 1316 14507 1337
rect 14565 1316 14625 1337
rect 14683 1316 14743 1337
rect 14447 1280 14743 1316
rect 14801 1317 14861 1337
rect 14919 1317 14979 1337
rect 15037 1317 15097 1337
rect 14801 1281 15097 1317
rect 15155 1317 15215 1337
rect 15273 1317 15333 1337
rect 15391 1317 15451 1337
rect 31649 1630 31709 2210
rect 31951 1831 32011 1857
rect 31919 1690 31986 1697
rect 32069 1690 32129 1857
rect 32187 1831 32247 1857
rect 32305 1831 32365 1857
rect 31919 1681 32129 1690
rect 31919 1647 31935 1681
rect 31969 1647 32129 1681
rect 31919 1631 32129 1647
rect 31649 1614 31800 1630
rect 31649 1580 31750 1614
rect 31784 1580 31800 1614
rect 31649 1564 31800 1580
rect 31649 1525 31709 1564
rect 32069 1525 32129 1631
rect 32423 1690 32483 1857
rect 32541 1831 32601 1857
rect 32566 1690 32633 1697
rect 32423 1681 32633 1690
rect 32423 1647 32583 1681
rect 32617 1647 32633 1681
rect 32423 1631 32633 1647
rect 32185 1597 32251 1613
rect 32185 1563 32201 1597
rect 32235 1563 32251 1597
rect 32185 1547 32251 1563
rect 32303 1598 32369 1613
rect 32303 1564 32319 1598
rect 32353 1564 32369 1598
rect 32303 1548 32369 1564
rect 32187 1525 32247 1547
rect 32305 1525 32365 1548
rect 32423 1525 32483 1631
rect 32947 1629 33007 2330
rect 33554 2310 33614 2336
rect 33672 2310 33732 2521
rect 34025 2515 34085 2547
rect 34143 2521 34203 2547
rect 34261 2521 34321 2547
rect 34022 2499 34088 2515
rect 34022 2465 34038 2499
rect 34072 2465 34088 2499
rect 34022 2449 34088 2465
rect 36697 2501 36736 2559
rect 36697 2441 36751 2501
rect 37151 2441 37626 2501
rect 33904 2382 33970 2398
rect 33904 2348 33920 2382
rect 33954 2348 33970 2382
rect 33904 2332 33970 2348
rect 36697 2383 36736 2441
rect 33907 2310 33967 2332
rect 36697 2323 36751 2383
rect 37151 2323 37177 2383
rect 33907 2084 33967 2110
rect 36697 2092 36751 2152
rect 37151 2092 37177 2152
rect 36697 2034 36736 2092
rect 36697 1974 36751 2034
rect 37151 2033 37177 2034
rect 37338 2033 37404 2036
rect 37151 2020 37404 2033
rect 37151 1986 37354 2020
rect 37388 1986 37404 2020
rect 37151 1974 37404 1986
rect 37569 2034 37626 2441
rect 37836 2226 37881 3000
rect 37836 2166 38084 2226
rect 38284 2166 38310 2226
rect 37725 2034 37804 2045
rect 37569 2032 38084 2034
rect 37569 1974 37738 2032
rect 37793 1974 38084 2032
rect 38484 1974 38510 2034
rect 33554 1888 33614 1910
rect 33672 1888 33732 1910
rect 33551 1872 33617 1888
rect 33551 1838 33567 1872
rect 33601 1838 33617 1872
rect 33551 1822 33617 1838
rect 33669 1872 33735 1888
rect 33669 1838 33685 1872
rect 33719 1838 33735 1872
rect 33669 1822 33735 1838
rect 36697 1916 36736 1974
rect 37337 1970 37404 1974
rect 37725 1964 37804 1974
rect 37438 1916 37525 1933
rect 36697 1856 36751 1916
rect 37151 1856 37177 1916
rect 37438 1914 38084 1916
rect 37438 1856 37453 1914
rect 37508 1856 38084 1914
rect 38484 1856 38510 1916
rect 37438 1838 37525 1856
rect 36697 1738 36751 1798
rect 37151 1738 37177 1798
rect 36697 1680 36736 1738
rect 37476 1680 37525 1838
rect 37958 1798 38024 1801
rect 38557 1843 38623 1859
rect 38557 1809 38573 1843
rect 38607 1809 38623 1843
rect 37958 1785 38084 1798
rect 37958 1751 37974 1785
rect 38008 1751 38084 1785
rect 37958 1738 38084 1751
rect 38484 1738 38510 1798
rect 38557 1793 38623 1809
rect 37958 1735 38024 1738
rect 32857 1613 33007 1629
rect 32857 1579 32873 1613
rect 32907 1579 33007 1613
rect 32857 1563 33007 1579
rect 32947 1525 33007 1563
rect 36697 1620 36751 1680
rect 37151 1620 37525 1680
rect 37567 1680 37636 1685
rect 37567 1666 38084 1680
rect 37567 1632 37584 1666
rect 37618 1632 38084 1666
rect 37567 1620 38084 1632
rect 38484 1620 38510 1680
rect 36697 1562 36736 1620
rect 37567 1616 37634 1620
rect 29784 1424 29844 1450
rect 29902 1424 29962 1450
rect 30020 1424 30080 1450
rect 30138 1430 30198 1450
rect 30138 1424 30199 1430
rect 30256 1424 30316 1450
rect 30374 1424 30434 1450
rect 15155 1281 15451 1317
rect 21096 1304 21156 1325
rect 21214 1304 21274 1325
rect 21332 1304 21392 1325
rect 21096 1268 21392 1304
rect 21450 1305 21510 1325
rect 21568 1305 21628 1325
rect 21686 1305 21746 1325
rect 21450 1269 21746 1305
rect 21804 1305 21864 1325
rect 21922 1305 21982 1325
rect 22040 1305 22100 1325
rect 21804 1269 22100 1305
rect -3874 1128 -3823 1186
rect -3198 1185 -3138 1243
rect -2548 1185 -2489 1268
rect 30021 1239 30079 1424
rect 30021 1213 30081 1239
rect 30139 1213 30199 1424
rect 30492 1418 30552 1450
rect 30610 1424 30670 1450
rect 30728 1424 30788 1450
rect 30489 1402 30555 1418
rect 30489 1368 30505 1402
rect 30539 1368 30555 1402
rect 30489 1352 30555 1368
rect 30371 1285 30437 1301
rect 31649 1299 31709 1325
rect 30371 1251 30387 1285
rect 30421 1251 30437 1285
rect 30371 1235 30437 1251
rect 30374 1213 30434 1235
rect -3874 1068 -3808 1128
rect -3408 1068 -3382 1128
rect -3198 1125 -3115 1185
rect -2715 1125 -2383 1185
rect -1983 1125 -1957 1185
rect -3874 1010 -3823 1068
rect -3198 1067 -3138 1125
rect -2471 1067 -2405 1069
rect -3874 950 -3808 1010
rect -3408 950 -3382 1010
rect -3198 1007 -3115 1067
rect -2715 1007 -2689 1067
rect -2471 1053 -2383 1067
rect -2471 1019 -2455 1053
rect -2421 1019 -2383 1053
rect -2471 1007 -2383 1019
rect -1983 1007 -1957 1067
rect -2471 1003 -2405 1007
rect -2471 949 -2406 951
rect -3834 832 -3808 892
rect -3408 832 -3338 892
rect -3389 774 -3338 832
rect -3834 714 -3808 774
rect -3408 714 -3338 774
rect -3389 656 -3338 714
rect -3834 596 -3808 656
rect -3408 596 -3338 656
rect -3199 889 -3115 949
rect -2715 889 -2689 949
rect -2471 935 -2383 949
rect -2471 901 -2456 935
rect -2422 901 -2383 935
rect -2471 889 -2383 901
rect -1983 889 -1957 949
rect -3199 831 -3139 889
rect -2471 885 -2406 889
rect -3199 771 -3115 831
rect -2715 771 -2383 831
rect -1983 771 -1957 831
rect 36697 1502 36751 1562
rect 37151 1502 37177 1562
rect 32947 1299 33007 1325
rect 36697 1265 36751 1325
rect 37151 1265 37177 1325
rect 36697 1207 36736 1265
rect 37567 1207 37624 1616
rect 38565 1484 38616 1793
rect 36697 1147 36751 1207
rect 37151 1147 37624 1207
rect 37836 1424 38084 1484
rect 38284 1424 38616 1484
rect 32069 1099 32129 1125
rect 32187 1099 32247 1125
rect 32305 1099 32365 1125
rect 32423 1099 32483 1125
rect 36697 1089 36736 1147
rect 36697 1029 36751 1089
rect 37151 1029 37177 1089
rect 30374 987 30434 1013
rect 30021 791 30081 813
rect 30139 791 30199 813
rect 36896 792 36951 852
rect 37151 792 37177 852
rect 30018 775 30084 791
rect -3199 713 -3139 771
rect -3199 653 -3115 713
rect -2715 653 -2689 713
rect -2548 688 -2489 771
rect 30018 741 30034 775
rect 30068 741 30084 775
rect 30018 725 30084 741
rect 30136 775 30202 791
rect 30136 741 30152 775
rect 30186 741 30202 775
rect 30136 725 30202 741
rect 36896 734 36935 792
rect -2555 671 -2489 688
rect -3389 409 -3338 596
rect -2555 637 -2539 671
rect -2505 637 -2489 671
rect -2555 621 -2489 637
rect 36896 674 36951 734
rect 37151 674 37177 734
rect 37297 710 37363 726
rect 37297 676 37313 710
rect 37347 676 37363 710
rect 36896 616 36935 674
rect 37297 660 37363 676
rect 37300 616 37360 660
rect 37836 616 37881 1424
rect 36896 556 36951 616
rect 37151 556 37881 616
rect -3676 349 -3608 409
rect -3408 349 -3338 409
rect -2487 381 -2421 397
rect -3251 359 -3197 375
rect -3676 291 -3625 349
rect -3251 325 -3241 359
rect -3207 325 -3197 359
rect -3251 307 -3197 325
rect -2487 347 -2471 381
rect -2437 347 -2421 381
rect -2487 307 -2421 347
rect -3389 291 -2383 307
rect -3676 231 -3608 291
rect -3408 247 -2383 291
rect -2183 247 -2157 307
rect -3408 232 -3338 247
rect -3408 231 -3382 232
rect -3676 173 -3625 231
rect -3676 113 -3608 173
rect -3408 113 -3382 173
<< polycont >>
rect 8052 27822 8086 27856
rect 9182 27828 9216 27862
rect 14565 27819 14599 27853
rect 15695 27825 15729 27859
rect 8052 27704 8086 27738
rect 9182 27708 9216 27742
rect 21099 27814 21133 27848
rect 22229 27820 22263 27854
rect 14565 27701 14599 27735
rect 6609 27338 6643 27372
rect 15695 27705 15729 27739
rect 27657 27818 27691 27852
rect 28787 27824 28821 27858
rect 21099 27696 21133 27730
rect 6491 27221 6525 27255
rect 8372 26948 8406 26982
rect 13122 27335 13156 27369
rect 22229 27700 22263 27734
rect 27657 27700 27691 27734
rect 13004 27218 13038 27252
rect 9514 26952 9548 26986
rect 6138 26711 6172 26745
rect 6256 26711 6290 26745
rect 14885 26945 14919 26979
rect 19656 27330 19690 27364
rect 28787 27704 28821 27738
rect 19538 27213 19572 27247
rect 16027 26949 16061 26983
rect 12651 26708 12685 26742
rect 12769 26708 12803 26742
rect 21419 26940 21453 26974
rect 26214 27334 26248 27368
rect 26096 27217 26130 27251
rect 22561 26944 22595 26978
rect 19185 26703 19219 26737
rect 19303 26703 19337 26737
rect 27977 26944 28011 26978
rect 29119 26948 29153 26982
rect 25743 26707 25777 26741
rect 25861 26707 25895 26741
rect 6623 25688 6657 25722
rect 6505 25571 6539 25605
rect 6152 25061 6186 25095
rect 6270 25061 6304 25095
rect 13136 25685 13170 25719
rect 13018 25568 13052 25602
rect 8784 24893 8818 24927
rect 7777 24250 7811 24284
rect 7592 24183 7626 24217
rect 8425 24250 8459 24284
rect 8043 24166 8077 24200
rect 8161 24167 8195 24201
rect 8715 24182 8749 24216
rect 12665 25058 12699 25092
rect 12783 25058 12817 25092
rect 19670 25680 19704 25714
rect 19552 25563 19586 25597
rect 10891 24872 10925 24906
rect 9405 24377 9439 24411
rect 9675 24250 9709 24284
rect 9490 24183 9524 24217
rect 10321 24251 10355 24285
rect 9941 24166 9975 24200
rect 10059 24167 10093 24201
rect 10613 24182 10647 24216
rect 15297 24890 15331 24924
rect 14290 24247 14324 24281
rect 14105 24180 14139 24214
rect 6618 24084 6652 24118
rect 6500 23967 6534 24001
rect 14938 24247 14972 24281
rect 14556 24163 14590 24197
rect 14674 24164 14708 24198
rect 15228 24179 15262 24213
rect 19199 25053 19233 25087
rect 19317 25053 19351 25087
rect 26228 25684 26262 25718
rect 26110 25567 26144 25601
rect 17404 24869 17438 24903
rect 15918 24374 15952 24408
rect 16188 24247 16222 24281
rect 16003 24180 16037 24214
rect 16834 24248 16868 24282
rect 16454 24163 16488 24197
rect 16572 24164 16606 24198
rect 17126 24179 17160 24213
rect 21831 24885 21865 24919
rect 20824 24242 20858 24276
rect 20639 24175 20673 24209
rect 13131 24081 13165 24115
rect 13013 23964 13047 23998
rect 6147 23457 6181 23491
rect 6265 23457 6299 23491
rect 21472 24242 21506 24276
rect 21090 24158 21124 24192
rect 21208 24159 21242 24193
rect 21762 24174 21796 24208
rect 25757 25057 25791 25091
rect 25875 25057 25909 25091
rect 23938 24864 23972 24898
rect 22452 24369 22486 24403
rect 22722 24242 22756 24276
rect 22537 24175 22571 24209
rect 23368 24243 23402 24277
rect 22988 24158 23022 24192
rect 23106 24159 23140 24193
rect 23660 24174 23694 24208
rect 28389 24889 28423 24923
rect 27382 24246 27416 24280
rect 27197 24179 27231 24213
rect 19665 24076 19699 24110
rect 19547 23959 19581 23993
rect 12660 23454 12694 23488
rect 12778 23454 12812 23488
rect 28030 24246 28064 24280
rect 27648 24162 27682 24196
rect 27766 24163 27800 24197
rect 28320 24178 28354 24212
rect 37458 24985 37513 25043
rect 30496 24868 30530 24902
rect 29010 24373 29044 24407
rect 29280 24246 29314 24280
rect 29095 24179 29129 24213
rect 29926 24247 29960 24281
rect 29546 24162 29580 24196
rect 29664 24163 29698 24197
rect 30218 24178 30252 24212
rect 26223 24080 26257 24114
rect 26105 23963 26139 23997
rect 19194 23449 19228 23483
rect 19312 23449 19346 23483
rect 37358 24028 37392 24062
rect 37742 24016 37797 24074
rect 37457 23898 37512 23956
rect 38577 23851 38611 23885
rect 37978 23793 38012 23827
rect 37588 23674 37622 23708
rect 25752 23453 25786 23487
rect 25870 23453 25904 23487
rect 37317 22718 37351 22752
rect 6688 22220 6722 22254
rect 7818 22214 7852 22248
rect 13246 22216 13280 22250
rect 14376 22210 14410 22244
rect 6688 22100 6722 22134
rect 7818 22096 7852 22130
rect 19780 22221 19814 22255
rect 20910 22215 20944 22249
rect 13246 22096 13280 22130
rect 9261 21730 9295 21764
rect 6356 21344 6390 21378
rect 9379 21613 9413 21647
rect 14376 22092 14410 22126
rect 7498 21340 7532 21374
rect 26293 22224 26327 22258
rect 27423 22218 27457 22252
rect 19780 22101 19814 22135
rect 15819 21726 15853 21760
rect 12914 21340 12948 21374
rect 15937 21609 15971 21643
rect 20910 22097 20944 22131
rect 14056 21336 14090 21370
rect 9614 21103 9648 21137
rect 9732 21103 9766 21137
rect 26293 22104 26327 22138
rect 22353 21731 22387 21765
rect 19448 21345 19482 21379
rect 22471 21614 22505 21648
rect 27423 22100 27457 22134
rect 20590 21341 20624 21375
rect 16172 21099 16206 21133
rect 16290 21099 16324 21133
rect 37458 21841 37513 21899
rect 28866 21734 28900 21768
rect 25961 21348 25995 21382
rect 28984 21617 29018 21651
rect 27103 21344 27137 21378
rect 22706 21104 22740 21138
rect 22824 21104 22858 21138
rect 29219 21107 29253 21141
rect 29337 21107 29371 21141
rect 37358 20884 37392 20918
rect 37742 20872 37797 20930
rect 37457 20754 37512 20812
rect 38577 20707 38611 20741
rect 37978 20649 38012 20683
rect 37588 20530 37622 20564
rect 9247 20080 9281 20114
rect 9365 19963 9399 19997
rect 15805 20076 15839 20110
rect 15923 19959 15957 19993
rect 4979 19264 5013 19298
rect 5549 18643 5583 18677
rect 5257 18574 5291 18608
rect 22339 20081 22373 20115
rect 22457 19964 22491 19998
rect 6465 18769 6499 18803
rect 6195 18642 6229 18676
rect 5811 18559 5845 18593
rect 5929 18558 5963 18592
rect 6380 18575 6414 18609
rect 9600 19453 9634 19487
rect 9718 19453 9752 19487
rect 7086 19285 7120 19319
rect 7445 18642 7479 18676
rect 7155 18574 7189 18608
rect 8093 18642 8127 18676
rect 7709 18559 7743 18593
rect 7827 18558 7861 18592
rect 11537 19260 11571 19294
rect 8278 18575 8312 18609
rect 12107 18639 12141 18673
rect 11815 18570 11849 18604
rect 9252 18476 9286 18510
rect 9370 18359 9404 18393
rect 28852 20084 28886 20118
rect 28970 19967 29004 20001
rect 13023 18765 13057 18799
rect 12753 18638 12787 18672
rect 12369 18555 12403 18589
rect 12487 18554 12521 18588
rect 12938 18571 12972 18605
rect 16158 19449 16192 19483
rect 16276 19449 16310 19483
rect 13644 19281 13678 19315
rect 14003 18638 14037 18672
rect 13713 18570 13747 18604
rect 14651 18638 14685 18672
rect 14267 18555 14301 18589
rect 14385 18554 14419 18588
rect 18071 19265 18105 19299
rect 14836 18571 14870 18605
rect 18641 18644 18675 18678
rect 18349 18575 18383 18609
rect 15810 18472 15844 18506
rect 15928 18355 15962 18389
rect 19557 18770 19591 18804
rect 19287 18643 19321 18677
rect 18903 18560 18937 18594
rect 19021 18559 19055 18593
rect 19472 18576 19506 18610
rect 22692 19454 22726 19488
rect 22810 19454 22844 19488
rect 20178 19286 20212 19320
rect 20537 18643 20571 18677
rect 20247 18575 20281 18609
rect 21185 18643 21219 18677
rect 20801 18560 20835 18594
rect 20919 18559 20953 18593
rect 24584 19268 24618 19302
rect 21370 18576 21404 18610
rect 25154 18647 25188 18681
rect 24862 18578 24896 18612
rect 9605 17849 9639 17883
rect 9723 17849 9757 17883
rect 22344 18477 22378 18511
rect 22462 18360 22496 18394
rect 37317 19574 37351 19608
rect 26070 18773 26104 18807
rect 25800 18646 25834 18680
rect 25416 18563 25450 18597
rect 25534 18562 25568 18596
rect 25985 18579 26019 18613
rect 29205 19457 29239 19491
rect 29323 19457 29357 19491
rect 26691 19289 26725 19323
rect 27050 18646 27084 18680
rect 26760 18578 26794 18612
rect 27698 18646 27732 18680
rect 27314 18563 27348 18597
rect 27432 18562 27466 18596
rect 27883 18579 27917 18613
rect 37454 18709 37509 18767
rect 16163 17845 16197 17879
rect 16281 17845 16315 17879
rect 28857 18480 28891 18514
rect 28975 18363 29009 18397
rect 22697 17850 22731 17884
rect 22815 17850 22849 17884
rect 29210 17853 29244 17887
rect 29328 17853 29362 17887
rect 37354 17752 37388 17786
rect 37738 17740 37793 17798
rect 37453 17622 37508 17680
rect 38573 17575 38607 17609
rect 37974 17517 38008 17551
rect 37584 17398 37618 17432
rect 37313 16442 37347 16476
rect -3043 16198 -3009 16232
rect -2468 15949 -2434 15983
rect -2535 15764 -2501 15798
rect -2451 15498 -2417 15532
rect 37454 15565 37509 15623
rect -2452 15380 -2418 15414
rect -2535 15116 -2501 15150
rect -3237 14804 -3203 14838
rect -2467 14826 -2433 14860
rect 8579 14954 8613 14988
rect 8461 14837 8495 14871
rect 15128 14953 15162 14987
rect 15010 14836 15044 14870
rect 21782 14974 21816 15008
rect 21664 14857 21698 14891
rect 30435 14807 30469 14841
rect 30317 14690 30351 14724
rect 8108 14327 8142 14361
rect 8226 14327 8260 14361
rect 14657 14326 14691 14360
rect 14775 14326 14809 14360
rect 21311 14347 21345 14381
rect 21429 14347 21463 14381
rect 29964 14180 29998 14214
rect 30082 14180 30116 14214
rect 37354 14608 37388 14642
rect 37738 14596 37793 14654
rect 33128 14280 33162 14314
rect -3045 14130 -3011 14164
rect 31728 14161 31762 14195
rect -2470 13881 -2436 13915
rect -2537 13696 -2503 13730
rect -2453 13430 -2419 13464
rect -2454 13312 -2420 13346
rect 6248 13271 6282 13305
rect 7378 13277 7412 13311
rect 12797 13359 12831 13393
rect 13927 13365 13961 13399
rect 12797 13241 12831 13275
rect 13927 13245 13961 13279
rect 19451 13291 19485 13325
rect 20581 13297 20615 13331
rect 26076 13359 26110 13393
rect 27206 13365 27240 13399
rect 31933 13581 31967 13615
rect 31748 13514 31782 13548
rect 32581 13581 32615 13615
rect 32199 13497 32233 13531
rect 32317 13498 32351 13532
rect 34036 14399 34070 14433
rect 37453 14478 37508 14536
rect 33918 14282 33952 14316
rect 38573 14431 38607 14465
rect 37974 14373 38008 14407
rect 37584 14254 37618 14288
rect 33565 13772 33599 13806
rect 33683 13772 33717 13806
rect 32871 13513 32905 13547
rect 6248 13153 6282 13187
rect 7378 13157 7412 13191
rect -2537 13048 -2503 13082
rect 1915 13054 1949 13088
rect 1797 12937 1831 12971
rect -3239 12736 -3205 12770
rect -2469 12758 -2435 12792
rect 4805 12787 4839 12821
rect 4687 12670 4721 12704
rect 1444 12427 1478 12461
rect 1562 12427 1596 12461
rect 6568 12397 6602 12431
rect 11354 12875 11388 12909
rect 26076 13241 26110 13275
rect 19451 13173 19485 13207
rect 20581 13177 20615 13211
rect 27206 13245 27240 13279
rect 11236 12758 11270 12792
rect 7710 12401 7744 12435
rect 4334 12160 4368 12194
rect 4452 12160 4486 12194
rect 13117 12485 13151 12519
rect 18008 12807 18042 12841
rect 17890 12690 17924 12724
rect 14259 12489 14293 12523
rect 10883 12248 10917 12282
rect 11001 12248 11035 12282
rect 19771 12417 19805 12451
rect 24633 12875 24667 12909
rect 37313 13298 37347 13332
rect 24515 12758 24549 12792
rect 20913 12421 20947 12455
rect 17537 12180 17571 12214
rect 17655 12180 17689 12214
rect 26396 12485 26430 12519
rect 27538 12489 27572 12523
rect 24162 12248 24196 12282
rect 24280 12248 24314 12282
rect 37458 12363 37513 12421
rect -3043 12061 -3009 12095
rect 30430 12236 30464 12270
rect 30312 12119 30346 12153
rect -2468 11812 -2434 11846
rect -2535 11627 -2501 11661
rect 29959 11609 29993 11643
rect -2451 11361 -2417 11395
rect -2452 11243 -2418 11277
rect 30077 11609 30111 11643
rect -2535 10979 -2501 11013
rect 4819 11137 4853 11171
rect 11368 11225 11402 11259
rect 37358 11406 37392 11440
rect 37742 11394 37797 11452
rect 11250 11108 11284 11142
rect 4701 11020 4735 11054
rect -3237 10667 -3203 10701
rect -2467 10689 -2433 10723
rect 1907 10469 1941 10503
rect 4348 10510 4382 10544
rect 4466 10510 4500 10544
rect 1789 10352 1823 10386
rect -3045 9993 -3011 10027
rect 1436 9842 1470 9876
rect 1554 9842 1588 9876
rect -2470 9744 -2436 9778
rect 6980 10342 7014 10376
rect 5973 9699 6007 9733
rect 5788 9632 5822 9666
rect -2537 9559 -2503 9593
rect 6621 9699 6655 9733
rect 6239 9615 6273 9649
rect 6357 9616 6391 9650
rect 6911 9631 6945 9665
rect 10897 10598 10931 10632
rect 11015 10598 11049 10632
rect 18022 11157 18056 11191
rect 17904 11040 17938 11074
rect 24647 11225 24681 11259
rect 24529 11108 24563 11142
rect 37457 11276 37512 11334
rect 38577 11229 38611 11263
rect 37978 11171 38012 11205
rect 9087 10321 9121 10355
rect 7601 9826 7635 9860
rect 7871 9699 7905 9733
rect 7686 9632 7720 9666
rect 8517 9700 8551 9734
rect 8137 9615 8171 9649
rect 8255 9616 8289 9650
rect 13529 10430 13563 10464
rect 12522 9787 12556 9821
rect 12337 9720 12371 9754
rect 8809 9631 8843 9665
rect 4814 9533 4848 9567
rect 4696 9416 4730 9450
rect -2453 9293 -2419 9327
rect -2454 9175 -2420 9209
rect 13170 9787 13204 9821
rect 12788 9703 12822 9737
rect 12906 9704 12940 9738
rect 13460 9719 13494 9753
rect 17551 10530 17585 10564
rect 17669 10530 17703 10564
rect 15636 10409 15670 10443
rect 14150 9914 14184 9948
rect 14420 9787 14454 9821
rect 14235 9720 14269 9754
rect 15066 9788 15100 9822
rect 14686 9703 14720 9737
rect 14804 9704 14838 9738
rect 15358 9719 15392 9753
rect 11363 9621 11397 9655
rect 11245 9504 11279 9538
rect 20183 10362 20217 10396
rect 19176 9719 19210 9753
rect 18991 9652 19025 9686
rect 19824 9719 19858 9753
rect 19442 9635 19476 9669
rect 19560 9636 19594 9670
rect 20114 9651 20148 9685
rect 24176 10598 24210 10632
rect 24294 10598 24328 10632
rect 37588 11052 37622 11086
rect 22290 10341 22324 10375
rect 20804 9846 20838 9880
rect 21074 9719 21108 9753
rect 20889 9652 20923 9686
rect 21720 9720 21754 9754
rect 21340 9635 21374 9669
rect 21458 9636 21492 9670
rect 26808 10430 26842 10464
rect 25801 9787 25835 9821
rect 25616 9720 25650 9754
rect 22012 9651 22046 9685
rect 18017 9553 18051 9587
rect 17899 9436 17933 9470
rect -2537 8911 -2503 8945
rect 4343 8906 4377 8940
rect 4461 8906 4495 8940
rect 10892 8994 10926 9028
rect 11010 8994 11044 9028
rect 26449 9787 26483 9821
rect 26067 9703 26101 9737
rect 26185 9704 26219 9738
rect 26739 9719 26773 9753
rect 28915 10409 28949 10443
rect 27429 9914 27463 9948
rect 27699 9787 27733 9821
rect 27514 9720 27548 9754
rect 28345 9788 28379 9822
rect 27965 9703 27999 9737
rect 28083 9704 28117 9738
rect 28637 9719 28671 9753
rect 33130 10189 33164 10223
rect 31730 10070 31764 10104
rect 24642 9621 24676 9655
rect 24524 9504 24558 9538
rect 31935 9490 31969 9524
rect 31750 9423 31784 9457
rect 32583 9490 32617 9524
rect 32201 9406 32235 9440
rect 32319 9407 32353 9441
rect 34038 10308 34072 10342
rect 33920 10191 33954 10225
rect 37317 10096 37351 10130
rect 33567 9681 33601 9715
rect 33685 9681 33719 9715
rect 32873 9422 32907 9456
rect 17546 8926 17580 8960
rect 17664 8926 17698 8960
rect 24171 8994 24205 9028
rect 24289 8994 24323 9028
rect 30430 9203 30464 9237
rect 30312 9086 30346 9120
rect -3239 8599 -3205 8633
rect -2469 8621 -2435 8655
rect 37458 9219 37513 9277
rect 29959 8576 29993 8610
rect 30077 8576 30111 8610
rect 37358 8262 37392 8296
rect 37742 8250 37797 8308
rect 37457 8132 37512 8190
rect -3045 7924 -3011 7958
rect 38577 8085 38611 8119
rect 37978 8027 38012 8061
rect 37588 7908 37622 7942
rect -2470 7675 -2436 7709
rect -2537 7490 -2503 7524
rect 6240 7491 6274 7525
rect 7370 7497 7404 7531
rect -2453 7224 -2419 7258
rect 12791 7489 12825 7523
rect 13921 7495 13955 7529
rect 6240 7373 6274 7407
rect 7370 7377 7404 7411
rect 19446 7490 19480 7524
rect 20576 7496 20610 7530
rect 12791 7371 12825 7405
rect -2454 7106 -2420 7140
rect 1888 7191 1922 7225
rect 1770 7074 1804 7108
rect -2537 6842 -2503 6876
rect 4797 7007 4831 7041
rect 13921 7375 13955 7409
rect 26068 7491 26102 7525
rect 27198 7497 27232 7531
rect 19446 7372 19480 7406
rect 4679 6890 4713 6924
rect -3239 6530 -3205 6564
rect -2469 6552 -2435 6586
rect 1417 6564 1451 6598
rect 1535 6564 1569 6598
rect 6560 6617 6594 6651
rect 11348 7005 11382 7039
rect 20576 7376 20610 7410
rect 26068 7373 26102 7407
rect 11230 6888 11264 6922
rect 7702 6621 7736 6655
rect 4326 6380 4360 6414
rect 4444 6380 4478 6414
rect 13111 6615 13145 6649
rect 18003 7006 18037 7040
rect 27198 7377 27232 7411
rect 17885 6889 17919 6923
rect 14253 6619 14287 6653
rect 10877 6378 10911 6412
rect 10995 6378 11029 6412
rect 19766 6616 19800 6650
rect 24625 7007 24659 7041
rect 30501 7283 30535 7317
rect 30383 7166 30417 7200
rect 24507 6890 24541 6924
rect 20908 6620 20942 6654
rect 17532 6379 17566 6413
rect 17650 6379 17684 6413
rect 26388 6617 26422 6651
rect 27530 6621 27564 6655
rect 30030 6656 30064 6690
rect 30148 6656 30182 6690
rect 37317 6952 37351 6986
rect 33130 6694 33164 6728
rect 24154 6380 24188 6414
rect 24272 6380 24306 6414
rect 31730 6575 31764 6609
rect -3047 5856 -3013 5890
rect 31935 5995 31969 6029
rect 31750 5928 31784 5962
rect 32583 5995 32617 6029
rect 32201 5911 32235 5945
rect 32319 5912 32353 5946
rect 34038 6813 34072 6847
rect 33920 6696 33954 6730
rect 33567 6186 33601 6220
rect 33685 6186 33719 6220
rect 37454 6087 37509 6145
rect 32873 5927 32907 5961
rect -2472 5607 -2438 5641
rect -2539 5422 -2505 5456
rect -2455 5156 -2421 5190
rect 4811 5357 4845 5391
rect 4693 5240 4727 5274
rect -2456 5038 -2422 5072
rect -2539 4774 -2505 4808
rect 4340 4730 4374 4764
rect 4458 4730 4492 4764
rect 11362 5355 11396 5389
rect 11244 5238 11278 5272
rect -3241 4462 -3207 4496
rect -2471 4484 -2437 4518
rect 1904 4431 1938 4465
rect 1786 4314 1820 4348
rect -3045 3787 -3011 3821
rect 1433 3804 1467 3838
rect 1551 3804 1585 3838
rect 6972 4562 7006 4596
rect 5965 3919 5999 3953
rect 5780 3852 5814 3886
rect -2470 3538 -2436 3572
rect 6613 3919 6647 3953
rect 6231 3835 6265 3869
rect 6349 3836 6383 3870
rect 6903 3851 6937 3885
rect 10891 4728 10925 4762
rect 11009 4728 11043 4762
rect 18017 5356 18051 5390
rect 17899 5239 17933 5273
rect 9079 4541 9113 4575
rect 7593 4046 7627 4080
rect 7863 3919 7897 3953
rect 7678 3852 7712 3886
rect 8509 3920 8543 3954
rect 8129 3835 8163 3869
rect 8247 3836 8281 3870
rect 8801 3851 8835 3885
rect 13523 4560 13557 4594
rect 12516 3917 12550 3951
rect 12331 3850 12365 3884
rect 4806 3753 4840 3787
rect 4688 3636 4722 3670
rect -2537 3353 -2503 3387
rect 13164 3917 13198 3951
rect 12782 3833 12816 3867
rect 12900 3834 12934 3868
rect 13454 3849 13488 3883
rect 17546 4729 17580 4763
rect 17664 4729 17698 4763
rect 24639 5357 24673 5391
rect 24521 5240 24555 5274
rect 15630 4539 15664 4573
rect 14144 4044 14178 4078
rect 14414 3917 14448 3951
rect 14229 3850 14263 3884
rect 15060 3918 15094 3952
rect 14680 3833 14714 3867
rect 14798 3834 14832 3868
rect 15352 3849 15386 3883
rect 20178 4561 20212 4595
rect 19171 3918 19205 3952
rect 18986 3851 19020 3885
rect 11357 3751 11391 3785
rect 11239 3634 11273 3668
rect -2453 3087 -2419 3121
rect 4335 3126 4369 3160
rect 4453 3126 4487 3160
rect 19819 3918 19853 3952
rect 19437 3834 19471 3868
rect 19555 3835 19589 3869
rect 20109 3850 20143 3884
rect 24168 4730 24202 4764
rect 24286 4730 24320 4764
rect 37354 5130 37388 5164
rect 37738 5118 37793 5176
rect 37453 5000 37508 5058
rect 22285 4540 22319 4574
rect 20799 4045 20833 4079
rect 21069 3918 21103 3952
rect 20884 3851 20918 3885
rect 21715 3919 21749 3953
rect 21335 3834 21369 3868
rect 21453 3835 21487 3869
rect 22007 3850 22041 3884
rect 26800 4562 26834 4596
rect 25793 3919 25827 3953
rect 25608 3852 25642 3886
rect 18012 3752 18046 3786
rect 17894 3635 17928 3669
rect -2454 2969 -2420 3003
rect 10886 3124 10920 3158
rect 11004 3124 11038 3158
rect 26441 3919 26475 3953
rect 26059 3835 26093 3869
rect 26177 3836 26211 3870
rect 26731 3851 26765 3885
rect 38573 4953 38607 4987
rect 37974 4895 38008 4929
rect 37584 4776 37618 4810
rect 28907 4541 28941 4575
rect 27421 4046 27455 4080
rect 27691 3919 27725 3953
rect 27506 3852 27540 3886
rect 28337 3920 28371 3954
rect 27957 3835 27991 3869
rect 28075 3836 28109 3870
rect 30498 4213 30532 4247
rect 30380 4096 30414 4130
rect 28629 3851 28663 3885
rect 24634 3753 24668 3787
rect 24516 3636 24550 3670
rect 17541 3125 17575 3159
rect 17659 3125 17693 3159
rect 37313 3820 37347 3854
rect 30027 3586 30061 3620
rect 30145 3586 30179 3620
rect 24163 3126 24197 3160
rect 24281 3126 24315 3160
rect -2537 2705 -2503 2739
rect 37454 2943 37509 3001
rect -3239 2393 -3205 2427
rect -2469 2415 -2435 2449
rect 33130 2346 33164 2380
rect 8143 2207 8177 2241
rect 8261 2207 8295 2241
rect 14697 2212 14731 2246
rect 14815 2212 14849 2246
rect 21346 2200 21380 2234
rect 21464 2200 21498 2234
rect 31730 2227 31764 2261
rect -3047 1719 -3013 1753
rect 8496 1697 8530 1731
rect 8614 1580 8648 1614
rect -2472 1470 -2438 1504
rect 15050 1702 15084 1736
rect 15168 1585 15202 1619
rect 21699 1690 21733 1724
rect 21817 1573 21851 1607
rect -2539 1285 -2505 1319
rect 31935 1647 31969 1681
rect 31750 1580 31784 1614
rect 32583 1647 32617 1681
rect 32201 1563 32235 1597
rect 32319 1564 32353 1598
rect 34038 2465 34072 2499
rect 33920 2348 33954 2382
rect 37354 1986 37388 2020
rect 37738 1974 37793 2032
rect 33567 1838 33601 1872
rect 33685 1838 33719 1872
rect 37453 1856 37508 1914
rect 38573 1809 38607 1843
rect 37974 1751 38008 1785
rect 32873 1579 32907 1613
rect 37584 1632 37618 1666
rect 30505 1368 30539 1402
rect 30387 1251 30421 1285
rect -2455 1019 -2421 1053
rect -2456 901 -2422 935
rect 30034 741 30068 775
rect 30152 741 30186 775
rect -2539 637 -2505 671
rect 37313 676 37347 710
rect -3241 325 -3207 359
rect -2471 347 -2437 381
<< locali >>
rect 6237 28022 6460 28098
rect 6237 27873 6316 28022
rect 6383 27873 6460 28022
rect 6237 27767 6460 27873
rect 8719 28076 8942 28152
rect 8719 27927 8798 28076
rect 8865 27927 8942 28076
rect 8052 27856 8086 27872
rect 8052 27806 8086 27822
rect 8719 27821 8942 27927
rect 9866 28076 10089 28152
rect 9866 27927 9945 28076
rect 10012 27927 10089 28076
rect 9182 27862 9216 27878
rect 9182 27812 9216 27828
rect 9866 27821 10089 27927
rect 12750 28019 12973 28095
rect 12750 27870 12829 28019
rect 12896 27870 12973 28019
rect 12750 27764 12973 27870
rect 15232 28073 15455 28149
rect 15232 27924 15311 28073
rect 15378 27924 15455 28073
rect 14565 27853 14599 27869
rect 14565 27803 14599 27819
rect 15232 27818 15455 27924
rect 16379 28073 16602 28149
rect 16379 27924 16458 28073
rect 16525 27924 16602 28073
rect 15695 27859 15729 27875
rect 15695 27809 15729 27825
rect 16379 27818 16602 27924
rect 19284 28014 19507 28090
rect 19284 27865 19363 28014
rect 19430 27865 19507 28014
rect 19284 27759 19507 27865
rect 21766 28068 21989 28144
rect 21766 27919 21845 28068
rect 21912 27919 21989 28068
rect 21099 27848 21133 27864
rect 21099 27798 21133 27814
rect 21766 27813 21989 27919
rect 22913 28068 23136 28144
rect 22913 27919 22992 28068
rect 23059 27919 23136 28068
rect 22229 27854 22263 27870
rect 22229 27804 22263 27820
rect 22913 27813 23136 27919
rect 25842 28018 26065 28094
rect 25842 27869 25921 28018
rect 25988 27869 26065 28018
rect 25842 27763 26065 27869
rect 28324 28072 28547 28148
rect 28324 27923 28403 28072
rect 28470 27923 28547 28072
rect 27657 27852 27691 27868
rect 27657 27802 27691 27818
rect 28324 27817 28547 27923
rect 29471 28072 29694 28148
rect 29471 27923 29550 28072
rect 29617 27923 29694 28072
rect 28787 27858 28821 27874
rect 28787 27808 28821 27824
rect 29471 27817 29694 27923
rect 8052 27738 8086 27754
rect 6668 27658 6938 27692
rect 8052 27688 8086 27704
rect 9182 27742 9216 27758
rect 5842 27608 5876 27624
rect 5842 27416 5876 27432
rect 5960 27608 5994 27624
rect 5960 27416 5994 27432
rect 6078 27608 6112 27624
rect 6078 27416 6112 27432
rect 6196 27608 6230 27624
rect 6196 27416 6230 27432
rect 6314 27608 6348 27624
rect 6314 27416 6348 27432
rect 6432 27608 6466 27624
rect 6432 27416 6466 27432
rect 6550 27608 6584 27624
rect 6550 27416 6584 27432
rect 6668 27608 6702 27658
rect 6668 27416 6702 27432
rect 6786 27608 6820 27624
rect 6786 27416 6820 27432
rect 6904 27608 6938 27658
rect 6904 27416 6938 27432
rect 8167 27680 8201 27696
rect 6593 27338 6609 27372
rect 6643 27338 6659 27372
rect 8167 27288 8201 27304
rect 8285 27680 8319 27696
rect 8285 27288 8319 27304
rect 8403 27680 8437 27696
rect 8403 27288 8437 27304
rect 8521 27680 8555 27696
rect 8521 27288 8555 27304
rect 8639 27680 8673 27696
rect 8639 27288 8673 27304
rect 8757 27680 8791 27696
rect 8757 27288 8791 27304
rect 8875 27680 8909 27696
rect 9182 27692 9216 27708
rect 14565 27735 14599 27751
rect 8875 27288 8909 27304
rect 9309 27684 9343 27700
rect 9309 27292 9343 27308
rect 9427 27684 9461 27700
rect 9427 27292 9461 27308
rect 9545 27684 9579 27700
rect 9545 27292 9579 27308
rect 9663 27684 9697 27700
rect 9663 27292 9697 27308
rect 9781 27684 9815 27700
rect 9781 27292 9815 27308
rect 9899 27684 9933 27700
rect 9899 27292 9933 27308
rect 10017 27684 10051 27700
rect 13181 27655 13451 27689
rect 14565 27685 14599 27701
rect 15695 27739 15729 27755
rect 12355 27605 12389 27621
rect 12355 27413 12389 27429
rect 12473 27605 12507 27621
rect 12473 27413 12507 27429
rect 12591 27605 12625 27621
rect 12591 27413 12625 27429
rect 12709 27605 12743 27621
rect 12709 27413 12743 27429
rect 12827 27605 12861 27621
rect 12827 27413 12861 27429
rect 12945 27605 12979 27621
rect 12945 27413 12979 27429
rect 13063 27605 13097 27621
rect 13063 27413 13097 27429
rect 13181 27605 13215 27655
rect 13181 27413 13215 27429
rect 13299 27605 13333 27621
rect 13299 27413 13333 27429
rect 13417 27605 13451 27655
rect 13417 27413 13451 27429
rect 14680 27677 14714 27693
rect 13106 27335 13122 27369
rect 13156 27335 13172 27369
rect 10017 27292 10051 27308
rect 14680 27285 14714 27301
rect 14798 27677 14832 27693
rect 14798 27285 14832 27301
rect 14916 27677 14950 27693
rect 14916 27285 14950 27301
rect 15034 27677 15068 27693
rect 15034 27285 15068 27301
rect 15152 27677 15186 27693
rect 15152 27285 15186 27301
rect 15270 27677 15304 27693
rect 15270 27285 15304 27301
rect 15388 27677 15422 27693
rect 15695 27689 15729 27705
rect 21099 27730 21133 27746
rect 15388 27285 15422 27301
rect 15822 27681 15856 27697
rect 15822 27289 15856 27305
rect 15940 27681 15974 27697
rect 15940 27289 15974 27305
rect 16058 27681 16092 27697
rect 16058 27289 16092 27305
rect 16176 27681 16210 27697
rect 16176 27289 16210 27305
rect 16294 27681 16328 27697
rect 16294 27289 16328 27305
rect 16412 27681 16446 27697
rect 16412 27289 16446 27305
rect 16530 27681 16564 27697
rect 19715 27650 19985 27684
rect 21099 27680 21133 27696
rect 22229 27734 22263 27750
rect 18889 27600 18923 27616
rect 18889 27408 18923 27424
rect 19007 27600 19041 27616
rect 19007 27408 19041 27424
rect 19125 27600 19159 27616
rect 19125 27408 19159 27424
rect 19243 27600 19277 27616
rect 19243 27408 19277 27424
rect 19361 27600 19395 27616
rect 19361 27408 19395 27424
rect 19479 27600 19513 27616
rect 19479 27408 19513 27424
rect 19597 27600 19631 27616
rect 19597 27408 19631 27424
rect 19715 27600 19749 27650
rect 19715 27408 19749 27424
rect 19833 27600 19867 27616
rect 19833 27408 19867 27424
rect 19951 27600 19985 27650
rect 19951 27408 19985 27424
rect 21214 27672 21248 27688
rect 19640 27330 19656 27364
rect 19690 27330 19706 27364
rect 16530 27289 16564 27305
rect 21214 27280 21248 27296
rect 21332 27672 21366 27688
rect 21332 27280 21366 27296
rect 21450 27672 21484 27688
rect 21450 27280 21484 27296
rect 21568 27672 21602 27688
rect 21568 27280 21602 27296
rect 21686 27672 21720 27688
rect 21686 27280 21720 27296
rect 21804 27672 21838 27688
rect 21804 27280 21838 27296
rect 21922 27672 21956 27688
rect 22229 27684 22263 27700
rect 27657 27734 27691 27750
rect 21922 27280 21956 27296
rect 22356 27676 22390 27692
rect 22356 27284 22390 27300
rect 22474 27676 22508 27692
rect 22474 27284 22508 27300
rect 22592 27676 22626 27692
rect 22592 27284 22626 27300
rect 22710 27676 22744 27692
rect 22710 27284 22744 27300
rect 22828 27676 22862 27692
rect 22828 27284 22862 27300
rect 22946 27676 22980 27692
rect 22946 27284 22980 27300
rect 23064 27676 23098 27692
rect 26273 27654 26543 27688
rect 27657 27684 27691 27700
rect 28787 27738 28821 27754
rect 25447 27604 25481 27620
rect 25447 27412 25481 27428
rect 25565 27604 25599 27620
rect 25565 27412 25599 27428
rect 25683 27604 25717 27620
rect 25683 27412 25717 27428
rect 25801 27604 25835 27620
rect 25801 27412 25835 27428
rect 25919 27604 25953 27620
rect 25919 27412 25953 27428
rect 26037 27604 26071 27620
rect 26037 27412 26071 27428
rect 26155 27604 26189 27620
rect 26155 27412 26189 27428
rect 26273 27604 26307 27654
rect 26273 27412 26307 27428
rect 26391 27604 26425 27620
rect 26391 27412 26425 27428
rect 26509 27604 26543 27654
rect 26509 27412 26543 27428
rect 27772 27676 27806 27692
rect 26198 27334 26214 27368
rect 26248 27334 26264 27368
rect 23064 27284 23098 27300
rect 27772 27284 27806 27300
rect 27890 27676 27924 27692
rect 27890 27284 27924 27300
rect 28008 27676 28042 27692
rect 28008 27284 28042 27300
rect 28126 27676 28160 27692
rect 28126 27284 28160 27300
rect 28244 27676 28278 27692
rect 28244 27284 28278 27300
rect 28362 27676 28396 27692
rect 28362 27284 28396 27300
rect 28480 27676 28514 27692
rect 28787 27688 28821 27704
rect 28480 27284 28514 27300
rect 28914 27680 28948 27696
rect 28914 27288 28948 27304
rect 29032 27680 29066 27696
rect 29032 27288 29066 27304
rect 29150 27680 29184 27696
rect 29150 27288 29184 27304
rect 29268 27680 29302 27696
rect 29268 27288 29302 27304
rect 29386 27680 29420 27696
rect 29386 27288 29420 27304
rect 29504 27680 29538 27696
rect 29504 27288 29538 27304
rect 29622 27680 29656 27696
rect 29622 27288 29656 27304
rect 6475 27221 6491 27255
rect 6525 27221 6541 27255
rect 12988 27218 13004 27252
rect 13038 27218 13054 27252
rect 19522 27213 19538 27247
rect 19572 27213 19588 27247
rect 26080 27217 26096 27251
rect 26130 27217 26146 27251
rect 6079 27171 6113 27187
rect 6079 26779 6113 26795
rect 6197 27171 6231 27187
rect 6197 26779 6231 26795
rect 6315 27171 6349 27187
rect 6432 27171 6466 27187
rect 6432 26979 6466 26995
rect 6550 27171 6584 27187
rect 6550 26979 6584 26995
rect 12592 27168 12626 27184
rect 8356 26948 8372 26982
rect 8406 26948 8422 26982
rect 9498 26952 9514 26986
rect 9548 26952 9564 26986
rect 8077 26897 8111 26913
rect 6315 26779 6349 26795
rect 6602 26845 6851 26888
rect 6602 26755 6649 26845
rect 6812 26755 6851 26845
rect 6122 26711 6138 26745
rect 6172 26711 6188 26745
rect 6240 26711 6256 26745
rect 6290 26711 6306 26745
rect 6602 26716 6851 26755
rect 8077 26705 8111 26721
rect 8195 26897 8229 26913
rect 8195 26705 8229 26721
rect 8313 26897 8347 26913
rect 8313 26705 8347 26721
rect 8431 26897 8465 26913
rect 8431 26705 8465 26721
rect 8596 26897 8630 26913
rect 8596 26705 8630 26721
rect 8714 26897 8748 26913
rect 8714 26705 8748 26721
rect 8832 26897 8866 26913
rect 8832 26705 8866 26721
rect 8950 26897 8984 26913
rect 8950 26705 8984 26721
rect 9219 26901 9253 26917
rect 9219 26709 9253 26725
rect 9337 26901 9371 26917
rect 9337 26709 9371 26725
rect 9455 26901 9489 26917
rect 9455 26709 9489 26725
rect 9573 26901 9607 26917
rect 9573 26709 9607 26725
rect 9738 26901 9772 26917
rect 9738 26709 9772 26725
rect 9856 26901 9890 26917
rect 9856 26709 9890 26725
rect 9974 26901 10008 26917
rect 9974 26709 10008 26725
rect 10092 26901 10126 26917
rect 12592 26776 12626 26792
rect 12710 27168 12744 27184
rect 12710 26776 12744 26792
rect 12828 27168 12862 27184
rect 12945 27168 12979 27184
rect 12945 26976 12979 26992
rect 13063 27168 13097 27184
rect 13063 26976 13097 26992
rect 19126 27163 19160 27179
rect 14869 26945 14885 26979
rect 14919 26945 14935 26979
rect 16011 26949 16027 26983
rect 16061 26949 16077 26983
rect 14590 26894 14624 26910
rect 12828 26776 12862 26792
rect 13115 26842 13364 26885
rect 13115 26752 13162 26842
rect 13325 26752 13364 26842
rect 10092 26709 10126 26725
rect 12635 26708 12651 26742
rect 12685 26708 12701 26742
rect 12753 26708 12769 26742
rect 12803 26708 12819 26742
rect 13115 26713 13364 26752
rect 14590 26702 14624 26718
rect 14708 26894 14742 26910
rect 14708 26702 14742 26718
rect 14826 26894 14860 26910
rect 14826 26702 14860 26718
rect 14944 26894 14978 26910
rect 14944 26702 14978 26718
rect 15109 26894 15143 26910
rect 15109 26702 15143 26718
rect 15227 26894 15261 26910
rect 15227 26702 15261 26718
rect 15345 26894 15379 26910
rect 15345 26702 15379 26718
rect 15463 26894 15497 26910
rect 15463 26702 15497 26718
rect 15732 26898 15766 26914
rect 15732 26706 15766 26722
rect 15850 26898 15884 26914
rect 15850 26706 15884 26722
rect 15968 26898 16002 26914
rect 15968 26706 16002 26722
rect 16086 26898 16120 26914
rect 16086 26706 16120 26722
rect 16251 26898 16285 26914
rect 16251 26706 16285 26722
rect 16369 26898 16403 26914
rect 16369 26706 16403 26722
rect 16487 26898 16521 26914
rect 16487 26706 16521 26722
rect 16605 26898 16639 26914
rect 19126 26771 19160 26787
rect 19244 27163 19278 27179
rect 19244 26771 19278 26787
rect 19362 27163 19396 27179
rect 19479 27163 19513 27179
rect 19479 26971 19513 26987
rect 19597 27163 19631 27179
rect 19597 26971 19631 26987
rect 25684 27167 25718 27183
rect 21403 26940 21419 26974
rect 21453 26940 21469 26974
rect 22545 26944 22561 26978
rect 22595 26944 22611 26978
rect 21124 26889 21158 26905
rect 19362 26771 19396 26787
rect 19649 26837 19898 26880
rect 19649 26747 19696 26837
rect 19859 26747 19898 26837
rect 16605 26706 16639 26722
rect 19169 26703 19185 26737
rect 19219 26703 19235 26737
rect 19287 26703 19303 26737
rect 19337 26703 19353 26737
rect 19649 26708 19898 26747
rect 21124 26697 21158 26713
rect 21242 26889 21276 26905
rect 21242 26697 21276 26713
rect 21360 26889 21394 26905
rect 21360 26697 21394 26713
rect 21478 26889 21512 26905
rect 21478 26697 21512 26713
rect 21643 26889 21677 26905
rect 21643 26697 21677 26713
rect 21761 26889 21795 26905
rect 21761 26697 21795 26713
rect 21879 26889 21913 26905
rect 21879 26697 21913 26713
rect 21997 26889 22031 26905
rect 21997 26697 22031 26713
rect 22266 26893 22300 26909
rect 22266 26701 22300 26717
rect 22384 26893 22418 26909
rect 22384 26701 22418 26717
rect 22502 26893 22536 26909
rect 22502 26701 22536 26717
rect 22620 26893 22654 26909
rect 22620 26701 22654 26717
rect 22785 26893 22819 26909
rect 22785 26701 22819 26717
rect 22903 26893 22937 26909
rect 22903 26701 22937 26717
rect 23021 26893 23055 26909
rect 23021 26701 23055 26717
rect 23139 26893 23173 26909
rect 25684 26775 25718 26791
rect 25802 27167 25836 27183
rect 25802 26775 25836 26791
rect 25920 27167 25954 27183
rect 26037 27167 26071 27183
rect 26037 26975 26071 26991
rect 26155 27167 26189 27183
rect 26155 26975 26189 26991
rect 27961 26944 27977 26978
rect 28011 26944 28027 26978
rect 29103 26948 29119 26982
rect 29153 26948 29169 26982
rect 27682 26893 27716 26909
rect 25920 26775 25954 26791
rect 26207 26841 26456 26884
rect 26207 26751 26254 26841
rect 26417 26751 26456 26841
rect 23139 26701 23173 26717
rect 25727 26707 25743 26741
rect 25777 26707 25793 26741
rect 25845 26707 25861 26741
rect 25895 26707 25911 26741
rect 26207 26712 26456 26751
rect 27682 26701 27716 26717
rect 27800 26893 27834 26909
rect 27800 26701 27834 26717
rect 27918 26893 27952 26909
rect 27918 26701 27952 26717
rect 28036 26893 28070 26909
rect 28036 26701 28070 26717
rect 28201 26893 28235 26909
rect 28201 26701 28235 26717
rect 28319 26893 28353 26909
rect 28319 26701 28353 26717
rect 28437 26893 28471 26909
rect 28437 26701 28471 26717
rect 28555 26893 28589 26909
rect 28555 26701 28589 26717
rect 28824 26897 28858 26913
rect 28824 26705 28858 26721
rect 28942 26897 28976 26913
rect 28942 26705 28976 26721
rect 29060 26897 29094 26913
rect 29060 26705 29094 26721
rect 29178 26897 29212 26913
rect 29178 26705 29212 26721
rect 29343 26897 29377 26913
rect 29343 26705 29377 26721
rect 29461 26897 29495 26913
rect 29461 26705 29495 26721
rect 29579 26897 29613 26913
rect 29579 26705 29613 26721
rect 29697 26897 29731 26913
rect 29697 26705 29731 26721
rect 8092 26474 8264 26521
rect 6251 26372 6474 26448
rect 6251 26223 6330 26372
rect 6397 26223 6474 26372
rect 8092 26311 8131 26474
rect 8221 26311 8264 26474
rect 8092 26272 8264 26311
rect 9234 26472 9406 26519
rect 9234 26309 9273 26472
rect 9363 26309 9406 26472
rect 14605 26471 14777 26518
rect 9234 26270 9406 26309
rect 12764 26369 12987 26445
rect 6251 26117 6474 26223
rect 12764 26220 12843 26369
rect 12910 26220 12987 26369
rect 14605 26308 14644 26471
rect 14734 26308 14777 26471
rect 14605 26269 14777 26308
rect 15747 26469 15919 26516
rect 15747 26306 15786 26469
rect 15876 26306 15919 26469
rect 21139 26466 21311 26513
rect 15747 26267 15919 26306
rect 19298 26364 19521 26440
rect 12764 26114 12987 26220
rect 19298 26215 19377 26364
rect 19444 26215 19521 26364
rect 21139 26303 21178 26466
rect 21268 26303 21311 26466
rect 21139 26264 21311 26303
rect 22281 26464 22453 26511
rect 22281 26301 22320 26464
rect 22410 26301 22453 26464
rect 27697 26470 27869 26517
rect 22281 26262 22453 26301
rect 25856 26368 26079 26444
rect 19298 26109 19521 26215
rect 25856 26219 25935 26368
rect 26002 26219 26079 26368
rect 27697 26307 27736 26470
rect 27826 26307 27869 26470
rect 27697 26268 27869 26307
rect 28839 26468 29011 26515
rect 28839 26305 28878 26468
rect 28968 26305 29011 26468
rect 28839 26266 29011 26305
rect 25856 26113 26079 26219
rect 6682 26008 6952 26042
rect 5856 25958 5890 25974
rect 54 25939 125 25946
rect 54 25890 64 25939
rect 118 25890 125 25939
rect -100 25518 -15 25527
rect -100 25447 -92 25518
rect -23 25447 -15 25518
rect -247 25094 -157 25103
rect -247 25023 -239 25094
rect -168 25023 -157 25094
rect -394 24634 -300 24647
rect -394 24573 -382 24634
rect -311 24573 -300 24634
rect -3681 16221 -3592 16255
rect -3416 16221 -3400 16255
rect -3681 16019 -3646 16221
rect -3608 16103 -3592 16137
rect -3416 16103 -3400 16137
rect -2383 16096 -2367 16130
rect -2191 16096 -2175 16130
rect -3681 15985 -3592 16019
rect -3416 15985 -3400 16019
rect -2484 15949 -2468 15983
rect -2434 15949 -2418 15983
rect -2383 15978 -2367 16012
rect -2191 15978 -2175 16012
rect -3608 15867 -3592 15901
rect -3416 15867 -3400 15901
rect -3115 15794 -3099 15828
rect -2723 15794 -2707 15828
rect -2551 15798 -2485 15814
rect -3808 15737 -3792 15771
rect -3416 15737 -3400 15771
rect -2551 15764 -2535 15798
rect -2501 15764 -2485 15798
rect -2551 15747 -2485 15764
rect -2770 15710 -2625 15711
rect -3115 15676 -3099 15710
rect -2723 15692 -2625 15710
rect -2723 15676 -2624 15692
rect -2383 15676 -2367 15710
rect -2770 15675 -2624 15676
rect -1991 15675 -1889 15710
rect -3808 15619 -3792 15653
rect -3416 15619 -3400 15653
rect -2665 15637 -2624 15675
rect -2665 15603 -2337 15637
rect -3115 15558 -3099 15592
rect -2723 15558 -2707 15592
rect -4083 15470 -3991 15504
rect -3808 15501 -3792 15535
rect -3416 15501 -3400 15535
rect -2665 15476 -2624 15603
rect -2383 15592 -2337 15603
rect -2383 15558 -2367 15592
rect -1991 15558 -1975 15592
rect -2451 15532 -2417 15548
rect -2451 15482 -2417 15498
rect -2770 15474 -2624 15476
rect -4083 15348 -4063 15470
rect -4019 15418 -3991 15470
rect -3115 15440 -3099 15474
rect -2723 15440 -2624 15474
rect -2383 15440 -2367 15474
rect -1991 15440 -1975 15474
rect -4009 15380 -3991 15418
rect -4019 15348 -3991 15380
rect -4083 15302 -3991 15348
rect -3880 15383 -3792 15417
rect -3416 15383 -3400 15417
rect -3880 15181 -3845 15383
rect -3115 15322 -3099 15356
rect -2723 15322 -2707 15356
rect -3808 15265 -3792 15299
rect -3416 15265 -3400 15299
rect -2665 15238 -2624 15440
rect -2452 15414 -2418 15430
rect -2452 15364 -2418 15380
rect -2383 15322 -2367 15356
rect -1991 15322 -1975 15356
rect -1924 15239 -1889 15675
rect -1819 15520 -1731 15536
rect -1819 15480 -1803 15520
rect -1819 15388 -1803 15430
rect -1747 15388 -1731 15520
rect -1819 15372 -1731 15388
rect -3115 15204 -3099 15238
rect -2723 15204 -2624 15238
rect -2383 15204 -2367 15238
rect -1991 15204 -1889 15239
rect -2769 15202 -2624 15204
rect -3880 15147 -3792 15181
rect -3416 15147 -3400 15181
rect -3115 15086 -3099 15120
rect -2723 15086 -2707 15120
rect -3808 15029 -3792 15063
rect -3416 15029 -3400 15063
rect -3608 14900 -3592 14934
rect -3416 14900 -3400 14934
rect -3237 14848 -3203 14854
rect -3608 14782 -3592 14816
rect -3416 14782 -3400 14816
rect -3237 14788 -3203 14794
rect -3608 14664 -3592 14698
rect -3416 14664 -3400 14698
rect -2665 14616 -2624 15202
rect -2551 15150 -2485 15167
rect -2551 15116 -2535 15150
rect -2501 15116 -2485 15150
rect -2551 15100 -2485 15116
rect -2483 14826 -2467 14860
rect -2433 14826 -2417 14860
rect -2383 14798 -2367 14832
rect -2191 14798 -2175 14832
rect -2383 14680 -2367 14714
rect -2191 14680 -2175 14714
rect -3608 14546 -3592 14580
rect -3416 14546 -3400 14580
rect -3683 14153 -3594 14187
rect -3418 14153 -3402 14187
rect -3683 13951 -3648 14153
rect -3610 14035 -3594 14069
rect -3418 14035 -3402 14069
rect -2385 14028 -2369 14062
rect -2193 14028 -2177 14062
rect -3683 13917 -3594 13951
rect -3418 13917 -3402 13951
rect -2486 13881 -2470 13915
rect -2436 13881 -2420 13915
rect -2385 13910 -2369 13944
rect -2193 13910 -2177 13944
rect -3610 13799 -3594 13833
rect -3418 13799 -3402 13833
rect -3117 13726 -3101 13760
rect -2725 13726 -2709 13760
rect -2553 13730 -2487 13746
rect -3810 13669 -3794 13703
rect -3418 13669 -3402 13703
rect -2553 13696 -2537 13730
rect -2503 13696 -2487 13730
rect -2553 13679 -2487 13696
rect -2772 13642 -2627 13643
rect -3117 13608 -3101 13642
rect -2725 13624 -2627 13642
rect -2725 13608 -2626 13624
rect -2385 13608 -2369 13642
rect -2772 13607 -2626 13608
rect -1993 13607 -1891 13642
rect -3810 13551 -3794 13585
rect -3418 13551 -3402 13585
rect -2667 13569 -2626 13607
rect -2667 13535 -2339 13569
rect -3117 13490 -3101 13524
rect -2725 13490 -2709 13524
rect -4085 13402 -3993 13436
rect -3810 13433 -3794 13467
rect -3418 13433 -3402 13467
rect -2667 13408 -2626 13535
rect -2385 13524 -2339 13535
rect -2385 13490 -2369 13524
rect -1993 13490 -1977 13524
rect -2453 13464 -2419 13480
rect -2453 13414 -2419 13430
rect -2772 13406 -2626 13408
rect -4085 13280 -4065 13402
rect -4021 13350 -3993 13402
rect -3117 13372 -3101 13406
rect -2725 13372 -2626 13406
rect -2385 13372 -2369 13406
rect -1993 13372 -1977 13406
rect -4011 13312 -3993 13350
rect -4021 13280 -3993 13312
rect -4085 13234 -3993 13280
rect -3882 13315 -3794 13349
rect -3418 13315 -3402 13349
rect -3882 13113 -3847 13315
rect -3117 13254 -3101 13288
rect -2725 13254 -2709 13288
rect -3810 13197 -3794 13231
rect -3418 13197 -3402 13231
rect -2667 13170 -2626 13372
rect -2454 13346 -2420 13362
rect -2454 13296 -2420 13312
rect -2385 13254 -2369 13288
rect -1993 13254 -1977 13288
rect -1926 13171 -1891 13607
rect -1821 13452 -1733 13468
rect -1821 13412 -1805 13452
rect -1821 13320 -1805 13362
rect -1749 13320 -1733 13452
rect -1821 13304 -1733 13320
rect -3117 13136 -3101 13170
rect -2725 13136 -2626 13170
rect -2385 13136 -2369 13170
rect -1993 13136 -1891 13171
rect -2771 13134 -2626 13136
rect -3882 13079 -3794 13113
rect -3418 13079 -3402 13113
rect -3117 13018 -3101 13052
rect -2725 13018 -2709 13052
rect -3810 12961 -3794 12995
rect -3418 12961 -3402 12995
rect -3610 12832 -3594 12866
rect -3418 12832 -3402 12866
rect -3239 12780 -3205 12786
rect -3610 12714 -3594 12748
rect -3418 12714 -3402 12748
rect -3239 12720 -3205 12726
rect -3610 12596 -3594 12630
rect -3418 12596 -3402 12630
rect -2667 12548 -2626 13134
rect -2553 13082 -2487 13099
rect -2553 13048 -2537 13082
rect -2503 13048 -2487 13082
rect -2553 13032 -2487 13048
rect -2485 12758 -2469 12792
rect -2435 12758 -2419 12792
rect -2385 12730 -2369 12764
rect -2193 12730 -2177 12764
rect -2385 12612 -2369 12646
rect -2193 12612 -2177 12646
rect -3610 12478 -3594 12512
rect -3418 12478 -3402 12512
rect -3681 12084 -3592 12118
rect -3416 12084 -3400 12118
rect -3681 11882 -3646 12084
rect -3608 11966 -3592 12000
rect -3416 11966 -3400 12000
rect -2383 11959 -2367 11993
rect -2191 11959 -2175 11993
rect -3681 11848 -3592 11882
rect -3416 11848 -3400 11882
rect -2484 11812 -2468 11846
rect -2434 11812 -2418 11846
rect -2383 11841 -2367 11875
rect -2191 11841 -2175 11875
rect -3608 11730 -3592 11764
rect -3416 11730 -3400 11764
rect -3115 11657 -3099 11691
rect -2723 11657 -2707 11691
rect -2551 11661 -2485 11677
rect -3808 11600 -3792 11634
rect -3416 11600 -3400 11634
rect -2551 11627 -2535 11661
rect -2501 11627 -2485 11661
rect -2551 11610 -2485 11627
rect -2770 11573 -2625 11574
rect -3115 11539 -3099 11573
rect -2723 11555 -2625 11573
rect -2723 11539 -2624 11555
rect -2383 11539 -2367 11573
rect -2770 11538 -2624 11539
rect -1991 11538 -1889 11573
rect -3808 11482 -3792 11516
rect -3416 11482 -3400 11516
rect -2665 11500 -2624 11538
rect -2665 11466 -2337 11500
rect -3115 11421 -3099 11455
rect -2723 11421 -2707 11455
rect -4083 11333 -3991 11367
rect -3808 11364 -3792 11398
rect -3416 11364 -3400 11398
rect -2665 11339 -2624 11466
rect -2383 11455 -2337 11466
rect -2383 11421 -2367 11455
rect -1991 11421 -1975 11455
rect -2451 11395 -2417 11411
rect -2451 11345 -2417 11361
rect -2770 11337 -2624 11339
rect -4083 11211 -4063 11333
rect -4019 11281 -3991 11333
rect -3115 11303 -3099 11337
rect -2723 11303 -2624 11337
rect -2383 11303 -2367 11337
rect -1991 11303 -1975 11337
rect -4009 11243 -3991 11281
rect -4019 11211 -3991 11243
rect -4083 11165 -3991 11211
rect -3880 11246 -3792 11280
rect -3416 11246 -3400 11280
rect -3880 11044 -3845 11246
rect -3115 11185 -3099 11219
rect -2723 11185 -2707 11219
rect -3808 11128 -3792 11162
rect -3416 11128 -3400 11162
rect -2665 11101 -2624 11303
rect -2452 11277 -2418 11293
rect -2452 11227 -2418 11243
rect -2383 11185 -2367 11219
rect -1991 11185 -1975 11219
rect -1924 11102 -1889 11538
rect -1819 11383 -1731 11399
rect -1819 11343 -1803 11383
rect -1819 11251 -1803 11293
rect -1747 11251 -1731 11383
rect -1819 11235 -1731 11251
rect -3115 11067 -3099 11101
rect -2723 11067 -2624 11101
rect -2383 11067 -2367 11101
rect -1991 11067 -1889 11102
rect -2769 11065 -2624 11067
rect -3880 11010 -3792 11044
rect -3416 11010 -3400 11044
rect -3115 10949 -3099 10983
rect -2723 10949 -2707 10983
rect -3808 10892 -3792 10926
rect -3416 10892 -3400 10926
rect -3608 10763 -3592 10797
rect -3416 10763 -3400 10797
rect -3237 10711 -3203 10717
rect -3608 10645 -3592 10679
rect -3416 10645 -3400 10679
rect -3237 10651 -3203 10657
rect -3608 10527 -3592 10561
rect -3416 10527 -3400 10561
rect -2665 10479 -2624 11065
rect -2551 11013 -2485 11030
rect -2551 10979 -2535 11013
rect -2501 10979 -2485 11013
rect -2551 10963 -2485 10979
rect -2483 10689 -2467 10723
rect -2433 10689 -2417 10723
rect -2383 10661 -2367 10695
rect -2191 10661 -2175 10695
rect -2383 10543 -2367 10577
rect -2191 10543 -2175 10577
rect -3608 10409 -3592 10443
rect -3416 10409 -3400 10443
rect -3683 10016 -3594 10050
rect -3418 10016 -3402 10050
rect -394 10028 -300 24573
rect -247 12564 -157 25023
rect -3683 9814 -3648 10016
rect -3610 9898 -3594 9932
rect -3418 9898 -3402 9932
rect -2385 9891 -2369 9925
rect -2193 9891 -2177 9925
rect -3683 9780 -3594 9814
rect -3418 9780 -3402 9814
rect -2486 9744 -2470 9778
rect -2436 9744 -2420 9778
rect -2385 9773 -2369 9807
rect -2193 9773 -2177 9807
rect -3610 9662 -3594 9696
rect -3418 9662 -3402 9696
rect -3117 9589 -3101 9623
rect -2725 9589 -2709 9623
rect -2553 9593 -2487 9609
rect -3810 9532 -3794 9566
rect -3418 9532 -3402 9566
rect -2553 9559 -2537 9593
rect -2503 9559 -2487 9593
rect -2553 9542 -2487 9559
rect -2772 9505 -2627 9506
rect -3117 9471 -3101 9505
rect -2725 9487 -2627 9505
rect -2725 9471 -2626 9487
rect -2385 9471 -2369 9505
rect -2772 9470 -2626 9471
rect -1993 9470 -1891 9505
rect -3810 9414 -3794 9448
rect -3418 9414 -3402 9448
rect -2667 9432 -2626 9470
rect -2667 9398 -2339 9432
rect -3117 9353 -3101 9387
rect -2725 9353 -2709 9387
rect -4085 9265 -3993 9299
rect -3810 9296 -3794 9330
rect -3418 9296 -3402 9330
rect -2667 9271 -2626 9398
rect -2385 9387 -2339 9398
rect -2385 9353 -2369 9387
rect -1993 9353 -1977 9387
rect -2453 9327 -2419 9343
rect -2453 9277 -2419 9293
rect -2772 9269 -2626 9271
rect -4085 9143 -4065 9265
rect -4021 9213 -3993 9265
rect -3117 9235 -3101 9269
rect -2725 9235 -2626 9269
rect -2385 9235 -2369 9269
rect -1993 9235 -1977 9269
rect -4011 9175 -3993 9213
rect -4021 9143 -3993 9175
rect -4085 9097 -3993 9143
rect -3882 9178 -3794 9212
rect -3418 9178 -3402 9212
rect -3882 8976 -3847 9178
rect -3117 9117 -3101 9151
rect -2725 9117 -2709 9151
rect -3810 9060 -3794 9094
rect -3418 9060 -3402 9094
rect -2667 9033 -2626 9235
rect -2454 9209 -2420 9225
rect -2454 9159 -2420 9175
rect -2385 9117 -2369 9151
rect -1993 9117 -1977 9151
rect -1926 9034 -1891 9470
rect -1821 9315 -1733 9331
rect -1821 9275 -1805 9315
rect -1821 9183 -1805 9225
rect -1749 9183 -1733 9315
rect -1821 9167 -1733 9183
rect -3117 8999 -3101 9033
rect -2725 8999 -2626 9033
rect -2385 8999 -2369 9033
rect -1993 8999 -1891 9034
rect -2771 8997 -2626 8999
rect -3882 8942 -3794 8976
rect -3418 8942 -3402 8976
rect -3117 8881 -3101 8915
rect -2725 8881 -2709 8915
rect -3810 8824 -3794 8858
rect -3418 8824 -3402 8858
rect -3610 8695 -3594 8729
rect -3418 8695 -3402 8729
rect -3239 8643 -3205 8649
rect -3610 8577 -3594 8611
rect -3418 8577 -3402 8611
rect -3239 8583 -3205 8589
rect -3610 8459 -3594 8493
rect -3418 8459 -3402 8493
rect -2667 8411 -2626 8997
rect -2553 8945 -2487 8962
rect -2553 8911 -2537 8945
rect -2503 8911 -2487 8945
rect -2553 8895 -2487 8911
rect -2485 8621 -2469 8655
rect -2435 8621 -2419 8655
rect -2385 8593 -2369 8627
rect -2193 8593 -2177 8627
rect -2385 8475 -2369 8509
rect -2193 8475 -2177 8509
rect -3610 8341 -3594 8375
rect -3418 8341 -3402 8375
rect -3683 7947 -3594 7981
rect -3418 7947 -3402 7981
rect -3683 7745 -3648 7947
rect -3610 7829 -3594 7863
rect -3418 7829 -3402 7863
rect -2385 7822 -2369 7856
rect -2193 7822 -2177 7856
rect -3683 7711 -3594 7745
rect -3418 7711 -3402 7745
rect -2486 7675 -2470 7709
rect -2436 7675 -2420 7709
rect -2385 7704 -2369 7738
rect -2193 7704 -2177 7738
rect -3610 7593 -3594 7627
rect -3418 7593 -3402 7627
rect -3117 7520 -3101 7554
rect -2725 7520 -2709 7554
rect -2553 7524 -2487 7540
rect -3810 7463 -3794 7497
rect -3418 7463 -3402 7497
rect -2553 7490 -2537 7524
rect -2503 7490 -2487 7524
rect -2553 7473 -2487 7490
rect -2772 7436 -2627 7437
rect -3117 7402 -3101 7436
rect -2725 7418 -2627 7436
rect -2725 7402 -2626 7418
rect -2385 7402 -2369 7436
rect -2772 7401 -2626 7402
rect -1993 7401 -1891 7436
rect -3810 7345 -3794 7379
rect -3418 7345 -3402 7379
rect -2667 7363 -2626 7401
rect -2667 7329 -2339 7363
rect -3117 7284 -3101 7318
rect -2725 7284 -2709 7318
rect -4085 7196 -3993 7230
rect -3810 7227 -3794 7261
rect -3418 7227 -3402 7261
rect -2667 7202 -2626 7329
rect -2385 7318 -2339 7329
rect -2385 7284 -2369 7318
rect -1993 7284 -1977 7318
rect -2453 7258 -2419 7274
rect -2453 7208 -2419 7224
rect -2772 7200 -2626 7202
rect -4085 7074 -4065 7196
rect -4021 7144 -3993 7196
rect -3117 7166 -3101 7200
rect -2725 7166 -2626 7200
rect -2385 7166 -2369 7200
rect -1993 7166 -1977 7200
rect -4011 7106 -3993 7144
rect -4021 7074 -3993 7106
rect -4085 7028 -3993 7074
rect -3882 7109 -3794 7143
rect -3418 7109 -3402 7143
rect -3882 6907 -3847 7109
rect -3117 7048 -3101 7082
rect -2725 7048 -2709 7082
rect -3810 6991 -3794 7025
rect -3418 6991 -3402 7025
rect -2667 6964 -2626 7166
rect -2454 7140 -2420 7156
rect -2454 7090 -2420 7106
rect -2385 7048 -2369 7082
rect -1993 7048 -1977 7082
rect -1926 6965 -1891 7401
rect -1821 7246 -1733 7262
rect -1821 7206 -1805 7246
rect -1821 7114 -1805 7156
rect -1749 7114 -1733 7246
rect -1821 7098 -1733 7114
rect -3117 6930 -3101 6964
rect -2725 6930 -2626 6964
rect -2385 6930 -2369 6964
rect -1993 6930 -1891 6965
rect -2771 6928 -2626 6930
rect -3882 6873 -3794 6907
rect -3418 6873 -3402 6907
rect -3117 6812 -3101 6846
rect -2725 6812 -2709 6846
rect -3810 6755 -3794 6789
rect -3418 6755 -3402 6789
rect -3610 6626 -3594 6660
rect -3418 6626 -3402 6660
rect -3239 6574 -3205 6580
rect -3610 6508 -3594 6542
rect -3418 6508 -3402 6542
rect -3239 6514 -3205 6520
rect -3610 6390 -3594 6424
rect -3418 6390 -3402 6424
rect -2667 6342 -2626 6928
rect -2553 6876 -2487 6893
rect -2553 6842 -2537 6876
rect -2503 6842 -2487 6876
rect -2553 6826 -2487 6842
rect -2485 6552 -2469 6586
rect -2435 6552 -2419 6586
rect -2385 6524 -2369 6558
rect -2193 6524 -2177 6558
rect -2385 6406 -2369 6440
rect -2193 6406 -2177 6440
rect -3610 6272 -3594 6306
rect -3418 6272 -3402 6306
rect -1078 6087 -998 6092
rect -1078 6025 -1077 6087
rect -1011 6025 -998 6087
rect -3685 5879 -3596 5913
rect -3420 5879 -3404 5913
rect -3685 5677 -3650 5879
rect -3612 5761 -3596 5795
rect -3420 5761 -3404 5795
rect -2387 5754 -2371 5788
rect -2195 5754 -2179 5788
rect -3685 5643 -3596 5677
rect -3420 5643 -3404 5677
rect -2488 5607 -2472 5641
rect -2438 5607 -2422 5641
rect -2387 5636 -2371 5670
rect -2195 5636 -2179 5670
rect -3612 5525 -3596 5559
rect -3420 5525 -3404 5559
rect -3119 5452 -3103 5486
rect -2727 5452 -2711 5486
rect -2555 5456 -2489 5472
rect -3812 5395 -3796 5429
rect -3420 5395 -3404 5429
rect -2555 5422 -2539 5456
rect -2505 5422 -2489 5456
rect -2555 5405 -2489 5422
rect -2774 5368 -2629 5369
rect -3119 5334 -3103 5368
rect -2727 5350 -2629 5368
rect -2727 5334 -2628 5350
rect -2387 5334 -2371 5368
rect -2774 5333 -2628 5334
rect -1995 5333 -1893 5368
rect -3812 5277 -3796 5311
rect -3420 5277 -3404 5311
rect -2669 5295 -2628 5333
rect -2669 5261 -2341 5295
rect -3119 5216 -3103 5250
rect -2727 5216 -2711 5250
rect -4087 5128 -3995 5162
rect -3812 5159 -3796 5193
rect -3420 5159 -3404 5193
rect -2669 5134 -2628 5261
rect -2387 5250 -2341 5261
rect -2387 5216 -2371 5250
rect -1995 5216 -1979 5250
rect -2455 5190 -2421 5206
rect -2455 5140 -2421 5156
rect -2774 5132 -2628 5134
rect -4087 5006 -4067 5128
rect -4023 5076 -3995 5128
rect -3119 5098 -3103 5132
rect -2727 5098 -2628 5132
rect -2387 5098 -2371 5132
rect -1995 5098 -1979 5132
rect -4013 5038 -3995 5076
rect -4023 5006 -3995 5038
rect -4087 4960 -3995 5006
rect -3884 5041 -3796 5075
rect -3420 5041 -3404 5075
rect -3884 4839 -3849 5041
rect -3119 4980 -3103 5014
rect -2727 4980 -2711 5014
rect -3812 4923 -3796 4957
rect -3420 4923 -3404 4957
rect -2669 4896 -2628 5098
rect -2456 5072 -2422 5088
rect -2456 5022 -2422 5038
rect -2387 4980 -2371 5014
rect -1995 4980 -1979 5014
rect -1928 4897 -1893 5333
rect -1823 5178 -1735 5194
rect -1823 5138 -1807 5178
rect -1823 5046 -1807 5088
rect -1751 5046 -1735 5178
rect -1823 5030 -1735 5046
rect -3119 4862 -3103 4896
rect -2727 4862 -2628 4896
rect -2387 4862 -2371 4896
rect -1995 4862 -1893 4897
rect -2773 4860 -2628 4862
rect -3884 4805 -3796 4839
rect -3420 4805 -3404 4839
rect -3119 4744 -3103 4778
rect -2727 4744 -2711 4778
rect -3812 4687 -3796 4721
rect -3420 4687 -3404 4721
rect -3612 4558 -3596 4592
rect -3420 4558 -3404 4592
rect -3241 4506 -3207 4512
rect -3612 4440 -3596 4474
rect -3420 4440 -3404 4474
rect -3241 4446 -3207 4452
rect -3612 4322 -3596 4356
rect -3420 4322 -3404 4356
rect -2669 4274 -2628 4860
rect -2555 4808 -2489 4825
rect -2555 4774 -2539 4808
rect -2505 4774 -2489 4808
rect -2555 4758 -2489 4774
rect -2487 4484 -2471 4518
rect -2437 4484 -2421 4518
rect -2387 4456 -2371 4490
rect -2195 4456 -2179 4490
rect -2387 4338 -2371 4372
rect -2195 4338 -2179 4372
rect -3612 4204 -3596 4238
rect -3420 4204 -3404 4238
rect -1230 4008 -1144 4020
rect -1230 3953 -1224 4008
rect -1154 3953 -1144 4008
rect -3683 3810 -3594 3844
rect -3418 3810 -3402 3844
rect -3683 3608 -3648 3810
rect -3610 3692 -3594 3726
rect -3418 3692 -3402 3726
rect -2385 3685 -2369 3719
rect -2193 3685 -2177 3719
rect -3683 3574 -3594 3608
rect -3418 3574 -3402 3608
rect -2486 3538 -2470 3572
rect -2436 3538 -2420 3572
rect -2385 3567 -2369 3601
rect -2193 3567 -2177 3601
rect -3610 3456 -3594 3490
rect -3418 3456 -3402 3490
rect -3117 3383 -3101 3417
rect -2725 3383 -2709 3417
rect -2553 3387 -2487 3403
rect -3810 3326 -3794 3360
rect -3418 3326 -3402 3360
rect -2553 3353 -2537 3387
rect -2503 3353 -2487 3387
rect -2553 3336 -2487 3353
rect -2772 3299 -2627 3300
rect -3117 3265 -3101 3299
rect -2725 3281 -2627 3299
rect -2725 3265 -2626 3281
rect -2385 3265 -2369 3299
rect -2772 3264 -2626 3265
rect -1993 3264 -1891 3299
rect -3810 3208 -3794 3242
rect -3418 3208 -3402 3242
rect -2667 3226 -2626 3264
rect -2667 3192 -2339 3226
rect -3117 3147 -3101 3181
rect -2725 3147 -2709 3181
rect -4085 3059 -3993 3093
rect -3810 3090 -3794 3124
rect -3418 3090 -3402 3124
rect -2667 3065 -2626 3192
rect -2385 3181 -2339 3192
rect -2385 3147 -2369 3181
rect -1993 3147 -1977 3181
rect -2453 3121 -2419 3137
rect -2453 3071 -2419 3087
rect -2772 3063 -2626 3065
rect -4085 2937 -4065 3059
rect -4021 3007 -3993 3059
rect -3117 3029 -3101 3063
rect -2725 3029 -2626 3063
rect -2385 3029 -2369 3063
rect -1993 3029 -1977 3063
rect -4011 2969 -3993 3007
rect -4021 2937 -3993 2969
rect -4085 2891 -3993 2937
rect -3882 2972 -3794 3006
rect -3418 2972 -3402 3006
rect -3882 2770 -3847 2972
rect -3117 2911 -3101 2945
rect -2725 2911 -2709 2945
rect -3810 2854 -3794 2888
rect -3418 2854 -3402 2888
rect -2667 2827 -2626 3029
rect -2454 3003 -2420 3019
rect -2454 2953 -2420 2969
rect -2385 2911 -2369 2945
rect -1993 2911 -1977 2945
rect -1926 2828 -1891 3264
rect -1821 3109 -1733 3125
rect -1821 3069 -1805 3109
rect -1821 2977 -1805 3019
rect -1749 2977 -1733 3109
rect -1821 2961 -1733 2977
rect -3117 2793 -3101 2827
rect -2725 2793 -2626 2827
rect -2385 2793 -2369 2827
rect -1993 2793 -1891 2828
rect -2771 2791 -2626 2793
rect -3882 2736 -3794 2770
rect -3418 2736 -3402 2770
rect -3117 2675 -3101 2709
rect -2725 2675 -2709 2709
rect -3810 2618 -3794 2652
rect -3418 2618 -3402 2652
rect -3610 2489 -3594 2523
rect -3418 2489 -3402 2523
rect -3239 2437 -3205 2443
rect -3610 2371 -3594 2405
rect -3418 2371 -3402 2405
rect -3239 2377 -3205 2383
rect -3610 2253 -3594 2287
rect -3418 2253 -3402 2287
rect -2667 2205 -2626 2791
rect -2553 2739 -2487 2756
rect -2553 2705 -2537 2739
rect -2503 2705 -2487 2739
rect -2553 2689 -2487 2705
rect -2485 2415 -2469 2449
rect -2435 2415 -2419 2449
rect -2385 2387 -2369 2421
rect -2193 2387 -2177 2421
rect -2385 2269 -2369 2303
rect -2193 2269 -2177 2303
rect -3610 2135 -3594 2169
rect -3418 2135 -3402 2169
rect -3685 1742 -3596 1776
rect -3420 1742 -3404 1776
rect -3685 1540 -3650 1742
rect -3612 1624 -3596 1658
rect -3420 1624 -3404 1658
rect -2387 1617 -2371 1651
rect -2195 1617 -2179 1651
rect -3685 1506 -3596 1540
rect -3420 1506 -3404 1540
rect -2488 1470 -2472 1504
rect -2438 1470 -2422 1504
rect -2387 1499 -2371 1533
rect -2195 1499 -2179 1533
rect -3612 1388 -3596 1422
rect -3420 1388 -3404 1422
rect -3119 1315 -3103 1349
rect -2727 1315 -2711 1349
rect -2555 1319 -2489 1335
rect -3812 1258 -3796 1292
rect -3420 1258 -3404 1292
rect -2555 1285 -2539 1319
rect -2505 1285 -2489 1319
rect -2555 1268 -2489 1285
rect -2774 1231 -2629 1232
rect -3119 1197 -3103 1231
rect -2727 1213 -2629 1231
rect -2727 1197 -2628 1213
rect -2387 1197 -2371 1231
rect -2774 1196 -2628 1197
rect -1995 1196 -1893 1231
rect -3812 1140 -3796 1174
rect -3420 1140 -3404 1174
rect -2669 1158 -2628 1196
rect -2669 1124 -2341 1158
rect -3119 1079 -3103 1113
rect -2727 1079 -2711 1113
rect -4087 991 -3995 1025
rect -3812 1022 -3796 1056
rect -3420 1022 -3404 1056
rect -2669 997 -2628 1124
rect -2387 1113 -2341 1124
rect -2387 1079 -2371 1113
rect -1995 1079 -1979 1113
rect -2455 1053 -2421 1069
rect -2455 1003 -2421 1019
rect -2774 995 -2628 997
rect -4087 869 -4067 991
rect -4023 939 -3995 991
rect -3119 961 -3103 995
rect -2727 961 -2628 995
rect -2387 961 -2371 995
rect -1995 961 -1979 995
rect -4013 901 -3995 939
rect -4023 869 -3995 901
rect -4087 823 -3995 869
rect -3884 904 -3796 938
rect -3420 904 -3404 938
rect -3884 702 -3849 904
rect -3119 843 -3103 877
rect -2727 843 -2711 877
rect -3812 786 -3796 820
rect -3420 786 -3404 820
rect -2669 759 -2628 961
rect -2456 935 -2422 951
rect -2456 885 -2422 901
rect -2387 843 -2371 877
rect -1995 843 -1979 877
rect -1928 760 -1893 1196
rect -1823 1041 -1735 1057
rect -1823 1001 -1807 1041
rect -1823 909 -1807 951
rect -1751 909 -1735 1041
rect -1823 893 -1735 909
rect -3119 725 -3103 759
rect -2727 725 -2628 759
rect -2387 725 -2371 759
rect -1995 725 -1893 760
rect -2773 723 -2628 725
rect -3884 668 -3796 702
rect -3420 668 -3404 702
rect -3119 607 -3103 641
rect -2727 607 -2711 641
rect -3812 550 -3796 584
rect -3420 550 -3404 584
rect -3612 421 -3596 455
rect -3420 421 -3404 455
rect -3241 369 -3207 375
rect -3612 303 -3596 337
rect -3420 303 -3404 337
rect -3241 309 -3207 315
rect -3612 185 -3596 219
rect -3420 185 -3404 219
rect -2669 137 -2628 723
rect -2555 671 -2489 688
rect -2555 637 -2539 671
rect -2505 637 -2489 671
rect -2555 621 -2489 637
rect -2487 347 -2471 381
rect -2437 347 -2421 381
rect -1230 371 -1144 3953
rect -1078 909 -998 6025
rect -393 4009 -300 10028
rect -248 9795 -157 12564
rect -100 12597 -15 25447
rect 54 13927 125 25890
rect 5856 25766 5890 25782
rect 5974 25958 6008 25974
rect 5974 25766 6008 25782
rect 6092 25958 6126 25974
rect 6092 25766 6126 25782
rect 6210 25958 6244 25974
rect 6210 25766 6244 25782
rect 6328 25958 6362 25974
rect 6328 25766 6362 25782
rect 6446 25958 6480 25974
rect 6446 25766 6480 25782
rect 6564 25958 6598 25974
rect 6564 25766 6598 25782
rect 6682 25958 6716 26008
rect 6682 25766 6716 25782
rect 6800 25958 6834 25974
rect 6800 25766 6834 25782
rect 6918 25958 6952 26008
rect 6918 25766 6952 25782
rect 9962 26029 10187 26105
rect 9962 25880 10041 26029
rect 10108 25880 10187 26029
rect 13195 26005 13465 26039
rect 9962 25774 10187 25880
rect 12369 25955 12403 25971
rect 12369 25763 12403 25779
rect 12487 25955 12521 25971
rect 12487 25763 12521 25779
rect 12605 25955 12639 25971
rect 12605 25763 12639 25779
rect 12723 25955 12757 25971
rect 12723 25763 12757 25779
rect 12841 25955 12875 25971
rect 12841 25763 12875 25779
rect 12959 25955 12993 25971
rect 12959 25763 12993 25779
rect 13077 25955 13111 25971
rect 13077 25763 13111 25779
rect 13195 25955 13229 26005
rect 13195 25763 13229 25779
rect 13313 25955 13347 25971
rect 13313 25763 13347 25779
rect 13431 25955 13465 26005
rect 13431 25763 13465 25779
rect 16475 26026 16700 26102
rect 16475 25877 16554 26026
rect 16621 25877 16700 26026
rect 19729 26000 19999 26034
rect 16475 25771 16700 25877
rect 18903 25950 18937 25966
rect 18903 25758 18937 25774
rect 19021 25950 19055 25966
rect 19021 25758 19055 25774
rect 19139 25950 19173 25966
rect 19139 25758 19173 25774
rect 19257 25950 19291 25966
rect 19257 25758 19291 25774
rect 19375 25950 19409 25966
rect 19375 25758 19409 25774
rect 19493 25950 19527 25966
rect 19493 25758 19527 25774
rect 19611 25950 19645 25966
rect 19611 25758 19645 25774
rect 19729 25950 19763 26000
rect 19729 25758 19763 25774
rect 19847 25950 19881 25966
rect 19847 25758 19881 25774
rect 19965 25950 19999 26000
rect 19965 25758 19999 25774
rect 23009 26021 23234 26097
rect 23009 25872 23088 26021
rect 23155 25872 23234 26021
rect 26287 26004 26557 26038
rect 23009 25766 23234 25872
rect 25461 25954 25495 25970
rect 25461 25762 25495 25778
rect 25579 25954 25613 25970
rect 25579 25762 25613 25778
rect 25697 25954 25731 25970
rect 25697 25762 25731 25778
rect 25815 25954 25849 25970
rect 25815 25762 25849 25778
rect 25933 25954 25967 25970
rect 25933 25762 25967 25778
rect 26051 25954 26085 25970
rect 26051 25762 26085 25778
rect 26169 25954 26203 25970
rect 26169 25762 26203 25778
rect 26287 25954 26321 26004
rect 26287 25762 26321 25778
rect 26405 25954 26439 25970
rect 26405 25762 26439 25778
rect 26523 25954 26557 26004
rect 26523 25762 26557 25778
rect 29567 26025 29792 26101
rect 29567 25876 29646 26025
rect 29713 25876 29792 26025
rect 29567 25770 29792 25876
rect 6607 25688 6623 25722
rect 6657 25688 6673 25722
rect 13120 25685 13136 25719
rect 13170 25685 13186 25719
rect 19654 25680 19670 25714
rect 19704 25680 19720 25714
rect 26212 25684 26228 25718
rect 26262 25684 26278 25718
rect 6489 25571 6505 25605
rect 6539 25571 6555 25605
rect 8158 25594 8428 25629
rect 7804 25541 7838 25557
rect 6093 25521 6127 25537
rect 6093 25129 6127 25145
rect 6211 25521 6245 25537
rect 6211 25129 6245 25145
rect 6329 25521 6363 25537
rect 6446 25521 6480 25537
rect 6446 25329 6480 25345
rect 6564 25521 6598 25537
rect 6564 25329 6598 25345
rect 7320 25395 7590 25430
rect 7320 25341 7354 25395
rect 6329 25129 6363 25145
rect 6616 25195 6865 25238
rect 6616 25105 6663 25195
rect 6826 25105 6865 25195
rect 7320 25149 7354 25165
rect 7438 25341 7472 25357
rect 7438 25149 7472 25165
rect 7556 25341 7590 25395
rect 7556 25149 7590 25165
rect 7674 25341 7708 25357
rect 7674 25149 7708 25165
rect 7804 25149 7838 25165
rect 7922 25541 7956 25557
rect 7922 25149 7956 25165
rect 8040 25541 8074 25557
rect 8040 25149 8074 25165
rect 8158 25541 8192 25594
rect 8158 25149 8192 25165
rect 8276 25541 8310 25557
rect 8276 25149 8310 25165
rect 8394 25541 8428 25594
rect 10056 25594 10326 25629
rect 8394 25149 8428 25165
rect 8512 25541 8546 25557
rect 9702 25541 9736 25557
rect 9218 25395 9488 25430
rect 8512 25149 8546 25165
rect 8641 25341 8675 25357
rect 8641 25149 8675 25165
rect 8759 25341 8793 25357
rect 8759 25149 8793 25165
rect 8877 25341 8911 25357
rect 8877 25149 8911 25165
rect 8995 25341 9029 25357
rect 8995 25149 9029 25165
rect 9218 25341 9252 25395
rect 9218 25149 9252 25165
rect 9336 25341 9370 25357
rect 9336 25149 9370 25165
rect 9454 25341 9488 25395
rect 9454 25149 9488 25165
rect 9572 25341 9606 25357
rect 9572 25149 9606 25165
rect 9702 25149 9736 25165
rect 9820 25541 9854 25557
rect 9820 25149 9854 25165
rect 9938 25541 9972 25557
rect 9938 25149 9972 25165
rect 10056 25541 10090 25594
rect 10056 25149 10090 25165
rect 10174 25541 10208 25557
rect 10174 25149 10208 25165
rect 10292 25541 10326 25594
rect 13002 25568 13018 25602
rect 13052 25568 13068 25602
rect 14671 25591 14941 25626
rect 10292 25149 10326 25165
rect 10410 25541 10444 25557
rect 14317 25538 14351 25554
rect 12606 25518 12640 25534
rect 10410 25149 10444 25165
rect 10539 25341 10573 25357
rect 10539 25149 10573 25165
rect 10657 25341 10691 25357
rect 10657 25149 10691 25165
rect 10775 25341 10809 25357
rect 10775 25149 10809 25165
rect 10893 25341 10927 25357
rect 10893 25149 10927 25165
rect 12606 25126 12640 25142
rect 12724 25518 12758 25534
rect 12724 25126 12758 25142
rect 12842 25518 12876 25534
rect 12959 25518 12993 25534
rect 12959 25326 12993 25342
rect 13077 25518 13111 25534
rect 13077 25326 13111 25342
rect 13833 25392 14103 25427
rect 13833 25338 13867 25392
rect 12842 25126 12876 25142
rect 13129 25192 13378 25235
rect 6136 25061 6152 25095
rect 6186 25061 6202 25095
rect 6254 25061 6270 25095
rect 6304 25061 6320 25095
rect 6616 25066 6865 25105
rect 13129 25102 13176 25192
rect 13339 25102 13378 25192
rect 13833 25146 13867 25162
rect 13951 25338 13985 25354
rect 13951 25146 13985 25162
rect 14069 25338 14103 25392
rect 14069 25146 14103 25162
rect 14187 25338 14221 25354
rect 14187 25146 14221 25162
rect 14317 25146 14351 25162
rect 14435 25538 14469 25554
rect 14435 25146 14469 25162
rect 14553 25538 14587 25554
rect 14553 25146 14587 25162
rect 14671 25538 14705 25591
rect 14671 25146 14705 25162
rect 14789 25538 14823 25554
rect 14789 25146 14823 25162
rect 14907 25538 14941 25591
rect 16569 25591 16839 25626
rect 14907 25146 14941 25162
rect 15025 25538 15059 25554
rect 16215 25538 16249 25554
rect 15731 25392 16001 25427
rect 15025 25146 15059 25162
rect 15154 25338 15188 25354
rect 15154 25146 15188 25162
rect 15272 25338 15306 25354
rect 15272 25146 15306 25162
rect 15390 25338 15424 25354
rect 15390 25146 15424 25162
rect 15508 25338 15542 25354
rect 15508 25146 15542 25162
rect 15731 25338 15765 25392
rect 15731 25146 15765 25162
rect 15849 25338 15883 25354
rect 15849 25146 15883 25162
rect 15967 25338 16001 25392
rect 15967 25146 16001 25162
rect 16085 25338 16119 25354
rect 16085 25146 16119 25162
rect 16215 25146 16249 25162
rect 16333 25538 16367 25554
rect 16333 25146 16367 25162
rect 16451 25538 16485 25554
rect 16451 25146 16485 25162
rect 16569 25538 16603 25591
rect 16569 25146 16603 25162
rect 16687 25538 16721 25554
rect 16687 25146 16721 25162
rect 16805 25538 16839 25591
rect 19536 25563 19552 25597
rect 19586 25563 19602 25597
rect 21205 25586 21475 25621
rect 16805 25146 16839 25162
rect 16923 25538 16957 25554
rect 20851 25533 20885 25549
rect 19140 25513 19174 25529
rect 16923 25146 16957 25162
rect 17052 25338 17086 25354
rect 17052 25146 17086 25162
rect 17170 25338 17204 25354
rect 17170 25146 17204 25162
rect 17288 25338 17322 25354
rect 17288 25146 17322 25162
rect 17406 25338 17440 25354
rect 17406 25146 17440 25162
rect 19140 25121 19174 25137
rect 19258 25513 19292 25529
rect 19258 25121 19292 25137
rect 19376 25513 19410 25529
rect 19493 25513 19527 25529
rect 19493 25321 19527 25337
rect 19611 25513 19645 25529
rect 19611 25321 19645 25337
rect 20367 25387 20637 25422
rect 20367 25333 20401 25387
rect 19376 25121 19410 25137
rect 19663 25187 19912 25230
rect 12649 25058 12665 25092
rect 12699 25058 12715 25092
rect 12767 25058 12783 25092
rect 12817 25058 12833 25092
rect 13129 25063 13378 25102
rect 19663 25097 19710 25187
rect 19873 25097 19912 25187
rect 20367 25141 20401 25157
rect 20485 25333 20519 25349
rect 20485 25141 20519 25157
rect 20603 25333 20637 25387
rect 20603 25141 20637 25157
rect 20721 25333 20755 25349
rect 20721 25141 20755 25157
rect 20851 25141 20885 25157
rect 20969 25533 21003 25549
rect 20969 25141 21003 25157
rect 21087 25533 21121 25549
rect 21087 25141 21121 25157
rect 21205 25533 21239 25586
rect 21205 25141 21239 25157
rect 21323 25533 21357 25549
rect 21323 25141 21357 25157
rect 21441 25533 21475 25586
rect 23103 25586 23373 25621
rect 21441 25141 21475 25157
rect 21559 25533 21593 25549
rect 22749 25533 22783 25549
rect 22265 25387 22535 25422
rect 21559 25141 21593 25157
rect 21688 25333 21722 25349
rect 21688 25141 21722 25157
rect 21806 25333 21840 25349
rect 21806 25141 21840 25157
rect 21924 25333 21958 25349
rect 21924 25141 21958 25157
rect 22042 25333 22076 25349
rect 22042 25141 22076 25157
rect 22265 25333 22299 25387
rect 22265 25141 22299 25157
rect 22383 25333 22417 25349
rect 22383 25141 22417 25157
rect 22501 25333 22535 25387
rect 22501 25141 22535 25157
rect 22619 25333 22653 25349
rect 22619 25141 22653 25157
rect 22749 25141 22783 25157
rect 22867 25533 22901 25549
rect 22867 25141 22901 25157
rect 22985 25533 23019 25549
rect 22985 25141 23019 25157
rect 23103 25533 23137 25586
rect 23103 25141 23137 25157
rect 23221 25533 23255 25549
rect 23221 25141 23255 25157
rect 23339 25533 23373 25586
rect 26094 25567 26110 25601
rect 26144 25567 26160 25601
rect 27763 25590 28033 25625
rect 23339 25141 23373 25157
rect 23457 25533 23491 25549
rect 27409 25537 27443 25553
rect 25698 25517 25732 25533
rect 23457 25141 23491 25157
rect 23586 25333 23620 25349
rect 23586 25141 23620 25157
rect 23704 25333 23738 25349
rect 23704 25141 23738 25157
rect 23822 25333 23856 25349
rect 23822 25141 23856 25157
rect 23940 25333 23974 25349
rect 23940 25141 23974 25157
rect 25698 25125 25732 25141
rect 25816 25517 25850 25533
rect 25816 25125 25850 25141
rect 25934 25517 25968 25533
rect 26051 25517 26085 25533
rect 26051 25325 26085 25341
rect 26169 25517 26203 25533
rect 26169 25325 26203 25341
rect 26925 25391 27195 25426
rect 26925 25337 26959 25391
rect 25934 25125 25968 25141
rect 26221 25191 26470 25234
rect 19183 25053 19199 25087
rect 19233 25053 19249 25087
rect 19301 25053 19317 25087
rect 19351 25053 19367 25087
rect 19663 25058 19912 25097
rect 26221 25101 26268 25191
rect 26431 25101 26470 25191
rect 26925 25145 26959 25161
rect 27043 25337 27077 25353
rect 27043 25145 27077 25161
rect 27161 25337 27195 25391
rect 27161 25145 27195 25161
rect 27279 25337 27313 25353
rect 27279 25145 27313 25161
rect 27409 25145 27443 25161
rect 27527 25537 27561 25553
rect 27527 25145 27561 25161
rect 27645 25537 27679 25553
rect 27645 25145 27679 25161
rect 27763 25537 27797 25590
rect 27763 25145 27797 25161
rect 27881 25537 27915 25553
rect 27881 25145 27915 25161
rect 27999 25537 28033 25590
rect 29661 25590 29931 25625
rect 27999 25145 28033 25161
rect 28117 25537 28151 25553
rect 29307 25537 29341 25553
rect 28823 25391 29093 25426
rect 28117 25145 28151 25161
rect 28246 25337 28280 25353
rect 28246 25145 28280 25161
rect 28364 25337 28398 25353
rect 28364 25145 28398 25161
rect 28482 25337 28516 25353
rect 28482 25145 28516 25161
rect 28600 25337 28634 25353
rect 28600 25145 28634 25161
rect 28823 25337 28857 25391
rect 28823 25145 28857 25161
rect 28941 25337 28975 25353
rect 28941 25145 28975 25161
rect 29059 25337 29093 25391
rect 29059 25145 29093 25161
rect 29177 25337 29211 25353
rect 29177 25145 29211 25161
rect 29307 25145 29341 25161
rect 29425 25537 29459 25553
rect 29425 25145 29459 25161
rect 29543 25537 29577 25553
rect 29543 25145 29577 25161
rect 29661 25537 29695 25590
rect 29661 25145 29695 25161
rect 29779 25537 29813 25553
rect 29779 25145 29813 25161
rect 29897 25537 29931 25590
rect 29897 25145 29931 25161
rect 30015 25537 30049 25553
rect 34841 25387 34964 25403
rect 30015 25145 30049 25161
rect 30144 25337 30178 25353
rect 30144 25145 30178 25161
rect 30262 25337 30296 25353
rect 30262 25145 30296 25161
rect 30380 25337 30414 25353
rect 30380 25145 30414 25161
rect 30498 25337 30532 25353
rect 30498 25145 30532 25161
rect 34841 25322 34860 25387
rect 34943 25322 34964 25387
rect 25741 25057 25757 25091
rect 25791 25057 25807 25091
rect 25859 25057 25875 25091
rect 25909 25057 25925 25091
rect 26221 25062 26470 25101
rect 8784 24927 8818 24943
rect 15297 24924 15331 24940
rect 8784 24877 8818 24893
rect 10874 24906 10941 24922
rect 10874 24872 10891 24906
rect 10925 24872 10941 24906
rect 21831 24919 21865 24935
rect 15297 24874 15331 24890
rect 17387 24903 17454 24919
rect 7747 24848 7781 24864
rect 6246 24768 6469 24844
rect 6246 24619 6325 24768
rect 6392 24619 6469 24768
rect 6246 24513 6469 24619
rect 7865 24848 7899 24864
rect 7747 24456 7781 24472
rect 7864 24472 7865 24519
rect 7983 24848 8017 24864
rect 7899 24472 7900 24519
rect 6677 24404 6947 24438
rect 5851 24354 5885 24370
rect 5851 24162 5885 24178
rect 5969 24354 6003 24370
rect 5969 24162 6003 24178
rect 6087 24354 6121 24370
rect 6087 24162 6121 24178
rect 6205 24354 6239 24370
rect 6205 24162 6239 24178
rect 6323 24354 6357 24370
rect 6323 24162 6357 24178
rect 6441 24354 6475 24370
rect 6441 24162 6475 24178
rect 6559 24354 6593 24370
rect 6559 24162 6593 24178
rect 6677 24354 6711 24404
rect 6677 24162 6711 24178
rect 6795 24354 6829 24370
rect 6795 24162 6829 24178
rect 6913 24354 6947 24404
rect 7864 24414 7900 24472
rect 8101 24848 8135 24864
rect 7983 24456 8017 24472
rect 8099 24472 8101 24519
rect 8099 24414 8135 24472
rect 8219 24848 8253 24864
rect 8219 24456 8253 24472
rect 8337 24848 8371 24864
rect 8455 24848 8489 24864
rect 8371 24472 8373 24518
rect 8337 24414 8373 24472
rect 8455 24456 8489 24472
rect 9645 24848 9679 24864
rect 9763 24848 9797 24864
rect 9645 24456 9679 24472
rect 9762 24472 9763 24519
rect 9881 24848 9915 24864
rect 9797 24472 9798 24519
rect 8960 24414 9457 24432
rect 7864 24411 9457 24414
rect 7864 24377 9405 24411
rect 9439 24377 9457 24411
rect 7864 24374 9457 24377
rect 9762 24414 9798 24472
rect 9999 24848 10033 24864
rect 9881 24456 9915 24472
rect 9997 24472 9999 24519
rect 9997 24414 10033 24472
rect 10117 24848 10151 24864
rect 10117 24456 10151 24472
rect 10235 24848 10269 24864
rect 10353 24848 10387 24864
rect 10874 24856 10941 24872
rect 17387 24869 17404 24903
rect 17438 24869 17454 24903
rect 28389 24923 28423 24939
rect 21831 24869 21865 24885
rect 23921 24898 23988 24914
rect 10269 24472 10271 24518
rect 10235 24414 10271 24472
rect 14260 24845 14294 24861
rect 12759 24765 12982 24841
rect 12759 24616 12838 24765
rect 12905 24616 12982 24765
rect 12759 24510 12982 24616
rect 10353 24456 10387 24472
rect 14378 24845 14412 24861
rect 14260 24453 14294 24469
rect 14377 24469 14378 24516
rect 14496 24845 14530 24861
rect 14412 24469 14413 24516
rect 10858 24443 10958 24444
rect 10858 24414 11146 24443
rect 9762 24374 11146 24414
rect 7883 24373 9457 24374
rect 9781 24373 11146 24374
rect 7761 24284 7828 24300
rect 7761 24250 7777 24284
rect 7811 24250 7828 24284
rect 7761 24234 7828 24250
rect 6913 24162 6947 24178
rect 7592 24217 7626 24233
rect 7592 24167 7626 24183
rect 7938 24132 7972 24373
rect 8960 24356 9457 24373
rect 8408 24284 8475 24300
rect 8408 24250 8425 24284
rect 8459 24250 8475 24284
rect 8408 24234 8475 24250
rect 9659 24284 9726 24300
rect 9659 24250 9675 24284
rect 9709 24250 9726 24284
rect 9659 24234 9726 24250
rect 8715 24216 8749 24232
rect 8027 24166 8043 24200
rect 8077 24166 8093 24200
rect 8145 24167 8161 24201
rect 8195 24167 8211 24201
rect 8715 24166 8749 24182
rect 9490 24217 9524 24233
rect 9490 24167 9524 24183
rect 9836 24132 9870 24373
rect 10858 24368 11146 24373
rect 13190 24401 13460 24435
rect 10858 24345 11148 24368
rect 10858 24344 10958 24345
rect 10304 24285 10371 24301
rect 10304 24251 10321 24285
rect 10355 24251 10371 24285
rect 10304 24235 10371 24251
rect 10613 24216 10647 24232
rect 9925 24166 9941 24200
rect 9975 24166 9991 24200
rect 10043 24167 10059 24201
rect 10093 24167 10109 24201
rect 10613 24166 10647 24182
rect 6602 24084 6618 24118
rect 6652 24084 6668 24118
rect 7445 24116 7479 24132
rect 6484 23967 6500 24001
rect 6534 23967 6550 24001
rect 6088 23917 6122 23933
rect 6088 23525 6122 23541
rect 6206 23917 6240 23933
rect 6206 23525 6240 23541
rect 6324 23917 6358 23933
rect 6441 23917 6475 23933
rect 6441 23725 6475 23741
rect 6559 23917 6593 23933
rect 7445 23924 7479 23940
rect 7563 24116 7597 24132
rect 7563 23924 7597 23940
rect 7865 24116 7899 24132
rect 6559 23725 6593 23741
rect 7938 24116 8017 24132
rect 7938 24086 7983 24116
rect 7865 23673 7900 23740
rect 7983 23724 8017 23740
rect 8101 24116 8135 24132
rect 8101 23724 8135 23740
rect 8219 24116 8253 24132
rect 8337 24116 8371 24132
rect 8743 24116 8777 24132
rect 8743 23924 8777 23940
rect 8861 24116 8895 24132
rect 8861 23924 8895 23940
rect 9343 24116 9377 24132
rect 9343 23924 9377 23940
rect 9461 24116 9495 24132
rect 9461 23924 9495 23940
rect 9763 24116 9797 24132
rect 8219 23724 8253 23740
rect 8336 23673 8371 23740
rect 7865 23638 8371 23673
rect 9836 24116 9915 24132
rect 9836 24086 9881 24116
rect 9763 23673 9798 23740
rect 9881 23724 9915 23740
rect 9999 24116 10033 24132
rect 9999 23724 10033 23740
rect 10117 24116 10151 24132
rect 10235 24116 10269 24132
rect 10641 24116 10675 24132
rect 10641 23924 10675 23940
rect 10759 24116 10793 24132
rect 10759 23924 10793 23940
rect 10117 23724 10151 23740
rect 10234 23673 10269 23740
rect 9763 23638 10269 23673
rect 6324 23525 6358 23541
rect 6611 23591 6860 23634
rect 6611 23501 6658 23591
rect 6821 23501 6860 23591
rect 6131 23457 6147 23491
rect 6181 23457 6197 23491
rect 6249 23457 6265 23491
rect 6299 23457 6315 23491
rect 6611 23462 6860 23501
rect 8036 23431 8208 23478
rect 8036 23268 8075 23431
rect 8165 23268 8208 23431
rect 8036 23228 8208 23268
rect 11007 22728 11148 24345
rect 12364 24351 12398 24367
rect 12364 24159 12398 24175
rect 12482 24351 12516 24367
rect 12482 24159 12516 24175
rect 12600 24351 12634 24367
rect 12600 24159 12634 24175
rect 12718 24351 12752 24367
rect 12718 24159 12752 24175
rect 12836 24351 12870 24367
rect 12836 24159 12870 24175
rect 12954 24351 12988 24367
rect 12954 24159 12988 24175
rect 13072 24351 13106 24367
rect 13072 24159 13106 24175
rect 13190 24351 13224 24401
rect 13190 24159 13224 24175
rect 13308 24351 13342 24367
rect 13308 24159 13342 24175
rect 13426 24351 13460 24401
rect 14377 24411 14413 24469
rect 14614 24845 14648 24861
rect 14496 24453 14530 24469
rect 14612 24469 14614 24516
rect 14612 24411 14648 24469
rect 14732 24845 14766 24861
rect 14732 24453 14766 24469
rect 14850 24845 14884 24861
rect 14968 24845 15002 24861
rect 14884 24469 14886 24515
rect 14850 24411 14886 24469
rect 14968 24453 15002 24469
rect 16158 24845 16192 24861
rect 16276 24845 16310 24861
rect 16158 24453 16192 24469
rect 16275 24469 16276 24516
rect 16394 24845 16428 24861
rect 16310 24469 16311 24516
rect 15473 24411 15970 24429
rect 14377 24408 15970 24411
rect 14377 24374 15918 24408
rect 15952 24374 15970 24408
rect 14377 24371 15970 24374
rect 16275 24411 16311 24469
rect 16512 24845 16546 24861
rect 16394 24453 16428 24469
rect 16510 24469 16512 24516
rect 16510 24411 16546 24469
rect 16630 24845 16664 24861
rect 16630 24453 16664 24469
rect 16748 24845 16782 24861
rect 16866 24845 16900 24861
rect 17387 24853 17454 24869
rect 23921 24864 23938 24898
rect 23972 24864 23988 24898
rect 28389 24873 28423 24889
rect 30479 24902 30546 24918
rect 16782 24469 16784 24515
rect 16748 24411 16784 24469
rect 20794 24840 20828 24856
rect 19293 24760 19516 24836
rect 19293 24611 19372 24760
rect 19439 24611 19516 24760
rect 19293 24505 19516 24611
rect 16866 24453 16900 24469
rect 20912 24840 20946 24856
rect 20794 24448 20828 24464
rect 20911 24464 20912 24511
rect 21030 24840 21064 24856
rect 20946 24464 20947 24511
rect 17371 24440 17471 24441
rect 17371 24411 17659 24440
rect 16275 24399 17659 24411
rect 16275 24371 17660 24399
rect 14396 24370 15970 24371
rect 16294 24370 17660 24371
rect 14274 24281 14341 24297
rect 14274 24247 14290 24281
rect 14324 24247 14341 24281
rect 14274 24231 14341 24247
rect 13426 24159 13460 24175
rect 14105 24214 14139 24230
rect 14105 24164 14139 24180
rect 14451 24129 14485 24370
rect 15473 24353 15970 24370
rect 14921 24281 14988 24297
rect 14921 24247 14938 24281
rect 14972 24247 14988 24281
rect 14921 24231 14988 24247
rect 16172 24281 16239 24297
rect 16172 24247 16188 24281
rect 16222 24247 16239 24281
rect 16172 24231 16239 24247
rect 15228 24213 15262 24229
rect 14540 24163 14556 24197
rect 14590 24163 14606 24197
rect 14658 24164 14674 24198
rect 14708 24164 14724 24198
rect 15228 24163 15262 24179
rect 16003 24214 16037 24230
rect 16003 24164 16037 24180
rect 16349 24129 16383 24370
rect 17371 24342 17660 24370
rect 19724 24396 19994 24430
rect 17371 24341 17471 24342
rect 16817 24282 16884 24298
rect 16817 24248 16834 24282
rect 16868 24248 16884 24282
rect 16817 24232 16884 24248
rect 17126 24213 17160 24229
rect 16438 24163 16454 24197
rect 16488 24163 16504 24197
rect 16556 24164 16572 24198
rect 16606 24164 16622 24198
rect 17126 24163 17160 24179
rect 13115 24081 13131 24115
rect 13165 24081 13181 24115
rect 13958 24113 13992 24129
rect 12997 23964 13013 23998
rect 13047 23964 13063 23998
rect 12601 23914 12635 23930
rect 12601 23522 12635 23538
rect 12719 23914 12753 23930
rect 12719 23522 12753 23538
rect 12837 23914 12871 23930
rect 12954 23914 12988 23930
rect 12954 23722 12988 23738
rect 13072 23914 13106 23930
rect 13958 23921 13992 23937
rect 14076 24113 14110 24129
rect 14076 23921 14110 23937
rect 14378 24113 14412 24129
rect 13072 23722 13106 23738
rect 14451 24113 14530 24129
rect 14451 24083 14496 24113
rect 14378 23670 14413 23737
rect 14496 23721 14530 23737
rect 14614 24113 14648 24129
rect 14614 23721 14648 23737
rect 14732 24113 14766 24129
rect 14850 24113 14884 24129
rect 15256 24113 15290 24129
rect 15256 23921 15290 23937
rect 15374 24113 15408 24129
rect 15374 23921 15408 23937
rect 15856 24113 15890 24129
rect 15856 23921 15890 23937
rect 15974 24113 16008 24129
rect 15974 23921 16008 23937
rect 16276 24113 16310 24129
rect 14732 23721 14766 23737
rect 14849 23670 14884 23737
rect 14378 23635 14884 23670
rect 16349 24113 16428 24129
rect 16349 24083 16394 24113
rect 16276 23670 16311 23737
rect 16394 23721 16428 23737
rect 16512 24113 16546 24129
rect 16512 23721 16546 23737
rect 16630 24113 16664 24129
rect 16748 24113 16782 24129
rect 17154 24113 17188 24129
rect 17154 23921 17188 23937
rect 17272 24113 17306 24129
rect 17272 23921 17306 23937
rect 16630 23721 16664 23737
rect 16747 23670 16782 23737
rect 16276 23635 16782 23670
rect 12837 23522 12871 23538
rect 13124 23588 13373 23631
rect 13124 23498 13171 23588
rect 13334 23498 13373 23588
rect 12644 23454 12660 23488
rect 12694 23454 12710 23488
rect 12762 23454 12778 23488
rect 12812 23454 12828 23488
rect 13124 23459 13373 23498
rect 14549 23428 14721 23475
rect 14549 23265 14588 23428
rect 14678 23265 14721 23428
rect 14549 23225 14721 23265
rect 17532 22915 17660 24342
rect 18898 24346 18932 24362
rect 18898 24154 18932 24170
rect 19016 24346 19050 24362
rect 19016 24154 19050 24170
rect 19134 24346 19168 24362
rect 19134 24154 19168 24170
rect 19252 24346 19286 24362
rect 19252 24154 19286 24170
rect 19370 24346 19404 24362
rect 19370 24154 19404 24170
rect 19488 24346 19522 24362
rect 19488 24154 19522 24170
rect 19606 24346 19640 24362
rect 19606 24154 19640 24170
rect 19724 24346 19758 24396
rect 19724 24154 19758 24170
rect 19842 24346 19876 24362
rect 19842 24154 19876 24170
rect 19960 24346 19994 24396
rect 20911 24406 20947 24464
rect 21148 24840 21182 24856
rect 21030 24448 21064 24464
rect 21146 24464 21148 24511
rect 21146 24406 21182 24464
rect 21266 24840 21300 24856
rect 21266 24448 21300 24464
rect 21384 24840 21418 24856
rect 21502 24840 21536 24856
rect 21418 24464 21420 24510
rect 21384 24406 21420 24464
rect 21502 24448 21536 24464
rect 22692 24840 22726 24856
rect 22810 24840 22844 24856
rect 22692 24448 22726 24464
rect 22809 24464 22810 24511
rect 22928 24840 22962 24856
rect 22844 24464 22845 24511
rect 22007 24406 22504 24424
rect 20911 24403 22504 24406
rect 20911 24369 22452 24403
rect 22486 24369 22504 24403
rect 20911 24366 22504 24369
rect 22809 24406 22845 24464
rect 23046 24840 23080 24856
rect 22928 24448 22962 24464
rect 23044 24464 23046 24511
rect 23044 24406 23080 24464
rect 23164 24840 23198 24856
rect 23164 24448 23198 24464
rect 23282 24840 23316 24856
rect 23400 24840 23434 24856
rect 23921 24848 23988 24864
rect 30479 24868 30496 24902
rect 30530 24868 30546 24902
rect 27352 24844 27386 24860
rect 23316 24464 23318 24510
rect 23282 24406 23318 24464
rect 25851 24764 26074 24840
rect 25851 24615 25930 24764
rect 25997 24615 26074 24764
rect 25851 24509 26074 24615
rect 23400 24448 23434 24464
rect 27470 24844 27504 24860
rect 27352 24452 27386 24468
rect 27469 24468 27470 24515
rect 27588 24844 27622 24860
rect 27504 24468 27505 24515
rect 23905 24435 24005 24436
rect 23905 24406 24193 24435
rect 22809 24382 24193 24406
rect 26282 24400 26552 24434
rect 22809 24366 24194 24382
rect 20930 24365 22504 24366
rect 22828 24365 24194 24366
rect 20808 24276 20875 24292
rect 20808 24242 20824 24276
rect 20858 24242 20875 24276
rect 20808 24226 20875 24242
rect 19960 24154 19994 24170
rect 20639 24209 20673 24225
rect 20639 24159 20673 24175
rect 20985 24124 21019 24365
rect 22007 24348 22504 24365
rect 21455 24276 21522 24292
rect 21455 24242 21472 24276
rect 21506 24242 21522 24276
rect 21455 24226 21522 24242
rect 22706 24276 22773 24292
rect 22706 24242 22722 24276
rect 22756 24242 22773 24276
rect 22706 24226 22773 24242
rect 21762 24208 21796 24224
rect 21074 24158 21090 24192
rect 21124 24158 21140 24192
rect 21192 24159 21208 24193
rect 21242 24159 21258 24193
rect 21762 24158 21796 24174
rect 22537 24209 22571 24225
rect 22537 24159 22571 24175
rect 22883 24124 22917 24365
rect 23905 24337 24194 24365
rect 23905 24336 24005 24337
rect 23351 24277 23418 24293
rect 23351 24243 23368 24277
rect 23402 24243 23418 24277
rect 23351 24227 23418 24243
rect 23660 24208 23694 24224
rect 22972 24158 22988 24192
rect 23022 24158 23038 24192
rect 23090 24159 23106 24193
rect 23140 24159 23156 24193
rect 23660 24158 23694 24174
rect 19649 24076 19665 24110
rect 19699 24076 19715 24110
rect 20492 24108 20526 24124
rect 19531 23959 19547 23993
rect 19581 23959 19597 23993
rect 19135 23909 19169 23925
rect 19135 23517 19169 23533
rect 19253 23909 19287 23925
rect 19253 23517 19287 23533
rect 19371 23909 19405 23925
rect 19488 23909 19522 23925
rect 19488 23717 19522 23733
rect 19606 23909 19640 23925
rect 20492 23916 20526 23932
rect 20610 24108 20644 24124
rect 20610 23916 20644 23932
rect 20912 24108 20946 24124
rect 19606 23717 19640 23733
rect 20985 24108 21064 24124
rect 20985 24078 21030 24108
rect 20912 23665 20947 23732
rect 21030 23716 21064 23732
rect 21148 24108 21182 24124
rect 21148 23716 21182 23732
rect 21266 24108 21300 24124
rect 21384 24108 21418 24124
rect 21790 24108 21824 24124
rect 21790 23916 21824 23932
rect 21908 24108 21942 24124
rect 21908 23916 21942 23932
rect 22390 24108 22424 24124
rect 22390 23916 22424 23932
rect 22508 24108 22542 24124
rect 22508 23916 22542 23932
rect 22810 24108 22844 24124
rect 21266 23716 21300 23732
rect 21383 23665 21418 23732
rect 20912 23630 21418 23665
rect 22883 24108 22962 24124
rect 22883 24078 22928 24108
rect 22810 23665 22845 23732
rect 22928 23716 22962 23732
rect 23046 24108 23080 24124
rect 23046 23716 23080 23732
rect 23164 24108 23198 24124
rect 23282 24108 23316 24124
rect 23688 24108 23722 24124
rect 23688 23916 23722 23932
rect 23806 24108 23840 24124
rect 23806 23916 23840 23932
rect 23164 23716 23198 23732
rect 23281 23665 23316 23732
rect 22810 23630 23316 23665
rect 19371 23517 19405 23533
rect 19658 23583 19907 23626
rect 19658 23493 19705 23583
rect 19868 23493 19907 23583
rect 19178 23449 19194 23483
rect 19228 23449 19244 23483
rect 19296 23449 19312 23483
rect 19346 23449 19362 23483
rect 19658 23454 19907 23493
rect 21083 23423 21255 23470
rect 21083 23260 21122 23423
rect 21212 23260 21255 23423
rect 21083 23220 21255 23260
rect 24060 23064 24194 24337
rect 25456 24350 25490 24366
rect 25456 24158 25490 24174
rect 25574 24350 25608 24366
rect 25574 24158 25608 24174
rect 25692 24350 25726 24366
rect 25692 24158 25726 24174
rect 25810 24350 25844 24366
rect 25810 24158 25844 24174
rect 25928 24350 25962 24366
rect 25928 24158 25962 24174
rect 26046 24350 26080 24366
rect 26046 24158 26080 24174
rect 26164 24350 26198 24366
rect 26164 24158 26198 24174
rect 26282 24350 26316 24400
rect 26282 24158 26316 24174
rect 26400 24350 26434 24366
rect 26400 24158 26434 24174
rect 26518 24350 26552 24400
rect 27469 24410 27505 24468
rect 27706 24844 27740 24860
rect 27588 24452 27622 24468
rect 27704 24468 27706 24515
rect 27704 24410 27740 24468
rect 27824 24844 27858 24860
rect 27824 24452 27858 24468
rect 27942 24844 27976 24860
rect 28060 24844 28094 24860
rect 27976 24468 27978 24514
rect 27942 24410 27978 24468
rect 28060 24452 28094 24468
rect 29250 24844 29284 24860
rect 29368 24844 29402 24860
rect 29250 24452 29284 24468
rect 29367 24468 29368 24515
rect 29486 24844 29520 24860
rect 29402 24468 29403 24515
rect 28565 24410 29062 24428
rect 27469 24407 29062 24410
rect 27469 24373 29010 24407
rect 29044 24373 29062 24407
rect 27469 24370 29062 24373
rect 29367 24410 29403 24468
rect 29604 24844 29638 24860
rect 29486 24452 29520 24468
rect 29602 24468 29604 24515
rect 29602 24410 29638 24468
rect 29722 24844 29756 24860
rect 29722 24452 29756 24468
rect 29840 24844 29874 24860
rect 29958 24844 29992 24860
rect 30479 24852 30546 24868
rect 29874 24468 29876 24514
rect 29840 24410 29876 24468
rect 29958 24452 29992 24468
rect 30463 24439 30563 24440
rect 30642 24439 32317 24440
rect 30463 24429 32317 24439
rect 30463 24410 32159 24429
rect 29367 24370 32159 24410
rect 27488 24369 29062 24370
rect 29386 24369 32159 24370
rect 27366 24280 27433 24296
rect 27366 24246 27382 24280
rect 27416 24246 27433 24280
rect 27366 24230 27433 24246
rect 26518 24158 26552 24174
rect 27197 24213 27231 24229
rect 27197 24163 27231 24179
rect 27543 24128 27577 24369
rect 28565 24352 29062 24369
rect 28013 24280 28080 24296
rect 28013 24246 28030 24280
rect 28064 24246 28080 24280
rect 28013 24230 28080 24246
rect 29264 24280 29331 24296
rect 29264 24246 29280 24280
rect 29314 24246 29331 24280
rect 29264 24230 29331 24246
rect 28320 24212 28354 24228
rect 27632 24162 27648 24196
rect 27682 24162 27698 24196
rect 27750 24163 27766 24197
rect 27800 24163 27816 24197
rect 28320 24162 28354 24178
rect 29095 24213 29129 24229
rect 29095 24163 29129 24179
rect 29441 24128 29475 24369
rect 30463 24351 32159 24369
rect 32304 24351 32317 24429
rect 30463 24343 32317 24351
rect 30463 24341 30751 24343
rect 30463 24340 30563 24341
rect 29909 24281 29976 24297
rect 29909 24247 29926 24281
rect 29960 24247 29976 24281
rect 29909 24231 29976 24247
rect 30218 24212 30252 24228
rect 29530 24162 29546 24196
rect 29580 24162 29596 24196
rect 29648 24163 29664 24197
rect 29698 24163 29714 24197
rect 30218 24162 30252 24178
rect 26207 24080 26223 24114
rect 26257 24080 26273 24114
rect 27050 24112 27084 24128
rect 26089 23963 26105 23997
rect 26139 23963 26155 23997
rect 25693 23913 25727 23929
rect 25693 23521 25727 23537
rect 25811 23913 25845 23929
rect 25811 23521 25845 23537
rect 25929 23913 25963 23929
rect 26046 23913 26080 23929
rect 26046 23721 26080 23737
rect 26164 23913 26198 23929
rect 27050 23920 27084 23936
rect 27168 24112 27202 24128
rect 27168 23920 27202 23936
rect 27470 24112 27504 24128
rect 26164 23721 26198 23737
rect 27543 24112 27622 24128
rect 27543 24082 27588 24112
rect 27470 23669 27505 23736
rect 27588 23720 27622 23736
rect 27706 24112 27740 24128
rect 27706 23720 27740 23736
rect 27824 24112 27858 24128
rect 27942 24112 27976 24128
rect 28348 24112 28382 24128
rect 28348 23920 28382 23936
rect 28466 24112 28500 24128
rect 28466 23920 28500 23936
rect 28948 24112 28982 24128
rect 28948 23920 28982 23936
rect 29066 24112 29100 24128
rect 29066 23920 29100 23936
rect 29368 24112 29402 24128
rect 27824 23720 27858 23736
rect 27941 23669 27976 23736
rect 27470 23634 27976 23669
rect 29441 24112 29520 24128
rect 29441 24082 29486 24112
rect 29368 23669 29403 23736
rect 29486 23720 29520 23736
rect 29604 24112 29638 24128
rect 29604 23720 29638 23736
rect 29722 24112 29756 24128
rect 29840 24112 29874 24128
rect 30246 24112 30280 24128
rect 30246 23920 30280 23936
rect 30364 24112 30398 24128
rect 30364 23920 30398 23936
rect 29722 23720 29756 23736
rect 29839 23669 29874 23736
rect 29368 23634 29874 23669
rect 25929 23521 25963 23537
rect 26216 23587 26465 23630
rect 26216 23497 26263 23587
rect 26426 23497 26465 23587
rect 25736 23453 25752 23487
rect 25786 23453 25802 23487
rect 25854 23453 25870 23487
rect 25904 23453 25920 23487
rect 26216 23458 26465 23497
rect 27641 23427 27813 23474
rect 27641 23264 27680 23427
rect 27770 23264 27813 23427
rect 27641 23224 27813 23264
rect 24060 23063 32825 23064
rect 24060 23049 32831 23063
rect 24060 22977 32676 23049
rect 32811 22977 32831 23049
rect 24060 22969 32831 22977
rect 24060 22965 32825 22969
rect 24060 22961 24194 22965
rect 17529 22899 33393 22915
rect 17529 22809 33244 22899
rect 33374 22809 33393 22899
rect 17529 22792 33393 22809
rect 34841 22728 34964 25322
rect 35178 25322 37815 25404
rect 35178 25178 35295 25322
rect 37727 25287 37815 25322
rect 37727 25238 37741 25287
rect 37801 25238 37815 25287
rect 37727 25222 37815 25238
rect 35178 23450 35297 25178
rect 36877 25114 36967 25148
rect 37143 25114 37159 25148
rect 36877 24912 36916 25114
rect 37441 25043 37526 25059
rect 36951 24996 36967 25030
rect 37143 24996 37233 25030
rect 36877 24878 36967 24912
rect 37143 24878 37159 24912
rect 37194 24794 37233 24996
rect 37441 24983 37458 25043
rect 37513 24983 37526 25043
rect 37441 24967 37526 24983
rect 36951 24760 36967 24794
rect 37143 24760 37233 24794
rect 36675 24673 36767 24707
rect 37143 24673 37159 24707
rect 36675 24471 36714 24673
rect 36751 24555 36767 24589
rect 37143 24555 37233 24589
rect 36675 24437 36767 24471
rect 37143 24437 37159 24471
rect 37194 24353 37233 24555
rect 36751 24319 36767 24353
rect 37143 24319 37233 24353
rect 36676 24206 36767 24240
rect 37143 24206 37159 24240
rect 36676 24004 36715 24206
rect 37194 24122 37233 24319
rect 38084 24280 38100 24314
rect 38276 24280 38292 24314
rect 38084 24162 38100 24196
rect 38276 24162 38292 24196
rect 38088 24122 38288 24162
rect 36751 24088 36767 24122
rect 37143 24088 37233 24122
rect 36479 23962 36589 23978
rect 36676 23970 36767 24004
rect 37143 23970 37159 24004
rect 36479 23766 36497 23962
rect 36573 23766 36589 23962
rect 37194 23886 37233 24088
rect 37729 24076 37814 24092
rect 38084 24088 38100 24122
rect 38476 24088 38492 24122
rect 37342 24028 37358 24062
rect 37392 24028 37408 24062
rect 37729 24016 37742 24076
rect 37797 24016 37814 24076
rect 37729 24000 37814 24016
rect 36751 23852 36767 23886
rect 37143 23852 37233 23886
rect 37444 23958 37529 23974
rect 38084 23970 38100 24004
rect 38476 23970 38492 24004
rect 37444 23898 37457 23958
rect 37512 23898 37529 23958
rect 38725 23904 38811 23920
rect 37444 23882 37529 23898
rect 38084 23852 38100 23886
rect 38476 23852 38492 23886
rect 38577 23885 38611 23901
rect 36479 23750 36589 23766
rect 36676 23734 36767 23768
rect 37143 23734 37159 23768
rect 36676 23532 36715 23734
rect 37194 23650 37233 23852
rect 38577 23835 38611 23851
rect 38725 23882 38743 23904
rect 37962 23793 37978 23827
rect 38012 23793 38028 23827
rect 38725 23824 38729 23882
rect 38725 23800 38743 23824
rect 38789 23800 38811 23904
rect 38725 23784 38811 23800
rect 38084 23734 38100 23768
rect 38476 23734 38492 23768
rect 37572 23674 37588 23708
rect 37622 23674 37638 23708
rect 36751 23616 36767 23650
rect 37143 23616 37233 23650
rect 38084 23616 38100 23650
rect 38476 23616 38492 23650
rect 36676 23498 36767 23532
rect 37143 23498 37159 23532
rect 35178 22934 35296 23450
rect 37194 23413 37233 23616
rect 38088 23572 38288 23616
rect 38084 23538 38100 23572
rect 38276 23538 38292 23572
rect 38084 23420 38100 23454
rect 38276 23420 38292 23454
rect 36751 23379 36767 23413
rect 37143 23379 37233 23413
rect 36676 23261 36767 23295
rect 37143 23261 37159 23295
rect 36676 23059 36715 23261
rect 37194 23177 37233 23379
rect 36751 23143 36767 23177
rect 37143 23143 37233 23177
rect 36676 23025 36767 23059
rect 37143 23025 37159 23059
rect 11007 22607 34964 22728
rect 11007 22606 34960 22607
rect 11007 22604 11146 22606
rect 35174 22570 35298 22934
rect 36951 22906 36967 22940
rect 37143 22906 37236 22940
rect 5815 22468 6038 22544
rect 5815 22319 5892 22468
rect 5959 22319 6038 22468
rect 5815 22213 6038 22319
rect 6962 22468 7185 22544
rect 6962 22319 7039 22468
rect 7106 22319 7185 22468
rect 6688 22254 6722 22270
rect 6688 22204 6722 22220
rect 6962 22213 7185 22319
rect 9444 22414 9667 22490
rect 9444 22265 9521 22414
rect 9588 22265 9667 22414
rect 7818 22248 7852 22264
rect 7818 22198 7852 22214
rect 9444 22159 9667 22265
rect 12373 22464 12596 22540
rect 12373 22315 12450 22464
rect 12517 22315 12596 22464
rect 12373 22209 12596 22315
rect 13520 22464 13743 22540
rect 13520 22315 13597 22464
rect 13664 22315 13743 22464
rect 13246 22250 13280 22266
rect 13246 22200 13280 22216
rect 13520 22209 13743 22315
rect 16002 22410 16225 22486
rect 16002 22261 16079 22410
rect 16146 22261 16225 22410
rect 14376 22244 14410 22260
rect 14376 22194 14410 22210
rect 16002 22155 16225 22261
rect 18907 22469 19130 22545
rect 18907 22320 18984 22469
rect 19051 22320 19130 22469
rect 18907 22214 19130 22320
rect 20054 22469 20277 22545
rect 20054 22320 20131 22469
rect 20198 22320 20277 22469
rect 19780 22255 19814 22271
rect 19780 22205 19814 22221
rect 20054 22214 20277 22320
rect 22536 22415 22759 22491
rect 22536 22266 22613 22415
rect 22680 22266 22759 22415
rect 20910 22249 20944 22265
rect 20910 22199 20944 22215
rect 22536 22160 22759 22266
rect 25420 22472 25643 22548
rect 25420 22323 25497 22472
rect 25564 22323 25643 22472
rect 25420 22217 25643 22323
rect 26567 22472 26790 22548
rect 30844 22528 35298 22570
rect 36880 22788 36967 22822
rect 37143 22788 37159 22822
rect 36880 22586 36917 22788
rect 37197 22704 37236 22906
rect 36951 22670 36967 22704
rect 37143 22670 37236 22704
rect 37317 22752 37351 22768
rect 37317 22702 37351 22718
rect 36880 22552 36967 22586
rect 37143 22552 37159 22586
rect 26567 22323 26644 22472
rect 26711 22323 26790 22472
rect 26293 22258 26327 22274
rect 26293 22208 26327 22224
rect 26567 22217 26790 22323
rect 29049 22418 29272 22494
rect 29049 22269 29126 22418
rect 29193 22269 29272 22418
rect 27423 22252 27457 22268
rect 27423 22202 27457 22218
rect 29049 22163 29272 22269
rect 30844 22445 35300 22528
rect 6688 22134 6722 22150
rect 5853 22076 5887 22092
rect 5853 21684 5887 21700
rect 5971 22076 6005 22092
rect 5971 21684 6005 21700
rect 6089 22076 6123 22092
rect 6089 21684 6123 21700
rect 6207 22076 6241 22092
rect 6207 21684 6241 21700
rect 6325 22076 6359 22092
rect 6325 21684 6359 21700
rect 6443 22076 6477 22092
rect 6443 21684 6477 21700
rect 6561 22076 6595 22092
rect 6688 22084 6722 22100
rect 7818 22130 7852 22146
rect 6561 21684 6595 21700
rect 6995 22072 7029 22088
rect 6995 21680 7029 21696
rect 7113 22072 7147 22088
rect 7113 21680 7147 21696
rect 7231 22072 7265 22088
rect 7231 21680 7265 21696
rect 7349 22072 7383 22088
rect 7349 21680 7383 21696
rect 7467 22072 7501 22088
rect 7467 21680 7501 21696
rect 7585 22072 7619 22088
rect 7585 21680 7619 21696
rect 7703 22072 7737 22088
rect 7818 22080 7852 22096
rect 13246 22130 13280 22146
rect 8966 22050 9236 22084
rect 8966 22000 9000 22050
rect 8966 21808 9000 21824
rect 9084 22000 9118 22016
rect 9084 21808 9118 21824
rect 9202 22000 9236 22050
rect 12411 22072 12445 22088
rect 9202 21808 9236 21824
rect 9320 22000 9354 22016
rect 9320 21808 9354 21824
rect 9438 22000 9472 22016
rect 9438 21808 9472 21824
rect 9556 22000 9590 22016
rect 9556 21808 9590 21824
rect 9674 22000 9708 22016
rect 9674 21808 9708 21824
rect 9792 22000 9826 22016
rect 9792 21808 9826 21824
rect 9910 22000 9944 22016
rect 9910 21808 9944 21824
rect 10028 22000 10062 22016
rect 10028 21808 10062 21824
rect 9245 21730 9261 21764
rect 9295 21730 9311 21764
rect 7703 21680 7737 21696
rect 12411 21680 12445 21696
rect 12529 22072 12563 22088
rect 12529 21680 12563 21696
rect 12647 22072 12681 22088
rect 12647 21680 12681 21696
rect 12765 22072 12799 22088
rect 12765 21680 12799 21696
rect 12883 22072 12917 22088
rect 12883 21680 12917 21696
rect 13001 22072 13035 22088
rect 13001 21680 13035 21696
rect 13119 22072 13153 22088
rect 13246 22080 13280 22096
rect 14376 22126 14410 22142
rect 19780 22135 19814 22151
rect 13119 21680 13153 21696
rect 13553 22068 13587 22084
rect 13553 21676 13587 21692
rect 13671 22068 13705 22084
rect 13671 21676 13705 21692
rect 13789 22068 13823 22084
rect 13789 21676 13823 21692
rect 13907 22068 13941 22084
rect 13907 21676 13941 21692
rect 14025 22068 14059 22084
rect 14025 21676 14059 21692
rect 14143 22068 14177 22084
rect 14143 21676 14177 21692
rect 14261 22068 14295 22084
rect 14376 22076 14410 22092
rect 15524 22046 15794 22080
rect 15524 21996 15558 22046
rect 15524 21804 15558 21820
rect 15642 21996 15676 22012
rect 15642 21804 15676 21820
rect 15760 21996 15794 22046
rect 18945 22077 18979 22093
rect 15760 21804 15794 21820
rect 15878 21996 15912 22012
rect 15878 21804 15912 21820
rect 15996 21996 16030 22012
rect 15996 21804 16030 21820
rect 16114 21996 16148 22012
rect 16114 21804 16148 21820
rect 16232 21996 16266 22012
rect 16232 21804 16266 21820
rect 16350 21996 16384 22012
rect 16350 21804 16384 21820
rect 16468 21996 16502 22012
rect 16468 21804 16502 21820
rect 16586 21996 16620 22012
rect 16586 21804 16620 21820
rect 15803 21726 15819 21760
rect 15853 21726 15869 21760
rect 14261 21676 14295 21692
rect 18945 21685 18979 21701
rect 19063 22077 19097 22093
rect 19063 21685 19097 21701
rect 19181 22077 19215 22093
rect 19181 21685 19215 21701
rect 19299 22077 19333 22093
rect 19299 21685 19333 21701
rect 19417 22077 19451 22093
rect 19417 21685 19451 21701
rect 19535 22077 19569 22093
rect 19535 21685 19569 21701
rect 19653 22077 19687 22093
rect 19780 22085 19814 22101
rect 20910 22131 20944 22147
rect 19653 21685 19687 21701
rect 20087 22073 20121 22089
rect 20087 21681 20121 21697
rect 20205 22073 20239 22089
rect 20205 21681 20239 21697
rect 20323 22073 20357 22089
rect 20323 21681 20357 21697
rect 20441 22073 20475 22089
rect 20441 21681 20475 21697
rect 20559 22073 20593 22089
rect 20559 21681 20593 21697
rect 20677 22073 20711 22089
rect 20677 21681 20711 21697
rect 20795 22073 20829 22089
rect 20910 22081 20944 22097
rect 26293 22138 26327 22154
rect 22058 22051 22328 22085
rect 22058 22001 22092 22051
rect 22058 21809 22092 21825
rect 22176 22001 22210 22017
rect 22176 21809 22210 21825
rect 22294 22001 22328 22051
rect 25458 22080 25492 22096
rect 22294 21809 22328 21825
rect 22412 22001 22446 22017
rect 22412 21809 22446 21825
rect 22530 22001 22564 22017
rect 22530 21809 22564 21825
rect 22648 22001 22682 22017
rect 22648 21809 22682 21825
rect 22766 22001 22800 22017
rect 22766 21809 22800 21825
rect 22884 22001 22918 22017
rect 22884 21809 22918 21825
rect 23002 22001 23036 22017
rect 23002 21809 23036 21825
rect 23120 22001 23154 22017
rect 23120 21809 23154 21825
rect 22337 21731 22353 21765
rect 22387 21731 22403 21765
rect 20795 21681 20829 21697
rect 25458 21688 25492 21704
rect 25576 22080 25610 22096
rect 25576 21688 25610 21704
rect 25694 22080 25728 22096
rect 25694 21688 25728 21704
rect 25812 22080 25846 22096
rect 25812 21688 25846 21704
rect 25930 22080 25964 22096
rect 25930 21688 25964 21704
rect 26048 22080 26082 22096
rect 26048 21688 26082 21704
rect 26166 22080 26200 22096
rect 26293 22088 26327 22104
rect 27423 22134 27457 22150
rect 26166 21688 26200 21704
rect 26600 22076 26634 22092
rect 26600 21684 26634 21700
rect 26718 22076 26752 22092
rect 26718 21684 26752 21700
rect 26836 22076 26870 22092
rect 26836 21684 26870 21700
rect 26954 22076 26988 22092
rect 26954 21684 26988 21700
rect 27072 22076 27106 22092
rect 27072 21684 27106 21700
rect 27190 22076 27224 22092
rect 27190 21684 27224 21700
rect 27308 22076 27342 22092
rect 27423 22084 27457 22100
rect 28571 22054 28841 22088
rect 28571 22004 28605 22054
rect 28571 21812 28605 21828
rect 28689 22004 28723 22020
rect 28689 21812 28723 21828
rect 28807 22004 28841 22054
rect 28807 21812 28841 21828
rect 28925 22004 28959 22020
rect 28925 21812 28959 21828
rect 29043 22004 29077 22020
rect 29043 21812 29077 21828
rect 29161 22004 29195 22020
rect 29161 21812 29195 21828
rect 29279 22004 29313 22020
rect 29279 21812 29313 21828
rect 29397 22004 29431 22020
rect 29397 21812 29431 21828
rect 29515 22004 29549 22020
rect 29515 21812 29549 21828
rect 29633 22004 29667 22020
rect 29633 21812 29667 21828
rect 28850 21734 28866 21768
rect 28900 21734 28916 21768
rect 27308 21684 27342 21700
rect 9363 21613 9379 21647
rect 9413 21613 9429 21647
rect 15921 21609 15937 21643
rect 15971 21609 15987 21643
rect 22455 21614 22471 21648
rect 22505 21614 22521 21648
rect 28968 21617 28984 21651
rect 29018 21617 29034 21651
rect 9320 21563 9354 21579
rect 6340 21344 6356 21378
rect 6390 21344 6406 21378
rect 7482 21340 7498 21374
rect 7532 21340 7548 21374
rect 9320 21371 9354 21387
rect 9438 21563 9472 21579
rect 9438 21371 9472 21387
rect 9555 21563 9589 21579
rect 5778 21293 5812 21309
rect 5778 21101 5812 21117
rect 5896 21293 5930 21309
rect 5896 21101 5930 21117
rect 6014 21293 6048 21309
rect 6014 21101 6048 21117
rect 6132 21293 6166 21309
rect 6132 21101 6166 21117
rect 6297 21293 6331 21309
rect 6297 21101 6331 21117
rect 6415 21293 6449 21309
rect 6415 21101 6449 21117
rect 6533 21293 6567 21309
rect 6533 21101 6567 21117
rect 6651 21293 6685 21309
rect 6651 21101 6685 21117
rect 6920 21289 6954 21305
rect 6920 21097 6954 21113
rect 7038 21289 7072 21305
rect 7038 21097 7072 21113
rect 7156 21289 7190 21305
rect 7156 21097 7190 21113
rect 7274 21289 7308 21305
rect 7274 21097 7308 21113
rect 7439 21289 7473 21305
rect 7439 21097 7473 21113
rect 7557 21289 7591 21305
rect 7557 21097 7591 21113
rect 7675 21289 7709 21305
rect 7675 21097 7709 21113
rect 7793 21289 7827 21305
rect 7793 21097 7827 21113
rect 9053 21237 9302 21280
rect 9053 21147 9092 21237
rect 9255 21147 9302 21237
rect 9555 21171 9589 21187
rect 9673 21563 9707 21579
rect 9673 21171 9707 21187
rect 9791 21563 9825 21579
rect 15878 21559 15912 21575
rect 12898 21340 12914 21374
rect 12948 21340 12964 21374
rect 14040 21336 14056 21370
rect 14090 21336 14106 21370
rect 15878 21367 15912 21383
rect 15996 21559 16030 21575
rect 15996 21367 16030 21383
rect 16113 21559 16147 21575
rect 9791 21171 9825 21187
rect 12336 21289 12370 21305
rect 9053 21108 9302 21147
rect 9598 21103 9614 21137
rect 9648 21103 9664 21137
rect 9716 21103 9732 21137
rect 9766 21103 9782 21137
rect 12336 21097 12370 21113
rect 12454 21289 12488 21305
rect 12454 21097 12488 21113
rect 12572 21289 12606 21305
rect 12572 21097 12606 21113
rect 12690 21289 12724 21305
rect 12690 21097 12724 21113
rect 12855 21289 12889 21305
rect 12855 21097 12889 21113
rect 12973 21289 13007 21305
rect 12973 21097 13007 21113
rect 13091 21289 13125 21305
rect 13091 21097 13125 21113
rect 13209 21289 13243 21305
rect 13209 21097 13243 21113
rect 13478 21285 13512 21301
rect 13478 21093 13512 21109
rect 13596 21285 13630 21301
rect 13596 21093 13630 21109
rect 13714 21285 13748 21301
rect 13714 21093 13748 21109
rect 13832 21285 13866 21301
rect 13832 21093 13866 21109
rect 13997 21285 14031 21301
rect 13997 21093 14031 21109
rect 14115 21285 14149 21301
rect 14115 21093 14149 21109
rect 14233 21285 14267 21301
rect 14233 21093 14267 21109
rect 14351 21285 14385 21301
rect 14351 21093 14385 21109
rect 15611 21233 15860 21276
rect 15611 21143 15650 21233
rect 15813 21143 15860 21233
rect 16113 21167 16147 21183
rect 16231 21559 16265 21575
rect 16231 21167 16265 21183
rect 16349 21559 16383 21575
rect 22412 21564 22446 21580
rect 19432 21345 19448 21379
rect 19482 21345 19498 21379
rect 20574 21341 20590 21375
rect 20624 21341 20640 21375
rect 22412 21372 22446 21388
rect 22530 21564 22564 21580
rect 22530 21372 22564 21388
rect 22647 21564 22681 21580
rect 16349 21167 16383 21183
rect 18870 21294 18904 21310
rect 15611 21104 15860 21143
rect 16156 21099 16172 21133
rect 16206 21099 16222 21133
rect 16274 21099 16290 21133
rect 16324 21099 16340 21133
rect 18870 21102 18904 21118
rect 18988 21294 19022 21310
rect 18988 21102 19022 21118
rect 19106 21294 19140 21310
rect 19106 21102 19140 21118
rect 19224 21294 19258 21310
rect 19224 21102 19258 21118
rect 19389 21294 19423 21310
rect 19389 21102 19423 21118
rect 19507 21294 19541 21310
rect 19507 21102 19541 21118
rect 19625 21294 19659 21310
rect 19625 21102 19659 21118
rect 19743 21294 19777 21310
rect 19743 21102 19777 21118
rect 20012 21290 20046 21306
rect 20012 21098 20046 21114
rect 20130 21290 20164 21306
rect 20130 21098 20164 21114
rect 20248 21290 20282 21306
rect 20248 21098 20282 21114
rect 20366 21290 20400 21306
rect 20366 21098 20400 21114
rect 20531 21290 20565 21306
rect 20531 21098 20565 21114
rect 20649 21290 20683 21306
rect 20649 21098 20683 21114
rect 20767 21290 20801 21306
rect 20767 21098 20801 21114
rect 20885 21290 20919 21306
rect 20885 21098 20919 21114
rect 22145 21238 22394 21281
rect 22145 21148 22184 21238
rect 22347 21148 22394 21238
rect 22647 21172 22681 21188
rect 22765 21564 22799 21580
rect 22765 21172 22799 21188
rect 22883 21564 22917 21580
rect 28925 21567 28959 21583
rect 25945 21348 25961 21382
rect 25995 21348 26011 21382
rect 27087 21344 27103 21378
rect 27137 21344 27153 21378
rect 28925 21375 28959 21391
rect 29043 21567 29077 21583
rect 29043 21375 29077 21391
rect 29160 21567 29194 21583
rect 22883 21172 22917 21188
rect 25383 21297 25417 21313
rect 22145 21109 22394 21148
rect 22690 21104 22706 21138
rect 22740 21104 22756 21138
rect 22808 21104 22824 21138
rect 22858 21104 22874 21138
rect 25383 21105 25417 21121
rect 25501 21297 25535 21313
rect 25501 21105 25535 21121
rect 25619 21297 25653 21313
rect 25619 21105 25653 21121
rect 25737 21297 25771 21313
rect 25737 21105 25771 21121
rect 25902 21297 25936 21313
rect 25902 21105 25936 21121
rect 26020 21297 26054 21313
rect 26020 21105 26054 21121
rect 26138 21297 26172 21313
rect 26138 21105 26172 21121
rect 26256 21297 26290 21313
rect 26256 21105 26290 21121
rect 26525 21293 26559 21309
rect 26525 21101 26559 21117
rect 26643 21293 26677 21309
rect 26643 21101 26677 21117
rect 26761 21293 26795 21309
rect 26761 21101 26795 21117
rect 26879 21293 26913 21309
rect 26879 21101 26913 21117
rect 27044 21293 27078 21309
rect 27044 21101 27078 21117
rect 27162 21293 27196 21309
rect 27162 21101 27196 21117
rect 27280 21293 27314 21309
rect 27280 21101 27314 21117
rect 27398 21293 27432 21309
rect 27398 21101 27432 21117
rect 28658 21241 28907 21284
rect 28658 21151 28697 21241
rect 28860 21151 28907 21241
rect 29160 21175 29194 21191
rect 29278 21567 29312 21583
rect 29278 21175 29312 21191
rect 29396 21567 29430 21583
rect 29396 21175 29430 21191
rect 28658 21112 28907 21151
rect 29203 21107 29219 21141
rect 29253 21107 29269 21141
rect 29321 21107 29337 21141
rect 29371 21107 29387 21141
rect 6498 20864 6670 20911
rect 6498 20701 6541 20864
rect 6631 20701 6670 20864
rect 6498 20662 6670 20701
rect 7640 20866 7812 20913
rect 7640 20703 7683 20866
rect 7773 20703 7812 20866
rect 13056 20860 13228 20907
rect 7640 20664 7812 20703
rect 9430 20764 9653 20840
rect 9430 20615 9507 20764
rect 9574 20615 9653 20764
rect 9430 20509 9653 20615
rect 10699 20658 10988 20705
rect 13056 20697 13099 20860
rect 13189 20697 13228 20860
rect 13056 20658 13228 20697
rect 14198 20862 14370 20909
rect 14198 20699 14241 20862
rect 14331 20699 14370 20862
rect 19590 20865 19762 20912
rect 14198 20660 14370 20699
rect 15988 20760 16211 20836
rect 10699 20549 10738 20658
rect 10849 20549 10988 20658
rect 10699 20537 10988 20549
rect 5717 20421 5942 20497
rect 5717 20272 5796 20421
rect 5863 20272 5942 20421
rect 5717 20166 5942 20272
rect 8952 20400 9222 20434
rect 8952 20350 8986 20400
rect 8952 20158 8986 20174
rect 9070 20350 9104 20366
rect 9070 20158 9104 20174
rect 9188 20350 9222 20400
rect 9188 20158 9222 20174
rect 9306 20350 9340 20366
rect 9306 20158 9340 20174
rect 9424 20350 9458 20366
rect 9424 20158 9458 20174
rect 9542 20350 9576 20366
rect 9542 20158 9576 20174
rect 9660 20350 9694 20366
rect 9660 20158 9694 20174
rect 9778 20350 9812 20366
rect 9778 20158 9812 20174
rect 9896 20350 9930 20366
rect 9896 20158 9930 20174
rect 10014 20350 10048 20366
rect 10014 20158 10048 20174
rect 9231 20080 9247 20114
rect 9281 20080 9297 20114
rect 5578 19986 5848 20021
rect 5460 19933 5494 19949
rect 4977 19733 5011 19749
rect 4977 19541 5011 19557
rect 5095 19733 5129 19749
rect 5095 19541 5129 19557
rect 5213 19733 5247 19749
rect 5213 19541 5247 19557
rect 5331 19733 5365 19749
rect 5331 19541 5365 19557
rect 5460 19541 5494 19557
rect 5578 19933 5612 19986
rect 5578 19541 5612 19557
rect 5696 19933 5730 19949
rect 5696 19541 5730 19557
rect 5814 19933 5848 19986
rect 7476 19986 7746 20021
rect 5814 19541 5848 19557
rect 5932 19933 5966 19949
rect 5932 19541 5966 19557
rect 6050 19933 6084 19949
rect 6050 19541 6084 19557
rect 6168 19933 6202 19949
rect 7358 19933 7392 19949
rect 6416 19787 6686 19822
rect 6168 19541 6202 19557
rect 6298 19733 6332 19749
rect 6298 19541 6332 19557
rect 6416 19733 6450 19787
rect 6416 19541 6450 19557
rect 6534 19733 6568 19749
rect 6534 19541 6568 19557
rect 6652 19733 6686 19787
rect 6652 19541 6686 19557
rect 6875 19733 6909 19749
rect 6875 19541 6909 19557
rect 6993 19733 7027 19749
rect 6993 19541 7027 19557
rect 7111 19733 7145 19749
rect 7111 19541 7145 19557
rect 7229 19733 7263 19749
rect 7229 19541 7263 19557
rect 7358 19541 7392 19557
rect 7476 19933 7510 19986
rect 7476 19541 7510 19557
rect 7594 19933 7628 19949
rect 7594 19541 7628 19557
rect 7712 19933 7746 19986
rect 9349 19963 9365 19997
rect 9399 19963 9415 19997
rect 7712 19541 7746 19557
rect 7830 19933 7864 19949
rect 7830 19541 7864 19557
rect 7948 19933 7982 19949
rect 7948 19541 7982 19557
rect 8066 19933 8100 19949
rect 9306 19913 9340 19929
rect 8314 19787 8584 19822
rect 8066 19541 8100 19557
rect 8196 19733 8230 19749
rect 8196 19541 8230 19557
rect 8314 19733 8348 19787
rect 8314 19541 8348 19557
rect 8432 19733 8466 19749
rect 8432 19541 8466 19557
rect 8550 19733 8584 19787
rect 9306 19721 9340 19737
rect 9424 19913 9458 19929
rect 9424 19721 9458 19737
rect 9541 19913 9575 19929
rect 8550 19541 8584 19557
rect 9039 19587 9288 19630
rect 9039 19497 9078 19587
rect 9241 19497 9288 19587
rect 9541 19521 9575 19537
rect 9659 19913 9693 19929
rect 9659 19521 9693 19537
rect 9777 19913 9811 19929
rect 9777 19521 9811 19537
rect 9039 19458 9288 19497
rect 9584 19453 9600 19487
rect 9634 19453 9650 19487
rect 9702 19453 9718 19487
rect 9752 19453 9768 19487
rect 7086 19319 7120 19335
rect 4963 19298 5030 19314
rect 4963 19264 4979 19298
rect 5013 19264 5030 19298
rect 7086 19269 7120 19285
rect 4963 19248 5030 19264
rect 5517 19240 5551 19256
rect 5635 19240 5669 19256
rect 5517 18848 5551 18864
rect 5633 18864 5635 18910
rect 4946 18835 5046 18836
rect 4890 18806 5046 18835
rect 5633 18806 5669 18864
rect 5753 19240 5787 19256
rect 5753 18848 5787 18864
rect 5871 19240 5905 19256
rect 5989 19240 6023 19256
rect 5905 18864 5907 18911
rect 5871 18806 5907 18864
rect 6107 19240 6141 19256
rect 5989 18848 6023 18864
rect 6106 18864 6107 18911
rect 6225 19240 6259 19256
rect 6141 18864 6142 18911
rect 6106 18806 6142 18864
rect 6225 18848 6259 18864
rect 7415 19240 7449 19256
rect 7533 19240 7567 19256
rect 7415 18848 7449 18864
rect 7531 18864 7533 18910
rect 4890 18766 6142 18806
rect 6447 18806 6944 18824
rect 7531 18806 7567 18864
rect 7651 19240 7685 19256
rect 7651 18848 7685 18864
rect 7769 19240 7803 19256
rect 7887 19240 7921 19256
rect 7803 18864 7805 18911
rect 7769 18806 7805 18864
rect 8005 19240 8039 19256
rect 7887 18848 7921 18864
rect 8004 18864 8005 18911
rect 8123 19240 8157 19256
rect 8039 18864 8040 18911
rect 8004 18806 8040 18864
rect 9435 19160 9658 19236
rect 9435 19011 9512 19160
rect 9579 19011 9658 19160
rect 9435 18905 9658 19011
rect 8123 18848 8157 18864
rect 6447 18803 8040 18806
rect 6447 18769 6465 18803
rect 6499 18769 8040 18803
rect 6447 18766 8040 18769
rect 8957 18796 9227 18830
rect 4890 18765 6123 18766
rect 6447 18765 8021 18766
rect 4890 18737 5046 18765
rect 4946 18736 5046 18737
rect 5533 18677 5600 18693
rect 5533 18643 5549 18677
rect 5583 18643 5600 18677
rect 5533 18627 5600 18643
rect 5257 18608 5291 18624
rect 5257 18558 5291 18574
rect 5795 18559 5811 18593
rect 5845 18559 5861 18593
rect 5913 18558 5929 18592
rect 5963 18558 5979 18592
rect 6034 18524 6068 18765
rect 6447 18748 6944 18765
rect 6178 18676 6245 18692
rect 6178 18642 6195 18676
rect 6229 18642 6245 18676
rect 6178 18626 6245 18642
rect 7429 18676 7496 18692
rect 7429 18642 7445 18676
rect 7479 18642 7496 18676
rect 7429 18626 7496 18642
rect 6380 18609 6414 18625
rect 6380 18559 6414 18575
rect 7155 18608 7189 18624
rect 7155 18558 7189 18574
rect 7693 18559 7709 18593
rect 7743 18559 7759 18593
rect 7811 18558 7827 18592
rect 7861 18558 7877 18592
rect 7932 18524 7966 18765
rect 8957 18746 8991 18796
rect 8076 18676 8143 18692
rect 8076 18642 8093 18676
rect 8127 18642 8143 18676
rect 8076 18626 8143 18642
rect 8278 18609 8312 18625
rect 8278 18559 8312 18575
rect 8957 18554 8991 18570
rect 9075 18746 9109 18762
rect 9075 18554 9109 18570
rect 9193 18746 9227 18796
rect 9193 18554 9227 18570
rect 9311 18746 9345 18762
rect 9311 18554 9345 18570
rect 9429 18746 9463 18762
rect 9429 18554 9463 18570
rect 9547 18746 9581 18762
rect 9547 18554 9581 18570
rect 9665 18746 9699 18762
rect 9665 18554 9699 18570
rect 9783 18746 9817 18762
rect 9783 18554 9817 18570
rect 9901 18746 9935 18762
rect 9901 18554 9935 18570
rect 10019 18746 10053 18762
rect 10019 18554 10053 18570
rect 5111 18508 5145 18524
rect 5111 18316 5145 18332
rect 5229 18508 5263 18524
rect 5229 18316 5263 18332
rect 5635 18508 5669 18524
rect 5753 18508 5787 18524
rect 5635 18065 5670 18132
rect 5753 18116 5787 18132
rect 5871 18508 5905 18524
rect 5871 18116 5905 18132
rect 5989 18508 6068 18524
rect 6023 18478 6068 18508
rect 6107 18508 6141 18524
rect 6409 18508 6443 18524
rect 6409 18316 6443 18332
rect 6527 18508 6561 18524
rect 6527 18316 6561 18332
rect 7009 18508 7043 18524
rect 7009 18316 7043 18332
rect 7127 18508 7161 18524
rect 7127 18316 7161 18332
rect 7533 18508 7567 18524
rect 5989 18116 6023 18132
rect 6106 18065 6141 18132
rect 5635 18030 6141 18065
rect 7651 18508 7685 18524
rect 7533 18065 7568 18132
rect 7651 18116 7685 18132
rect 7769 18508 7803 18524
rect 7769 18116 7803 18132
rect 7887 18508 7966 18524
rect 7921 18478 7966 18508
rect 8005 18508 8039 18524
rect 8307 18508 8341 18524
rect 8307 18316 8341 18332
rect 8425 18508 8459 18524
rect 9236 18476 9252 18510
rect 9286 18476 9302 18510
rect 9354 18359 9370 18393
rect 9404 18359 9420 18393
rect 8425 18316 8459 18332
rect 7887 18116 7921 18132
rect 8004 18065 8039 18132
rect 9311 18309 9345 18325
rect 9311 18117 9345 18133
rect 9429 18309 9463 18325
rect 9429 18117 9463 18133
rect 9546 18309 9580 18325
rect 7533 18030 8039 18065
rect 9044 17983 9293 18026
rect 9044 17893 9083 17983
rect 9246 17893 9293 17983
rect 9546 17917 9580 17933
rect 9664 18309 9698 18325
rect 9664 17917 9698 17933
rect 9782 18309 9816 18325
rect 9782 17917 9816 17933
rect 7696 17823 7868 17870
rect 9044 17854 9293 17893
rect 9589 17849 9605 17883
rect 9639 17849 9655 17883
rect 9707 17849 9723 17883
rect 9757 17849 9773 17883
rect 7696 17660 7739 17823
rect 7829 17660 7868 17823
rect 7696 17620 7868 17660
rect 10851 15790 10988 20537
rect 15988 20611 16065 20760
rect 16132 20611 16211 20760
rect 15988 20505 16211 20611
rect 17255 20646 17552 20704
rect 19590 20702 19633 20865
rect 19723 20702 19762 20865
rect 19590 20663 19762 20702
rect 20732 20867 20904 20914
rect 20732 20704 20775 20867
rect 20865 20704 20904 20867
rect 26103 20868 26275 20915
rect 20732 20665 20904 20704
rect 22522 20765 22745 20841
rect 17255 20549 17301 20646
rect 17404 20549 17552 20646
rect 17255 20533 17552 20549
rect 12275 20417 12500 20493
rect 12275 20268 12354 20417
rect 12421 20268 12500 20417
rect 12275 20162 12500 20268
rect 15510 20396 15780 20430
rect 15510 20346 15544 20396
rect 15510 20154 15544 20170
rect 15628 20346 15662 20362
rect 15628 20154 15662 20170
rect 15746 20346 15780 20396
rect 15746 20154 15780 20170
rect 15864 20346 15898 20362
rect 15864 20154 15898 20170
rect 15982 20346 16016 20362
rect 15982 20154 16016 20170
rect 16100 20346 16134 20362
rect 16100 20154 16134 20170
rect 16218 20346 16252 20362
rect 16218 20154 16252 20170
rect 16336 20346 16370 20362
rect 16336 20154 16370 20170
rect 16454 20346 16488 20362
rect 16454 20154 16488 20170
rect 16572 20346 16606 20362
rect 16572 20154 16606 20170
rect 15789 20076 15805 20110
rect 15839 20076 15855 20110
rect 12136 19982 12406 20017
rect 12018 19929 12052 19945
rect 11535 19729 11569 19745
rect 11535 19537 11569 19553
rect 11653 19729 11687 19745
rect 11653 19537 11687 19553
rect 11771 19729 11805 19745
rect 11771 19537 11805 19553
rect 11889 19729 11923 19745
rect 11889 19537 11923 19553
rect 12018 19537 12052 19553
rect 12136 19929 12170 19982
rect 12136 19537 12170 19553
rect 12254 19929 12288 19945
rect 12254 19537 12288 19553
rect 12372 19929 12406 19982
rect 14034 19982 14304 20017
rect 12372 19537 12406 19553
rect 12490 19929 12524 19945
rect 12490 19537 12524 19553
rect 12608 19929 12642 19945
rect 12608 19537 12642 19553
rect 12726 19929 12760 19945
rect 13916 19929 13950 19945
rect 12974 19783 13244 19818
rect 12726 19537 12760 19553
rect 12856 19729 12890 19745
rect 12856 19537 12890 19553
rect 12974 19729 13008 19783
rect 12974 19537 13008 19553
rect 13092 19729 13126 19745
rect 13092 19537 13126 19553
rect 13210 19729 13244 19783
rect 13210 19537 13244 19553
rect 13433 19729 13467 19745
rect 13433 19537 13467 19553
rect 13551 19729 13585 19745
rect 13551 19537 13585 19553
rect 13669 19729 13703 19745
rect 13669 19537 13703 19553
rect 13787 19729 13821 19745
rect 13787 19537 13821 19553
rect 13916 19537 13950 19553
rect 14034 19929 14068 19982
rect 14034 19537 14068 19553
rect 14152 19929 14186 19945
rect 14152 19537 14186 19553
rect 14270 19929 14304 19982
rect 15907 19959 15923 19993
rect 15957 19959 15973 19993
rect 14270 19537 14304 19553
rect 14388 19929 14422 19945
rect 14388 19537 14422 19553
rect 14506 19929 14540 19945
rect 14506 19537 14540 19553
rect 14624 19929 14658 19945
rect 15864 19909 15898 19925
rect 14872 19783 15142 19818
rect 14624 19537 14658 19553
rect 14754 19729 14788 19745
rect 14754 19537 14788 19553
rect 14872 19729 14906 19783
rect 14872 19537 14906 19553
rect 14990 19729 15024 19745
rect 14990 19537 15024 19553
rect 15108 19729 15142 19783
rect 15864 19717 15898 19733
rect 15982 19909 16016 19925
rect 15982 19717 16016 19733
rect 16099 19909 16133 19925
rect 15108 19537 15142 19553
rect 15597 19583 15846 19626
rect 15597 19493 15636 19583
rect 15799 19493 15846 19583
rect 16099 19517 16133 19533
rect 16217 19909 16251 19925
rect 16217 19517 16251 19533
rect 16335 19909 16369 19925
rect 16335 19517 16369 19533
rect 15597 19454 15846 19493
rect 16142 19449 16158 19483
rect 16192 19449 16208 19483
rect 16260 19449 16276 19483
rect 16310 19449 16326 19483
rect 13644 19315 13678 19331
rect 11521 19294 11588 19310
rect 11521 19260 11537 19294
rect 11571 19260 11588 19294
rect 13644 19265 13678 19281
rect 11521 19244 11588 19260
rect 12075 19236 12109 19252
rect 12193 19236 12227 19252
rect 12075 18844 12109 18860
rect 12191 18860 12193 18906
rect 11504 18831 11604 18832
rect 11448 18802 11604 18831
rect 12191 18802 12227 18860
rect 12311 19236 12345 19252
rect 12311 18844 12345 18860
rect 12429 19236 12463 19252
rect 12547 19236 12581 19252
rect 12463 18860 12465 18907
rect 12429 18802 12465 18860
rect 12665 19236 12699 19252
rect 12547 18844 12581 18860
rect 12664 18860 12665 18907
rect 12783 19236 12817 19252
rect 12699 18860 12700 18907
rect 12664 18802 12700 18860
rect 12783 18844 12817 18860
rect 13973 19236 14007 19252
rect 14091 19236 14125 19252
rect 13973 18844 14007 18860
rect 14089 18860 14091 18906
rect 11448 18762 12700 18802
rect 13005 18802 13502 18820
rect 14089 18802 14125 18860
rect 14209 19236 14243 19252
rect 14209 18844 14243 18860
rect 14327 19236 14361 19252
rect 14445 19236 14479 19252
rect 14361 18860 14363 18907
rect 14327 18802 14363 18860
rect 14563 19236 14597 19252
rect 14445 18844 14479 18860
rect 14562 18860 14563 18907
rect 14681 19236 14715 19252
rect 14597 18860 14598 18907
rect 14562 18802 14598 18860
rect 15993 19156 16216 19232
rect 15993 19007 16070 19156
rect 16137 19007 16216 19156
rect 15993 18901 16216 19007
rect 14681 18844 14715 18860
rect 13005 18799 14598 18802
rect 13005 18765 13023 18799
rect 13057 18765 14598 18799
rect 13005 18762 14598 18765
rect 15515 18792 15785 18826
rect 11448 18761 12681 18762
rect 13005 18761 14579 18762
rect 11448 18733 11604 18761
rect 11504 18732 11604 18733
rect 12091 18673 12158 18689
rect 12091 18639 12107 18673
rect 12141 18639 12158 18673
rect 12091 18623 12158 18639
rect 11815 18604 11849 18620
rect 11815 18554 11849 18570
rect 12353 18555 12369 18589
rect 12403 18555 12419 18589
rect 12471 18554 12487 18588
rect 12521 18554 12537 18588
rect 12592 18520 12626 18761
rect 13005 18744 13502 18761
rect 12736 18672 12803 18688
rect 12736 18638 12753 18672
rect 12787 18638 12803 18672
rect 12736 18622 12803 18638
rect 13987 18672 14054 18688
rect 13987 18638 14003 18672
rect 14037 18638 14054 18672
rect 13987 18622 14054 18638
rect 12938 18605 12972 18621
rect 12938 18555 12972 18571
rect 13713 18604 13747 18620
rect 13713 18554 13747 18570
rect 14251 18555 14267 18589
rect 14301 18555 14317 18589
rect 14369 18554 14385 18588
rect 14419 18554 14435 18588
rect 14490 18520 14524 18761
rect 15515 18742 15549 18792
rect 14634 18672 14701 18688
rect 14634 18638 14651 18672
rect 14685 18638 14701 18672
rect 14634 18622 14701 18638
rect 14836 18605 14870 18621
rect 14836 18555 14870 18571
rect 15515 18550 15549 18566
rect 15633 18742 15667 18758
rect 15633 18550 15667 18566
rect 15751 18742 15785 18792
rect 15751 18550 15785 18566
rect 15869 18742 15903 18758
rect 15869 18550 15903 18566
rect 15987 18742 16021 18758
rect 15987 18550 16021 18566
rect 16105 18742 16139 18758
rect 16105 18550 16139 18566
rect 16223 18742 16257 18758
rect 16223 18550 16257 18566
rect 16341 18742 16375 18758
rect 16341 18550 16375 18566
rect 16459 18742 16493 18758
rect 16459 18550 16493 18566
rect 16577 18742 16611 18758
rect 16577 18550 16611 18566
rect 11669 18504 11703 18520
rect 11669 18312 11703 18328
rect 11787 18504 11821 18520
rect 11787 18312 11821 18328
rect 12193 18504 12227 18520
rect 12311 18504 12345 18520
rect 12193 18061 12228 18128
rect 12311 18112 12345 18128
rect 12429 18504 12463 18520
rect 12429 18112 12463 18128
rect 12547 18504 12626 18520
rect 12581 18474 12626 18504
rect 12665 18504 12699 18520
rect 12967 18504 13001 18520
rect 12967 18312 13001 18328
rect 13085 18504 13119 18520
rect 13085 18312 13119 18328
rect 13567 18504 13601 18520
rect 13567 18312 13601 18328
rect 13685 18504 13719 18520
rect 13685 18312 13719 18328
rect 14091 18504 14125 18520
rect 12547 18112 12581 18128
rect 12664 18061 12699 18128
rect 12193 18026 12699 18061
rect 14209 18504 14243 18520
rect 14091 18061 14126 18128
rect 14209 18112 14243 18128
rect 14327 18504 14361 18520
rect 14327 18112 14361 18128
rect 14445 18504 14524 18520
rect 14479 18474 14524 18504
rect 14563 18504 14597 18520
rect 14865 18504 14899 18520
rect 14865 18312 14899 18328
rect 14983 18504 15017 18520
rect 15794 18472 15810 18506
rect 15844 18472 15860 18506
rect 15912 18355 15928 18389
rect 15962 18355 15978 18389
rect 14983 18312 15017 18328
rect 14445 18112 14479 18128
rect 14562 18061 14597 18128
rect 15869 18305 15903 18321
rect 15869 18113 15903 18129
rect 15987 18305 16021 18321
rect 15987 18113 16021 18129
rect 16104 18305 16138 18321
rect 14091 18026 14597 18061
rect 15602 17979 15851 18022
rect 15602 17889 15641 17979
rect 15804 17889 15851 17979
rect 16104 17913 16138 17929
rect 16222 18305 16256 18321
rect 16222 17913 16256 17929
rect 16340 18305 16374 18321
rect 16340 17913 16374 17929
rect 14254 17819 14426 17866
rect 15602 17850 15851 17889
rect 16147 17845 16163 17879
rect 16197 17845 16213 17879
rect 16265 17845 16281 17879
rect 16315 17845 16331 17879
rect 14254 17656 14297 17819
rect 14387 17656 14426 17819
rect 14254 17616 14426 17656
rect 17431 16123 17552 20533
rect 22522 20616 22599 20765
rect 22666 20616 22745 20765
rect 26103 20705 26146 20868
rect 26236 20705 26275 20868
rect 22522 20510 22745 20616
rect 23789 20650 24075 20704
rect 26103 20666 26275 20705
rect 27245 20870 27417 20917
rect 27245 20707 27288 20870
rect 27378 20707 27417 20870
rect 27245 20668 27417 20707
rect 29035 20768 29258 20844
rect 23789 20558 23837 20650
rect 23935 20558 24075 20650
rect 23789 20539 24075 20558
rect 18809 20422 19034 20498
rect 18809 20273 18888 20422
rect 18955 20273 19034 20422
rect 18809 20167 19034 20273
rect 22044 20401 22314 20435
rect 22044 20351 22078 20401
rect 22044 20159 22078 20175
rect 22162 20351 22196 20367
rect 22162 20159 22196 20175
rect 22280 20351 22314 20401
rect 22280 20159 22314 20175
rect 22398 20351 22432 20367
rect 22398 20159 22432 20175
rect 22516 20351 22550 20367
rect 22516 20159 22550 20175
rect 22634 20351 22668 20367
rect 22634 20159 22668 20175
rect 22752 20351 22786 20367
rect 22752 20159 22786 20175
rect 22870 20351 22904 20367
rect 22870 20159 22904 20175
rect 22988 20351 23022 20367
rect 22988 20159 23022 20175
rect 23106 20351 23140 20367
rect 23106 20159 23140 20175
rect 22323 20081 22339 20115
rect 22373 20081 22389 20115
rect 18670 19987 18940 20022
rect 18552 19934 18586 19950
rect 18069 19734 18103 19750
rect 18069 19542 18103 19558
rect 18187 19734 18221 19750
rect 18187 19542 18221 19558
rect 18305 19734 18339 19750
rect 18305 19542 18339 19558
rect 18423 19734 18457 19750
rect 18423 19542 18457 19558
rect 18552 19542 18586 19558
rect 18670 19934 18704 19987
rect 18670 19542 18704 19558
rect 18788 19934 18822 19950
rect 18788 19542 18822 19558
rect 18906 19934 18940 19987
rect 20568 19987 20838 20022
rect 18906 19542 18940 19558
rect 19024 19934 19058 19950
rect 19024 19542 19058 19558
rect 19142 19934 19176 19950
rect 19142 19542 19176 19558
rect 19260 19934 19294 19950
rect 20450 19934 20484 19950
rect 19508 19788 19778 19823
rect 19260 19542 19294 19558
rect 19390 19734 19424 19750
rect 19390 19542 19424 19558
rect 19508 19734 19542 19788
rect 19508 19542 19542 19558
rect 19626 19734 19660 19750
rect 19626 19542 19660 19558
rect 19744 19734 19778 19788
rect 19744 19542 19778 19558
rect 19967 19734 20001 19750
rect 19967 19542 20001 19558
rect 20085 19734 20119 19750
rect 20085 19542 20119 19558
rect 20203 19734 20237 19750
rect 20203 19542 20237 19558
rect 20321 19734 20355 19750
rect 20321 19542 20355 19558
rect 20450 19542 20484 19558
rect 20568 19934 20602 19987
rect 20568 19542 20602 19558
rect 20686 19934 20720 19950
rect 20686 19542 20720 19558
rect 20804 19934 20838 19987
rect 22441 19964 22457 19998
rect 22491 19964 22507 19998
rect 20804 19542 20838 19558
rect 20922 19934 20956 19950
rect 20922 19542 20956 19558
rect 21040 19934 21074 19950
rect 21040 19542 21074 19558
rect 21158 19934 21192 19950
rect 22398 19914 22432 19930
rect 21406 19788 21676 19823
rect 21158 19542 21192 19558
rect 21288 19734 21322 19750
rect 21288 19542 21322 19558
rect 21406 19734 21440 19788
rect 21406 19542 21440 19558
rect 21524 19734 21558 19750
rect 21524 19542 21558 19558
rect 21642 19734 21676 19788
rect 22398 19722 22432 19738
rect 22516 19914 22550 19930
rect 22516 19722 22550 19738
rect 22633 19914 22667 19930
rect 21642 19542 21676 19558
rect 22131 19588 22380 19631
rect 22131 19498 22170 19588
rect 22333 19498 22380 19588
rect 22633 19522 22667 19538
rect 22751 19914 22785 19930
rect 22751 19522 22785 19538
rect 22869 19914 22903 19930
rect 22869 19522 22903 19538
rect 22131 19459 22380 19498
rect 22676 19454 22692 19488
rect 22726 19454 22742 19488
rect 22794 19454 22810 19488
rect 22844 19454 22860 19488
rect 20178 19320 20212 19336
rect 18055 19299 18122 19315
rect 18055 19265 18071 19299
rect 18105 19265 18122 19299
rect 20178 19270 20212 19286
rect 18055 19249 18122 19265
rect 18609 19241 18643 19257
rect 18727 19241 18761 19257
rect 18609 18849 18643 18865
rect 18725 18865 18727 18911
rect 18038 18836 18138 18837
rect 17982 18807 18138 18836
rect 18725 18807 18761 18865
rect 18845 19241 18879 19257
rect 18845 18849 18879 18865
rect 18963 19241 18997 19257
rect 19081 19241 19115 19257
rect 18997 18865 18999 18912
rect 18963 18807 18999 18865
rect 19199 19241 19233 19257
rect 19081 18849 19115 18865
rect 19198 18865 19199 18912
rect 19317 19241 19351 19257
rect 19233 18865 19234 18912
rect 19198 18807 19234 18865
rect 19317 18849 19351 18865
rect 20507 19241 20541 19257
rect 20625 19241 20659 19257
rect 20507 18849 20541 18865
rect 20623 18865 20625 18911
rect 17982 18767 19234 18807
rect 19539 18807 20036 18825
rect 20623 18807 20659 18865
rect 20743 19241 20777 19257
rect 20743 18849 20777 18865
rect 20861 19241 20895 19257
rect 20979 19241 21013 19257
rect 20895 18865 20897 18912
rect 20861 18807 20897 18865
rect 21097 19241 21131 19257
rect 20979 18849 21013 18865
rect 21096 18865 21097 18912
rect 21215 19241 21249 19257
rect 21131 18865 21132 18912
rect 21096 18807 21132 18865
rect 22527 19161 22750 19237
rect 22527 19012 22604 19161
rect 22671 19012 22750 19161
rect 22527 18906 22750 19012
rect 21215 18849 21249 18865
rect 19539 18804 21132 18807
rect 19539 18770 19557 18804
rect 19591 18770 21132 18804
rect 19539 18767 21132 18770
rect 22049 18797 22319 18831
rect 17982 18766 19215 18767
rect 19539 18766 21113 18767
rect 17982 18738 18138 18766
rect 18038 18737 18138 18738
rect 18625 18678 18692 18694
rect 18625 18644 18641 18678
rect 18675 18644 18692 18678
rect 18625 18628 18692 18644
rect 18349 18609 18383 18625
rect 18349 18559 18383 18575
rect 18887 18560 18903 18594
rect 18937 18560 18953 18594
rect 19005 18559 19021 18593
rect 19055 18559 19071 18593
rect 19126 18525 19160 18766
rect 19539 18749 20036 18766
rect 19270 18677 19337 18693
rect 19270 18643 19287 18677
rect 19321 18643 19337 18677
rect 19270 18627 19337 18643
rect 20521 18677 20588 18693
rect 20521 18643 20537 18677
rect 20571 18643 20588 18677
rect 20521 18627 20588 18643
rect 19472 18610 19506 18626
rect 19472 18560 19506 18576
rect 20247 18609 20281 18625
rect 20247 18559 20281 18575
rect 20785 18560 20801 18594
rect 20835 18560 20851 18594
rect 20903 18559 20919 18593
rect 20953 18559 20969 18593
rect 21024 18525 21058 18766
rect 22049 18747 22083 18797
rect 21168 18677 21235 18693
rect 21168 18643 21185 18677
rect 21219 18643 21235 18677
rect 21168 18627 21235 18643
rect 21370 18610 21404 18626
rect 21370 18560 21404 18576
rect 22049 18555 22083 18571
rect 22167 18747 22201 18763
rect 22167 18555 22201 18571
rect 22285 18747 22319 18797
rect 22285 18555 22319 18571
rect 22403 18747 22437 18763
rect 22403 18555 22437 18571
rect 22521 18747 22555 18763
rect 22521 18555 22555 18571
rect 22639 18747 22673 18763
rect 22639 18555 22673 18571
rect 22757 18747 22791 18763
rect 22757 18555 22791 18571
rect 22875 18747 22909 18763
rect 22875 18555 22909 18571
rect 22993 18747 23027 18763
rect 22993 18555 23027 18571
rect 23111 18747 23145 18763
rect 23111 18555 23145 18571
rect 18203 18509 18237 18525
rect 18203 18317 18237 18333
rect 18321 18509 18355 18525
rect 18321 18317 18355 18333
rect 18727 18509 18761 18525
rect 18845 18509 18879 18525
rect 18727 18066 18762 18133
rect 18845 18117 18879 18133
rect 18963 18509 18997 18525
rect 18963 18117 18997 18133
rect 19081 18509 19160 18525
rect 19115 18479 19160 18509
rect 19199 18509 19233 18525
rect 19501 18509 19535 18525
rect 19501 18317 19535 18333
rect 19619 18509 19653 18525
rect 19619 18317 19653 18333
rect 20101 18509 20135 18525
rect 20101 18317 20135 18333
rect 20219 18509 20253 18525
rect 20219 18317 20253 18333
rect 20625 18509 20659 18525
rect 19081 18117 19115 18133
rect 19198 18066 19233 18133
rect 18727 18031 19233 18066
rect 20743 18509 20777 18525
rect 20625 18066 20660 18133
rect 20743 18117 20777 18133
rect 20861 18509 20895 18525
rect 20861 18117 20895 18133
rect 20979 18509 21058 18525
rect 21013 18479 21058 18509
rect 21097 18509 21131 18525
rect 21399 18509 21433 18525
rect 21399 18317 21433 18333
rect 21517 18509 21551 18525
rect 22328 18477 22344 18511
rect 22378 18477 22394 18511
rect 22446 18360 22462 18394
rect 22496 18360 22512 18394
rect 21517 18317 21551 18333
rect 20979 18117 21013 18133
rect 21096 18066 21131 18133
rect 22403 18310 22437 18326
rect 22403 18118 22437 18134
rect 22521 18310 22555 18326
rect 22521 18118 22555 18134
rect 22638 18310 22672 18326
rect 20625 18031 21131 18066
rect 22136 17984 22385 18027
rect 22136 17894 22175 17984
rect 22338 17894 22385 17984
rect 22638 17918 22672 17934
rect 22756 18310 22790 18326
rect 22756 17918 22790 17934
rect 22874 18310 22908 18326
rect 22874 17918 22908 17934
rect 20788 17824 20960 17871
rect 22136 17855 22385 17894
rect 22681 17850 22697 17884
rect 22731 17850 22747 17884
rect 22799 17850 22815 17884
rect 22849 17850 22865 17884
rect 20788 17661 20831 17824
rect 20921 17661 20960 17824
rect 20788 17621 20960 17661
rect 23951 16648 24075 20539
rect 29035 20619 29112 20768
rect 29179 20619 29258 20768
rect 29035 20513 29258 20619
rect 25322 20425 25547 20501
rect 25322 20276 25401 20425
rect 25468 20276 25547 20425
rect 25322 20170 25547 20276
rect 28557 20404 28827 20438
rect 28557 20354 28591 20404
rect 28557 20162 28591 20178
rect 28675 20354 28709 20370
rect 28675 20162 28709 20178
rect 28793 20354 28827 20404
rect 28793 20162 28827 20178
rect 28911 20354 28945 20370
rect 28911 20162 28945 20178
rect 29029 20354 29063 20370
rect 29029 20162 29063 20178
rect 29147 20354 29181 20370
rect 29147 20162 29181 20178
rect 29265 20354 29299 20370
rect 29265 20162 29299 20178
rect 29383 20354 29417 20370
rect 29383 20162 29417 20178
rect 29501 20354 29535 20370
rect 29501 20162 29535 20178
rect 29619 20354 29653 20370
rect 29619 20162 29653 20178
rect 28836 20084 28852 20118
rect 28886 20084 28902 20118
rect 25183 19990 25453 20025
rect 25065 19937 25099 19953
rect 24582 19737 24616 19753
rect 24582 19545 24616 19561
rect 24700 19737 24734 19753
rect 24700 19545 24734 19561
rect 24818 19737 24852 19753
rect 24818 19545 24852 19561
rect 24936 19737 24970 19753
rect 24936 19545 24970 19561
rect 25065 19545 25099 19561
rect 25183 19937 25217 19990
rect 25183 19545 25217 19561
rect 25301 19937 25335 19953
rect 25301 19545 25335 19561
rect 25419 19937 25453 19990
rect 27081 19990 27351 20025
rect 25419 19545 25453 19561
rect 25537 19937 25571 19953
rect 25537 19545 25571 19561
rect 25655 19937 25689 19953
rect 25655 19545 25689 19561
rect 25773 19937 25807 19953
rect 26963 19937 26997 19953
rect 26021 19791 26291 19826
rect 25773 19545 25807 19561
rect 25903 19737 25937 19753
rect 25903 19545 25937 19561
rect 26021 19737 26055 19791
rect 26021 19545 26055 19561
rect 26139 19737 26173 19753
rect 26139 19545 26173 19561
rect 26257 19737 26291 19791
rect 26257 19545 26291 19561
rect 26480 19737 26514 19753
rect 26480 19545 26514 19561
rect 26598 19737 26632 19753
rect 26598 19545 26632 19561
rect 26716 19737 26750 19753
rect 26716 19545 26750 19561
rect 26834 19737 26868 19753
rect 26834 19545 26868 19561
rect 26963 19545 26997 19561
rect 27081 19937 27115 19990
rect 27081 19545 27115 19561
rect 27199 19937 27233 19953
rect 27199 19545 27233 19561
rect 27317 19937 27351 19990
rect 28954 19967 28970 20001
rect 29004 19967 29020 20001
rect 27317 19545 27351 19561
rect 27435 19937 27469 19953
rect 27435 19545 27469 19561
rect 27553 19937 27587 19953
rect 27553 19545 27587 19561
rect 27671 19937 27705 19953
rect 28911 19917 28945 19933
rect 27919 19791 28189 19826
rect 27671 19545 27705 19561
rect 27801 19737 27835 19753
rect 27801 19545 27835 19561
rect 27919 19737 27953 19791
rect 27919 19545 27953 19561
rect 28037 19737 28071 19753
rect 28037 19545 28071 19561
rect 28155 19737 28189 19791
rect 28911 19725 28945 19741
rect 29029 19917 29063 19933
rect 29029 19725 29063 19741
rect 29146 19917 29180 19933
rect 28155 19545 28189 19561
rect 28644 19591 28893 19634
rect 28644 19501 28683 19591
rect 28846 19501 28893 19591
rect 29146 19525 29180 19541
rect 29264 19917 29298 19933
rect 29264 19525 29298 19541
rect 29382 19917 29416 19933
rect 29382 19525 29416 19541
rect 28644 19462 28893 19501
rect 29189 19457 29205 19491
rect 29239 19457 29255 19491
rect 29307 19457 29323 19491
rect 29357 19457 29373 19491
rect 26691 19323 26725 19339
rect 24568 19302 24635 19318
rect 24568 19268 24584 19302
rect 24618 19268 24635 19302
rect 26691 19273 26725 19289
rect 24568 19252 24635 19268
rect 25122 19244 25156 19260
rect 25240 19244 25274 19260
rect 25122 18852 25156 18868
rect 25238 18868 25240 18914
rect 24551 18839 24651 18840
rect 24495 18810 24651 18839
rect 25238 18810 25274 18868
rect 25358 19244 25392 19260
rect 25358 18852 25392 18868
rect 25476 19244 25510 19260
rect 25594 19244 25628 19260
rect 25510 18868 25512 18915
rect 25476 18810 25512 18868
rect 25712 19244 25746 19260
rect 25594 18852 25628 18868
rect 25711 18868 25712 18915
rect 25830 19244 25864 19260
rect 25746 18868 25747 18915
rect 25711 18810 25747 18868
rect 25830 18852 25864 18868
rect 27020 19244 27054 19260
rect 27138 19244 27172 19260
rect 27020 18852 27054 18868
rect 27136 18868 27138 18914
rect 24495 18770 25747 18810
rect 26052 18810 26549 18828
rect 27136 18810 27172 18868
rect 27256 19244 27290 19260
rect 27256 18852 27290 18868
rect 27374 19244 27408 19260
rect 27492 19244 27526 19260
rect 27408 18868 27410 18915
rect 27374 18810 27410 18868
rect 27610 19244 27644 19260
rect 27492 18852 27526 18868
rect 27609 18868 27610 18915
rect 27728 19244 27762 19260
rect 27644 18868 27645 18915
rect 27609 18810 27645 18868
rect 29040 19164 29263 19240
rect 29040 19015 29117 19164
rect 29184 19015 29263 19164
rect 29040 18909 29263 19015
rect 27728 18852 27762 18868
rect 26052 18807 27645 18810
rect 26052 18773 26070 18807
rect 26104 18773 27645 18807
rect 26052 18770 27645 18773
rect 28562 18800 28832 18834
rect 24495 18769 25728 18770
rect 26052 18769 27626 18770
rect 24495 18741 24651 18769
rect 24551 18740 24651 18741
rect 25138 18681 25205 18697
rect 25138 18647 25154 18681
rect 25188 18647 25205 18681
rect 25138 18631 25205 18647
rect 24862 18612 24896 18628
rect 24862 18562 24896 18578
rect 25400 18563 25416 18597
rect 25450 18563 25466 18597
rect 25518 18562 25534 18596
rect 25568 18562 25584 18596
rect 25639 18528 25673 18769
rect 26052 18752 26549 18769
rect 25783 18680 25850 18696
rect 25783 18646 25800 18680
rect 25834 18646 25850 18680
rect 25783 18630 25850 18646
rect 27034 18680 27101 18696
rect 27034 18646 27050 18680
rect 27084 18646 27101 18680
rect 27034 18630 27101 18646
rect 25985 18613 26019 18629
rect 25985 18563 26019 18579
rect 26760 18612 26794 18628
rect 26760 18562 26794 18578
rect 27298 18563 27314 18597
rect 27348 18563 27364 18597
rect 27416 18562 27432 18596
rect 27466 18562 27482 18596
rect 27537 18528 27571 18769
rect 28562 18750 28596 18800
rect 27681 18680 27748 18696
rect 27681 18646 27698 18680
rect 27732 18646 27748 18680
rect 27681 18630 27748 18646
rect 27883 18613 27917 18629
rect 27883 18563 27917 18579
rect 28562 18558 28596 18574
rect 28680 18750 28714 18766
rect 28680 18558 28714 18574
rect 28798 18750 28832 18800
rect 28798 18558 28832 18574
rect 28916 18750 28950 18766
rect 28916 18558 28950 18574
rect 29034 18750 29068 18766
rect 29034 18558 29068 18574
rect 29152 18750 29186 18766
rect 29152 18558 29186 18574
rect 29270 18750 29304 18766
rect 29270 18558 29304 18574
rect 29388 18750 29422 18766
rect 29388 18558 29422 18574
rect 29506 18750 29540 18766
rect 29506 18558 29540 18574
rect 29624 18750 29658 18766
rect 29624 18558 29658 18574
rect 24716 18512 24750 18528
rect 24716 18320 24750 18336
rect 24834 18512 24868 18528
rect 24834 18320 24868 18336
rect 25240 18512 25274 18528
rect 25358 18512 25392 18528
rect 25240 18069 25275 18136
rect 25358 18120 25392 18136
rect 25476 18512 25510 18528
rect 25476 18120 25510 18136
rect 25594 18512 25673 18528
rect 25628 18482 25673 18512
rect 25712 18512 25746 18528
rect 26014 18512 26048 18528
rect 26014 18320 26048 18336
rect 26132 18512 26166 18528
rect 26132 18320 26166 18336
rect 26614 18512 26648 18528
rect 26614 18320 26648 18336
rect 26732 18512 26766 18528
rect 26732 18320 26766 18336
rect 27138 18512 27172 18528
rect 25594 18120 25628 18136
rect 25711 18069 25746 18136
rect 25240 18034 25746 18069
rect 27256 18512 27290 18528
rect 27138 18069 27173 18136
rect 27256 18120 27290 18136
rect 27374 18512 27408 18528
rect 27374 18120 27408 18136
rect 27492 18512 27571 18528
rect 27526 18482 27571 18512
rect 27610 18512 27644 18528
rect 27912 18512 27946 18528
rect 27912 18320 27946 18336
rect 28030 18512 28064 18528
rect 28841 18480 28857 18514
rect 28891 18480 28907 18514
rect 28959 18363 28975 18397
rect 29009 18363 29025 18397
rect 28030 18320 28064 18336
rect 27492 18120 27526 18136
rect 27609 18069 27644 18136
rect 28916 18313 28950 18329
rect 28916 18121 28950 18137
rect 29034 18313 29068 18329
rect 29034 18121 29068 18137
rect 29151 18313 29185 18329
rect 27138 18034 27644 18069
rect 28649 17987 28898 18030
rect 28649 17897 28688 17987
rect 28851 17897 28898 17987
rect 29151 17921 29185 17937
rect 29269 18313 29303 18329
rect 29269 17921 29303 17937
rect 29387 18313 29421 18329
rect 29387 17921 29421 17937
rect 27301 17827 27473 17874
rect 28649 17858 28898 17897
rect 29194 17853 29210 17887
rect 29244 17853 29260 17887
rect 29312 17853 29328 17887
rect 29362 17853 29378 17887
rect 27301 17664 27344 17827
rect 27434 17664 27473 17827
rect 27301 17624 27473 17664
rect 23950 16242 24076 16648
rect 23950 16184 23984 16242
rect 24052 16184 24076 16242
rect 23950 16153 24076 16184
rect 17431 16067 17459 16123
rect 17530 16067 17552 16123
rect 17431 16041 17552 16067
rect 30844 16012 30942 22445
rect 34475 22236 37815 22257
rect 34475 22173 34502 22236
rect 34551 22173 37815 22236
rect 34475 22171 37815 22173
rect 37728 22143 37815 22171
rect 37728 22094 37741 22143
rect 37801 22094 37815 22143
rect 37728 22072 37815 22094
rect 36877 21970 36967 22004
rect 37143 21970 37159 22004
rect 36877 21768 36916 21970
rect 37441 21899 37526 21915
rect 36951 21852 36967 21886
rect 37143 21852 37233 21886
rect 36877 21734 36967 21768
rect 37143 21734 37159 21768
rect 37194 21650 37233 21852
rect 37441 21839 37458 21899
rect 37513 21839 37526 21899
rect 37441 21823 37526 21839
rect 36951 21616 36967 21650
rect 37143 21616 37233 21650
rect 36675 21529 36767 21563
rect 37143 21529 37159 21563
rect 36675 21327 36714 21529
rect 36751 21411 36767 21445
rect 37143 21411 37233 21445
rect 36675 21293 36767 21327
rect 37143 21293 37159 21327
rect 37194 21209 37233 21411
rect 36751 21175 36767 21209
rect 37143 21175 37233 21209
rect 36676 21062 36767 21096
rect 37143 21062 37159 21096
rect 36676 20860 36715 21062
rect 37194 20978 37233 21175
rect 38084 21136 38100 21170
rect 38276 21136 38292 21170
rect 38084 21018 38100 21052
rect 38276 21018 38292 21052
rect 38088 20978 38288 21018
rect 36751 20944 36767 20978
rect 37143 20944 37233 20978
rect 36479 20818 36589 20834
rect 36676 20826 36767 20860
rect 37143 20826 37159 20860
rect 36479 20622 36497 20818
rect 36573 20622 36589 20818
rect 37194 20742 37233 20944
rect 37729 20932 37814 20948
rect 38084 20944 38100 20978
rect 38476 20944 38492 20978
rect 37342 20884 37358 20918
rect 37392 20884 37408 20918
rect 37729 20872 37742 20932
rect 37797 20872 37814 20932
rect 37729 20856 37814 20872
rect 36751 20708 36767 20742
rect 37143 20708 37233 20742
rect 37444 20814 37529 20830
rect 38084 20826 38100 20860
rect 38476 20826 38492 20860
rect 37444 20754 37457 20814
rect 37512 20754 37529 20814
rect 38725 20760 38811 20776
rect 37444 20738 37529 20754
rect 38084 20708 38100 20742
rect 38476 20708 38492 20742
rect 38577 20741 38611 20757
rect 36479 20606 36589 20622
rect 36676 20590 36767 20624
rect 37143 20590 37159 20624
rect 36676 20388 36715 20590
rect 37194 20506 37233 20708
rect 38577 20691 38611 20707
rect 38725 20738 38743 20760
rect 37962 20649 37978 20683
rect 38012 20649 38028 20683
rect 38725 20680 38729 20738
rect 38725 20656 38743 20680
rect 38789 20656 38811 20760
rect 38725 20640 38811 20656
rect 38084 20590 38100 20624
rect 38476 20590 38492 20624
rect 37572 20530 37588 20564
rect 37622 20530 37638 20564
rect 36751 20472 36767 20506
rect 37143 20472 37233 20506
rect 38084 20472 38100 20506
rect 38476 20472 38492 20506
rect 36676 20354 36767 20388
rect 37143 20354 37159 20388
rect 37194 20269 37233 20472
rect 38088 20428 38288 20472
rect 38084 20394 38100 20428
rect 38276 20394 38292 20428
rect 38084 20276 38100 20310
rect 38276 20276 38292 20310
rect 36751 20235 36767 20269
rect 37143 20235 37233 20269
rect 36676 20117 36767 20151
rect 37143 20117 37159 20151
rect 36676 19915 36715 20117
rect 37194 20033 37233 20235
rect 36751 19999 36767 20033
rect 37143 19999 37233 20033
rect 36676 19881 36767 19915
rect 37143 19881 37159 19915
rect 36951 19762 36967 19796
rect 37143 19762 37236 19796
rect 36880 19644 36967 19678
rect 37143 19644 37159 19678
rect 36880 19442 36917 19644
rect 37197 19560 37236 19762
rect 36951 19526 36967 19560
rect 37143 19526 37236 19560
rect 37317 19608 37351 19624
rect 37317 19558 37351 19574
rect 36880 19408 36967 19442
rect 37143 19408 37159 19442
rect 34779 19035 37812 19116
rect 10851 15745 10883 15790
rect 10962 15745 10988 15790
rect 10851 15722 10988 15745
rect 21304 15484 21472 15500
rect 8101 15464 8269 15480
rect 8101 15394 8117 15464
rect 8253 15394 8269 15464
rect 8101 15378 8269 15394
rect 14650 15463 14818 15479
rect 14650 15393 14666 15463
rect 14802 15393 14818 15463
rect 21304 15414 21320 15484
rect 21456 15414 21472 15484
rect 21304 15398 21472 15414
rect 30846 15452 30940 16012
rect 14650 15377 14818 15393
rect 30846 15380 30852 15452
rect 30930 15380 30940 15452
rect 30846 15375 30940 15380
rect 32099 15410 32543 15416
rect 8638 15274 8908 15308
rect 7812 15224 7846 15240
rect 7812 15032 7846 15048
rect 7930 15224 7964 15240
rect 7930 15032 7964 15048
rect 8048 15224 8082 15240
rect 8048 15032 8082 15048
rect 8166 15224 8200 15240
rect 8166 15032 8200 15048
rect 8284 15224 8318 15240
rect 8284 15032 8318 15048
rect 8402 15224 8436 15240
rect 8402 15032 8436 15048
rect 8520 15224 8554 15240
rect 8520 15032 8554 15048
rect 8638 15224 8672 15274
rect 8638 15032 8672 15048
rect 8756 15224 8790 15240
rect 8756 15032 8790 15048
rect 8874 15224 8908 15274
rect 15187 15273 15457 15307
rect 8874 15032 8908 15048
rect 14361 15223 14395 15239
rect 14361 15031 14395 15047
rect 14479 15223 14513 15239
rect 14479 15031 14513 15047
rect 14597 15223 14631 15239
rect 14597 15031 14631 15047
rect 14715 15223 14749 15239
rect 14715 15031 14749 15047
rect 14833 15223 14867 15239
rect 14833 15031 14867 15047
rect 14951 15223 14985 15239
rect 14951 15031 14985 15047
rect 15069 15223 15103 15239
rect 15069 15031 15103 15047
rect 15187 15223 15221 15273
rect 15187 15031 15221 15047
rect 15305 15223 15339 15239
rect 15305 15031 15339 15047
rect 15423 15223 15457 15273
rect 21841 15294 22111 15328
rect 21015 15244 21049 15260
rect 21015 15052 21049 15068
rect 21133 15244 21167 15260
rect 21133 15052 21167 15068
rect 21251 15244 21285 15260
rect 21251 15052 21285 15068
rect 21369 15244 21403 15260
rect 21369 15052 21403 15068
rect 21487 15244 21521 15260
rect 21487 15052 21521 15068
rect 21605 15244 21639 15260
rect 21605 15052 21639 15068
rect 21723 15244 21757 15260
rect 21723 15052 21757 15068
rect 21841 15244 21875 15294
rect 21841 15052 21875 15068
rect 21959 15244 21993 15260
rect 21959 15052 21993 15068
rect 22077 15244 22111 15294
rect 29957 15317 30125 15333
rect 29957 15247 29973 15317
rect 30109 15247 30125 15317
rect 29957 15231 30125 15247
rect 32099 15210 32110 15410
rect 32531 15210 32543 15410
rect 32099 15204 32543 15210
rect 30494 15127 30764 15161
rect 22077 15052 22111 15068
rect 29668 15077 29702 15093
rect 15423 15031 15457 15047
rect 8563 14954 8579 14988
rect 8613 14954 8629 14988
rect 15112 14953 15128 14987
rect 15162 14953 15178 14987
rect 21766 14974 21782 15008
rect 21816 14974 21832 15008
rect 8445 14837 8461 14871
rect 8495 14837 8511 14871
rect 14994 14836 15010 14870
rect 15044 14836 15060 14870
rect 21648 14857 21664 14891
rect 21698 14857 21714 14891
rect 29668 14885 29702 14901
rect 29786 15077 29820 15093
rect 29786 14885 29820 14901
rect 29904 15077 29938 15093
rect 29904 14885 29938 14901
rect 30022 15077 30056 15093
rect 30022 14885 30056 14901
rect 30140 15077 30174 15093
rect 30140 14885 30174 14901
rect 30258 15077 30292 15093
rect 30258 14885 30292 14901
rect 30376 15077 30410 15093
rect 30376 14885 30410 14901
rect 30494 15077 30528 15127
rect 30494 14885 30528 14901
rect 30612 15077 30646 15093
rect 30612 14885 30646 14901
rect 30730 15077 30764 15127
rect 30730 14885 30764 14901
rect 32314 14925 32584 14960
rect 31960 14872 31994 14888
rect 21252 14807 21286 14823
rect 8049 14787 8083 14803
rect 8049 14395 8083 14411
rect 8167 14787 8201 14803
rect 8167 14395 8201 14411
rect 8285 14787 8319 14803
rect 8402 14787 8436 14803
rect 8402 14595 8436 14611
rect 8520 14787 8554 14803
rect 8520 14595 8554 14611
rect 14598 14786 14632 14802
rect 8285 14395 8319 14411
rect 14598 14394 14632 14410
rect 14716 14786 14750 14802
rect 14716 14394 14750 14410
rect 14834 14786 14868 14802
rect 14951 14786 14985 14802
rect 14951 14594 14985 14610
rect 15069 14786 15103 14802
rect 15069 14594 15103 14610
rect 21252 14415 21286 14431
rect 21370 14807 21404 14823
rect 21370 14415 21404 14431
rect 21488 14807 21522 14823
rect 21605 14807 21639 14823
rect 21605 14615 21639 14631
rect 21723 14807 21757 14823
rect 30419 14807 30435 14841
rect 30469 14807 30485 14841
rect 31476 14726 31746 14761
rect 30301 14690 30317 14724
rect 30351 14690 30367 14724
rect 31476 14672 31510 14726
rect 21723 14615 21757 14631
rect 29905 14640 29939 14656
rect 21488 14415 21522 14431
rect 14834 14394 14868 14410
rect 21114 14383 21185 14385
rect 14283 14361 14563 14366
rect 8092 14327 8108 14361
rect 8142 14327 8158 14361
rect 8210 14327 8226 14361
rect 8260 14327 8276 14361
rect 14283 14315 14511 14361
rect 14560 14315 14563 14361
rect 14641 14326 14657 14360
rect 14691 14326 14707 14360
rect 14759 14326 14775 14360
rect 14809 14326 14825 14360
rect 21114 14335 21118 14383
rect 21179 14335 21185 14383
rect 21295 14347 21311 14381
rect 21345 14347 21361 14381
rect 21413 14347 21429 14381
rect 21463 14347 21479 14381
rect 14283 14310 14563 14315
rect 21114 14322 21185 14335
rect 8325 14256 8493 14274
rect 8325 14200 8341 14256
rect 8475 14200 8493 14256
rect 8325 14184 8493 14200
rect 54 13871 66 13927
rect 54 13864 125 13871
rect 203 14109 311 14112
rect 203 14059 227 14109
rect 288 14059 311 14109
rect -100 12582 127 12597
rect -100 12512 23 12582
rect 97 12512 127 12582
rect -100 12497 127 12512
rect -97 12496 127 12497
rect 203 12417 311 14059
rect 14283 14028 14336 14310
rect 14874 14255 15042 14273
rect 14874 14199 14890 14255
rect 15024 14199 15042 14255
rect 14874 14183 15042 14199
rect 362 13975 14336 14028
rect 362 13536 453 13975
rect 21114 13940 21177 14322
rect 492 13936 21177 13940
rect 492 13882 7930 13936
rect 7979 13882 21177 13936
rect 492 13874 21177 13882
rect 21211 14293 21272 14298
rect 21211 14255 21220 14293
rect 21265 14255 21272 14293
rect 492 13710 602 13874
rect 21211 13829 21272 14255
rect 21528 14276 21696 14294
rect 21528 14220 21544 14276
rect 21678 14220 21696 14276
rect 29905 14248 29939 14264
rect 30023 14640 30057 14656
rect 30023 14248 30057 14264
rect 30141 14640 30175 14656
rect 30258 14640 30292 14656
rect 30258 14448 30292 14464
rect 30376 14640 30410 14656
rect 31476 14480 31510 14496
rect 31594 14672 31628 14688
rect 31594 14480 31628 14496
rect 31712 14672 31746 14726
rect 31712 14480 31746 14496
rect 31830 14672 31864 14688
rect 31830 14480 31864 14496
rect 31960 14480 31994 14496
rect 32078 14872 32112 14888
rect 32078 14480 32112 14496
rect 32196 14872 32230 14888
rect 32196 14480 32230 14496
rect 32314 14872 32348 14925
rect 32314 14480 32348 14496
rect 32432 14872 32466 14888
rect 32432 14480 32466 14496
rect 32550 14872 32584 14925
rect 33558 14909 33726 14925
rect 32550 14480 32584 14496
rect 32668 14872 32702 14888
rect 33558 14839 33574 14909
rect 33710 14839 33726 14909
rect 33558 14823 33726 14839
rect 34095 14719 34365 14753
rect 32668 14480 32702 14496
rect 32797 14672 32831 14688
rect 32797 14480 32831 14496
rect 32915 14672 32949 14688
rect 32915 14480 32949 14496
rect 33033 14672 33067 14688
rect 33033 14480 33067 14496
rect 33151 14672 33185 14688
rect 33151 14480 33185 14496
rect 33269 14669 33303 14685
rect 33269 14477 33303 14493
rect 33387 14669 33421 14685
rect 33387 14477 33421 14493
rect 33505 14669 33539 14685
rect 33505 14477 33539 14493
rect 33623 14669 33657 14685
rect 33623 14477 33657 14493
rect 33741 14669 33775 14685
rect 33741 14477 33775 14493
rect 33859 14669 33893 14685
rect 33859 14477 33893 14493
rect 33977 14669 34011 14685
rect 33977 14477 34011 14493
rect 34095 14669 34129 14719
rect 34095 14477 34129 14493
rect 34213 14669 34247 14685
rect 34213 14477 34247 14493
rect 34331 14669 34365 14719
rect 34331 14477 34365 14493
rect 30376 14448 30410 14464
rect 34020 14399 34036 14433
rect 34070 14399 34086 14433
rect 33128 14314 33162 14330
rect 33902 14282 33918 14316
rect 33952 14282 33968 14316
rect 33128 14264 33162 14280
rect 30141 14248 30175 14264
rect 21528 14204 21696 14220
rect 33506 14232 33540 14248
rect 29948 14180 29964 14214
rect 29998 14180 30014 14214
rect 30066 14180 30082 14214
rect 30116 14180 30132 14214
rect 31205 14208 31547 14214
rect 31205 14140 31455 14208
rect 31535 14140 31547 14208
rect 31722 14195 31778 14212
rect 31722 14161 31728 14195
rect 31762 14161 31778 14195
rect 31722 14144 31778 14161
rect 31903 14179 31937 14195
rect 31205 14134 31547 14140
rect 30181 14109 30349 14127
rect 30181 14053 30197 14109
rect 30331 14053 30349 14109
rect 30181 14037 30349 14053
rect 362 13491 380 13536
rect 437 13491 453 13536
rect 362 13484 453 13491
rect 203 12416 331 12417
rect 192 12402 331 12416
rect 192 12335 207 12402
rect 193 12318 207 12335
rect 320 12318 331 12402
rect -248 9775 125 9795
rect -248 9694 20 9775
rect 114 9694 125 9775
rect -248 9678 125 9694
rect -393 4001 118 4009
rect -393 3919 21 4001
rect 103 3919 118 4001
rect -393 3908 118 3919
rect -1078 897 122 909
rect -1078 821 15 897
rect 109 821 122 897
rect -1078 813 122 821
rect 193 493 331 12318
rect 491 4000 602 13710
rect 2748 13763 21272 13829
rect 1437 13564 1605 13580
rect 1437 13494 1453 13564
rect 1589 13494 1605 13564
rect 1437 13478 1605 13494
rect 1974 13374 2244 13408
rect 1148 13324 1182 13340
rect 1148 13132 1182 13148
rect 1266 13324 1300 13340
rect 1266 13132 1300 13148
rect 1384 13324 1418 13340
rect 1384 13132 1418 13148
rect 1502 13324 1536 13340
rect 1502 13132 1536 13148
rect 1620 13324 1654 13340
rect 1620 13132 1654 13148
rect 1738 13324 1772 13340
rect 1738 13132 1772 13148
rect 1856 13324 1890 13340
rect 1856 13132 1890 13148
rect 1974 13324 2008 13374
rect 1974 13132 2008 13148
rect 2092 13324 2126 13340
rect 2092 13132 2126 13148
rect 2210 13324 2244 13374
rect 2210 13132 2244 13148
rect 1899 13054 1915 13088
rect 1949 13054 1965 13088
rect 1781 12937 1797 12971
rect 1831 12937 1847 12971
rect 1385 12887 1419 12903
rect 491 3919 499 4000
rect 601 3919 602 4000
rect 491 3908 602 3919
rect 637 12580 740 12588
rect 637 12504 645 12580
rect 734 12504 740 12580
rect 637 642 740 12504
rect 1385 12495 1419 12511
rect 1503 12887 1537 12903
rect 1503 12495 1537 12511
rect 1621 12887 1655 12903
rect 1738 12887 1772 12903
rect 1738 12695 1772 12711
rect 1856 12887 1890 12903
rect 1856 12695 1890 12711
rect 1621 12495 1655 12511
rect 1428 12427 1444 12461
rect 1478 12427 1494 12461
rect 1546 12427 1562 12461
rect 1596 12427 1612 12461
rect 883 12386 1198 12391
rect 883 12342 1139 12386
rect 1195 12342 1198 12386
rect 883 12338 1198 12342
rect 1661 12356 1829 12374
rect 883 6532 965 12338
rect 1661 12300 1677 12356
rect 1811 12300 1829 12356
rect 1661 12284 1829 12300
rect 1429 10979 1597 10995
rect 1429 10909 1445 10979
rect 1581 10909 1597 10979
rect 1429 10893 1597 10909
rect 1966 10789 2236 10823
rect 1140 10739 1174 10755
rect 1140 10547 1174 10563
rect 1258 10739 1292 10755
rect 1258 10547 1292 10563
rect 1376 10739 1410 10755
rect 1376 10547 1410 10563
rect 1494 10739 1528 10755
rect 1494 10547 1528 10563
rect 1612 10739 1646 10755
rect 1612 10547 1646 10563
rect 1730 10739 1764 10755
rect 1730 10547 1764 10563
rect 1848 10739 1882 10755
rect 1848 10547 1882 10563
rect 1966 10739 2000 10789
rect 1966 10547 2000 10563
rect 2084 10739 2118 10755
rect 2084 10547 2118 10563
rect 2202 10739 2236 10789
rect 2202 10547 2236 10563
rect 1891 10469 1907 10503
rect 1941 10469 1957 10503
rect 1773 10352 1789 10386
rect 1823 10352 1839 10386
rect 1377 10302 1411 10318
rect 1377 9910 1411 9926
rect 1495 10302 1529 10318
rect 1495 9910 1529 9926
rect 1613 10302 1647 10318
rect 1730 10302 1764 10318
rect 1730 10110 1764 10126
rect 1848 10302 1882 10318
rect 1848 10110 1882 10126
rect 1613 9910 1647 9926
rect 1420 9842 1436 9876
rect 1470 9842 1486 9876
rect 1538 9842 1554 9876
rect 1588 9842 1604 9876
rect 1653 9771 1821 9789
rect 1653 9715 1669 9771
rect 1803 9715 1821 9771
rect 1653 9699 1821 9715
rect 1410 7701 1578 7717
rect 1410 7631 1426 7701
rect 1562 7631 1578 7701
rect 1410 7615 1578 7631
rect 1947 7511 2217 7545
rect 1121 7461 1155 7477
rect 1121 7269 1155 7285
rect 1239 7461 1273 7477
rect 1239 7269 1273 7285
rect 1357 7461 1391 7477
rect 1357 7269 1391 7285
rect 1475 7461 1509 7477
rect 1475 7269 1509 7285
rect 1593 7461 1627 7477
rect 1593 7269 1627 7285
rect 1711 7461 1745 7477
rect 1711 7269 1745 7285
rect 1829 7461 1863 7477
rect 1829 7269 1863 7285
rect 1947 7461 1981 7511
rect 1947 7269 1981 7285
rect 2065 7461 2099 7477
rect 2065 7269 2099 7285
rect 2183 7461 2217 7511
rect 2183 7269 2217 7285
rect 1872 7191 1888 7225
rect 1922 7191 1938 7225
rect 1754 7074 1770 7108
rect 1804 7074 1820 7108
rect 1358 7024 1392 7040
rect 1358 6632 1392 6648
rect 1476 7024 1510 7040
rect 1476 6632 1510 6648
rect 1594 7024 1628 7040
rect 1711 7024 1745 7040
rect 1711 6832 1745 6848
rect 1829 7024 1863 7040
rect 1829 6832 1863 6848
rect 1594 6632 1628 6648
rect 1401 6564 1417 6598
rect 1451 6564 1467 6598
rect 1519 6564 1535 6598
rect 1569 6564 1585 6598
rect 883 6527 1148 6532
rect 883 6474 1083 6527
rect 1143 6474 1148 6527
rect 883 6470 1148 6474
rect 1634 6493 1802 6511
rect 1634 6437 1650 6493
rect 1784 6437 1802 6493
rect 1634 6421 1802 6437
rect 1426 4941 1594 4957
rect 1426 4871 1442 4941
rect 1578 4871 1594 4941
rect 1426 4855 1594 4871
rect 1963 4751 2233 4785
rect 1137 4701 1171 4717
rect 1137 4509 1171 4525
rect 1255 4701 1289 4717
rect 1255 4509 1289 4525
rect 1373 4701 1407 4717
rect 1373 4509 1407 4525
rect 1491 4701 1525 4717
rect 1491 4509 1525 4525
rect 1609 4701 1643 4717
rect 1609 4509 1643 4525
rect 1727 4701 1761 4717
rect 1727 4509 1761 4525
rect 1845 4701 1879 4717
rect 1845 4509 1879 4525
rect 1963 4701 1997 4751
rect 1963 4509 1997 4525
rect 2081 4701 2115 4717
rect 2081 4509 2115 4525
rect 2199 4701 2233 4751
rect 2199 4509 2233 4525
rect 1888 4431 1904 4465
rect 1938 4431 1954 4465
rect 1770 4314 1786 4348
rect 1820 4314 1836 4348
rect 1374 4264 1408 4280
rect 1374 3872 1408 3888
rect 1492 4264 1526 4280
rect 1492 3872 1526 3888
rect 1610 4264 1644 4280
rect 1727 4264 1761 4280
rect 1727 4072 1761 4088
rect 1845 4264 1879 4280
rect 1845 4072 1879 4088
rect 1610 3872 1644 3888
rect 1417 3804 1433 3838
rect 1467 3804 1483 3838
rect 1535 3804 1551 3838
rect 1585 3804 1601 3838
rect 1650 3733 1818 3751
rect 1650 3677 1666 3733
rect 1800 3677 1818 3733
rect 1650 3661 1818 3677
rect 594 633 785 642
rect 594 567 619 633
rect 763 567 785 633
rect 594 559 785 567
rect 193 422 204 493
rect 318 422 331 493
rect 193 405 331 422
rect -1230 361 136 371
rect 2748 370 2875 13763
rect 4433 13472 4656 13547
rect 4433 13471 4513 13472
rect 4433 13322 4512 13471
rect 4580 13323 4656 13472
rect 4579 13322 4656 13323
rect 4433 13216 4656 13322
rect 6915 13525 7138 13601
rect 6915 13376 6994 13525
rect 7061 13522 7138 13525
rect 6915 13373 6995 13376
rect 7062 13373 7138 13522
rect 6248 13305 6282 13321
rect 6248 13255 6282 13271
rect 6915 13270 7138 13373
rect 8062 13525 8285 13601
rect 8062 13524 8141 13525
rect 8062 13375 8137 13524
rect 8208 13376 8285 13525
rect 8204 13375 8285 13376
rect 7378 13311 7412 13327
rect 7378 13261 7412 13277
rect 8062 13270 8285 13375
rect 10982 13560 11205 13635
rect 10982 13559 11062 13560
rect 10982 13410 11061 13559
rect 11129 13411 11205 13560
rect 11128 13410 11205 13411
rect 10982 13304 11205 13410
rect 13464 13613 13687 13689
rect 13464 13464 13543 13613
rect 13610 13611 13687 13613
rect 13464 13462 13545 13464
rect 13612 13462 13687 13611
rect 12797 13393 12831 13409
rect 12797 13343 12831 13359
rect 13464 13358 13687 13462
rect 14611 13613 14834 13689
rect 14611 13464 14689 13613
rect 14757 13464 14834 13613
rect 13927 13399 13961 13415
rect 13927 13349 13961 13365
rect 14611 13358 14834 13464
rect 17636 13491 17859 13567
rect 17636 13341 17715 13491
rect 17782 13341 17859 13491
rect 20118 13546 20341 13621
rect 20118 13397 20196 13546
rect 20263 13545 20341 13546
rect 20118 13396 20197 13397
rect 20264 13396 20341 13545
rect 12797 13275 12831 13291
rect 6248 13187 6282 13203
rect 4864 13107 5134 13141
rect 6248 13137 6282 13153
rect 7378 13191 7412 13207
rect 11413 13195 11683 13229
rect 12797 13225 12831 13241
rect 13927 13279 13961 13295
rect 4038 13057 4072 13073
rect 4038 12865 4072 12881
rect 4156 13057 4190 13073
rect 4156 12865 4190 12881
rect 4274 13057 4308 13073
rect 4274 12865 4308 12881
rect 4392 13057 4426 13073
rect 4392 12865 4426 12881
rect 4510 13057 4544 13073
rect 4510 12865 4544 12881
rect 4628 13057 4662 13073
rect 4628 12865 4662 12881
rect 4746 13057 4780 13073
rect 4746 12865 4780 12881
rect 4864 13057 4898 13107
rect 4864 12865 4898 12881
rect 4982 13057 5016 13073
rect 4982 12865 5016 12881
rect 5100 13057 5134 13107
rect 5100 12865 5134 12881
rect 6363 13129 6397 13145
rect 4789 12787 4805 12821
rect 4839 12787 4855 12821
rect 6363 12737 6397 12753
rect 6481 13129 6515 13145
rect 6481 12737 6515 12753
rect 6599 13129 6633 13145
rect 6599 12737 6633 12753
rect 6717 13129 6751 13145
rect 6717 12737 6751 12753
rect 6835 13129 6869 13145
rect 6835 12737 6869 12753
rect 6953 13129 6987 13145
rect 6953 12737 6987 12753
rect 7071 13129 7105 13145
rect 7378 13141 7412 13157
rect 7071 12737 7105 12753
rect 7505 13133 7539 13149
rect 7505 12741 7539 12757
rect 7623 13133 7657 13149
rect 7623 12741 7657 12757
rect 7741 13133 7775 13149
rect 7741 12741 7775 12757
rect 7859 13133 7893 13149
rect 7859 12741 7893 12757
rect 7977 13133 8011 13149
rect 7977 12741 8011 12757
rect 8095 13133 8129 13149
rect 8095 12741 8129 12757
rect 8213 13133 8247 13149
rect 10587 13145 10621 13161
rect 10587 12953 10621 12969
rect 10705 13145 10739 13161
rect 10705 12953 10739 12969
rect 10823 13145 10857 13161
rect 10823 12953 10857 12969
rect 10941 13145 10975 13161
rect 10941 12953 10975 12969
rect 11059 13145 11093 13161
rect 11059 12953 11093 12969
rect 11177 13145 11211 13161
rect 11177 12953 11211 12969
rect 11295 13145 11329 13161
rect 11295 12953 11329 12969
rect 11413 13145 11447 13195
rect 11413 12953 11447 12969
rect 11531 13145 11565 13161
rect 11531 12953 11565 12969
rect 11649 13145 11683 13195
rect 11649 12953 11683 12969
rect 12912 13217 12946 13233
rect 11338 12875 11354 12909
rect 11388 12875 11404 12909
rect 12912 12825 12946 12841
rect 13030 13217 13064 13233
rect 13030 12825 13064 12841
rect 13148 13217 13182 13233
rect 13148 12825 13182 12841
rect 13266 13217 13300 13233
rect 13266 12825 13300 12841
rect 13384 13217 13418 13233
rect 13384 12825 13418 12841
rect 13502 13217 13536 13233
rect 13502 12825 13536 12841
rect 13620 13217 13654 13233
rect 13927 13229 13961 13245
rect 13620 12825 13654 12841
rect 14054 13221 14088 13237
rect 14054 12829 14088 12845
rect 14172 13221 14206 13237
rect 14172 12829 14206 12845
rect 14290 13221 14324 13237
rect 14290 12829 14324 12845
rect 14408 13221 14442 13237
rect 14408 12829 14442 12845
rect 14526 13221 14560 13237
rect 14526 12829 14560 12845
rect 14644 13221 14678 13237
rect 14644 12829 14678 12845
rect 14762 13221 14796 13237
rect 17636 13236 17859 13341
rect 19451 13325 19485 13341
rect 19451 13275 19485 13291
rect 20118 13290 20341 13396
rect 21265 13545 21488 13621
rect 21265 13396 21343 13545
rect 21411 13396 21488 13545
rect 20581 13331 20615 13347
rect 20581 13281 20615 13297
rect 21265 13290 21488 13396
rect 24261 13559 24484 13635
rect 24261 13410 24335 13559
rect 24407 13410 24484 13559
rect 24261 13304 24484 13410
rect 26743 13613 26966 13689
rect 26743 13611 26822 13613
rect 26743 13462 26819 13611
rect 26889 13464 26966 13613
rect 26886 13462 26966 13464
rect 26076 13393 26110 13409
rect 26076 13343 26110 13359
rect 26743 13358 26966 13462
rect 27890 13617 28113 13689
rect 27890 13468 27968 13617
rect 28035 13613 28113 13617
rect 27890 13464 27969 13468
rect 28036 13464 28113 13613
rect 27206 13399 27240 13415
rect 27206 13349 27240 13365
rect 27890 13358 28113 13464
rect 26076 13275 26110 13291
rect 19451 13207 19485 13223
rect 18067 13127 18337 13161
rect 19451 13157 19485 13173
rect 20581 13211 20615 13227
rect 17241 13077 17275 13093
rect 17241 12885 17275 12901
rect 17359 13077 17393 13093
rect 17359 12885 17393 12901
rect 17477 13077 17511 13093
rect 17477 12885 17511 12901
rect 17595 13077 17629 13093
rect 17595 12885 17629 12901
rect 17713 13077 17747 13093
rect 17713 12885 17747 12901
rect 17831 13077 17865 13093
rect 17831 12885 17865 12901
rect 17949 13077 17983 13093
rect 17949 12885 17983 12901
rect 18067 13077 18101 13127
rect 18067 12885 18101 12901
rect 18185 13077 18219 13093
rect 18185 12885 18219 12901
rect 18303 13077 18337 13127
rect 18303 12885 18337 12901
rect 19566 13149 19600 13165
rect 14762 12829 14796 12845
rect 17992 12807 18008 12841
rect 18042 12807 18058 12841
rect 11220 12758 11236 12792
rect 11270 12758 11286 12792
rect 19566 12757 19600 12773
rect 19684 13149 19718 13165
rect 19684 12757 19718 12773
rect 19802 13149 19836 13165
rect 19802 12757 19836 12773
rect 19920 13149 19954 13165
rect 19920 12757 19954 12773
rect 20038 13149 20072 13165
rect 20038 12757 20072 12773
rect 20156 13149 20190 13165
rect 20156 12757 20190 12773
rect 20274 13149 20308 13165
rect 20581 13161 20615 13177
rect 24692 13195 24962 13229
rect 26076 13225 26110 13241
rect 27206 13279 27240 13295
rect 20274 12757 20308 12773
rect 20708 13153 20742 13169
rect 20708 12761 20742 12777
rect 20826 13153 20860 13169
rect 20826 12761 20860 12777
rect 20944 13153 20978 13169
rect 20944 12761 20978 12777
rect 21062 13153 21096 13169
rect 21062 12761 21096 12777
rect 21180 13153 21214 13169
rect 21180 12761 21214 12777
rect 21298 13153 21332 13169
rect 21298 12761 21332 12777
rect 21416 13153 21450 13169
rect 23866 13145 23900 13161
rect 23866 12953 23900 12969
rect 23984 13145 24018 13161
rect 23984 12953 24018 12969
rect 24102 13145 24136 13161
rect 24102 12953 24136 12969
rect 24220 13145 24254 13161
rect 24220 12953 24254 12969
rect 24338 13145 24372 13161
rect 24338 12953 24372 12969
rect 24456 13145 24490 13161
rect 24456 12953 24490 12969
rect 24574 13145 24608 13161
rect 24574 12953 24608 12969
rect 24692 13145 24726 13195
rect 24692 12953 24726 12969
rect 24810 13145 24844 13161
rect 24810 12953 24844 12969
rect 24928 13145 24962 13195
rect 24928 12953 24962 12969
rect 26191 13217 26225 13233
rect 24617 12875 24633 12909
rect 24667 12875 24683 12909
rect 26191 12825 26225 12841
rect 26309 13217 26343 13233
rect 26309 12825 26343 12841
rect 26427 13217 26461 13233
rect 26427 12825 26461 12841
rect 26545 13217 26579 13233
rect 26545 12825 26579 12841
rect 26663 13217 26697 13233
rect 26663 12825 26697 12841
rect 26781 13217 26815 13233
rect 26781 12825 26815 12841
rect 26899 13217 26933 13233
rect 27206 13229 27240 13245
rect 26899 12825 26933 12841
rect 27333 13221 27367 13237
rect 27333 12829 27367 12845
rect 27451 13221 27485 13237
rect 27451 12829 27485 12845
rect 27569 13221 27603 13237
rect 27569 12829 27603 12845
rect 27687 13221 27721 13237
rect 27687 12829 27721 12845
rect 27805 13221 27839 13237
rect 27805 12829 27839 12845
rect 27923 13221 27957 13237
rect 27923 12829 27957 12845
rect 28041 13221 28075 13237
rect 28041 12829 28075 12845
rect 21416 12761 21450 12777
rect 24499 12758 24515 12792
rect 24549 12758 24565 12792
rect 8213 12741 8247 12757
rect 29952 12746 30120 12762
rect 10824 12708 10858 12724
rect 4671 12670 4687 12704
rect 4721 12670 4737 12704
rect 4275 12620 4309 12636
rect 4275 12228 4309 12244
rect 4393 12620 4427 12636
rect 4393 12228 4427 12244
rect 4511 12620 4545 12636
rect 4628 12620 4662 12636
rect 4628 12428 4662 12444
rect 4746 12620 4780 12636
rect 4746 12428 4780 12444
rect 6552 12397 6568 12431
rect 6602 12397 6618 12431
rect 7694 12401 7710 12435
rect 7744 12401 7760 12435
rect 6273 12346 6307 12362
rect 4511 12228 4545 12244
rect 4798 12294 5047 12337
rect 4798 12204 4845 12294
rect 5008 12204 5047 12294
rect 4318 12160 4334 12194
rect 4368 12160 4384 12194
rect 4436 12160 4452 12194
rect 4486 12160 4502 12194
rect 4798 12165 5047 12204
rect 6273 12154 6307 12170
rect 6391 12346 6425 12362
rect 6391 12154 6425 12170
rect 6509 12346 6543 12362
rect 6509 12154 6543 12170
rect 6627 12346 6661 12362
rect 6627 12154 6661 12170
rect 6792 12346 6826 12362
rect 6792 12154 6826 12170
rect 6910 12346 6944 12362
rect 6910 12154 6944 12170
rect 7028 12346 7062 12362
rect 7028 12154 7062 12170
rect 7146 12346 7180 12362
rect 7146 12154 7180 12170
rect 7415 12350 7449 12366
rect 7415 12158 7449 12174
rect 7533 12350 7567 12366
rect 7533 12158 7567 12174
rect 7651 12350 7685 12366
rect 7651 12158 7685 12174
rect 7769 12350 7803 12366
rect 7769 12158 7803 12174
rect 7934 12350 7968 12366
rect 7934 12158 7968 12174
rect 8052 12350 8086 12366
rect 8052 12158 8086 12174
rect 8170 12350 8204 12366
rect 8170 12158 8204 12174
rect 8288 12350 8322 12366
rect 10824 12316 10858 12332
rect 10942 12708 10976 12724
rect 10942 12316 10976 12332
rect 11060 12708 11094 12724
rect 11177 12708 11211 12724
rect 11177 12516 11211 12532
rect 11295 12708 11329 12724
rect 17874 12690 17890 12724
rect 17924 12690 17940 12724
rect 24103 12708 24137 12724
rect 11295 12516 11329 12532
rect 17478 12640 17512 12656
rect 13101 12485 13117 12519
rect 13151 12485 13167 12519
rect 14243 12489 14259 12523
rect 14293 12489 14309 12523
rect 12822 12434 12856 12450
rect 11060 12316 11094 12332
rect 11347 12382 11596 12425
rect 11347 12292 11394 12382
rect 11557 12292 11596 12382
rect 10867 12248 10883 12282
rect 10917 12248 10933 12282
rect 10985 12248 11001 12282
rect 11035 12248 11051 12282
rect 11347 12253 11596 12292
rect 12822 12242 12856 12258
rect 12940 12434 12974 12450
rect 12940 12242 12974 12258
rect 13058 12434 13092 12450
rect 13058 12242 13092 12258
rect 13176 12434 13210 12450
rect 13176 12242 13210 12258
rect 13341 12434 13375 12450
rect 13341 12242 13375 12258
rect 13459 12434 13493 12450
rect 13459 12242 13493 12258
rect 13577 12434 13611 12450
rect 13577 12242 13611 12258
rect 13695 12434 13729 12450
rect 13695 12242 13729 12258
rect 13964 12438 13998 12454
rect 13964 12246 13998 12262
rect 14082 12438 14116 12454
rect 14082 12246 14116 12262
rect 14200 12438 14234 12454
rect 14200 12246 14234 12262
rect 14318 12438 14352 12454
rect 14318 12246 14352 12262
rect 14483 12438 14517 12454
rect 14483 12246 14517 12262
rect 14601 12438 14635 12454
rect 14601 12246 14635 12262
rect 14719 12438 14753 12454
rect 14719 12246 14753 12262
rect 14837 12438 14871 12454
rect 14837 12246 14871 12262
rect 17478 12248 17512 12264
rect 17596 12640 17630 12656
rect 17596 12248 17630 12264
rect 17714 12640 17748 12656
rect 17831 12640 17865 12656
rect 17831 12448 17865 12464
rect 17949 12640 17983 12656
rect 17949 12448 17983 12464
rect 19755 12417 19771 12451
rect 19805 12417 19821 12451
rect 20897 12421 20913 12455
rect 20947 12421 20963 12455
rect 19476 12366 19510 12382
rect 17714 12248 17748 12264
rect 18001 12314 18250 12357
rect 18001 12224 18048 12314
rect 18211 12224 18250 12314
rect 17521 12180 17537 12214
rect 17571 12180 17587 12214
rect 17639 12180 17655 12214
rect 17689 12180 17705 12214
rect 18001 12185 18250 12224
rect 19476 12174 19510 12190
rect 19594 12366 19628 12382
rect 19594 12174 19628 12190
rect 19712 12366 19746 12382
rect 19712 12174 19746 12190
rect 19830 12366 19864 12382
rect 19830 12174 19864 12190
rect 19995 12366 20029 12382
rect 19995 12174 20029 12190
rect 20113 12366 20147 12382
rect 20113 12174 20147 12190
rect 20231 12366 20265 12382
rect 20231 12174 20265 12190
rect 20349 12366 20383 12382
rect 20349 12174 20383 12190
rect 20618 12370 20652 12386
rect 20618 12178 20652 12194
rect 20736 12370 20770 12386
rect 20736 12178 20770 12194
rect 20854 12370 20888 12386
rect 20854 12178 20888 12194
rect 20972 12370 21006 12386
rect 20972 12178 21006 12194
rect 21137 12370 21171 12386
rect 21137 12178 21171 12194
rect 21255 12370 21289 12386
rect 21255 12178 21289 12194
rect 21373 12370 21407 12386
rect 21373 12178 21407 12194
rect 21491 12370 21525 12386
rect 24103 12316 24137 12332
rect 24221 12708 24255 12724
rect 24221 12316 24255 12332
rect 24339 12708 24373 12724
rect 24456 12708 24490 12724
rect 24456 12516 24490 12532
rect 24574 12708 24608 12724
rect 29952 12676 29968 12746
rect 30104 12676 30120 12746
rect 29952 12660 30120 12676
rect 24574 12516 24608 12532
rect 30489 12556 30759 12590
rect 26380 12485 26396 12519
rect 26430 12485 26446 12519
rect 27522 12489 27538 12523
rect 27572 12489 27588 12523
rect 29663 12506 29697 12522
rect 26101 12434 26135 12450
rect 24339 12316 24373 12332
rect 24626 12382 24875 12425
rect 24626 12292 24673 12382
rect 24836 12292 24875 12382
rect 24146 12248 24162 12282
rect 24196 12248 24212 12282
rect 24264 12248 24280 12282
rect 24314 12248 24330 12282
rect 24626 12253 24875 12292
rect 26101 12242 26135 12258
rect 26219 12434 26253 12450
rect 26219 12242 26253 12258
rect 26337 12434 26371 12450
rect 26337 12242 26371 12258
rect 26455 12434 26489 12450
rect 26455 12242 26489 12258
rect 26620 12434 26654 12450
rect 26620 12242 26654 12258
rect 26738 12434 26772 12450
rect 26738 12242 26772 12258
rect 26856 12434 26890 12450
rect 26856 12242 26890 12258
rect 26974 12434 27008 12450
rect 26974 12242 27008 12258
rect 27243 12438 27277 12454
rect 27243 12246 27277 12262
rect 27361 12438 27395 12454
rect 27361 12246 27395 12262
rect 27479 12438 27513 12454
rect 27479 12246 27513 12262
rect 27597 12438 27631 12454
rect 27597 12246 27631 12262
rect 27762 12438 27796 12454
rect 27762 12246 27796 12262
rect 27880 12438 27914 12454
rect 27880 12246 27914 12262
rect 27998 12438 28032 12454
rect 27998 12246 28032 12262
rect 28116 12438 28150 12454
rect 29663 12314 29697 12330
rect 29781 12506 29815 12522
rect 29781 12314 29815 12330
rect 29899 12506 29933 12522
rect 29899 12314 29933 12330
rect 30017 12506 30051 12522
rect 30017 12314 30051 12330
rect 30135 12506 30169 12522
rect 30135 12314 30169 12330
rect 30253 12506 30287 12522
rect 30253 12314 30287 12330
rect 30371 12506 30405 12522
rect 30371 12314 30405 12330
rect 30489 12506 30523 12556
rect 30489 12314 30523 12330
rect 30607 12506 30641 12522
rect 30607 12314 30641 12330
rect 30725 12506 30759 12556
rect 30725 12314 30759 12330
rect 28116 12246 28150 12262
rect 30414 12236 30430 12270
rect 30464 12236 30480 12270
rect 21491 12178 21525 12194
rect 8288 12158 8322 12174
rect 30296 12119 30312 12153
rect 30346 12119 30362 12153
rect 29900 12069 29934 12085
rect 12837 12011 13009 12058
rect 6288 11923 6460 11970
rect 4447 11821 4670 11897
rect 4447 11672 4525 11821
rect 4593 11672 4670 11821
rect 6288 11760 6327 11923
rect 6417 11760 6460 11923
rect 6288 11721 6460 11760
rect 7430 11921 7602 11968
rect 7430 11758 7469 11921
rect 7559 11758 7602 11921
rect 7430 11719 7602 11758
rect 10996 11909 11219 11985
rect 10996 11760 11075 11909
rect 11142 11908 11219 11909
rect 10996 11759 11076 11760
rect 11143 11759 11219 11908
rect 12837 11848 12876 12011
rect 12966 11848 13009 12011
rect 12837 11809 13009 11848
rect 13979 12009 14151 12056
rect 13979 11846 14018 12009
rect 14108 11846 14151 12009
rect 26116 12011 26288 12058
rect 19491 11943 19663 11990
rect 13979 11807 14151 11846
rect 17650 11842 17873 11917
rect 17650 11841 17730 11842
rect 4447 11566 4670 11672
rect 10996 11654 11219 11759
rect 17650 11692 17729 11841
rect 17797 11693 17873 11842
rect 19491 11780 19530 11943
rect 19620 11780 19663 11943
rect 19491 11741 19663 11780
rect 20633 11941 20805 11988
rect 20633 11778 20672 11941
rect 20762 11778 20805 11941
rect 20633 11739 20805 11778
rect 24275 11909 24498 11985
rect 24275 11760 24354 11909
rect 24421 11908 24498 11909
rect 24275 11759 24358 11760
rect 24425 11759 24498 11908
rect 26116 11848 26155 12011
rect 26245 11848 26288 12011
rect 26116 11846 26159 11848
rect 26226 11846 26288 11848
rect 26116 11809 26288 11846
rect 27258 12009 27430 12056
rect 27258 11846 27297 12009
rect 27387 11846 27430 12009
rect 27258 11807 27430 11846
rect 17796 11692 17873 11693
rect 4878 11457 5148 11491
rect 4052 11407 4086 11423
rect 4052 11215 4086 11231
rect 4170 11407 4204 11423
rect 4170 11215 4204 11231
rect 4288 11407 4322 11423
rect 4288 11215 4322 11231
rect 4406 11407 4440 11423
rect 4406 11215 4440 11231
rect 4524 11407 4558 11423
rect 4524 11215 4558 11231
rect 4642 11407 4676 11423
rect 4642 11215 4676 11231
rect 4760 11407 4794 11423
rect 4760 11215 4794 11231
rect 4878 11407 4912 11457
rect 4878 11215 4912 11231
rect 4996 11407 5030 11423
rect 4996 11215 5030 11231
rect 5114 11407 5148 11457
rect 5114 11215 5148 11231
rect 8158 11479 8383 11554
rect 11427 11545 11697 11579
rect 8158 11329 8237 11479
rect 8304 11329 8383 11479
rect 8158 11223 8383 11329
rect 10601 11495 10635 11511
rect 10601 11303 10635 11319
rect 10719 11495 10753 11511
rect 10719 11303 10753 11319
rect 10837 11495 10871 11511
rect 10837 11303 10871 11319
rect 10955 11495 10989 11511
rect 10955 11303 10989 11319
rect 11073 11495 11107 11511
rect 11073 11303 11107 11319
rect 11191 11495 11225 11511
rect 11191 11303 11225 11319
rect 11309 11495 11343 11511
rect 11309 11303 11343 11319
rect 11427 11495 11461 11545
rect 11427 11303 11461 11319
rect 11545 11495 11579 11511
rect 11545 11303 11579 11319
rect 11663 11495 11697 11545
rect 11663 11303 11697 11319
rect 14707 11566 14932 11642
rect 17650 11586 17873 11692
rect 24275 11654 24498 11759
rect 29900 11677 29934 11693
rect 30018 12069 30052 12085
rect 30018 11677 30052 11693
rect 30136 12069 30170 12085
rect 30253 12069 30287 12085
rect 30253 11877 30287 11893
rect 30371 12069 30405 12085
rect 30371 11877 30405 11893
rect 30136 11677 30170 11693
rect 14707 11417 14786 11566
rect 14858 11417 14932 11566
rect 18081 11477 18351 11511
rect 14707 11311 14932 11417
rect 17255 11427 17289 11443
rect 11352 11225 11368 11259
rect 11402 11225 11418 11259
rect 17255 11235 17289 11251
rect 17373 11427 17407 11443
rect 17373 11235 17407 11251
rect 17491 11427 17525 11443
rect 17491 11235 17525 11251
rect 17609 11427 17643 11443
rect 17609 11235 17643 11251
rect 17727 11427 17761 11443
rect 17727 11235 17761 11251
rect 17845 11427 17879 11443
rect 17845 11235 17879 11251
rect 17963 11427 17997 11443
rect 17963 11235 17997 11251
rect 18081 11427 18115 11477
rect 18081 11235 18115 11251
rect 18199 11427 18233 11443
rect 18199 11235 18233 11251
rect 18317 11427 18351 11477
rect 18317 11235 18351 11251
rect 21361 11498 21586 11574
rect 24706 11545 24976 11579
rect 21361 11494 21440 11498
rect 21361 11345 21437 11494
rect 21507 11349 21586 11498
rect 21504 11345 21586 11349
rect 21361 11243 21586 11345
rect 23880 11495 23914 11511
rect 23880 11303 23914 11319
rect 23998 11495 24032 11511
rect 23998 11303 24032 11319
rect 24116 11495 24150 11511
rect 24116 11303 24150 11319
rect 24234 11495 24268 11511
rect 24234 11303 24268 11319
rect 24352 11495 24386 11511
rect 24352 11303 24386 11319
rect 24470 11495 24504 11511
rect 24470 11303 24504 11319
rect 24588 11495 24622 11511
rect 24588 11303 24622 11319
rect 24706 11495 24740 11545
rect 24706 11303 24740 11319
rect 24824 11495 24858 11511
rect 24824 11303 24858 11319
rect 24942 11495 24976 11545
rect 24942 11303 24976 11319
rect 27986 11566 28211 11642
rect 29943 11609 29959 11643
rect 29993 11609 30009 11643
rect 30061 11609 30077 11643
rect 30111 11609 30127 11643
rect 27986 11414 28065 11566
rect 28132 11414 28211 11566
rect 30176 11538 30344 11556
rect 30176 11482 30192 11538
rect 30326 11482 30344 11538
rect 30176 11466 30344 11482
rect 27986 11311 28211 11414
rect 24631 11225 24647 11259
rect 24681 11225 24697 11259
rect 4803 11137 4819 11171
rect 4853 11137 4869 11171
rect 11234 11108 11250 11142
rect 11284 11108 11300 11142
rect 12903 11131 13173 11166
rect 12549 11078 12583 11094
rect 4685 11020 4701 11054
rect 4735 11020 4751 11054
rect 6354 11043 6624 11078
rect 6000 10990 6034 11006
rect 4289 10970 4323 10986
rect 3143 10630 3403 10632
rect 3141 10601 3403 10630
rect 3141 10491 3250 10601
rect 3368 10491 3403 10601
rect 4289 10578 4323 10594
rect 4407 10970 4441 10986
rect 4407 10578 4441 10594
rect 4525 10970 4559 10986
rect 4642 10970 4676 10986
rect 4642 10778 4676 10794
rect 4760 10970 4794 10986
rect 4760 10778 4794 10794
rect 5516 10844 5786 10879
rect 5516 10790 5550 10844
rect 4525 10578 4559 10594
rect 4812 10644 5061 10687
rect 4812 10554 4859 10644
rect 5022 10554 5061 10644
rect 5516 10598 5550 10614
rect 5634 10790 5668 10806
rect 5634 10598 5668 10614
rect 5752 10790 5786 10844
rect 5752 10598 5786 10614
rect 5870 10790 5904 10806
rect 5870 10598 5904 10614
rect 6000 10598 6034 10614
rect 6118 10990 6152 11006
rect 6118 10598 6152 10614
rect 6236 10990 6270 11006
rect 6236 10598 6270 10614
rect 6354 10990 6388 11043
rect 6354 10598 6388 10614
rect 6472 10990 6506 11006
rect 6472 10598 6506 10614
rect 6590 10990 6624 11043
rect 8252 11043 8522 11078
rect 6590 10598 6624 10614
rect 6708 10990 6742 11006
rect 7898 10990 7932 11006
rect 7414 10844 7684 10879
rect 6708 10598 6742 10614
rect 6837 10790 6871 10806
rect 6837 10598 6871 10614
rect 6955 10790 6989 10806
rect 6955 10598 6989 10614
rect 7073 10790 7107 10806
rect 7073 10598 7107 10614
rect 7191 10790 7225 10806
rect 7191 10598 7225 10614
rect 7414 10790 7448 10844
rect 7414 10598 7448 10614
rect 7532 10790 7566 10806
rect 7532 10598 7566 10614
rect 7650 10790 7684 10844
rect 7650 10598 7684 10614
rect 7768 10790 7802 10806
rect 7768 10598 7802 10614
rect 7898 10598 7932 10614
rect 8016 10990 8050 11006
rect 8016 10598 8050 10614
rect 8134 10990 8168 11006
rect 8134 10598 8168 10614
rect 8252 10990 8286 11043
rect 8252 10598 8286 10614
rect 8370 10990 8404 11006
rect 8370 10598 8404 10614
rect 8488 10990 8522 11043
rect 10838 11058 10872 11074
rect 8488 10598 8522 10614
rect 8606 10990 8640 11006
rect 8606 10598 8640 10614
rect 8735 10790 8769 10806
rect 8735 10598 8769 10614
rect 8853 10790 8887 10806
rect 8853 10598 8887 10614
rect 8971 10790 9005 10806
rect 8971 10598 9005 10614
rect 9089 10790 9123 10806
rect 10838 10666 10872 10682
rect 10956 11058 10990 11074
rect 10956 10666 10990 10682
rect 11074 11058 11108 11074
rect 11191 11058 11225 11074
rect 11191 10866 11225 10882
rect 11309 11058 11343 11074
rect 11309 10866 11343 10882
rect 12065 10932 12335 10967
rect 12065 10878 12099 10932
rect 11074 10666 11108 10682
rect 11361 10732 11610 10775
rect 11361 10642 11408 10732
rect 11571 10642 11610 10732
rect 12065 10686 12099 10702
rect 12183 10878 12217 10894
rect 12183 10686 12217 10702
rect 12301 10878 12335 10932
rect 12301 10686 12335 10702
rect 12419 10878 12453 10894
rect 12419 10686 12453 10702
rect 12549 10686 12583 10702
rect 12667 11078 12701 11094
rect 12667 10686 12701 10702
rect 12785 11078 12819 11094
rect 12785 10686 12819 10702
rect 12903 11078 12937 11131
rect 12903 10686 12937 10702
rect 13021 11078 13055 11094
rect 13021 10686 13055 10702
rect 13139 11078 13173 11131
rect 14801 11131 15071 11166
rect 18006 11157 18022 11191
rect 18056 11157 18072 11191
rect 13139 10686 13173 10702
rect 13257 11078 13291 11094
rect 14447 11078 14481 11094
rect 13963 10932 14233 10967
rect 13257 10686 13291 10702
rect 13386 10878 13420 10894
rect 13386 10686 13420 10702
rect 13504 10878 13538 10894
rect 13504 10686 13538 10702
rect 13622 10878 13656 10894
rect 13622 10686 13656 10702
rect 13740 10878 13774 10894
rect 13740 10686 13774 10702
rect 13963 10878 13997 10932
rect 13963 10686 13997 10702
rect 14081 10878 14115 10894
rect 14081 10686 14115 10702
rect 14199 10878 14233 10932
rect 14199 10686 14233 10702
rect 14317 10878 14351 10894
rect 14317 10686 14351 10702
rect 14447 10686 14481 10702
rect 14565 11078 14599 11094
rect 14565 10686 14599 10702
rect 14683 11078 14717 11094
rect 14683 10686 14717 10702
rect 14801 11078 14835 11131
rect 14801 10686 14835 10702
rect 14919 11078 14953 11094
rect 14919 10686 14953 10702
rect 15037 11078 15071 11131
rect 24513 11108 24529 11142
rect 24563 11108 24579 11142
rect 26182 11131 26452 11166
rect 15037 10686 15071 10702
rect 15155 11078 15189 11094
rect 17888 11040 17904 11074
rect 17938 11040 17954 11074
rect 19557 11063 19827 11098
rect 19203 11010 19237 11026
rect 17492 10990 17526 11006
rect 15155 10686 15189 10702
rect 15284 10878 15318 10894
rect 15284 10686 15318 10702
rect 15402 10878 15436 10894
rect 15402 10686 15436 10702
rect 15520 10878 15554 10894
rect 15520 10686 15554 10702
rect 15638 10878 15672 10894
rect 15638 10686 15672 10702
rect 9089 10598 9123 10614
rect 10881 10598 10897 10632
rect 10931 10598 10947 10632
rect 10999 10598 11015 10632
rect 11049 10598 11065 10632
rect 11361 10603 11610 10642
rect 16386 10630 16612 10652
rect 4332 10510 4348 10544
rect 4382 10510 4398 10544
rect 4450 10510 4466 10544
rect 4500 10510 4516 10544
rect 4812 10515 5061 10554
rect 16386 10513 16452 10630
rect 16591 10513 16612 10630
rect 17492 10598 17526 10614
rect 17610 10990 17644 11006
rect 17610 10598 17644 10614
rect 17728 10990 17762 11006
rect 17845 10990 17879 11006
rect 17845 10798 17879 10814
rect 17963 10990 17997 11006
rect 17963 10798 17997 10814
rect 18719 10864 18989 10899
rect 18719 10810 18753 10864
rect 17728 10598 17762 10614
rect 18015 10664 18264 10707
rect 18015 10574 18062 10664
rect 18225 10574 18264 10664
rect 18719 10618 18753 10634
rect 18837 10810 18871 10826
rect 18837 10618 18871 10634
rect 18955 10810 18989 10864
rect 18955 10618 18989 10634
rect 19073 10810 19107 10826
rect 19073 10618 19107 10634
rect 19203 10618 19237 10634
rect 19321 11010 19355 11026
rect 19321 10618 19355 10634
rect 19439 11010 19473 11026
rect 19439 10618 19473 10634
rect 19557 11010 19591 11063
rect 19557 10618 19591 10634
rect 19675 11010 19709 11026
rect 19675 10618 19709 10634
rect 19793 11010 19827 11063
rect 21455 11063 21725 11098
rect 25828 11078 25862 11094
rect 19793 10618 19827 10634
rect 19911 11010 19945 11026
rect 21101 11010 21135 11026
rect 20617 10864 20887 10899
rect 19911 10618 19945 10634
rect 20040 10810 20074 10826
rect 20040 10618 20074 10634
rect 20158 10810 20192 10826
rect 20158 10618 20192 10634
rect 20276 10810 20310 10826
rect 20276 10618 20310 10634
rect 20394 10810 20428 10826
rect 20394 10618 20428 10634
rect 20617 10810 20651 10864
rect 20617 10618 20651 10634
rect 20735 10810 20769 10826
rect 20735 10618 20769 10634
rect 20853 10810 20887 10864
rect 20853 10618 20887 10634
rect 20971 10810 21005 10826
rect 20971 10618 21005 10634
rect 21101 10618 21135 10634
rect 21219 11010 21253 11026
rect 21219 10618 21253 10634
rect 21337 11010 21371 11026
rect 21337 10618 21371 10634
rect 21455 11010 21489 11063
rect 21455 10618 21489 10634
rect 21573 11010 21607 11026
rect 21573 10618 21607 10634
rect 21691 11010 21725 11063
rect 24117 11058 24151 11074
rect 21691 10618 21725 10634
rect 21809 11010 21843 11026
rect 21809 10618 21843 10634
rect 21938 10810 21972 10826
rect 21938 10618 21972 10634
rect 22056 10810 22090 10826
rect 22056 10618 22090 10634
rect 22174 10810 22208 10826
rect 22174 10618 22208 10634
rect 22292 10810 22326 10826
rect 24117 10666 24151 10682
rect 24235 11058 24269 11074
rect 24235 10666 24269 10682
rect 24353 11058 24387 11074
rect 24470 11058 24504 11074
rect 24470 10866 24504 10882
rect 24588 11058 24622 11074
rect 24588 10866 24622 10882
rect 25344 10932 25614 10967
rect 25344 10878 25378 10932
rect 24353 10666 24387 10682
rect 24640 10732 24889 10775
rect 22292 10618 22326 10634
rect 24640 10642 24687 10732
rect 24850 10642 24889 10732
rect 25344 10686 25378 10702
rect 25462 10878 25496 10894
rect 25462 10686 25496 10702
rect 25580 10878 25614 10932
rect 25580 10686 25614 10702
rect 25698 10878 25732 10894
rect 25698 10686 25732 10702
rect 25828 10686 25862 10702
rect 25946 11078 25980 11094
rect 25946 10686 25980 10702
rect 26064 11078 26098 11094
rect 26064 10686 26098 10702
rect 26182 11078 26216 11131
rect 26182 10686 26216 10702
rect 26300 11078 26334 11094
rect 26300 10686 26334 10702
rect 26418 11078 26452 11131
rect 28080 11131 28350 11166
rect 26418 10686 26452 10702
rect 26536 11078 26570 11094
rect 27726 11078 27760 11094
rect 27242 10932 27512 10967
rect 26536 10686 26570 10702
rect 26665 10878 26699 10894
rect 26665 10686 26699 10702
rect 26783 10878 26817 10894
rect 26783 10686 26817 10702
rect 26901 10878 26935 10894
rect 26901 10686 26935 10702
rect 27019 10878 27053 10894
rect 27019 10686 27053 10702
rect 27242 10878 27276 10932
rect 27242 10686 27276 10702
rect 27360 10878 27394 10894
rect 27360 10686 27394 10702
rect 27478 10878 27512 10932
rect 27478 10686 27512 10702
rect 27596 10878 27630 10894
rect 27596 10686 27630 10702
rect 27726 10686 27760 10702
rect 27844 11078 27878 11094
rect 27844 10686 27878 10702
rect 27962 11078 27996 11094
rect 27962 10686 27996 10702
rect 28080 11078 28114 11131
rect 28080 10686 28114 10702
rect 28198 11078 28232 11094
rect 28198 10686 28232 10702
rect 28316 11078 28350 11131
rect 28316 10686 28350 10702
rect 28434 11078 28468 11094
rect 28434 10686 28468 10702
rect 28563 10878 28597 10894
rect 28563 10686 28597 10702
rect 28681 10878 28715 10894
rect 28681 10686 28715 10702
rect 28799 10878 28833 10894
rect 28799 10686 28833 10702
rect 28917 10878 28951 10894
rect 28917 10686 28951 10702
rect 24160 10598 24176 10632
rect 24210 10598 24226 10632
rect 24278 10598 24294 10632
rect 24328 10598 24344 10632
rect 24640 10603 24889 10642
rect 17535 10530 17551 10564
rect 17585 10530 17601 10564
rect 17653 10530 17669 10564
rect 17703 10530 17719 10564
rect 18015 10535 18264 10574
rect 16386 10501 16612 10513
rect 3141 10481 3403 10491
rect 3141 8083 3305 10481
rect 13529 10464 13563 10480
rect 13529 10414 13563 10430
rect 15619 10443 15686 10459
rect 15619 10409 15636 10443
rect 15670 10409 15686 10443
rect 6980 10376 7014 10392
rect 12492 10385 12526 10401
rect 6980 10326 7014 10342
rect 9070 10355 9137 10371
rect 9070 10321 9087 10355
rect 9121 10321 9137 10355
rect 5943 10297 5977 10313
rect 4442 10217 4665 10293
rect 4442 10068 4521 10217
rect 4588 10215 4665 10217
rect 4442 10066 4523 10068
rect 4590 10066 4665 10215
rect 4442 9962 4665 10066
rect 6061 10297 6095 10313
rect 5943 9905 5977 9921
rect 6060 9921 6061 9968
rect 6179 10297 6213 10313
rect 6095 9921 6096 9968
rect 4873 9853 5143 9887
rect 4047 9803 4081 9819
rect 4047 9611 4081 9627
rect 4165 9803 4199 9819
rect 4165 9611 4199 9627
rect 4283 9803 4317 9819
rect 4283 9611 4317 9627
rect 4401 9803 4435 9819
rect 4401 9611 4435 9627
rect 4519 9803 4553 9819
rect 4519 9611 4553 9627
rect 4637 9803 4671 9819
rect 4637 9611 4671 9627
rect 4755 9803 4789 9819
rect 4755 9611 4789 9627
rect 4873 9803 4907 9853
rect 4873 9611 4907 9627
rect 4991 9803 5025 9819
rect 4991 9611 5025 9627
rect 5109 9803 5143 9853
rect 6060 9863 6096 9921
rect 6297 10297 6331 10313
rect 6179 9905 6213 9921
rect 6295 9921 6297 9968
rect 6295 9863 6331 9921
rect 6415 10297 6449 10313
rect 6415 9905 6449 9921
rect 6533 10297 6567 10313
rect 6651 10297 6685 10313
rect 6567 9921 6569 9967
rect 6533 9863 6569 9921
rect 6651 9905 6685 9921
rect 7841 10297 7875 10313
rect 7959 10297 7993 10313
rect 7841 9905 7875 9921
rect 7958 9921 7959 9968
rect 8077 10297 8111 10313
rect 7993 9921 7994 9968
rect 7156 9863 7653 9881
rect 6060 9860 7653 9863
rect 6060 9826 7601 9860
rect 7635 9826 7653 9860
rect 6060 9823 7653 9826
rect 7958 9863 7994 9921
rect 8195 10297 8229 10313
rect 8077 9905 8111 9921
rect 8193 9921 8195 9968
rect 8193 9863 8229 9921
rect 8313 10297 8347 10313
rect 8313 9905 8347 9921
rect 8431 10297 8465 10313
rect 8549 10297 8583 10313
rect 9070 10305 9137 10321
rect 10991 10308 11214 10381
rect 8465 9921 8467 9967
rect 8431 9863 8467 9921
rect 10991 10159 11068 10308
rect 11135 10305 11214 10308
rect 10991 10156 11070 10159
rect 11137 10156 11214 10305
rect 10991 10050 11214 10156
rect 12610 10385 12644 10401
rect 12492 9993 12526 10009
rect 12609 10009 12610 10056
rect 12728 10385 12762 10401
rect 12644 10009 12645 10056
rect 8549 9905 8583 9921
rect 11422 9941 11692 9975
rect 9054 9863 9317 9893
rect 7958 9823 9317 9863
rect 6079 9822 7653 9823
rect 7977 9822 9317 9823
rect 5957 9733 6024 9749
rect 5957 9699 5973 9733
rect 6007 9699 6024 9733
rect 5957 9683 6024 9699
rect 5109 9611 5143 9627
rect 5788 9666 5822 9682
rect 5788 9616 5822 9632
rect 6134 9581 6168 9822
rect 7156 9805 7653 9822
rect 6604 9733 6671 9749
rect 6604 9699 6621 9733
rect 6655 9699 6671 9733
rect 6604 9683 6671 9699
rect 7855 9733 7922 9749
rect 7855 9699 7871 9733
rect 7905 9699 7922 9733
rect 7855 9683 7922 9699
rect 6911 9665 6945 9681
rect 6223 9615 6239 9649
rect 6273 9615 6289 9649
rect 6341 9616 6357 9650
rect 6391 9616 6407 9650
rect 6911 9615 6945 9631
rect 7686 9666 7720 9682
rect 7686 9616 7720 9632
rect 8032 9581 8066 9822
rect 9054 9793 9317 9822
rect 8500 9734 8567 9750
rect 8500 9700 8517 9734
rect 8551 9700 8567 9734
rect 8500 9684 8567 9700
rect 8809 9665 8843 9681
rect 8121 9615 8137 9649
rect 8171 9615 8187 9649
rect 8239 9616 8255 9650
rect 8289 9616 8305 9650
rect 8809 9615 8843 9631
rect 4798 9533 4814 9567
rect 4848 9533 4864 9567
rect 5641 9565 5675 9581
rect 4680 9416 4696 9450
rect 4730 9416 4746 9450
rect 4284 9366 4318 9382
rect 4284 8974 4318 8990
rect 4402 9366 4436 9382
rect 4402 8974 4436 8990
rect 4520 9366 4554 9382
rect 4637 9366 4671 9382
rect 4637 9174 4671 9190
rect 4755 9366 4789 9382
rect 5641 9373 5675 9389
rect 5759 9565 5793 9581
rect 5759 9373 5793 9389
rect 6061 9565 6095 9581
rect 4755 9174 4789 9190
rect 6134 9565 6213 9581
rect 6134 9535 6179 9565
rect 6061 9122 6096 9189
rect 6179 9173 6213 9189
rect 6297 9565 6331 9581
rect 6297 9173 6331 9189
rect 6415 9565 6449 9581
rect 6533 9565 6567 9581
rect 6939 9565 6973 9581
rect 6939 9373 6973 9389
rect 7057 9565 7091 9581
rect 7057 9373 7091 9389
rect 7539 9565 7573 9581
rect 7539 9373 7573 9389
rect 7657 9565 7691 9581
rect 7657 9373 7691 9389
rect 7959 9565 7993 9581
rect 6415 9173 6449 9189
rect 6532 9122 6567 9189
rect 6061 9087 6567 9122
rect 8032 9565 8111 9581
rect 8032 9535 8077 9565
rect 7959 9122 7994 9189
rect 8077 9173 8111 9189
rect 8195 9565 8229 9581
rect 8195 9173 8229 9189
rect 8313 9565 8347 9581
rect 8431 9565 8465 9581
rect 8837 9565 8871 9581
rect 8837 9373 8871 9389
rect 8955 9565 8989 9581
rect 8955 9373 8989 9389
rect 8313 9173 8347 9189
rect 8430 9122 8465 9189
rect 7959 9087 8465 9122
rect 4520 8974 4554 8990
rect 4807 9040 5056 9083
rect 4807 8950 4854 9040
rect 5017 8950 5056 9040
rect 4327 8906 4343 8940
rect 4377 8906 4393 8940
rect 4445 8906 4461 8940
rect 4495 8906 4511 8940
rect 4807 8911 5056 8950
rect 6232 8880 6404 8927
rect 6232 8717 6271 8880
rect 6361 8717 6404 8880
rect 6232 8677 6404 8717
rect 9185 8335 9317 9793
rect 10596 9891 10630 9907
rect 10596 9699 10630 9715
rect 10714 9891 10748 9907
rect 10714 9699 10748 9715
rect 10832 9891 10866 9907
rect 10832 9699 10866 9715
rect 10950 9891 10984 9907
rect 10950 9699 10984 9715
rect 11068 9891 11102 9907
rect 11068 9699 11102 9715
rect 11186 9891 11220 9907
rect 11186 9699 11220 9715
rect 11304 9891 11338 9907
rect 11304 9699 11338 9715
rect 11422 9891 11456 9941
rect 11422 9699 11456 9715
rect 11540 9891 11574 9907
rect 11540 9699 11574 9715
rect 11658 9891 11692 9941
rect 12609 9951 12645 10009
rect 12846 10385 12880 10401
rect 12728 9993 12762 10009
rect 12844 10009 12846 10056
rect 12844 9951 12880 10009
rect 12964 10385 12998 10401
rect 12964 9993 12998 10009
rect 13082 10385 13116 10401
rect 13200 10385 13234 10401
rect 13116 10009 13118 10055
rect 13082 9951 13118 10009
rect 13200 9993 13234 10009
rect 14390 10385 14424 10401
rect 14508 10385 14542 10401
rect 14390 9993 14424 10009
rect 14507 10009 14508 10056
rect 14626 10385 14660 10401
rect 14542 10009 14543 10056
rect 13705 9951 14202 9969
rect 12609 9948 14202 9951
rect 12609 9914 14150 9948
rect 14184 9914 14202 9948
rect 12609 9911 14202 9914
rect 14507 9951 14543 10009
rect 14744 10385 14778 10401
rect 14626 9993 14660 10009
rect 14742 10009 14744 10056
rect 14742 9951 14778 10009
rect 14862 10385 14896 10401
rect 14862 9993 14896 10009
rect 14980 10385 15014 10401
rect 15098 10385 15132 10401
rect 15619 10393 15686 10409
rect 15014 10009 15016 10055
rect 14980 9951 15016 10009
rect 15098 9993 15132 10009
rect 15603 9980 15703 9981
rect 15603 9951 15759 9980
rect 14507 9911 15759 9951
rect 12628 9910 14202 9911
rect 14526 9910 15759 9911
rect 12506 9821 12573 9837
rect 12506 9787 12522 9821
rect 12556 9787 12573 9821
rect 12506 9771 12573 9787
rect 11658 9699 11692 9715
rect 12337 9754 12371 9770
rect 12337 9704 12371 9720
rect 12683 9669 12717 9910
rect 13705 9893 14202 9910
rect 13153 9821 13220 9837
rect 13153 9787 13170 9821
rect 13204 9787 13220 9821
rect 13153 9771 13220 9787
rect 14404 9821 14471 9837
rect 14404 9787 14420 9821
rect 14454 9787 14471 9821
rect 14404 9771 14471 9787
rect 13460 9753 13494 9769
rect 12772 9703 12788 9737
rect 12822 9703 12838 9737
rect 12890 9704 12906 9738
rect 12940 9704 12956 9738
rect 13460 9703 13494 9719
rect 14235 9754 14269 9770
rect 14235 9704 14269 9720
rect 14581 9669 14615 9910
rect 15603 9882 15759 9910
rect 15603 9881 15703 9882
rect 15049 9822 15116 9838
rect 15049 9788 15066 9822
rect 15100 9788 15116 9822
rect 15049 9772 15116 9788
rect 15358 9753 15392 9769
rect 14670 9703 14686 9737
rect 14720 9703 14736 9737
rect 14788 9704 14804 9738
rect 14838 9704 14854 9738
rect 15358 9703 15392 9719
rect 11347 9621 11363 9655
rect 11397 9621 11413 9655
rect 12190 9653 12224 9669
rect 11229 9504 11245 9538
rect 11279 9504 11295 9538
rect 10833 9454 10867 9470
rect 10833 9062 10867 9078
rect 10951 9454 10985 9470
rect 10951 9062 10985 9078
rect 11069 9454 11103 9470
rect 11186 9454 11220 9470
rect 11186 9262 11220 9278
rect 11304 9454 11338 9470
rect 12190 9461 12224 9477
rect 12308 9653 12342 9669
rect 12308 9461 12342 9477
rect 12610 9653 12644 9669
rect 11304 9262 11338 9278
rect 12683 9653 12762 9669
rect 12683 9623 12728 9653
rect 12610 9210 12645 9277
rect 12728 9261 12762 9277
rect 12846 9653 12880 9669
rect 12846 9261 12880 9277
rect 12964 9653 12998 9669
rect 13082 9653 13116 9669
rect 13488 9653 13522 9669
rect 13488 9461 13522 9477
rect 13606 9653 13640 9669
rect 13606 9461 13640 9477
rect 14088 9653 14122 9669
rect 14088 9461 14122 9477
rect 14206 9653 14240 9669
rect 14206 9461 14240 9477
rect 14508 9653 14542 9669
rect 12964 9261 12998 9277
rect 13081 9210 13116 9277
rect 12610 9175 13116 9210
rect 14581 9653 14660 9669
rect 14581 9623 14626 9653
rect 14508 9210 14543 9277
rect 14626 9261 14660 9277
rect 14744 9653 14778 9669
rect 14744 9261 14778 9277
rect 14862 9653 14896 9669
rect 14980 9653 15014 9669
rect 15386 9653 15420 9669
rect 15386 9461 15420 9477
rect 15504 9653 15538 9669
rect 15504 9461 15538 9477
rect 14862 9261 14896 9277
rect 14979 9210 15014 9277
rect 14508 9175 15014 9210
rect 11069 9062 11103 9078
rect 11356 9128 11605 9171
rect 11356 9038 11403 9128
rect 11566 9038 11605 9128
rect 10876 8994 10892 9028
rect 10926 8994 10942 9028
rect 10994 8994 11010 9028
rect 11044 8994 11060 9028
rect 11356 8999 11605 9038
rect 12781 8968 12953 9015
rect 12781 8805 12820 8968
rect 12910 8805 12953 8968
rect 12781 8765 12953 8805
rect 16387 8565 16550 10501
rect 26808 10464 26842 10480
rect 26808 10414 26842 10430
rect 28898 10443 28965 10459
rect 20183 10396 20217 10412
rect 28898 10409 28915 10443
rect 28949 10409 28965 10443
rect 20183 10346 20217 10362
rect 22273 10375 22340 10391
rect 25771 10385 25805 10401
rect 22273 10341 22290 10375
rect 22324 10341 22340 10375
rect 19146 10317 19180 10333
rect 17645 10239 17868 10313
rect 17645 10237 17725 10239
rect 17645 10088 17724 10237
rect 17792 10090 17868 10239
rect 17791 10088 17868 10090
rect 17645 9982 17868 10088
rect 19264 10317 19298 10333
rect 19146 9925 19180 9941
rect 19263 9941 19264 9988
rect 19382 10317 19416 10333
rect 19298 9941 19299 9988
rect 18076 9873 18346 9907
rect 17250 9823 17284 9839
rect 17250 9631 17284 9647
rect 17368 9823 17402 9839
rect 17368 9631 17402 9647
rect 17486 9823 17520 9839
rect 17486 9631 17520 9647
rect 17604 9823 17638 9839
rect 17604 9631 17638 9647
rect 17722 9823 17756 9839
rect 17722 9631 17756 9647
rect 17840 9823 17874 9839
rect 17840 9631 17874 9647
rect 17958 9823 17992 9839
rect 17958 9631 17992 9647
rect 18076 9823 18110 9873
rect 18076 9631 18110 9647
rect 18194 9823 18228 9839
rect 18194 9631 18228 9647
rect 18312 9823 18346 9873
rect 19263 9883 19299 9941
rect 19500 10317 19534 10333
rect 19382 9925 19416 9941
rect 19498 9941 19500 9988
rect 19498 9883 19534 9941
rect 19618 10317 19652 10333
rect 19618 9925 19652 9941
rect 19736 10317 19770 10333
rect 19854 10317 19888 10333
rect 19770 9941 19772 9987
rect 19736 9883 19772 9941
rect 19854 9925 19888 9941
rect 21044 10317 21078 10333
rect 21162 10317 21196 10333
rect 21044 9925 21078 9941
rect 21161 9941 21162 9988
rect 21280 10317 21314 10333
rect 21196 9941 21197 9988
rect 20359 9883 20856 9901
rect 19263 9880 20856 9883
rect 19263 9846 20804 9880
rect 20838 9846 20856 9880
rect 19263 9843 20856 9846
rect 21161 9883 21197 9941
rect 21398 10317 21432 10333
rect 21280 9925 21314 9941
rect 21396 9941 21398 9988
rect 21396 9883 21432 9941
rect 21516 10317 21550 10333
rect 21516 9925 21550 9941
rect 21634 10317 21668 10333
rect 21752 10317 21786 10333
rect 22273 10325 22340 10341
rect 21668 9941 21670 9987
rect 21634 9883 21670 9941
rect 24270 10305 24493 10381
rect 24270 10156 24349 10305
rect 24416 10300 24493 10305
rect 24270 10151 24350 10156
rect 24417 10151 24493 10300
rect 24270 10050 24493 10151
rect 25889 10385 25923 10401
rect 25771 9993 25805 10009
rect 25888 10009 25889 10056
rect 26007 10385 26041 10401
rect 25923 10009 25924 10056
rect 21752 9925 21786 9941
rect 24701 9941 24971 9975
rect 22867 9914 22976 9920
rect 22343 9913 22976 9914
rect 22257 9911 22976 9913
rect 22257 9883 22874 9911
rect 21161 9843 22874 9883
rect 19282 9842 20856 9843
rect 21180 9842 22874 9843
rect 19160 9753 19227 9769
rect 19160 9719 19176 9753
rect 19210 9719 19227 9753
rect 19160 9703 19227 9719
rect 18312 9631 18346 9647
rect 18991 9686 19025 9702
rect 18991 9636 19025 9652
rect 19337 9601 19371 9842
rect 20359 9825 20856 9842
rect 19807 9753 19874 9769
rect 19807 9719 19824 9753
rect 19858 9719 19874 9753
rect 19807 9703 19874 9719
rect 21058 9753 21125 9769
rect 21058 9719 21074 9753
rect 21108 9719 21125 9753
rect 21058 9703 21125 9719
rect 20114 9685 20148 9701
rect 19426 9635 19442 9669
rect 19476 9635 19492 9669
rect 19544 9636 19560 9670
rect 19594 9636 19610 9670
rect 20114 9635 20148 9651
rect 20889 9686 20923 9702
rect 20889 9636 20923 9652
rect 21235 9601 21269 9842
rect 22257 9813 22874 9842
rect 22343 9812 22874 9813
rect 22867 9811 22874 9812
rect 22970 9811 22976 9911
rect 22867 9805 22976 9811
rect 23875 9891 23909 9907
rect 21703 9754 21770 9770
rect 21703 9720 21720 9754
rect 21754 9720 21770 9754
rect 21703 9704 21770 9720
rect 22012 9685 22046 9701
rect 23875 9699 23909 9715
rect 23993 9891 24027 9907
rect 23993 9699 24027 9715
rect 24111 9891 24145 9907
rect 24111 9699 24145 9715
rect 24229 9891 24263 9907
rect 24229 9699 24263 9715
rect 24347 9891 24381 9907
rect 24347 9699 24381 9715
rect 24465 9891 24499 9907
rect 24465 9699 24499 9715
rect 24583 9891 24617 9907
rect 24583 9699 24617 9715
rect 24701 9891 24735 9941
rect 24701 9699 24735 9715
rect 24819 9891 24853 9907
rect 24819 9699 24853 9715
rect 24937 9891 24971 9941
rect 25888 9951 25924 10009
rect 26125 10385 26159 10401
rect 26007 9993 26041 10009
rect 26123 10009 26125 10056
rect 26123 9951 26159 10009
rect 26243 10385 26277 10401
rect 26243 9993 26277 10009
rect 26361 10385 26395 10401
rect 26479 10385 26513 10401
rect 26395 10009 26397 10055
rect 26361 9951 26397 10009
rect 26479 9993 26513 10009
rect 27669 10385 27703 10401
rect 27787 10385 27821 10401
rect 27669 9993 27703 10009
rect 27786 10009 27787 10056
rect 27905 10385 27939 10401
rect 27821 10009 27822 10056
rect 26984 9951 27481 9969
rect 25888 9948 27481 9951
rect 25888 9914 27429 9948
rect 27463 9914 27481 9948
rect 25888 9911 27481 9914
rect 27786 9951 27822 10009
rect 28023 10385 28057 10401
rect 27905 9993 27939 10009
rect 28021 10009 28023 10056
rect 28021 9951 28057 10009
rect 28141 10385 28175 10401
rect 28141 9993 28175 10009
rect 28259 10385 28293 10401
rect 28377 10385 28411 10401
rect 28898 10393 28965 10409
rect 28293 10009 28295 10055
rect 28259 9951 28295 10009
rect 28377 9993 28411 10009
rect 28882 9980 28982 9981
rect 28882 9951 29038 9980
rect 27786 9911 29038 9951
rect 25907 9910 27481 9911
rect 27805 9910 29038 9911
rect 25785 9821 25852 9837
rect 25785 9787 25801 9821
rect 25835 9787 25852 9821
rect 25785 9771 25852 9787
rect 24937 9699 24971 9715
rect 25616 9754 25650 9770
rect 25616 9704 25650 9720
rect 21324 9635 21340 9669
rect 21374 9635 21390 9669
rect 21442 9636 21458 9670
rect 21492 9636 21508 9670
rect 25962 9669 25996 9910
rect 26984 9893 27481 9910
rect 26432 9821 26499 9837
rect 26432 9787 26449 9821
rect 26483 9787 26499 9821
rect 26432 9771 26499 9787
rect 27683 9821 27750 9837
rect 27683 9787 27699 9821
rect 27733 9787 27750 9821
rect 27683 9771 27750 9787
rect 26739 9753 26773 9769
rect 26051 9703 26067 9737
rect 26101 9703 26117 9737
rect 26169 9704 26185 9738
rect 26219 9704 26235 9738
rect 26739 9703 26773 9719
rect 27514 9754 27548 9770
rect 27514 9704 27548 9720
rect 27860 9669 27894 9910
rect 28882 9882 29038 9910
rect 28882 9881 28982 9882
rect 28328 9822 28395 9838
rect 28328 9788 28345 9822
rect 28379 9788 28395 9822
rect 28328 9772 28395 9788
rect 28637 9753 28671 9769
rect 27949 9703 27965 9737
rect 27999 9703 28015 9737
rect 28067 9704 28083 9738
rect 28117 9704 28133 9738
rect 28637 9703 28671 9719
rect 29952 9713 30120 9729
rect 22012 9635 22046 9651
rect 24626 9621 24642 9655
rect 24676 9621 24692 9655
rect 25469 9653 25503 9669
rect 18001 9553 18017 9587
rect 18051 9553 18067 9587
rect 18844 9585 18878 9601
rect 17883 9436 17899 9470
rect 17933 9436 17949 9470
rect 17487 9386 17521 9402
rect 17487 8994 17521 9010
rect 17605 9386 17639 9402
rect 17605 8994 17639 9010
rect 17723 9386 17757 9402
rect 17840 9386 17874 9402
rect 17840 9194 17874 9210
rect 17958 9386 17992 9402
rect 18844 9393 18878 9409
rect 18962 9585 18996 9601
rect 18962 9393 18996 9409
rect 19264 9585 19298 9601
rect 17958 9194 17992 9210
rect 19337 9585 19416 9601
rect 19337 9555 19382 9585
rect 19264 9142 19299 9209
rect 19382 9193 19416 9209
rect 19500 9585 19534 9601
rect 19500 9193 19534 9209
rect 19618 9585 19652 9601
rect 19736 9585 19770 9601
rect 20142 9585 20176 9601
rect 20142 9393 20176 9409
rect 20260 9585 20294 9601
rect 20260 9393 20294 9409
rect 20742 9585 20776 9601
rect 20742 9393 20776 9409
rect 20860 9585 20894 9601
rect 20860 9393 20894 9409
rect 21162 9585 21196 9601
rect 19618 9193 19652 9209
rect 19735 9142 19770 9209
rect 19264 9107 19770 9142
rect 21235 9585 21314 9601
rect 21235 9555 21280 9585
rect 21162 9142 21197 9209
rect 21280 9193 21314 9209
rect 21398 9585 21432 9601
rect 21398 9193 21432 9209
rect 21516 9585 21550 9601
rect 21634 9585 21668 9601
rect 22040 9585 22074 9601
rect 22040 9393 22074 9409
rect 22158 9585 22192 9601
rect 24508 9504 24524 9538
rect 24558 9504 24574 9538
rect 22158 9393 22192 9409
rect 24112 9454 24146 9470
rect 21516 9193 21550 9209
rect 21633 9142 21668 9209
rect 21162 9107 21668 9142
rect 17723 8994 17757 9010
rect 18010 9060 18259 9103
rect 24112 9062 24146 9078
rect 24230 9454 24264 9470
rect 24230 9062 24264 9078
rect 24348 9454 24382 9470
rect 24465 9454 24499 9470
rect 24465 9262 24499 9278
rect 24583 9454 24617 9470
rect 25469 9461 25503 9477
rect 25587 9653 25621 9669
rect 25587 9461 25621 9477
rect 25889 9653 25923 9669
rect 24583 9262 24617 9278
rect 25962 9653 26041 9669
rect 25962 9623 26007 9653
rect 25889 9210 25924 9277
rect 26007 9261 26041 9277
rect 26125 9653 26159 9669
rect 26125 9261 26159 9277
rect 26243 9653 26277 9669
rect 26361 9653 26395 9669
rect 26767 9653 26801 9669
rect 26767 9461 26801 9477
rect 26885 9653 26919 9669
rect 26885 9461 26919 9477
rect 27367 9653 27401 9669
rect 27367 9461 27401 9477
rect 27485 9653 27519 9669
rect 27485 9461 27519 9477
rect 27787 9653 27821 9669
rect 26243 9261 26277 9277
rect 26360 9210 26395 9277
rect 25889 9175 26395 9210
rect 27860 9653 27939 9669
rect 27860 9623 27905 9653
rect 27787 9210 27822 9277
rect 27905 9261 27939 9277
rect 28023 9653 28057 9669
rect 28023 9261 28057 9277
rect 28141 9653 28175 9669
rect 28259 9653 28293 9669
rect 28665 9653 28699 9669
rect 28665 9461 28699 9477
rect 28783 9653 28817 9669
rect 29952 9643 29968 9713
rect 30104 9643 30120 9713
rect 29952 9627 30120 9643
rect 30489 9523 30759 9557
rect 28783 9461 28817 9477
rect 29663 9473 29697 9489
rect 29663 9281 29697 9297
rect 29781 9473 29815 9489
rect 29781 9281 29815 9297
rect 29899 9473 29933 9489
rect 29899 9281 29933 9297
rect 30017 9473 30051 9489
rect 30017 9281 30051 9297
rect 30135 9473 30169 9489
rect 30135 9281 30169 9297
rect 30253 9473 30287 9489
rect 30253 9281 30287 9297
rect 30371 9473 30405 9489
rect 30371 9281 30405 9297
rect 30489 9473 30523 9523
rect 30489 9281 30523 9297
rect 30607 9473 30641 9489
rect 30607 9281 30641 9297
rect 30725 9473 30759 9523
rect 30725 9281 30759 9297
rect 28141 9261 28175 9277
rect 28258 9210 28293 9277
rect 27787 9175 28293 9210
rect 30414 9203 30430 9237
rect 30464 9203 30480 9237
rect 24348 9062 24382 9078
rect 24635 9128 24884 9171
rect 18010 8970 18057 9060
rect 18220 8970 18259 9060
rect 24635 9038 24682 9128
rect 24845 9038 24884 9128
rect 30296 9086 30312 9120
rect 30346 9086 30362 9120
rect 24155 8994 24171 9028
rect 24205 8994 24221 9028
rect 24273 8994 24289 9028
rect 24323 8994 24339 9028
rect 24635 8999 24884 9038
rect 29900 9036 29934 9052
rect 17530 8926 17546 8960
rect 17580 8926 17596 8960
rect 17648 8926 17664 8960
rect 17698 8926 17714 8960
rect 18010 8931 18259 8970
rect 26060 8968 26232 9015
rect 19435 8900 19607 8947
rect 19435 8737 19474 8900
rect 19564 8737 19607 8900
rect 26060 8805 26099 8968
rect 26189 8805 26232 8968
rect 26060 8765 26232 8805
rect 19435 8697 19607 8737
rect 29900 8644 29934 8660
rect 30018 9036 30052 9052
rect 30018 8644 30052 8660
rect 30136 9036 30170 9052
rect 30253 9036 30287 9052
rect 30253 8844 30287 8860
rect 30371 9036 30405 9052
rect 30371 8844 30405 8860
rect 30136 8644 30170 8660
rect 16387 8497 16431 8565
rect 16501 8497 16550 8565
rect 16387 8481 16550 8497
rect 22383 8590 23655 8617
rect 22383 8491 22414 8590
rect 22520 8491 23523 8590
rect 23629 8491 23655 8590
rect 29943 8576 29959 8610
rect 29993 8576 30009 8610
rect 30061 8576 30077 8610
rect 30111 8576 30127 8610
rect 22383 8464 23655 8491
rect 30176 8505 30344 8523
rect 30176 8449 30192 8505
rect 30326 8449 30344 8505
rect 30176 8433 30344 8449
rect 16405 8337 28677 8338
rect 31205 8337 31324 14134
rect 32021 14179 32055 14195
rect 31903 13787 31937 13803
rect 32020 13803 32021 13850
rect 32139 14179 32173 14195
rect 32055 13803 32056 13850
rect 32020 13745 32056 13803
rect 32257 14179 32291 14195
rect 32139 13787 32173 13803
rect 32255 13803 32257 13850
rect 32255 13745 32291 13803
rect 32375 14179 32409 14195
rect 32375 13787 32409 13803
rect 32493 14179 32527 14195
rect 32611 14179 32645 14195
rect 32527 13803 32529 13849
rect 32493 13745 32529 13803
rect 32773 13974 32843 13978
rect 32773 13883 32777 13974
rect 32839 13883 32843 13974
rect 32773 13878 32843 13883
rect 32611 13787 32645 13803
rect 32788 13745 32829 13878
rect 33506 13840 33540 13856
rect 33624 14232 33658 14248
rect 33624 13840 33658 13856
rect 33742 14232 33776 14248
rect 33859 14232 33893 14248
rect 33859 14040 33893 14056
rect 33977 14232 34011 14248
rect 33977 14040 34011 14056
rect 34779 13985 34897 19035
rect 37723 19011 37812 19035
rect 37723 18962 37737 19011
rect 37797 18962 37812 19011
rect 37723 18946 37812 18962
rect 36873 18838 36963 18872
rect 37139 18838 37155 18872
rect 36873 18636 36912 18838
rect 37437 18767 37522 18783
rect 36947 18720 36963 18754
rect 37139 18720 37229 18754
rect 36873 18602 36963 18636
rect 37139 18602 37155 18636
rect 37190 18518 37229 18720
rect 37437 18707 37454 18767
rect 37509 18707 37522 18767
rect 37437 18691 37522 18707
rect 36947 18484 36963 18518
rect 37139 18484 37229 18518
rect 36671 18397 36763 18431
rect 37139 18397 37155 18431
rect 36671 18195 36710 18397
rect 36747 18279 36763 18313
rect 37139 18279 37229 18313
rect 36671 18161 36763 18195
rect 37139 18161 37155 18195
rect 37190 18077 37229 18279
rect 36747 18043 36763 18077
rect 37139 18043 37229 18077
rect 36672 17930 36763 17964
rect 37139 17930 37155 17964
rect 36672 17728 36711 17930
rect 37190 17846 37229 18043
rect 38080 18004 38096 18038
rect 38272 18004 38288 18038
rect 38080 17886 38096 17920
rect 38272 17886 38288 17920
rect 38084 17846 38284 17886
rect 36747 17812 36763 17846
rect 37139 17812 37229 17846
rect 36475 17686 36585 17702
rect 36672 17694 36763 17728
rect 37139 17694 37155 17728
rect 36475 17490 36493 17686
rect 36569 17490 36585 17686
rect 37190 17610 37229 17812
rect 37725 17800 37810 17816
rect 38080 17812 38096 17846
rect 38472 17812 38488 17846
rect 37338 17752 37354 17786
rect 37388 17752 37404 17786
rect 37725 17740 37738 17800
rect 37793 17740 37810 17800
rect 37725 17724 37810 17740
rect 36747 17576 36763 17610
rect 37139 17576 37229 17610
rect 37440 17682 37525 17698
rect 38080 17694 38096 17728
rect 38472 17694 38488 17728
rect 37440 17622 37453 17682
rect 37508 17622 37525 17682
rect 38721 17628 38807 17644
rect 37440 17606 37525 17622
rect 38080 17576 38096 17610
rect 38472 17576 38488 17610
rect 38573 17609 38607 17625
rect 36475 17474 36585 17490
rect 36672 17458 36763 17492
rect 37139 17458 37155 17492
rect 36672 17256 36711 17458
rect 37190 17374 37229 17576
rect 38573 17559 38607 17575
rect 38721 17606 38739 17628
rect 37958 17517 37974 17551
rect 38008 17517 38024 17551
rect 38721 17548 38725 17606
rect 38721 17524 38739 17548
rect 38785 17524 38807 17628
rect 38721 17508 38807 17524
rect 38080 17458 38096 17492
rect 38472 17458 38488 17492
rect 37568 17398 37584 17432
rect 37618 17398 37634 17432
rect 36747 17340 36763 17374
rect 37139 17340 37229 17374
rect 38080 17340 38096 17374
rect 38472 17340 38488 17374
rect 36672 17222 36763 17256
rect 37139 17222 37155 17256
rect 37190 17137 37229 17340
rect 38084 17296 38284 17340
rect 38080 17262 38096 17296
rect 38272 17262 38288 17296
rect 38080 17144 38096 17178
rect 38272 17144 38288 17178
rect 36747 17103 36763 17137
rect 37139 17103 37229 17137
rect 36672 16985 36763 17019
rect 37139 16985 37155 17019
rect 36672 16783 36711 16985
rect 37190 16901 37229 17103
rect 36747 16867 36763 16901
rect 37139 16867 37229 16901
rect 36672 16749 36763 16783
rect 37139 16749 37155 16783
rect 36947 16630 36963 16664
rect 37139 16630 37232 16664
rect 36876 16512 36963 16546
rect 37139 16512 37155 16546
rect 36876 16310 36913 16512
rect 37193 16428 37232 16630
rect 36947 16394 36963 16428
rect 37139 16394 37232 16428
rect 37313 16476 37347 16492
rect 37313 16426 37347 16442
rect 36876 16276 36963 16310
rect 37139 16276 37155 16310
rect 36873 15694 36963 15728
rect 37139 15694 37155 15728
rect 36873 15492 36912 15694
rect 37437 15623 37522 15639
rect 36947 15576 36963 15610
rect 37139 15576 37229 15610
rect 36873 15458 36963 15492
rect 37139 15458 37155 15492
rect 37190 15374 37229 15576
rect 37437 15563 37454 15623
rect 37509 15563 37522 15623
rect 37437 15547 37522 15563
rect 36947 15340 36963 15374
rect 37139 15340 37229 15374
rect 36671 15253 36763 15287
rect 37139 15253 37155 15287
rect 36671 15051 36710 15253
rect 36747 15135 36763 15169
rect 37139 15135 37229 15169
rect 36671 15017 36763 15051
rect 37139 15017 37155 15051
rect 37190 14933 37229 15135
rect 36747 14899 36763 14933
rect 37139 14899 37229 14933
rect 36672 14786 36763 14820
rect 37139 14786 37155 14820
rect 36672 14584 36711 14786
rect 37190 14702 37229 14899
rect 38080 14860 38096 14894
rect 38272 14860 38288 14894
rect 38080 14742 38096 14776
rect 38272 14742 38288 14776
rect 38084 14702 38284 14742
rect 36747 14668 36763 14702
rect 37139 14668 37229 14702
rect 36475 14542 36585 14558
rect 36672 14550 36763 14584
rect 37139 14550 37155 14584
rect 36475 14346 36493 14542
rect 36569 14346 36585 14542
rect 37190 14466 37229 14668
rect 37725 14656 37810 14672
rect 38080 14668 38096 14702
rect 38472 14668 38488 14702
rect 37338 14608 37354 14642
rect 37388 14608 37404 14642
rect 37725 14596 37738 14656
rect 37793 14596 37810 14656
rect 37725 14580 37810 14596
rect 36747 14432 36763 14466
rect 37139 14432 37229 14466
rect 37440 14538 37525 14554
rect 38080 14550 38096 14584
rect 38472 14550 38488 14584
rect 37440 14478 37453 14538
rect 37508 14478 37525 14538
rect 38721 14484 38807 14500
rect 37440 14462 37525 14478
rect 38080 14432 38096 14466
rect 38472 14432 38488 14466
rect 38573 14465 38607 14481
rect 36475 14330 36585 14346
rect 36672 14314 36763 14348
rect 37139 14314 37155 14348
rect 36672 14112 36711 14314
rect 37190 14230 37229 14432
rect 38573 14415 38607 14431
rect 38721 14462 38739 14484
rect 37958 14373 37974 14407
rect 38008 14373 38024 14407
rect 38721 14404 38725 14462
rect 38721 14380 38739 14404
rect 38785 14380 38807 14484
rect 38721 14364 38807 14380
rect 38080 14314 38096 14348
rect 38472 14314 38488 14348
rect 37568 14254 37584 14288
rect 37618 14254 37634 14288
rect 36747 14196 36763 14230
rect 37139 14196 37229 14230
rect 38080 14196 38096 14230
rect 38472 14196 38488 14230
rect 36672 14078 36763 14112
rect 37139 14078 37155 14112
rect 37190 13993 37229 14196
rect 38084 14152 38284 14196
rect 38080 14118 38096 14152
rect 38272 14118 38288 14152
rect 38080 14000 38096 14034
rect 38272 14000 38288 14034
rect 34250 13977 34897 13985
rect 34250 13883 34254 13977
rect 34377 13883 34897 13977
rect 36747 13959 36763 13993
rect 37139 13959 37229 13993
rect 34250 13870 34897 13883
rect 33742 13840 33776 13856
rect 36672 13841 36763 13875
rect 37139 13841 37155 13875
rect 33549 13772 33565 13806
rect 33599 13772 33615 13806
rect 33667 13772 33683 13806
rect 33717 13772 33733 13806
rect 32020 13705 32829 13745
rect 32039 13704 32829 13705
rect 31917 13615 31984 13631
rect 31917 13581 31933 13615
rect 31967 13581 31984 13615
rect 31917 13565 31984 13581
rect 31748 13548 31782 13564
rect 31748 13498 31782 13514
rect 32094 13463 32128 13704
rect 33782 13701 33950 13719
rect 33782 13645 33798 13701
rect 33932 13645 33950 13701
rect 32564 13615 32631 13631
rect 33782 13629 33950 13645
rect 36672 13639 36711 13841
rect 37190 13757 37229 13959
rect 36747 13723 36763 13757
rect 37139 13723 37229 13757
rect 32564 13581 32581 13615
rect 32615 13581 32631 13615
rect 36672 13605 36763 13639
rect 37139 13605 37155 13639
rect 32564 13565 32631 13581
rect 32871 13547 32905 13563
rect 32183 13497 32199 13531
rect 32233 13497 32249 13531
rect 32301 13498 32317 13532
rect 32351 13498 32367 13532
rect 32871 13497 32905 13513
rect 36947 13486 36963 13520
rect 37139 13486 37232 13520
rect 31601 13447 31635 13463
rect 31601 13255 31635 13271
rect 31719 13447 31753 13463
rect 31719 13255 31753 13271
rect 32021 13447 32055 13463
rect 32094 13447 32173 13463
rect 32094 13417 32139 13447
rect 32021 13004 32056 13071
rect 32139 13055 32173 13071
rect 32257 13447 32291 13463
rect 32257 13055 32291 13071
rect 32375 13447 32409 13463
rect 32493 13447 32527 13463
rect 32899 13447 32933 13463
rect 32899 13255 32933 13271
rect 33017 13447 33051 13463
rect 33017 13255 33051 13271
rect 36876 13368 36963 13402
rect 37139 13368 37155 13402
rect 36876 13166 36913 13368
rect 37193 13284 37232 13486
rect 36947 13250 36963 13284
rect 37139 13250 37232 13284
rect 37313 13332 37347 13348
rect 37313 13282 37347 13298
rect 36876 13132 36963 13166
rect 37139 13132 37155 13166
rect 32375 13055 32409 13071
rect 32492 13004 32527 13071
rect 32021 12969 32527 13004
rect 32168 12900 32410 12912
rect 32168 12798 32215 12900
rect 32350 12798 32410 12900
rect 32168 12781 32410 12798
rect 34451 12700 37813 12787
rect 34451 12563 34580 12700
rect 37727 12665 37813 12700
rect 37727 12616 37741 12665
rect 37801 12616 37813 12665
rect 37727 12597 37813 12616
rect 32101 11319 32545 11325
rect 32101 11119 32112 11319
rect 32533 11119 32545 11319
rect 32101 11113 32545 11119
rect 32316 10834 32586 10869
rect 31962 10781 31996 10797
rect 31478 10635 31748 10670
rect 31478 10581 31512 10635
rect 31478 10389 31512 10405
rect 31596 10581 31630 10597
rect 31596 10389 31630 10405
rect 31714 10581 31748 10635
rect 31714 10389 31748 10405
rect 31832 10581 31866 10597
rect 31832 10389 31866 10405
rect 31962 10389 31996 10405
rect 32080 10781 32114 10797
rect 32080 10389 32114 10405
rect 32198 10781 32232 10797
rect 32198 10389 32232 10405
rect 32316 10781 32350 10834
rect 32316 10389 32350 10405
rect 32434 10781 32468 10797
rect 32434 10389 32468 10405
rect 32552 10781 32586 10834
rect 33560 10818 33728 10834
rect 32552 10389 32586 10405
rect 32670 10781 32704 10797
rect 33560 10748 33576 10818
rect 33712 10748 33728 10818
rect 33560 10732 33728 10748
rect 34097 10628 34367 10662
rect 32670 10389 32704 10405
rect 32799 10581 32833 10597
rect 32799 10389 32833 10405
rect 32917 10581 32951 10597
rect 32917 10389 32951 10405
rect 33035 10581 33069 10597
rect 33035 10389 33069 10405
rect 33153 10581 33187 10597
rect 33153 10389 33187 10405
rect 33271 10578 33305 10594
rect 33271 10386 33305 10402
rect 33389 10578 33423 10594
rect 33389 10386 33423 10402
rect 33507 10578 33541 10594
rect 33507 10386 33541 10402
rect 33625 10578 33659 10594
rect 33625 10386 33659 10402
rect 33743 10578 33777 10594
rect 33743 10386 33777 10402
rect 33861 10578 33895 10594
rect 33861 10386 33895 10402
rect 33979 10578 34013 10594
rect 33979 10386 34013 10402
rect 34097 10578 34131 10628
rect 34097 10386 34131 10402
rect 34215 10578 34249 10594
rect 34215 10386 34249 10402
rect 34333 10578 34367 10628
rect 34333 10386 34367 10402
rect 34022 10308 34038 10342
rect 34072 10308 34088 10342
rect 33130 10223 33164 10239
rect 33904 10191 33920 10225
rect 33954 10191 33970 10225
rect 33130 10173 33164 10189
rect 33508 10141 33542 10157
rect 31724 10104 31780 10121
rect 31724 10070 31730 10104
rect 31764 10070 31780 10104
rect 31724 10053 31780 10070
rect 31905 10088 31939 10104
rect 32023 10088 32057 10104
rect 31905 9696 31939 9712
rect 32022 9712 32023 9759
rect 32141 10088 32175 10104
rect 32057 9712 32058 9759
rect 32022 9654 32058 9712
rect 32259 10088 32293 10104
rect 32141 9696 32175 9712
rect 32257 9712 32259 9759
rect 32257 9654 32293 9712
rect 32377 10088 32411 10104
rect 32377 9696 32411 9712
rect 32495 10088 32529 10104
rect 32613 10088 32647 10104
rect 32529 9712 32531 9758
rect 32495 9654 32531 9712
rect 32775 9883 32845 9887
rect 32775 9792 32779 9883
rect 32841 9792 32845 9883
rect 32775 9787 32845 9792
rect 32613 9696 32647 9712
rect 32790 9654 32831 9787
rect 33508 9749 33542 9765
rect 33626 10141 33660 10157
rect 33626 9749 33660 9765
rect 33744 10141 33778 10157
rect 33861 10141 33895 10157
rect 33861 9949 33895 9965
rect 33979 10141 34013 10157
rect 34211 10131 34367 10137
rect 34211 10060 34226 10131
rect 34353 10060 34367 10131
rect 34211 10050 34367 10060
rect 33979 9949 34013 9965
rect 33744 9749 33778 9765
rect 33551 9681 33567 9715
rect 33601 9681 33617 9715
rect 33669 9681 33685 9715
rect 33719 9681 33735 9715
rect 32022 9614 32831 9654
rect 32041 9613 32831 9614
rect 31919 9524 31986 9540
rect 31919 9490 31935 9524
rect 31969 9490 31986 9524
rect 31919 9474 31986 9490
rect 31750 9457 31784 9473
rect 31750 9407 31784 9423
rect 32096 9372 32130 9613
rect 33784 9610 33952 9628
rect 33784 9554 33800 9610
rect 33934 9554 33952 9610
rect 32566 9524 32633 9540
rect 33784 9538 33952 9554
rect 32566 9490 32583 9524
rect 32617 9490 32633 9524
rect 32566 9474 32633 9490
rect 32873 9456 32907 9472
rect 32185 9406 32201 9440
rect 32235 9406 32251 9440
rect 32303 9407 32319 9441
rect 32353 9407 32369 9441
rect 32873 9406 32907 9422
rect 31603 9356 31637 9372
rect 31603 9164 31637 9180
rect 31721 9356 31755 9372
rect 31721 9164 31755 9180
rect 32023 9356 32057 9372
rect 32096 9356 32175 9372
rect 32096 9326 32141 9356
rect 32023 8913 32058 8980
rect 32141 8964 32175 8980
rect 32259 9356 32293 9372
rect 32259 8964 32293 8980
rect 32377 9356 32411 9372
rect 32495 9356 32529 9372
rect 32901 9356 32935 9372
rect 32901 9164 32935 9180
rect 33019 9356 33053 9372
rect 33019 9164 33053 9180
rect 32377 8964 32411 8980
rect 32494 8913 32529 8980
rect 32023 8878 32529 8913
rect 32170 8809 32412 8821
rect 32170 8707 32217 8809
rect 32352 8707 32412 8809
rect 32170 8690 32412 8707
rect 16405 8336 31324 8337
rect 13940 8335 31324 8336
rect 9185 8226 31324 8335
rect 9185 8224 19612 8226
rect 28663 8225 31324 8226
rect 9185 8223 16189 8224
rect 3140 8081 31165 8083
rect 34274 8081 34367 10050
rect 3140 7954 34367 8081
rect 14531 7952 34367 7954
rect 32101 7824 32545 7830
rect 4425 7692 4648 7767
rect 4425 7543 4501 7692
rect 4568 7691 4648 7692
rect 4425 7542 4504 7543
rect 4571 7542 4648 7691
rect 4425 7436 4648 7542
rect 6907 7747 7130 7821
rect 6907 7598 6981 7747
rect 7048 7745 7130 7747
rect 6907 7596 6986 7598
rect 7053 7596 7130 7745
rect 6240 7525 6274 7541
rect 6240 7475 6274 7491
rect 6907 7490 7130 7596
rect 8054 7745 8277 7821
rect 8054 7596 8133 7745
rect 8200 7744 8277 7745
rect 8054 7595 8137 7596
rect 8204 7595 8277 7744
rect 7370 7531 7404 7547
rect 7370 7481 7404 7497
rect 8054 7490 8277 7595
rect 10976 7690 11199 7765
rect 10976 7689 11056 7690
rect 10976 7540 11055 7689
rect 11123 7541 11199 7690
rect 11122 7540 11199 7541
rect 10976 7434 11199 7540
rect 13458 7743 13681 7819
rect 13458 7594 13537 7743
rect 13604 7594 13681 7743
rect 12791 7523 12825 7539
rect 12791 7473 12825 7489
rect 13458 7488 13681 7594
rect 14605 7743 14828 7819
rect 14605 7594 14684 7743
rect 14752 7594 14828 7743
rect 13921 7529 13955 7545
rect 13921 7479 13955 7495
rect 14605 7488 14828 7594
rect 16387 7748 16549 7764
rect 16387 7680 16430 7748
rect 16500 7680 16549 7748
rect 6240 7407 6274 7423
rect 4856 7327 5126 7361
rect 6240 7357 6274 7373
rect 7370 7411 7404 7427
rect 4030 7277 4064 7293
rect 4030 7085 4064 7101
rect 4148 7277 4182 7293
rect 4148 7085 4182 7101
rect 4266 7277 4300 7293
rect 4266 7085 4300 7101
rect 4384 7277 4418 7293
rect 4384 7085 4418 7101
rect 4502 7277 4536 7293
rect 4502 7085 4536 7101
rect 4620 7277 4654 7293
rect 4620 7085 4654 7101
rect 4738 7277 4772 7293
rect 4738 7085 4772 7101
rect 4856 7277 4890 7327
rect 4856 7085 4890 7101
rect 4974 7277 5008 7293
rect 4974 7085 5008 7101
rect 5092 7277 5126 7327
rect 5092 7085 5126 7101
rect 6355 7349 6389 7365
rect 4781 7007 4797 7041
rect 4831 7007 4847 7041
rect 6355 6957 6389 6973
rect 6473 7349 6507 7365
rect 6473 6957 6507 6973
rect 6591 7349 6625 7365
rect 6591 6957 6625 6973
rect 6709 7349 6743 7365
rect 6709 6957 6743 6973
rect 6827 7349 6861 7365
rect 6827 6957 6861 6973
rect 6945 7349 6979 7365
rect 6945 6957 6979 6973
rect 7063 7349 7097 7365
rect 7370 7361 7404 7377
rect 12791 7405 12825 7421
rect 7063 6957 7097 6973
rect 7497 7353 7531 7369
rect 7497 6961 7531 6977
rect 7615 7353 7649 7369
rect 7615 6961 7649 6977
rect 7733 7353 7767 7369
rect 7733 6961 7767 6977
rect 7851 7353 7885 7369
rect 7851 6961 7885 6977
rect 7969 7353 8003 7369
rect 7969 6961 8003 6977
rect 8087 7353 8121 7369
rect 8087 6961 8121 6977
rect 8205 7353 8239 7369
rect 11407 7325 11677 7359
rect 12791 7355 12825 7371
rect 13921 7409 13955 7425
rect 10581 7275 10615 7291
rect 10581 7083 10615 7099
rect 10699 7275 10733 7291
rect 10699 7083 10733 7099
rect 10817 7275 10851 7291
rect 10817 7083 10851 7099
rect 10935 7275 10969 7291
rect 10935 7083 10969 7099
rect 11053 7275 11087 7291
rect 11053 7083 11087 7099
rect 11171 7275 11205 7291
rect 11171 7083 11205 7099
rect 11289 7275 11323 7291
rect 11289 7083 11323 7099
rect 11407 7275 11441 7325
rect 11407 7083 11441 7099
rect 11525 7275 11559 7291
rect 11525 7083 11559 7099
rect 11643 7275 11677 7325
rect 11643 7083 11677 7099
rect 12906 7347 12940 7363
rect 11332 7005 11348 7039
rect 11382 7005 11398 7039
rect 8205 6961 8239 6977
rect 12906 6955 12940 6971
rect 13024 7347 13058 7363
rect 13024 6955 13058 6971
rect 13142 7347 13176 7363
rect 13142 6955 13176 6971
rect 13260 7347 13294 7363
rect 13260 6955 13294 6971
rect 13378 7347 13412 7363
rect 13378 6955 13412 6971
rect 13496 7347 13530 7363
rect 13496 6955 13530 6971
rect 13614 7347 13648 7363
rect 13921 7359 13955 7375
rect 13614 6955 13648 6971
rect 14048 7351 14082 7367
rect 14048 6959 14082 6975
rect 14166 7351 14200 7367
rect 14166 6959 14200 6975
rect 14284 7351 14318 7367
rect 14284 6959 14318 6975
rect 14402 7351 14436 7367
rect 14402 6959 14436 6975
rect 14520 7351 14554 7367
rect 14520 6959 14554 6975
rect 14638 7351 14672 7367
rect 14638 6959 14672 6975
rect 14756 7351 14790 7367
rect 16387 7162 16549 7680
rect 17631 7690 17854 7766
rect 17631 7687 17710 7690
rect 17631 7538 17707 7687
rect 17777 7541 17854 7690
rect 17774 7538 17854 7541
rect 20113 7747 20336 7820
rect 20113 7595 20192 7747
rect 20259 7595 20336 7747
rect 17631 7435 17854 7538
rect 19446 7524 19480 7540
rect 19446 7474 19480 7490
rect 20113 7489 20336 7595
rect 21260 7744 21483 7820
rect 21260 7595 21339 7744
rect 21408 7595 21483 7744
rect 20576 7530 20610 7546
rect 20576 7480 20610 7496
rect 21260 7489 21483 7595
rect 24253 7692 24476 7767
rect 24253 7543 24331 7692
rect 24398 7691 24476 7692
rect 24253 7542 24332 7543
rect 24399 7542 24476 7691
rect 24253 7436 24476 7542
rect 26735 7745 26958 7821
rect 26735 7740 26814 7745
rect 26735 7591 26810 7740
rect 26881 7596 26958 7745
rect 26877 7591 26958 7596
rect 26068 7525 26102 7541
rect 26068 7475 26102 7491
rect 26735 7490 26958 7591
rect 27882 7746 28105 7821
rect 27882 7597 27958 7746
rect 28025 7745 28105 7746
rect 27882 7596 27961 7597
rect 28028 7596 28105 7745
rect 30023 7793 30191 7809
rect 30023 7723 30039 7793
rect 30175 7723 30191 7793
rect 30023 7707 30191 7723
rect 27198 7531 27232 7547
rect 27198 7481 27232 7497
rect 27882 7490 28105 7596
rect 30560 7603 30830 7637
rect 32101 7624 32112 7824
rect 32533 7624 32545 7824
rect 32101 7618 32545 7624
rect 29734 7553 29768 7569
rect 19446 7406 19480 7422
rect 18062 7326 18332 7360
rect 19446 7356 19480 7372
rect 20576 7410 20610 7426
rect 17236 7276 17270 7292
rect 14756 6959 14790 6975
rect 4663 6890 4679 6924
rect 4713 6890 4729 6924
rect 11214 6888 11230 6922
rect 11264 6888 11280 6922
rect 4267 6840 4301 6856
rect 4267 6448 4301 6464
rect 4385 6840 4419 6856
rect 4385 6448 4419 6464
rect 4503 6840 4537 6856
rect 4620 6840 4654 6856
rect 4620 6648 4654 6664
rect 4738 6840 4772 6856
rect 4738 6648 4772 6664
rect 10818 6838 10852 6854
rect 6544 6617 6560 6651
rect 6594 6617 6610 6651
rect 7686 6621 7702 6655
rect 7736 6621 7752 6655
rect 6265 6566 6299 6582
rect 4503 6448 4537 6464
rect 4790 6514 5039 6557
rect 4790 6424 4837 6514
rect 5000 6424 5039 6514
rect 4310 6380 4326 6414
rect 4360 6380 4376 6414
rect 4428 6380 4444 6414
rect 4478 6380 4494 6414
rect 4790 6385 5039 6424
rect 6265 6374 6299 6390
rect 6383 6566 6417 6582
rect 6383 6374 6417 6390
rect 6501 6566 6535 6582
rect 6501 6374 6535 6390
rect 6619 6566 6653 6582
rect 6619 6374 6653 6390
rect 6784 6566 6818 6582
rect 6784 6374 6818 6390
rect 6902 6566 6936 6582
rect 6902 6374 6936 6390
rect 7020 6566 7054 6582
rect 7020 6374 7054 6390
rect 7138 6566 7172 6582
rect 7138 6374 7172 6390
rect 7407 6570 7441 6586
rect 7407 6378 7441 6394
rect 7525 6570 7559 6586
rect 7525 6378 7559 6394
rect 7643 6570 7677 6586
rect 7643 6378 7677 6394
rect 7761 6570 7795 6586
rect 7761 6378 7795 6394
rect 7926 6570 7960 6586
rect 7926 6378 7960 6394
rect 8044 6570 8078 6586
rect 8044 6378 8078 6394
rect 8162 6570 8196 6586
rect 8162 6378 8196 6394
rect 8280 6570 8314 6586
rect 10818 6446 10852 6462
rect 10936 6838 10970 6854
rect 10936 6446 10970 6462
rect 11054 6838 11088 6854
rect 11171 6838 11205 6854
rect 11171 6646 11205 6662
rect 11289 6838 11323 6854
rect 11289 6646 11323 6662
rect 13095 6615 13111 6649
rect 13145 6615 13161 6649
rect 14237 6619 14253 6653
rect 14287 6619 14303 6653
rect 12816 6564 12850 6580
rect 11054 6446 11088 6462
rect 11341 6512 11590 6555
rect 11341 6422 11388 6512
rect 11551 6422 11590 6512
rect 8280 6378 8314 6394
rect 10861 6378 10877 6412
rect 10911 6378 10927 6412
rect 10979 6378 10995 6412
rect 11029 6378 11045 6412
rect 11341 6383 11590 6422
rect 12816 6372 12850 6388
rect 12934 6564 12968 6580
rect 12934 6372 12968 6388
rect 13052 6564 13086 6580
rect 13052 6372 13086 6388
rect 13170 6564 13204 6580
rect 13170 6372 13204 6388
rect 13335 6564 13369 6580
rect 13335 6372 13369 6388
rect 13453 6564 13487 6580
rect 13453 6372 13487 6388
rect 13571 6564 13605 6580
rect 13571 6372 13605 6388
rect 13689 6564 13723 6580
rect 13689 6372 13723 6388
rect 13958 6568 13992 6584
rect 13958 6376 13992 6392
rect 14076 6568 14110 6584
rect 14076 6376 14110 6392
rect 14194 6568 14228 6584
rect 14194 6376 14228 6392
rect 14312 6568 14346 6584
rect 14312 6376 14346 6392
rect 14477 6568 14511 6584
rect 14477 6376 14511 6392
rect 14595 6568 14629 6584
rect 14595 6376 14629 6392
rect 14713 6568 14747 6584
rect 14713 6376 14747 6392
rect 14831 6568 14865 6584
rect 14831 6376 14865 6392
rect 6280 6143 6452 6190
rect 4439 6041 4662 6117
rect 4439 5892 4518 6041
rect 4585 6039 4662 6041
rect 4439 5890 4522 5892
rect 4589 5890 4662 6039
rect 6280 5980 6319 6143
rect 6409 5980 6452 6143
rect 6280 5941 6452 5980
rect 7422 6141 7594 6188
rect 7422 5978 7461 6141
rect 7551 5978 7594 6141
rect 12831 6141 13003 6188
rect 7422 5939 7594 5978
rect 10990 6046 11213 6115
rect 4439 5786 4662 5890
rect 10990 5897 11067 6046
rect 11134 6039 11213 6046
rect 10990 5890 11069 5897
rect 11136 5890 11213 6039
rect 12831 5978 12870 6141
rect 12960 5978 13003 6141
rect 12831 5939 13003 5978
rect 13973 6139 14145 6186
rect 13973 5976 14012 6139
rect 14102 5976 14145 6139
rect 13973 5972 14020 5976
rect 14087 5972 14145 5976
rect 13973 5937 14145 5972
rect 10990 5784 11213 5890
rect 4870 5677 5140 5711
rect 4044 5627 4078 5643
rect 4044 5435 4078 5451
rect 4162 5627 4196 5643
rect 4162 5435 4196 5451
rect 4280 5627 4314 5643
rect 4280 5435 4314 5451
rect 4398 5627 4432 5643
rect 4398 5435 4432 5451
rect 4516 5627 4550 5643
rect 4516 5435 4550 5451
rect 4634 5627 4668 5643
rect 4634 5435 4668 5451
rect 4752 5627 4786 5643
rect 4752 5435 4786 5451
rect 4870 5627 4904 5677
rect 4870 5435 4904 5451
rect 4988 5627 5022 5643
rect 4988 5435 5022 5451
rect 5106 5627 5140 5677
rect 5106 5435 5140 5451
rect 8150 5698 8375 5774
rect 8150 5549 8228 5698
rect 8296 5549 8375 5698
rect 11421 5675 11691 5709
rect 8150 5443 8375 5549
rect 10595 5625 10629 5641
rect 10595 5433 10629 5449
rect 10713 5625 10747 5641
rect 10713 5433 10747 5449
rect 10831 5625 10865 5641
rect 10831 5433 10865 5449
rect 10949 5625 10983 5641
rect 10949 5433 10983 5449
rect 11067 5625 11101 5641
rect 11067 5433 11101 5449
rect 11185 5625 11219 5641
rect 11185 5433 11219 5449
rect 11303 5625 11337 5641
rect 11303 5433 11337 5449
rect 11421 5625 11455 5675
rect 11421 5433 11455 5449
rect 11539 5625 11573 5641
rect 11539 5433 11573 5449
rect 11657 5625 11691 5675
rect 11657 5433 11691 5449
rect 14701 5697 14926 5772
rect 14701 5696 14784 5697
rect 14701 5547 14780 5696
rect 14851 5548 14926 5697
rect 14847 5547 14926 5548
rect 14701 5441 14926 5547
rect 4795 5357 4811 5391
rect 4845 5357 4861 5391
rect 11346 5355 11362 5389
rect 11396 5355 11412 5389
rect 4677 5240 4693 5274
rect 4727 5240 4743 5274
rect 6346 5263 6616 5298
rect 5992 5210 6026 5226
rect 4281 5190 4315 5206
rect 4281 4798 4315 4814
rect 4399 5190 4433 5206
rect 4399 4798 4433 4814
rect 4517 5190 4551 5206
rect 4634 5190 4668 5206
rect 4634 4998 4668 5014
rect 4752 5190 4786 5206
rect 4752 4998 4786 5014
rect 5508 5064 5778 5099
rect 5508 5010 5542 5064
rect 4517 4798 4551 4814
rect 4804 4864 5053 4907
rect 4804 4774 4851 4864
rect 5014 4774 5053 4864
rect 5508 4818 5542 4834
rect 5626 5010 5660 5026
rect 5626 4818 5660 4834
rect 5744 5010 5778 5064
rect 5744 4818 5778 4834
rect 5862 5010 5896 5026
rect 5862 4818 5896 4834
rect 5992 4818 6026 4834
rect 6110 5210 6144 5226
rect 6110 4818 6144 4834
rect 6228 5210 6262 5226
rect 6228 4818 6262 4834
rect 6346 5210 6380 5263
rect 6346 4818 6380 4834
rect 6464 5210 6498 5226
rect 6464 4818 6498 4834
rect 6582 5210 6616 5263
rect 8244 5263 8514 5298
rect 6582 4818 6616 4834
rect 6700 5210 6734 5226
rect 7890 5210 7924 5226
rect 7406 5064 7676 5099
rect 6700 4818 6734 4834
rect 6829 5010 6863 5026
rect 6829 4818 6863 4834
rect 6947 5010 6981 5026
rect 6947 4818 6981 4834
rect 7065 5010 7099 5026
rect 7065 4818 7099 4834
rect 7183 5010 7217 5026
rect 7183 4818 7217 4834
rect 7406 5010 7440 5064
rect 7406 4818 7440 4834
rect 7524 5010 7558 5026
rect 7524 4818 7558 4834
rect 7642 5010 7676 5064
rect 7642 4818 7676 4834
rect 7760 5010 7794 5026
rect 7760 4818 7794 4834
rect 7890 4818 7924 4834
rect 8008 5210 8042 5226
rect 8008 4818 8042 4834
rect 8126 5210 8160 5226
rect 8126 4818 8160 4834
rect 8244 5210 8278 5263
rect 8244 4818 8278 4834
rect 8362 5210 8396 5226
rect 8362 4818 8396 4834
rect 8480 5210 8514 5263
rect 11228 5238 11244 5272
rect 11278 5238 11294 5272
rect 12897 5261 13167 5296
rect 8480 4818 8514 4834
rect 8598 5210 8632 5226
rect 12543 5208 12577 5224
rect 10832 5188 10866 5204
rect 8598 4818 8632 4834
rect 8727 5010 8761 5026
rect 8727 4818 8761 4834
rect 8845 5010 8879 5026
rect 8845 4818 8879 4834
rect 8963 5010 8997 5026
rect 8963 4818 8997 4834
rect 9081 5010 9115 5026
rect 9081 4818 9115 4834
rect 10832 4796 10866 4812
rect 10950 5188 10984 5204
rect 10950 4796 10984 4812
rect 11068 5188 11102 5204
rect 11185 5188 11219 5204
rect 11185 4996 11219 5012
rect 11303 5188 11337 5204
rect 11303 4996 11337 5012
rect 12059 5062 12329 5097
rect 12059 5008 12093 5062
rect 11068 4796 11102 4812
rect 11355 4862 11604 4905
rect 4324 4730 4340 4764
rect 4374 4730 4390 4764
rect 4442 4730 4458 4764
rect 4492 4730 4508 4764
rect 4804 4735 5053 4774
rect 11355 4772 11402 4862
rect 11565 4772 11604 4862
rect 12059 4816 12093 4832
rect 12177 5008 12211 5024
rect 12177 4816 12211 4832
rect 12295 5008 12329 5062
rect 12295 4816 12329 4832
rect 12413 5008 12447 5024
rect 12413 4816 12447 4832
rect 12543 4816 12577 4832
rect 12661 5208 12695 5224
rect 12661 4816 12695 4832
rect 12779 5208 12813 5224
rect 12779 4816 12813 4832
rect 12897 5208 12931 5261
rect 12897 4816 12931 4832
rect 13015 5208 13049 5224
rect 13015 4816 13049 4832
rect 13133 5208 13167 5261
rect 14795 5261 15065 5296
rect 13133 4816 13167 4832
rect 13251 5208 13285 5224
rect 14441 5208 14475 5224
rect 13957 5062 14227 5097
rect 13251 4816 13285 4832
rect 13380 5008 13414 5024
rect 13380 4816 13414 4832
rect 13498 5008 13532 5024
rect 13498 4816 13532 4832
rect 13616 5008 13650 5024
rect 13616 4816 13650 4832
rect 13734 5008 13768 5024
rect 13734 4816 13768 4832
rect 13957 5008 13991 5062
rect 13957 4816 13991 4832
rect 14075 5008 14109 5024
rect 14075 4816 14109 4832
rect 14193 5008 14227 5062
rect 14193 4816 14227 4832
rect 14311 5008 14345 5024
rect 14311 4816 14345 4832
rect 14441 4816 14475 4832
rect 14559 5208 14593 5224
rect 14559 4816 14593 4832
rect 14677 5208 14711 5224
rect 14677 4816 14711 4832
rect 14795 5208 14829 5261
rect 14795 4816 14829 4832
rect 14913 5208 14947 5224
rect 14913 4816 14947 4832
rect 15031 5208 15065 5261
rect 15031 4816 15065 4832
rect 15149 5208 15183 5224
rect 15149 4816 15183 4832
rect 15278 5008 15312 5024
rect 15278 4816 15312 4832
rect 15396 5008 15430 5024
rect 15396 4816 15430 4832
rect 15514 5008 15548 5024
rect 15514 4816 15548 4832
rect 15632 5008 15666 5024
rect 15632 4816 15666 4832
rect 10875 4728 10891 4762
rect 10925 4728 10941 4762
rect 10993 4728 11009 4762
rect 11043 4728 11059 4762
rect 11355 4733 11604 4772
rect 6972 4596 7006 4612
rect 13523 4594 13557 4610
rect 6972 4546 7006 4562
rect 9062 4575 9129 4591
rect 9062 4541 9079 4575
rect 9113 4541 9129 4575
rect 13523 4544 13557 4560
rect 15613 4573 15680 4589
rect 5935 4517 5969 4533
rect 4434 4440 4657 4513
rect 4434 4291 4511 4440
rect 4578 4437 4657 4440
rect 4434 4288 4513 4291
rect 4580 4288 4657 4437
rect 4434 4182 4657 4288
rect 6053 4517 6087 4533
rect 5935 4125 5969 4141
rect 6052 4141 6053 4188
rect 6171 4517 6205 4533
rect 6087 4141 6088 4188
rect 4865 4073 5135 4107
rect 4039 4023 4073 4039
rect 4039 3831 4073 3847
rect 4157 4023 4191 4039
rect 4157 3831 4191 3847
rect 4275 4023 4309 4039
rect 4275 3831 4309 3847
rect 4393 4023 4427 4039
rect 4393 3831 4427 3847
rect 4511 4023 4545 4039
rect 4511 3831 4545 3847
rect 4629 4023 4663 4039
rect 4629 3831 4663 3847
rect 4747 4023 4781 4039
rect 4747 3831 4781 3847
rect 4865 4023 4899 4073
rect 4865 3831 4899 3847
rect 4983 4023 5017 4039
rect 4983 3831 5017 3847
rect 5101 4023 5135 4073
rect 6052 4083 6088 4141
rect 6289 4517 6323 4533
rect 6171 4125 6205 4141
rect 6287 4141 6289 4188
rect 6287 4083 6323 4141
rect 6407 4517 6441 4533
rect 6407 4125 6441 4141
rect 6525 4517 6559 4533
rect 6643 4517 6677 4533
rect 6559 4141 6561 4187
rect 6525 4083 6561 4141
rect 6643 4125 6677 4141
rect 7833 4517 7867 4533
rect 7951 4517 7985 4533
rect 7833 4125 7867 4141
rect 7950 4141 7951 4188
rect 8069 4517 8103 4533
rect 7985 4141 7986 4188
rect 7148 4083 7645 4101
rect 6052 4080 7645 4083
rect 6052 4046 7593 4080
rect 7627 4046 7645 4080
rect 6052 4043 7645 4046
rect 7950 4083 7986 4141
rect 8187 4517 8221 4533
rect 8069 4125 8103 4141
rect 8185 4141 8187 4188
rect 8185 4083 8221 4141
rect 8305 4517 8339 4533
rect 8305 4125 8339 4141
rect 8423 4517 8457 4533
rect 8541 4517 8575 4533
rect 9062 4525 9129 4541
rect 15613 4539 15630 4573
rect 15664 4539 15680 4573
rect 8457 4141 8459 4187
rect 8423 4083 8459 4141
rect 12486 4515 12520 4531
rect 10985 4435 11208 4511
rect 10985 4286 11064 4435
rect 11134 4286 11208 4435
rect 10985 4180 11208 4286
rect 8541 4125 8575 4141
rect 12604 4515 12638 4531
rect 12486 4123 12520 4139
rect 12603 4139 12604 4186
rect 12722 4515 12756 4531
rect 12638 4139 12639 4186
rect 9046 4112 9146 4113
rect 9046 4083 9202 4112
rect 7950 4043 9202 4083
rect 6071 4042 7645 4043
rect 7969 4042 9202 4043
rect 5949 3953 6016 3969
rect 5949 3919 5965 3953
rect 5999 3919 6016 3953
rect 5949 3903 6016 3919
rect 5101 3831 5135 3847
rect 5780 3886 5814 3902
rect 5780 3836 5814 3852
rect 6126 3801 6160 4042
rect 7148 4025 7645 4042
rect 6596 3953 6663 3969
rect 6596 3919 6613 3953
rect 6647 3919 6663 3953
rect 6596 3903 6663 3919
rect 7847 3953 7914 3969
rect 7847 3919 7863 3953
rect 7897 3919 7914 3953
rect 7847 3903 7914 3919
rect 6903 3885 6937 3901
rect 6215 3835 6231 3869
rect 6265 3835 6281 3869
rect 6333 3836 6349 3870
rect 6383 3836 6399 3870
rect 6903 3835 6937 3851
rect 7678 3886 7712 3902
rect 7678 3836 7712 3852
rect 8024 3801 8058 4042
rect 9046 4014 9202 4042
rect 11416 4071 11686 4105
rect 10590 4021 10624 4037
rect 9046 4013 9146 4014
rect 8492 3954 8559 3970
rect 8492 3920 8509 3954
rect 8543 3920 8559 3954
rect 8492 3904 8559 3920
rect 8801 3885 8835 3901
rect 8113 3835 8129 3869
rect 8163 3835 8179 3869
rect 8231 3836 8247 3870
rect 8281 3836 8297 3870
rect 8801 3835 8835 3851
rect 10590 3829 10624 3845
rect 10708 4021 10742 4037
rect 10708 3829 10742 3845
rect 10826 4021 10860 4037
rect 10826 3829 10860 3845
rect 10944 4021 10978 4037
rect 10944 3829 10978 3845
rect 11062 4021 11096 4037
rect 11062 3829 11096 3845
rect 11180 4021 11214 4037
rect 11180 3829 11214 3845
rect 11298 4021 11332 4037
rect 11298 3829 11332 3845
rect 11416 4021 11450 4071
rect 11416 3829 11450 3845
rect 11534 4021 11568 4037
rect 11534 3829 11568 3845
rect 11652 4021 11686 4071
rect 12603 4081 12639 4139
rect 12840 4515 12874 4531
rect 12722 4123 12756 4139
rect 12838 4139 12840 4186
rect 12838 4081 12874 4139
rect 12958 4515 12992 4531
rect 12958 4123 12992 4139
rect 13076 4515 13110 4531
rect 13194 4515 13228 4531
rect 13110 4139 13112 4185
rect 13076 4081 13112 4139
rect 13194 4123 13228 4139
rect 14384 4515 14418 4531
rect 14502 4515 14536 4531
rect 14384 4123 14418 4139
rect 14501 4139 14502 4186
rect 14620 4515 14654 4531
rect 14536 4139 14537 4186
rect 13699 4081 14196 4099
rect 12603 4078 14196 4081
rect 12603 4044 14144 4078
rect 14178 4044 14196 4078
rect 12603 4041 14196 4044
rect 14501 4081 14537 4139
rect 14738 4515 14772 4531
rect 14620 4123 14654 4139
rect 14736 4139 14738 4186
rect 14736 4081 14772 4139
rect 14856 4515 14890 4531
rect 14856 4123 14890 4139
rect 14974 4515 15008 4531
rect 15092 4515 15126 4531
rect 15613 4523 15680 4539
rect 15008 4139 15010 4185
rect 14974 4081 15010 4139
rect 15092 4123 15126 4139
rect 15597 4081 15904 4111
rect 14501 4041 15904 4081
rect 12622 4040 14196 4041
rect 14520 4040 15904 4041
rect 12500 3951 12567 3967
rect 12500 3917 12516 3951
rect 12550 3917 12567 3951
rect 12500 3901 12567 3917
rect 11652 3829 11686 3845
rect 12331 3884 12365 3900
rect 12331 3834 12365 3850
rect 4790 3753 4806 3787
rect 4840 3753 4856 3787
rect 5633 3785 5667 3801
rect 4672 3636 4688 3670
rect 4722 3636 4738 3670
rect 4276 3586 4310 3602
rect 4276 3194 4310 3210
rect 4394 3586 4428 3602
rect 4394 3194 4428 3210
rect 4512 3586 4546 3602
rect 4629 3586 4663 3602
rect 4629 3394 4663 3410
rect 4747 3586 4781 3602
rect 5633 3593 5667 3609
rect 5751 3785 5785 3801
rect 5751 3593 5785 3609
rect 6053 3785 6087 3801
rect 4747 3394 4781 3410
rect 6126 3785 6205 3801
rect 6126 3755 6171 3785
rect 6053 3342 6088 3409
rect 6171 3393 6205 3409
rect 6289 3785 6323 3801
rect 6289 3393 6323 3409
rect 6407 3785 6441 3801
rect 6525 3785 6559 3801
rect 6931 3785 6965 3801
rect 6931 3593 6965 3609
rect 7049 3785 7083 3801
rect 7049 3593 7083 3609
rect 7531 3785 7565 3801
rect 7531 3593 7565 3609
rect 7649 3785 7683 3801
rect 7649 3593 7683 3609
rect 7951 3785 7985 3801
rect 6407 3393 6441 3409
rect 6524 3342 6559 3409
rect 6053 3307 6559 3342
rect 8024 3785 8103 3801
rect 8024 3755 8069 3785
rect 7951 3342 7986 3409
rect 8069 3393 8103 3409
rect 8187 3785 8221 3801
rect 8187 3393 8221 3409
rect 8305 3785 8339 3801
rect 8423 3785 8457 3801
rect 8829 3785 8863 3801
rect 8829 3593 8863 3609
rect 8947 3785 8981 3801
rect 12677 3799 12711 4040
rect 13699 4023 14196 4040
rect 13147 3951 13214 3967
rect 13147 3917 13164 3951
rect 13198 3917 13214 3951
rect 13147 3901 13214 3917
rect 14398 3951 14465 3967
rect 14398 3917 14414 3951
rect 14448 3917 14465 3951
rect 14398 3901 14465 3917
rect 13454 3883 13488 3899
rect 12766 3833 12782 3867
rect 12816 3833 12832 3867
rect 12884 3834 12900 3868
rect 12934 3834 12950 3868
rect 13454 3833 13488 3849
rect 14229 3884 14263 3900
rect 14229 3834 14263 3850
rect 14575 3799 14609 4040
rect 15597 4011 15904 4040
rect 15669 4010 15904 4011
rect 15043 3952 15110 3968
rect 15043 3918 15060 3952
rect 15094 3918 15110 3952
rect 15043 3902 15110 3918
rect 15352 3883 15386 3899
rect 14664 3833 14680 3867
rect 14714 3833 14730 3867
rect 14782 3834 14798 3868
rect 14832 3834 14848 3868
rect 15352 3833 15386 3849
rect 11341 3751 11357 3785
rect 11391 3751 11407 3785
rect 12184 3783 12218 3799
rect 11223 3634 11239 3668
rect 11273 3634 11289 3668
rect 8947 3593 8981 3609
rect 8305 3393 8339 3409
rect 8422 3342 8457 3409
rect 7951 3307 8457 3342
rect 10827 3584 10861 3600
rect 4512 3194 4546 3210
rect 4799 3260 5048 3303
rect 4799 3170 4846 3260
rect 5009 3170 5048 3260
rect 10827 3192 10861 3208
rect 10945 3584 10979 3600
rect 10945 3192 10979 3208
rect 11063 3584 11097 3600
rect 11180 3584 11214 3600
rect 11180 3392 11214 3408
rect 11298 3584 11332 3600
rect 12184 3591 12218 3607
rect 12302 3783 12336 3799
rect 12302 3591 12336 3607
rect 12604 3783 12638 3799
rect 11298 3392 11332 3408
rect 12677 3783 12756 3799
rect 12677 3753 12722 3783
rect 12604 3340 12639 3407
rect 12722 3391 12756 3407
rect 12840 3783 12874 3799
rect 12840 3391 12874 3407
rect 12958 3783 12992 3799
rect 13076 3783 13110 3799
rect 13482 3783 13516 3799
rect 13482 3591 13516 3607
rect 13600 3783 13634 3799
rect 13600 3591 13634 3607
rect 14082 3783 14116 3799
rect 14082 3591 14116 3607
rect 14200 3783 14234 3799
rect 14200 3591 14234 3607
rect 14502 3783 14536 3799
rect 12958 3391 12992 3407
rect 13075 3340 13110 3407
rect 12604 3305 13110 3340
rect 14575 3783 14654 3799
rect 14575 3753 14620 3783
rect 14502 3340 14537 3407
rect 14620 3391 14654 3407
rect 14738 3783 14772 3799
rect 14738 3391 14772 3407
rect 14856 3783 14890 3799
rect 14974 3783 15008 3799
rect 15380 3783 15414 3799
rect 15380 3591 15414 3607
rect 15498 3783 15532 3799
rect 15498 3591 15532 3607
rect 14856 3391 14890 3407
rect 14973 3340 15008 3407
rect 14502 3305 15008 3340
rect 11063 3192 11097 3208
rect 11350 3258 11599 3301
rect 4319 3126 4335 3160
rect 4369 3126 4385 3160
rect 4437 3126 4453 3160
rect 4487 3126 4503 3160
rect 4799 3131 5048 3170
rect 11350 3168 11397 3258
rect 11560 3168 11599 3258
rect 6224 3100 6396 3147
rect 10870 3124 10886 3158
rect 10920 3124 10936 3158
rect 10988 3124 11004 3158
rect 11038 3124 11054 3158
rect 11350 3129 11599 3168
rect 6224 2937 6263 3100
rect 6353 2937 6396 3100
rect 6224 2897 6396 2937
rect 12775 3098 12947 3145
rect 12775 2935 12814 3098
rect 12904 2935 12947 3098
rect 12775 2895 12947 2935
rect 15770 2655 15904 4010
rect 16384 2990 16552 7162
rect 17236 7084 17270 7100
rect 17354 7276 17388 7292
rect 17354 7084 17388 7100
rect 17472 7276 17506 7292
rect 17472 7084 17506 7100
rect 17590 7276 17624 7292
rect 17590 7084 17624 7100
rect 17708 7276 17742 7292
rect 17708 7084 17742 7100
rect 17826 7276 17860 7292
rect 17826 7084 17860 7100
rect 17944 7276 17978 7292
rect 17944 7084 17978 7100
rect 18062 7276 18096 7326
rect 18062 7084 18096 7100
rect 18180 7276 18214 7292
rect 18180 7084 18214 7100
rect 18298 7276 18332 7326
rect 18298 7084 18332 7100
rect 19561 7348 19595 7364
rect 17987 7006 18003 7040
rect 18037 7006 18053 7040
rect 19561 6956 19595 6972
rect 19679 7348 19713 7364
rect 19679 6956 19713 6972
rect 19797 7348 19831 7364
rect 19797 6956 19831 6972
rect 19915 7348 19949 7364
rect 19915 6956 19949 6972
rect 20033 7348 20067 7364
rect 20033 6956 20067 6972
rect 20151 7348 20185 7364
rect 20151 6956 20185 6972
rect 20269 7348 20303 7364
rect 20576 7360 20610 7376
rect 26068 7407 26102 7423
rect 20269 6956 20303 6972
rect 20703 7352 20737 7368
rect 20703 6960 20737 6976
rect 20821 7352 20855 7368
rect 20821 6960 20855 6976
rect 20939 7352 20973 7368
rect 20939 6960 20973 6976
rect 21057 7352 21091 7368
rect 21057 6960 21091 6976
rect 21175 7352 21209 7368
rect 21175 6960 21209 6976
rect 21293 7352 21327 7368
rect 21293 6960 21327 6976
rect 21411 7352 21445 7368
rect 24684 7327 24954 7361
rect 26068 7357 26102 7373
rect 27198 7411 27232 7427
rect 23858 7277 23892 7293
rect 23858 7085 23892 7101
rect 23976 7277 24010 7293
rect 23976 7085 24010 7101
rect 24094 7277 24128 7293
rect 24094 7085 24128 7101
rect 24212 7277 24246 7293
rect 24212 7085 24246 7101
rect 24330 7277 24364 7293
rect 24330 7085 24364 7101
rect 24448 7277 24482 7293
rect 24448 7085 24482 7101
rect 24566 7277 24600 7293
rect 24566 7085 24600 7101
rect 24684 7277 24718 7327
rect 24684 7085 24718 7101
rect 24802 7277 24836 7293
rect 24802 7085 24836 7101
rect 24920 7277 24954 7327
rect 24920 7085 24954 7101
rect 26183 7349 26217 7365
rect 24609 7007 24625 7041
rect 24659 7007 24675 7041
rect 21411 6960 21445 6976
rect 26183 6957 26217 6973
rect 26301 7349 26335 7365
rect 26301 6957 26335 6973
rect 26419 7349 26453 7365
rect 26419 6957 26453 6973
rect 26537 7349 26571 7365
rect 26537 6957 26571 6973
rect 26655 7349 26689 7365
rect 26655 6957 26689 6973
rect 26773 7349 26807 7365
rect 26773 6957 26807 6973
rect 26891 7349 26925 7365
rect 27198 7361 27232 7377
rect 26891 6957 26925 6973
rect 27325 7353 27359 7369
rect 27325 6961 27359 6977
rect 27443 7353 27477 7369
rect 27443 6961 27477 6977
rect 27561 7353 27595 7369
rect 27561 6961 27595 6977
rect 27679 7353 27713 7369
rect 27679 6961 27713 6977
rect 27797 7353 27831 7369
rect 27797 6961 27831 6977
rect 27915 7353 27949 7369
rect 27915 6961 27949 6977
rect 28033 7353 28067 7369
rect 29734 7361 29768 7377
rect 29852 7553 29886 7569
rect 29852 7361 29886 7377
rect 29970 7553 30004 7569
rect 29970 7361 30004 7377
rect 30088 7553 30122 7569
rect 30088 7361 30122 7377
rect 30206 7553 30240 7569
rect 30206 7361 30240 7377
rect 30324 7553 30358 7569
rect 30324 7361 30358 7377
rect 30442 7553 30476 7569
rect 30442 7361 30476 7377
rect 30560 7553 30594 7603
rect 30560 7361 30594 7377
rect 30678 7553 30712 7569
rect 30678 7361 30712 7377
rect 30796 7553 30830 7603
rect 30796 7361 30830 7377
rect 32316 7339 32586 7374
rect 30485 7283 30501 7317
rect 30535 7283 30551 7317
rect 31962 7286 31996 7302
rect 30367 7166 30383 7200
rect 30417 7166 30433 7200
rect 31478 7140 31748 7175
rect 28033 6961 28067 6977
rect 29971 7116 30005 7132
rect 17869 6889 17885 6923
rect 17919 6889 17935 6923
rect 24491 6890 24507 6924
rect 24541 6890 24557 6924
rect 17473 6839 17507 6855
rect 17473 6447 17507 6463
rect 17591 6839 17625 6855
rect 17591 6447 17625 6463
rect 17709 6839 17743 6855
rect 17826 6839 17860 6855
rect 17826 6647 17860 6663
rect 17944 6839 17978 6855
rect 17944 6647 17978 6663
rect 24095 6840 24129 6856
rect 19750 6616 19766 6650
rect 19800 6616 19816 6650
rect 20892 6620 20908 6654
rect 20942 6620 20958 6654
rect 19471 6565 19505 6581
rect 17709 6447 17743 6463
rect 17996 6513 18245 6556
rect 17996 6423 18043 6513
rect 18206 6423 18245 6513
rect 17516 6379 17532 6413
rect 17566 6379 17582 6413
rect 17634 6379 17650 6413
rect 17684 6379 17700 6413
rect 17996 6384 18245 6423
rect 19471 6373 19505 6389
rect 19589 6565 19623 6581
rect 19589 6373 19623 6389
rect 19707 6565 19741 6581
rect 19707 6373 19741 6389
rect 19825 6565 19859 6581
rect 19825 6373 19859 6389
rect 19990 6565 20024 6581
rect 19990 6373 20024 6389
rect 20108 6565 20142 6581
rect 20108 6373 20142 6389
rect 20226 6565 20260 6581
rect 20226 6373 20260 6389
rect 20344 6565 20378 6581
rect 20344 6373 20378 6389
rect 20613 6569 20647 6585
rect 20613 6377 20647 6393
rect 20731 6569 20765 6585
rect 20731 6377 20765 6393
rect 20849 6569 20883 6585
rect 20849 6377 20883 6393
rect 20967 6569 21001 6585
rect 20967 6377 21001 6393
rect 21132 6569 21166 6585
rect 21132 6377 21166 6393
rect 21250 6569 21284 6585
rect 21250 6377 21284 6393
rect 21368 6569 21402 6585
rect 21368 6377 21402 6393
rect 21486 6569 21520 6585
rect 24095 6448 24129 6464
rect 24213 6840 24247 6856
rect 24213 6448 24247 6464
rect 24331 6840 24365 6856
rect 24448 6840 24482 6856
rect 24448 6648 24482 6664
rect 24566 6840 24600 6856
rect 29971 6724 30005 6740
rect 30089 7116 30123 7132
rect 30089 6724 30123 6740
rect 30207 7116 30241 7132
rect 30324 7116 30358 7132
rect 30324 6924 30358 6940
rect 30442 7116 30476 7132
rect 30442 6924 30476 6940
rect 31478 7086 31512 7140
rect 31478 6894 31512 6910
rect 31596 7086 31630 7102
rect 31596 6894 31630 6910
rect 31714 7086 31748 7140
rect 31714 6894 31748 6910
rect 31832 7086 31866 7102
rect 31832 6894 31866 6910
rect 31962 6894 31996 6910
rect 32080 7286 32114 7302
rect 32080 6894 32114 6910
rect 32198 7286 32232 7302
rect 32198 6894 32232 6910
rect 32316 7286 32350 7339
rect 32316 6894 32350 6910
rect 32434 7286 32468 7302
rect 32434 6894 32468 6910
rect 32552 7286 32586 7339
rect 33560 7323 33728 7339
rect 32552 6894 32586 6910
rect 32670 7286 32704 7302
rect 33560 7253 33576 7323
rect 33712 7253 33728 7323
rect 33560 7237 33728 7253
rect 34097 7133 34367 7167
rect 32670 6894 32704 6910
rect 32799 7086 32833 7102
rect 32799 6894 32833 6910
rect 32917 7086 32951 7102
rect 32917 6894 32951 6910
rect 33035 7086 33069 7102
rect 33035 6894 33069 6910
rect 33153 7086 33187 7102
rect 33153 6894 33187 6910
rect 33271 7083 33305 7099
rect 33271 6891 33305 6907
rect 33389 7083 33423 7099
rect 33389 6891 33423 6907
rect 33507 7083 33541 7099
rect 33507 6891 33541 6907
rect 33625 7083 33659 7099
rect 33625 6891 33659 6907
rect 33743 7083 33777 7099
rect 33743 6891 33777 6907
rect 33861 7083 33895 7099
rect 33861 6891 33895 6907
rect 33979 7083 34013 7099
rect 33979 6891 34013 6907
rect 34097 7083 34131 7133
rect 34097 6891 34131 6907
rect 34215 7083 34249 7099
rect 34215 6891 34249 6907
rect 34333 7083 34367 7133
rect 34333 6891 34367 6907
rect 34022 6813 34038 6847
rect 34072 6813 34088 6847
rect 30207 6724 30241 6740
rect 33130 6728 33164 6744
rect 33904 6696 33920 6730
rect 33954 6696 33970 6730
rect 24566 6648 24600 6664
rect 30014 6656 30030 6690
rect 30064 6656 30080 6690
rect 30132 6656 30148 6690
rect 30182 6656 30198 6690
rect 33130 6678 33164 6694
rect 26372 6617 26388 6651
rect 26422 6617 26438 6651
rect 27514 6621 27530 6655
rect 27564 6621 27580 6655
rect 33508 6646 33542 6662
rect 31724 6609 31780 6626
rect 26093 6566 26127 6582
rect 24331 6448 24365 6464
rect 24618 6514 24867 6557
rect 24618 6424 24665 6514
rect 24828 6424 24867 6514
rect 21486 6377 21520 6393
rect 24138 6380 24154 6414
rect 24188 6380 24204 6414
rect 24256 6380 24272 6414
rect 24306 6380 24322 6414
rect 24618 6385 24867 6424
rect 26093 6374 26127 6390
rect 26211 6566 26245 6582
rect 26211 6374 26245 6390
rect 26329 6566 26363 6582
rect 26329 6374 26363 6390
rect 26447 6566 26481 6582
rect 26447 6374 26481 6390
rect 26612 6566 26646 6582
rect 26612 6374 26646 6390
rect 26730 6566 26764 6582
rect 26730 6374 26764 6390
rect 26848 6566 26882 6582
rect 26848 6374 26882 6390
rect 26966 6566 27000 6582
rect 26966 6374 27000 6390
rect 27235 6570 27269 6586
rect 27235 6378 27269 6394
rect 27353 6570 27387 6586
rect 27353 6378 27387 6394
rect 27471 6570 27505 6586
rect 27471 6378 27505 6394
rect 27589 6570 27623 6586
rect 27589 6378 27623 6394
rect 27754 6570 27788 6586
rect 27754 6378 27788 6394
rect 27872 6570 27906 6586
rect 27872 6378 27906 6394
rect 27990 6570 28024 6586
rect 27990 6378 28024 6394
rect 28108 6570 28142 6586
rect 30247 6585 30415 6603
rect 30247 6529 30263 6585
rect 30397 6529 30415 6585
rect 31724 6575 31730 6609
rect 31764 6575 31780 6609
rect 31724 6558 31780 6575
rect 31905 6593 31939 6609
rect 30247 6513 30415 6529
rect 28108 6378 28142 6394
rect 32023 6593 32057 6609
rect 31905 6201 31939 6217
rect 32022 6217 32023 6264
rect 32141 6593 32175 6609
rect 32057 6217 32058 6264
rect 19486 6142 19658 6189
rect 17645 6041 17868 6116
rect 17645 6040 17727 6041
rect 17645 5891 17724 6040
rect 17794 5892 17868 6041
rect 19486 5979 19525 6142
rect 19615 5979 19658 6142
rect 19486 5940 19658 5979
rect 20628 6140 20800 6187
rect 20628 5977 20667 6140
rect 20757 5977 20800 6140
rect 26108 6143 26280 6190
rect 20628 5938 20800 5977
rect 24267 6042 24490 6117
rect 17791 5891 17868 5892
rect 17645 5785 17868 5891
rect 24267 5892 24346 6042
rect 24413 5892 24490 6042
rect 26108 5980 26147 6143
rect 26237 5980 26280 6143
rect 26108 5941 26280 5980
rect 27250 6141 27422 6188
rect 27250 5978 27289 6141
rect 27379 5978 27422 6141
rect 32022 6159 32058 6217
rect 32259 6593 32293 6609
rect 32141 6201 32175 6217
rect 32257 6217 32259 6264
rect 32257 6159 32293 6217
rect 32377 6593 32411 6609
rect 32377 6201 32411 6217
rect 32495 6593 32529 6609
rect 32613 6593 32647 6609
rect 32529 6217 32531 6263
rect 32495 6159 32531 6217
rect 32775 6388 32845 6392
rect 32775 6297 32779 6388
rect 32841 6297 32845 6388
rect 32775 6292 32845 6297
rect 32613 6201 32647 6217
rect 32790 6159 32831 6292
rect 33508 6254 33542 6270
rect 33626 6646 33660 6662
rect 33626 6254 33660 6270
rect 33744 6646 33778 6662
rect 33861 6646 33895 6662
rect 33861 6454 33895 6470
rect 33979 6646 34013 6662
rect 33979 6454 34013 6470
rect 34451 6400 34581 12563
rect 36877 12492 36967 12526
rect 37143 12492 37159 12526
rect 36877 12290 36916 12492
rect 37441 12421 37526 12437
rect 36951 12374 36967 12408
rect 37143 12374 37233 12408
rect 36877 12256 36967 12290
rect 37143 12256 37159 12290
rect 37194 12172 37233 12374
rect 37441 12361 37458 12421
rect 37513 12361 37526 12421
rect 37441 12345 37526 12361
rect 36951 12138 36967 12172
rect 37143 12138 37233 12172
rect 36675 12051 36767 12085
rect 37143 12051 37159 12085
rect 36675 11849 36714 12051
rect 36751 11933 36767 11967
rect 37143 11933 37233 11967
rect 36675 11815 36767 11849
rect 37143 11815 37159 11849
rect 37194 11731 37233 11933
rect 36751 11697 36767 11731
rect 37143 11697 37233 11731
rect 36676 11584 36767 11618
rect 37143 11584 37159 11618
rect 36676 11382 36715 11584
rect 37194 11500 37233 11697
rect 38084 11658 38100 11692
rect 38276 11658 38292 11692
rect 38084 11540 38100 11574
rect 38276 11540 38292 11574
rect 38088 11500 38288 11540
rect 36751 11466 36767 11500
rect 37143 11466 37233 11500
rect 36479 11340 36589 11356
rect 36676 11348 36767 11382
rect 37143 11348 37159 11382
rect 36479 11144 36497 11340
rect 36573 11144 36589 11340
rect 37194 11264 37233 11466
rect 37729 11454 37814 11470
rect 38084 11466 38100 11500
rect 38476 11466 38492 11500
rect 37342 11406 37358 11440
rect 37392 11406 37408 11440
rect 37729 11394 37742 11454
rect 37797 11394 37814 11454
rect 37729 11378 37814 11394
rect 36751 11230 36767 11264
rect 37143 11230 37233 11264
rect 37444 11336 37529 11352
rect 38084 11348 38100 11382
rect 38476 11348 38492 11382
rect 37444 11276 37457 11336
rect 37512 11276 37529 11336
rect 38725 11282 38811 11298
rect 37444 11260 37529 11276
rect 38084 11230 38100 11264
rect 38476 11230 38492 11264
rect 38577 11263 38611 11279
rect 36479 11128 36589 11144
rect 36676 11112 36767 11146
rect 37143 11112 37159 11146
rect 36676 10910 36715 11112
rect 37194 11028 37233 11230
rect 38577 11213 38611 11229
rect 38725 11260 38743 11282
rect 37962 11171 37978 11205
rect 38012 11171 38028 11205
rect 38725 11202 38729 11260
rect 38725 11178 38743 11202
rect 38789 11178 38811 11282
rect 38725 11162 38811 11178
rect 38084 11112 38100 11146
rect 38476 11112 38492 11146
rect 37572 11052 37588 11086
rect 37622 11052 37638 11086
rect 36751 10994 36767 11028
rect 37143 10994 37233 11028
rect 38084 10994 38100 11028
rect 38476 10994 38492 11028
rect 36676 10876 36767 10910
rect 37143 10876 37159 10910
rect 37194 10791 37233 10994
rect 38088 10950 38288 10994
rect 38084 10916 38100 10950
rect 38276 10916 38292 10950
rect 38084 10798 38100 10832
rect 38276 10798 38292 10832
rect 36751 10757 36767 10791
rect 37143 10757 37233 10791
rect 36676 10639 36767 10673
rect 37143 10639 37159 10673
rect 36676 10437 36715 10639
rect 37194 10555 37233 10757
rect 36751 10521 36767 10555
rect 37143 10521 37233 10555
rect 36676 10403 36767 10437
rect 37143 10403 37159 10437
rect 36951 10284 36967 10318
rect 37143 10284 37236 10318
rect 36880 10166 36967 10200
rect 37143 10166 37159 10200
rect 36880 9964 36917 10166
rect 37197 10082 37236 10284
rect 36951 10048 36967 10082
rect 37143 10048 37236 10082
rect 37317 10130 37351 10146
rect 37317 10080 37351 10096
rect 36880 9930 36967 9964
rect 37143 9930 37159 9964
rect 36877 9348 36967 9382
rect 37143 9348 37159 9382
rect 36877 9146 36916 9348
rect 37441 9277 37526 9293
rect 36951 9230 36967 9264
rect 37143 9230 37233 9264
rect 36877 9112 36967 9146
rect 37143 9112 37159 9146
rect 37194 9028 37233 9230
rect 37441 9217 37458 9277
rect 37513 9217 37526 9277
rect 37441 9201 37526 9217
rect 36951 8994 36967 9028
rect 37143 8994 37233 9028
rect 36675 8907 36767 8941
rect 37143 8907 37159 8941
rect 36675 8705 36714 8907
rect 36751 8789 36767 8823
rect 37143 8789 37233 8823
rect 36675 8671 36767 8705
rect 37143 8671 37159 8705
rect 37194 8587 37233 8789
rect 36751 8553 36767 8587
rect 37143 8553 37233 8587
rect 36676 8440 36767 8474
rect 37143 8440 37159 8474
rect 36676 8238 36715 8440
rect 37194 8356 37233 8553
rect 38084 8514 38100 8548
rect 38276 8514 38292 8548
rect 38084 8396 38100 8430
rect 38276 8396 38292 8430
rect 38088 8356 38288 8396
rect 36751 8322 36767 8356
rect 37143 8322 37233 8356
rect 36479 8196 36589 8212
rect 36676 8204 36767 8238
rect 37143 8204 37159 8238
rect 36479 8000 36497 8196
rect 36573 8000 36589 8196
rect 37194 8120 37233 8322
rect 37729 8310 37814 8326
rect 38084 8322 38100 8356
rect 38476 8322 38492 8356
rect 37342 8262 37358 8296
rect 37392 8262 37408 8296
rect 37729 8250 37742 8310
rect 37797 8250 37814 8310
rect 37729 8234 37814 8250
rect 36751 8086 36767 8120
rect 37143 8086 37233 8120
rect 37444 8192 37529 8208
rect 38084 8204 38100 8238
rect 38476 8204 38492 8238
rect 37444 8132 37457 8192
rect 37512 8132 37529 8192
rect 38725 8138 38811 8154
rect 37444 8116 37529 8132
rect 38084 8086 38100 8120
rect 38476 8086 38492 8120
rect 38577 8119 38611 8135
rect 36479 7984 36589 8000
rect 36676 7968 36767 8002
rect 37143 7968 37159 8002
rect 36676 7766 36715 7968
rect 37194 7884 37233 8086
rect 38577 8069 38611 8085
rect 38725 8116 38743 8138
rect 37962 8027 37978 8061
rect 38012 8027 38028 8061
rect 38725 8058 38729 8116
rect 38725 8034 38743 8058
rect 38789 8034 38811 8138
rect 38725 8018 38811 8034
rect 38084 7968 38100 8002
rect 38476 7968 38492 8002
rect 37572 7908 37588 7942
rect 37622 7908 37638 7942
rect 36751 7850 36767 7884
rect 37143 7850 37233 7884
rect 38084 7850 38100 7884
rect 38476 7850 38492 7884
rect 36676 7732 36767 7766
rect 37143 7732 37159 7766
rect 37194 7647 37233 7850
rect 38088 7806 38288 7850
rect 38084 7772 38100 7806
rect 38276 7772 38292 7806
rect 38084 7654 38100 7688
rect 38276 7654 38292 7688
rect 36751 7613 36767 7647
rect 37143 7613 37233 7647
rect 36676 7495 36767 7529
rect 37143 7495 37159 7529
rect 36676 7293 36715 7495
rect 37194 7411 37233 7613
rect 36751 7377 36767 7411
rect 37143 7377 37233 7411
rect 36676 7259 36767 7293
rect 37143 7259 37159 7293
rect 36951 7140 36967 7174
rect 37143 7140 37236 7174
rect 36880 7022 36967 7056
rect 37143 7022 37159 7056
rect 36880 6820 36917 7022
rect 37197 6938 37236 7140
rect 36951 6904 36967 6938
rect 37143 6904 37236 6938
rect 37317 6986 37351 7002
rect 37317 6936 37351 6952
rect 36880 6786 36967 6820
rect 37143 6786 37159 6820
rect 34651 6486 37812 6503
rect 34651 6418 34662 6486
rect 34728 6418 37812 6486
rect 34651 6408 37812 6418
rect 34404 6375 34581 6400
rect 34404 6303 34434 6375
rect 34529 6303 34581 6375
rect 37723 6389 37812 6408
rect 37723 6340 37737 6389
rect 37797 6340 37812 6389
rect 37723 6320 37812 6340
rect 34404 6287 34581 6303
rect 33744 6254 33778 6270
rect 33551 6186 33567 6220
rect 33601 6186 33617 6220
rect 33669 6186 33685 6220
rect 33719 6186 33735 6220
rect 36873 6216 36963 6250
rect 37139 6216 37155 6250
rect 32022 6119 32831 6159
rect 32041 6118 32831 6119
rect 31919 6029 31986 6045
rect 31919 5995 31935 6029
rect 31969 5995 31986 6029
rect 31919 5979 31986 5995
rect 27250 5939 27422 5978
rect 31750 5962 31784 5978
rect 31750 5912 31784 5928
rect 24267 5786 24490 5892
rect 32096 5877 32130 6118
rect 33784 6115 33952 6133
rect 33784 6059 33800 6115
rect 33934 6059 33952 6115
rect 32566 6029 32633 6045
rect 33784 6043 33952 6059
rect 32566 5995 32583 6029
rect 32617 5995 32633 6029
rect 32566 5979 32633 5995
rect 36873 6014 36912 6216
rect 37437 6145 37522 6161
rect 36947 6098 36963 6132
rect 37139 6098 37229 6132
rect 36873 5980 36963 6014
rect 37139 5980 37155 6014
rect 32873 5961 32907 5977
rect 32185 5911 32201 5945
rect 32235 5911 32251 5945
rect 32303 5912 32319 5946
rect 32353 5912 32369 5946
rect 32873 5911 32907 5927
rect 37190 5896 37229 6098
rect 37437 6085 37454 6145
rect 37509 6085 37522 6145
rect 37437 6069 37522 6085
rect 31603 5861 31637 5877
rect 18076 5676 18346 5710
rect 17250 5626 17284 5642
rect 17250 5434 17284 5450
rect 17368 5626 17402 5642
rect 17368 5434 17402 5450
rect 17486 5626 17520 5642
rect 17486 5434 17520 5450
rect 17604 5626 17638 5642
rect 17604 5434 17638 5450
rect 17722 5626 17756 5642
rect 17722 5434 17756 5450
rect 17840 5626 17874 5642
rect 17840 5434 17874 5450
rect 17958 5626 17992 5642
rect 17958 5434 17992 5450
rect 18076 5626 18110 5676
rect 18076 5434 18110 5450
rect 18194 5626 18228 5642
rect 18194 5434 18228 5450
rect 18312 5626 18346 5676
rect 18312 5434 18346 5450
rect 21356 5699 21581 5773
rect 21356 5697 21438 5699
rect 21356 5548 21435 5697
rect 21505 5550 21581 5699
rect 24698 5677 24968 5711
rect 21502 5548 21581 5550
rect 21356 5442 21581 5548
rect 23872 5627 23906 5643
rect 23872 5435 23906 5451
rect 23990 5627 24024 5643
rect 23990 5435 24024 5451
rect 24108 5627 24142 5643
rect 24108 5435 24142 5451
rect 24226 5627 24260 5643
rect 24226 5435 24260 5451
rect 24344 5627 24378 5643
rect 24344 5435 24378 5451
rect 24462 5627 24496 5643
rect 24462 5435 24496 5451
rect 24580 5627 24614 5643
rect 24580 5435 24614 5451
rect 24698 5627 24732 5677
rect 24698 5435 24732 5451
rect 24816 5627 24850 5643
rect 24816 5435 24850 5451
rect 24934 5627 24968 5677
rect 24934 5435 24968 5451
rect 27978 5698 28203 5774
rect 27978 5549 28057 5698
rect 28124 5697 28203 5698
rect 27978 5548 28059 5549
rect 28126 5548 28203 5697
rect 31603 5669 31637 5685
rect 31721 5861 31755 5877
rect 31721 5669 31755 5685
rect 32023 5861 32057 5877
rect 27978 5443 28203 5548
rect 32096 5861 32175 5877
rect 32096 5831 32141 5861
rect 32023 5418 32058 5485
rect 32141 5469 32175 5485
rect 32259 5861 32293 5877
rect 32259 5469 32293 5485
rect 32377 5861 32411 5877
rect 32495 5861 32529 5877
rect 32901 5861 32935 5877
rect 32901 5669 32935 5685
rect 33019 5861 33053 5877
rect 36947 5862 36963 5896
rect 37139 5862 37229 5896
rect 33019 5669 33053 5685
rect 36671 5775 36763 5809
rect 37139 5775 37155 5809
rect 36671 5573 36710 5775
rect 36747 5657 36763 5691
rect 37139 5657 37229 5691
rect 36671 5539 36763 5573
rect 37139 5539 37155 5573
rect 32377 5469 32411 5485
rect 32494 5418 32529 5485
rect 37190 5455 37229 5657
rect 36747 5421 36763 5455
rect 37139 5421 37229 5455
rect 18001 5356 18017 5390
rect 18051 5356 18067 5390
rect 24623 5357 24639 5391
rect 24673 5357 24689 5391
rect 32023 5383 32529 5418
rect 32170 5314 32412 5326
rect 17883 5239 17899 5273
rect 17933 5239 17949 5273
rect 19552 5262 19822 5297
rect 19198 5209 19232 5225
rect 17487 5189 17521 5205
rect 17487 4797 17521 4813
rect 17605 5189 17639 5205
rect 17605 4797 17639 4813
rect 17723 5189 17757 5205
rect 17840 5189 17874 5205
rect 17840 4997 17874 5013
rect 17958 5189 17992 5205
rect 17958 4997 17992 5013
rect 18714 5063 18984 5098
rect 18714 5009 18748 5063
rect 17723 4797 17757 4813
rect 18010 4863 18259 4906
rect 18010 4773 18057 4863
rect 18220 4773 18259 4863
rect 18714 4817 18748 4833
rect 18832 5009 18866 5025
rect 18832 4817 18866 4833
rect 18950 5009 18984 5063
rect 18950 4817 18984 4833
rect 19068 5009 19102 5025
rect 19068 4817 19102 4833
rect 19198 4817 19232 4833
rect 19316 5209 19350 5225
rect 19316 4817 19350 4833
rect 19434 5209 19468 5225
rect 19434 4817 19468 4833
rect 19552 5209 19586 5262
rect 19552 4817 19586 4833
rect 19670 5209 19704 5225
rect 19670 4817 19704 4833
rect 19788 5209 19822 5262
rect 21450 5262 21720 5297
rect 19788 4817 19822 4833
rect 19906 5209 19940 5225
rect 21096 5209 21130 5225
rect 20612 5063 20882 5098
rect 19906 4817 19940 4833
rect 20035 5009 20069 5025
rect 20035 4817 20069 4833
rect 20153 5009 20187 5025
rect 20153 4817 20187 4833
rect 20271 5009 20305 5025
rect 20271 4817 20305 4833
rect 20389 5009 20423 5025
rect 20389 4817 20423 4833
rect 20612 5009 20646 5063
rect 20612 4817 20646 4833
rect 20730 5009 20764 5025
rect 20730 4817 20764 4833
rect 20848 5009 20882 5063
rect 20848 4817 20882 4833
rect 20966 5009 21000 5025
rect 20966 4817 21000 4833
rect 21096 4817 21130 4833
rect 21214 5209 21248 5225
rect 21214 4817 21248 4833
rect 21332 5209 21366 5225
rect 21332 4817 21366 4833
rect 21450 5209 21484 5262
rect 21450 4817 21484 4833
rect 21568 5209 21602 5225
rect 21568 4817 21602 4833
rect 21686 5209 21720 5262
rect 24505 5240 24521 5274
rect 24555 5240 24571 5274
rect 26174 5263 26444 5298
rect 21686 4817 21720 4833
rect 21804 5209 21838 5225
rect 25820 5210 25854 5226
rect 24109 5190 24143 5206
rect 21804 4817 21838 4833
rect 21933 5009 21967 5025
rect 21933 4817 21967 4833
rect 22051 5009 22085 5025
rect 22051 4817 22085 4833
rect 22169 5009 22203 5025
rect 22169 4817 22203 4833
rect 22287 5009 22321 5025
rect 22287 4817 22321 4833
rect 24109 4798 24143 4814
rect 24227 5190 24261 5206
rect 24227 4798 24261 4814
rect 24345 5190 24379 5206
rect 24462 5190 24496 5206
rect 24462 4998 24496 5014
rect 24580 5190 24614 5206
rect 24580 4998 24614 5014
rect 25336 5064 25606 5099
rect 25336 5010 25370 5064
rect 24345 4798 24379 4814
rect 24632 4864 24881 4907
rect 17530 4729 17546 4763
rect 17580 4729 17596 4763
rect 17648 4729 17664 4763
rect 17698 4729 17714 4763
rect 18010 4734 18259 4773
rect 24632 4774 24679 4864
rect 24842 4774 24881 4864
rect 25336 4818 25370 4834
rect 25454 5010 25488 5026
rect 25454 4818 25488 4834
rect 25572 5010 25606 5064
rect 25572 4818 25606 4834
rect 25690 5010 25724 5026
rect 25690 4818 25724 4834
rect 25820 4818 25854 4834
rect 25938 5210 25972 5226
rect 25938 4818 25972 4834
rect 26056 5210 26090 5226
rect 26056 4818 26090 4834
rect 26174 5210 26208 5263
rect 26174 4818 26208 4834
rect 26292 5210 26326 5226
rect 26292 4818 26326 4834
rect 26410 5210 26444 5263
rect 28072 5263 28342 5298
rect 26410 4818 26444 4834
rect 26528 5210 26562 5226
rect 27718 5210 27752 5226
rect 27234 5064 27504 5099
rect 26528 4818 26562 4834
rect 26657 5010 26691 5026
rect 26657 4818 26691 4834
rect 26775 5010 26809 5026
rect 26775 4818 26809 4834
rect 26893 5010 26927 5026
rect 26893 4818 26927 4834
rect 27011 5010 27045 5026
rect 27011 4818 27045 4834
rect 27234 5010 27268 5064
rect 27234 4818 27268 4834
rect 27352 5010 27386 5026
rect 27352 4818 27386 4834
rect 27470 5010 27504 5064
rect 27470 4818 27504 4834
rect 27588 5010 27622 5026
rect 27588 4818 27622 4834
rect 27718 4818 27752 4834
rect 27836 5210 27870 5226
rect 27836 4818 27870 4834
rect 27954 5210 27988 5226
rect 27954 4818 27988 4834
rect 28072 5210 28106 5263
rect 28072 4818 28106 4834
rect 28190 5210 28224 5226
rect 28190 4818 28224 4834
rect 28308 5210 28342 5263
rect 28308 4818 28342 4834
rect 28426 5210 28460 5226
rect 32170 5212 32217 5314
rect 32352 5212 32412 5314
rect 32170 5195 32412 5212
rect 36672 5308 36763 5342
rect 37139 5308 37155 5342
rect 36672 5106 36711 5308
rect 37190 5224 37229 5421
rect 38080 5382 38096 5416
rect 38272 5382 38288 5416
rect 38080 5264 38096 5298
rect 38272 5264 38288 5298
rect 38084 5224 38284 5264
rect 36747 5190 36763 5224
rect 37139 5190 37229 5224
rect 36475 5064 36585 5080
rect 36672 5072 36763 5106
rect 37139 5072 37155 5106
rect 28426 4818 28460 4834
rect 28555 5010 28589 5026
rect 28555 4818 28589 4834
rect 28673 5010 28707 5026
rect 28673 4818 28707 4834
rect 28791 5010 28825 5026
rect 28791 4818 28825 4834
rect 28909 5010 28943 5026
rect 36475 4868 36493 5064
rect 36569 4868 36585 5064
rect 37190 4988 37229 5190
rect 37725 5178 37810 5194
rect 38080 5190 38096 5224
rect 38472 5190 38488 5224
rect 37338 5130 37354 5164
rect 37388 5130 37404 5164
rect 37725 5118 37738 5178
rect 37793 5118 37810 5178
rect 37725 5102 37810 5118
rect 36747 4954 36763 4988
rect 37139 4954 37229 4988
rect 37440 5060 37525 5076
rect 38080 5072 38096 5106
rect 38472 5072 38488 5106
rect 37440 5000 37453 5060
rect 37508 5000 37525 5060
rect 38721 5006 38807 5022
rect 37440 4984 37525 5000
rect 38080 4954 38096 4988
rect 38472 4954 38488 4988
rect 38573 4987 38607 5003
rect 36475 4852 36585 4868
rect 28909 4818 28943 4834
rect 36672 4836 36763 4870
rect 37139 4836 37155 4870
rect 24152 4730 24168 4764
rect 24202 4730 24218 4764
rect 24270 4730 24286 4764
rect 24320 4730 24336 4764
rect 24632 4735 24881 4774
rect 30020 4723 30188 4739
rect 30020 4653 30036 4723
rect 30172 4653 30188 4723
rect 30020 4637 30188 4653
rect 36672 4634 36711 4836
rect 37190 4752 37229 4954
rect 38573 4937 38607 4953
rect 38721 4984 38739 5006
rect 37958 4895 37974 4929
rect 38008 4895 38024 4929
rect 38721 4926 38725 4984
rect 38721 4902 38739 4926
rect 38785 4902 38807 5006
rect 38721 4886 38807 4902
rect 38080 4836 38096 4870
rect 38472 4836 38488 4870
rect 37568 4776 37584 4810
rect 37618 4776 37634 4810
rect 36747 4718 36763 4752
rect 37139 4718 37229 4752
rect 38080 4718 38096 4752
rect 38472 4718 38488 4752
rect 20178 4595 20212 4611
rect 26800 4596 26834 4612
rect 36672 4600 36763 4634
rect 37139 4600 37155 4634
rect 20178 4545 20212 4561
rect 22268 4574 22335 4590
rect 22268 4540 22285 4574
rect 22319 4540 22335 4574
rect 26800 4546 26834 4562
rect 28890 4575 28957 4591
rect 19141 4516 19175 4532
rect 17640 4436 17863 4512
rect 17640 4287 17719 4436
rect 17786 4433 17863 4436
rect 17640 4284 17722 4287
rect 17789 4284 17863 4433
rect 17640 4181 17863 4284
rect 19259 4516 19293 4532
rect 19141 4124 19175 4140
rect 19258 4140 19259 4187
rect 19377 4516 19411 4532
rect 19293 4140 19294 4187
rect 18071 4072 18341 4106
rect 17245 4022 17279 4038
rect 17245 3830 17279 3846
rect 17363 4022 17397 4038
rect 17363 3830 17397 3846
rect 17481 4022 17515 4038
rect 17481 3830 17515 3846
rect 17599 4022 17633 4038
rect 17599 3830 17633 3846
rect 17717 4022 17751 4038
rect 17717 3830 17751 3846
rect 17835 4022 17869 4038
rect 17835 3830 17869 3846
rect 17953 4022 17987 4038
rect 17953 3830 17987 3846
rect 18071 4022 18105 4072
rect 18071 3830 18105 3846
rect 18189 4022 18223 4038
rect 18189 3830 18223 3846
rect 18307 4022 18341 4072
rect 19258 4082 19294 4140
rect 19495 4516 19529 4532
rect 19377 4124 19411 4140
rect 19493 4140 19495 4187
rect 19493 4082 19529 4140
rect 19613 4516 19647 4532
rect 19613 4124 19647 4140
rect 19731 4516 19765 4532
rect 19849 4516 19883 4532
rect 19765 4140 19767 4186
rect 19731 4082 19767 4140
rect 19849 4124 19883 4140
rect 21039 4516 21073 4532
rect 21157 4516 21191 4532
rect 21039 4124 21073 4140
rect 21156 4140 21157 4187
rect 21275 4516 21309 4532
rect 21191 4140 21192 4187
rect 20354 4082 20851 4100
rect 19258 4079 20851 4082
rect 19258 4045 20799 4079
rect 20833 4045 20851 4079
rect 19258 4042 20851 4045
rect 21156 4082 21192 4140
rect 21393 4516 21427 4532
rect 21275 4124 21309 4140
rect 21391 4140 21393 4187
rect 21391 4082 21427 4140
rect 21511 4516 21545 4532
rect 21511 4124 21545 4140
rect 21629 4516 21663 4532
rect 21747 4516 21781 4532
rect 22268 4524 22335 4540
rect 28890 4541 28907 4575
rect 28941 4541 28957 4575
rect 21663 4140 21665 4186
rect 21629 4082 21665 4140
rect 25763 4517 25797 4533
rect 24262 4437 24485 4513
rect 24262 4288 24341 4437
rect 24408 4433 24485 4437
rect 24262 4284 24343 4288
rect 24410 4284 24485 4433
rect 24262 4182 24485 4284
rect 21747 4124 21781 4140
rect 25881 4517 25915 4533
rect 25763 4125 25797 4141
rect 25880 4141 25881 4188
rect 25999 4517 26033 4533
rect 25915 4141 25916 4188
rect 22252 4111 22352 4112
rect 22252 4082 22408 4111
rect 21156 4042 22408 4082
rect 19277 4041 20851 4042
rect 21175 4041 22408 4042
rect 19155 3952 19222 3968
rect 19155 3918 19171 3952
rect 19205 3918 19222 3952
rect 19155 3902 19222 3918
rect 18307 3830 18341 3846
rect 18986 3885 19020 3901
rect 18986 3835 19020 3851
rect 19332 3800 19366 4041
rect 20354 4024 20851 4041
rect 19802 3952 19869 3968
rect 19802 3918 19819 3952
rect 19853 3918 19869 3952
rect 19802 3902 19869 3918
rect 21053 3952 21120 3968
rect 21053 3918 21069 3952
rect 21103 3918 21120 3952
rect 21053 3902 21120 3918
rect 20109 3884 20143 3900
rect 19421 3834 19437 3868
rect 19471 3834 19487 3868
rect 19539 3835 19555 3869
rect 19589 3835 19605 3869
rect 20109 3834 20143 3850
rect 20884 3885 20918 3901
rect 20884 3835 20918 3851
rect 21230 3800 21264 4041
rect 22252 4013 22408 4041
rect 24693 4073 24963 4107
rect 23867 4023 23901 4039
rect 22252 4012 22352 4013
rect 21698 3953 21765 3969
rect 21698 3919 21715 3953
rect 21749 3919 21765 3953
rect 21698 3903 21765 3919
rect 22007 3884 22041 3900
rect 21319 3834 21335 3868
rect 21369 3834 21385 3868
rect 21437 3835 21453 3869
rect 21487 3835 21503 3869
rect 22007 3834 22041 3850
rect 23867 3831 23901 3847
rect 23985 4023 24019 4039
rect 23985 3831 24019 3847
rect 24103 4023 24137 4039
rect 24103 3831 24137 3847
rect 24221 4023 24255 4039
rect 24221 3831 24255 3847
rect 24339 4023 24373 4039
rect 24339 3831 24373 3847
rect 24457 4023 24491 4039
rect 24457 3831 24491 3847
rect 24575 4023 24609 4039
rect 24575 3831 24609 3847
rect 24693 4023 24727 4073
rect 24693 3831 24727 3847
rect 24811 4023 24845 4039
rect 24811 3831 24845 3847
rect 24929 4023 24963 4073
rect 25880 4083 25916 4141
rect 26117 4517 26151 4533
rect 25999 4125 26033 4141
rect 26115 4141 26117 4188
rect 26115 4083 26151 4141
rect 26235 4517 26269 4533
rect 26235 4125 26269 4141
rect 26353 4517 26387 4533
rect 26471 4517 26505 4533
rect 26387 4141 26389 4187
rect 26353 4083 26389 4141
rect 26471 4125 26505 4141
rect 27661 4517 27695 4533
rect 27779 4517 27813 4533
rect 27661 4125 27695 4141
rect 27778 4141 27779 4188
rect 27897 4517 27931 4533
rect 27813 4141 27814 4188
rect 26976 4083 27473 4101
rect 25880 4080 27473 4083
rect 25880 4046 27421 4080
rect 27455 4046 27473 4080
rect 25880 4043 27473 4046
rect 27778 4083 27814 4141
rect 28015 4517 28049 4533
rect 27897 4125 27931 4141
rect 28013 4141 28015 4188
rect 28013 4083 28049 4141
rect 28133 4517 28167 4533
rect 28133 4125 28167 4141
rect 28251 4517 28285 4533
rect 28369 4517 28403 4533
rect 28890 4525 28957 4541
rect 30557 4533 30827 4567
rect 28285 4141 28287 4187
rect 28251 4083 28287 4141
rect 29731 4483 29765 4499
rect 29731 4291 29765 4307
rect 29849 4483 29883 4499
rect 29849 4291 29883 4307
rect 29967 4483 30001 4499
rect 29967 4291 30001 4307
rect 30085 4483 30119 4499
rect 30085 4291 30119 4307
rect 30203 4483 30237 4499
rect 30203 4291 30237 4307
rect 30321 4483 30355 4499
rect 30321 4291 30355 4307
rect 30439 4483 30473 4499
rect 30439 4291 30473 4307
rect 30557 4483 30591 4533
rect 30557 4291 30591 4307
rect 30675 4483 30709 4499
rect 30675 4291 30709 4307
rect 30793 4483 30827 4533
rect 37190 4515 37229 4718
rect 38084 4674 38284 4718
rect 38080 4640 38096 4674
rect 38272 4640 38288 4674
rect 38080 4522 38096 4556
rect 38272 4522 38288 4556
rect 36747 4481 36763 4515
rect 37139 4481 37229 4515
rect 30793 4291 30827 4307
rect 36672 4363 36763 4397
rect 37139 4363 37155 4397
rect 30482 4213 30498 4247
rect 30532 4213 30548 4247
rect 28369 4125 28403 4141
rect 36672 4161 36711 4363
rect 37190 4279 37229 4481
rect 36747 4245 36763 4279
rect 37139 4245 37229 4279
rect 28874 4112 28974 4113
rect 28874 4083 29030 4112
rect 27778 4043 29030 4083
rect 25899 4042 27473 4043
rect 27797 4042 29030 4043
rect 25777 3953 25844 3969
rect 25777 3919 25793 3953
rect 25827 3919 25844 3953
rect 25777 3903 25844 3919
rect 24929 3831 24963 3847
rect 25608 3886 25642 3902
rect 25608 3836 25642 3852
rect 25954 3801 25988 4042
rect 26976 4025 27473 4042
rect 26424 3953 26491 3969
rect 26424 3919 26441 3953
rect 26475 3919 26491 3953
rect 26424 3903 26491 3919
rect 27675 3953 27742 3969
rect 27675 3919 27691 3953
rect 27725 3919 27742 3953
rect 27675 3903 27742 3919
rect 26731 3885 26765 3901
rect 26043 3835 26059 3869
rect 26093 3835 26109 3869
rect 26161 3836 26177 3870
rect 26211 3836 26227 3870
rect 26731 3835 26765 3851
rect 27506 3886 27540 3902
rect 27506 3836 27540 3852
rect 27852 3801 27886 4042
rect 28874 4014 29030 4042
rect 30364 4096 30380 4130
rect 30414 4096 30430 4130
rect 36672 4127 36763 4161
rect 37139 4127 37155 4161
rect 29968 4046 30002 4062
rect 28874 4013 28974 4014
rect 28320 3954 28387 3970
rect 28320 3920 28337 3954
rect 28371 3920 28387 3954
rect 28320 3904 28387 3920
rect 28629 3885 28663 3901
rect 27941 3835 27957 3869
rect 27991 3835 28007 3869
rect 28059 3836 28075 3870
rect 28109 3836 28125 3870
rect 28629 3835 28663 3851
rect 17996 3752 18012 3786
rect 18046 3752 18062 3786
rect 18839 3784 18873 3800
rect 17878 3635 17894 3669
rect 17928 3635 17944 3669
rect 17482 3585 17516 3601
rect 17482 3193 17516 3209
rect 17600 3585 17634 3601
rect 17600 3193 17634 3209
rect 17718 3585 17752 3601
rect 17835 3585 17869 3601
rect 17835 3393 17869 3409
rect 17953 3585 17987 3601
rect 18839 3592 18873 3608
rect 18957 3784 18991 3800
rect 18957 3592 18991 3608
rect 19259 3784 19293 3800
rect 17953 3393 17987 3409
rect 19332 3784 19411 3800
rect 19332 3754 19377 3784
rect 19259 3341 19294 3408
rect 19377 3392 19411 3408
rect 19495 3784 19529 3800
rect 19495 3392 19529 3408
rect 19613 3784 19647 3800
rect 19731 3784 19765 3800
rect 20137 3784 20171 3800
rect 20137 3592 20171 3608
rect 20255 3784 20289 3800
rect 20255 3592 20289 3608
rect 20737 3784 20771 3800
rect 20737 3592 20771 3608
rect 20855 3784 20889 3800
rect 20855 3592 20889 3608
rect 21157 3784 21191 3800
rect 19613 3392 19647 3408
rect 19730 3341 19765 3408
rect 19259 3306 19765 3341
rect 21230 3784 21309 3800
rect 21230 3754 21275 3784
rect 21157 3341 21192 3408
rect 21275 3392 21309 3408
rect 21393 3784 21427 3800
rect 21393 3392 21427 3408
rect 21511 3784 21545 3800
rect 21629 3784 21663 3800
rect 22035 3784 22069 3800
rect 22035 3592 22069 3608
rect 22153 3784 22187 3800
rect 24618 3753 24634 3787
rect 24668 3753 24684 3787
rect 25461 3785 25495 3801
rect 24500 3636 24516 3670
rect 24550 3636 24566 3670
rect 22153 3592 22187 3608
rect 21511 3392 21545 3408
rect 21628 3341 21663 3408
rect 21157 3306 21663 3341
rect 24104 3586 24138 3602
rect 17718 3193 17752 3209
rect 18005 3259 18254 3302
rect 18005 3169 18052 3259
rect 18215 3239 18254 3259
rect 18218 3172 18254 3239
rect 24104 3194 24138 3210
rect 24222 3586 24256 3602
rect 24222 3194 24256 3210
rect 24340 3586 24374 3602
rect 24457 3586 24491 3602
rect 24457 3394 24491 3410
rect 24575 3586 24609 3602
rect 25461 3593 25495 3609
rect 25579 3785 25613 3801
rect 25579 3593 25613 3609
rect 25881 3785 25915 3801
rect 24575 3394 24609 3410
rect 25954 3785 26033 3801
rect 25954 3755 25999 3785
rect 25881 3342 25916 3409
rect 25999 3393 26033 3409
rect 26117 3785 26151 3801
rect 26117 3393 26151 3409
rect 26235 3785 26269 3801
rect 26353 3785 26387 3801
rect 26759 3785 26793 3801
rect 26759 3593 26793 3609
rect 26877 3785 26911 3801
rect 26877 3593 26911 3609
rect 27359 3785 27393 3801
rect 27359 3593 27393 3609
rect 27477 3785 27511 3801
rect 27477 3593 27511 3609
rect 27779 3785 27813 3801
rect 26235 3393 26269 3409
rect 26352 3342 26387 3409
rect 25881 3307 26387 3342
rect 27852 3785 27931 3801
rect 27852 3755 27897 3785
rect 27779 3342 27814 3409
rect 27897 3393 27931 3409
rect 28015 3785 28049 3801
rect 28015 3393 28049 3409
rect 28133 3785 28167 3801
rect 28251 3785 28285 3801
rect 28657 3785 28691 3801
rect 28657 3593 28691 3609
rect 28775 3785 28809 3801
rect 29968 3654 30002 3670
rect 30086 4046 30120 4062
rect 30086 3654 30120 3670
rect 30204 4046 30238 4062
rect 30321 4046 30355 4062
rect 30321 3854 30355 3870
rect 30439 4046 30473 4062
rect 36947 4008 36963 4042
rect 37139 4008 37232 4042
rect 30439 3854 30473 3870
rect 36876 3890 36963 3924
rect 37139 3890 37155 3924
rect 30204 3654 30238 3670
rect 36876 3688 36913 3890
rect 37193 3806 37232 4008
rect 36947 3772 36963 3806
rect 37139 3772 37232 3806
rect 37313 3854 37347 3870
rect 37313 3804 37347 3820
rect 36876 3654 36963 3688
rect 37139 3654 37155 3688
rect 28775 3593 28809 3609
rect 30011 3586 30027 3620
rect 30061 3586 30077 3620
rect 30129 3586 30145 3620
rect 30179 3586 30195 3620
rect 30244 3515 30412 3533
rect 30244 3459 30260 3515
rect 30394 3459 30412 3515
rect 30244 3443 30412 3459
rect 32101 3476 32545 3482
rect 28133 3393 28167 3409
rect 28250 3342 28285 3409
rect 27779 3307 28285 3342
rect 24340 3194 24374 3210
rect 24627 3260 24876 3303
rect 32101 3276 32112 3476
rect 32533 3276 32545 3476
rect 32101 3270 32545 3276
rect 34779 3349 34897 3361
rect 34779 3341 37809 3349
rect 34779 3275 34797 3341
rect 34890 3297 37809 3341
rect 34890 3275 37810 3297
rect 34779 3268 37810 3275
rect 18215 3169 18254 3172
rect 17525 3125 17541 3159
rect 17575 3125 17591 3159
rect 17643 3125 17659 3159
rect 17693 3125 17709 3159
rect 18005 3130 18254 3169
rect 24627 3170 24674 3260
rect 24837 3170 24876 3260
rect 16384 2922 16430 2990
rect 16500 2922 16552 2990
rect 16384 2909 16552 2922
rect 19430 3099 19602 3146
rect 24147 3126 24163 3160
rect 24197 3126 24213 3160
rect 24265 3126 24281 3160
rect 24315 3126 24331 3160
rect 24627 3131 24876 3170
rect 37724 3245 37810 3268
rect 37724 3196 37737 3245
rect 37797 3196 37810 3245
rect 37724 3165 37810 3196
rect 19430 2936 19469 3099
rect 19559 2936 19602 3099
rect 19430 2896 19602 2936
rect 26052 3100 26224 3147
rect 26052 2937 26091 3100
rect 26181 2937 26224 3100
rect 36873 3072 36963 3106
rect 37139 3072 37155 3106
rect 32316 2991 32586 3026
rect 26052 2897 26224 2937
rect 31962 2938 31996 2954
rect 31478 2792 31748 2827
rect 31478 2738 31512 2792
rect 15770 2503 31116 2655
rect 31478 2546 31512 2562
rect 31596 2738 31630 2754
rect 31596 2546 31630 2562
rect 31714 2738 31748 2792
rect 31714 2546 31748 2562
rect 31832 2738 31866 2754
rect 31832 2546 31866 2562
rect 31962 2546 31996 2562
rect 32080 2938 32114 2954
rect 32080 2546 32114 2562
rect 32198 2938 32232 2954
rect 32198 2546 32232 2562
rect 32316 2938 32350 2991
rect 32316 2546 32350 2562
rect 32434 2938 32468 2954
rect 32434 2546 32468 2562
rect 32552 2938 32586 2991
rect 33560 2975 33728 2991
rect 32552 2546 32586 2562
rect 32670 2938 32704 2954
rect 33560 2905 33576 2975
rect 33712 2905 33728 2975
rect 33560 2889 33728 2905
rect 36873 2870 36912 3072
rect 37437 3001 37522 3017
rect 36947 2954 36963 2988
rect 37139 2954 37229 2988
rect 36873 2836 36963 2870
rect 37139 2836 37155 2870
rect 34097 2785 34367 2819
rect 32670 2546 32704 2562
rect 32799 2738 32833 2754
rect 32799 2546 32833 2562
rect 32917 2738 32951 2754
rect 32917 2546 32951 2562
rect 33035 2738 33069 2754
rect 33035 2546 33069 2562
rect 33153 2738 33187 2754
rect 33153 2546 33187 2562
rect 33271 2735 33305 2751
rect 33271 2543 33305 2559
rect 33389 2735 33423 2751
rect 33389 2543 33423 2559
rect 33507 2735 33541 2751
rect 33507 2543 33541 2559
rect 33625 2735 33659 2751
rect 33625 2543 33659 2559
rect 33743 2735 33777 2751
rect 33743 2543 33777 2559
rect 33861 2735 33895 2751
rect 33861 2543 33895 2559
rect 33979 2735 34013 2751
rect 33979 2543 34013 2559
rect 34097 2735 34131 2785
rect 34097 2543 34131 2559
rect 34215 2735 34249 2751
rect 34215 2543 34249 2559
rect 34333 2735 34367 2785
rect 37190 2752 37229 2954
rect 37437 2941 37454 3001
rect 37509 2941 37522 3001
rect 37437 2925 37522 2941
rect 36947 2718 36963 2752
rect 37139 2718 37229 2752
rect 34333 2543 34367 2559
rect 36671 2631 36763 2665
rect 37139 2631 37155 2665
rect 31024 2406 31116 2503
rect 34022 2465 34038 2499
rect 34072 2465 34088 2499
rect 36671 2429 36710 2631
rect 36747 2513 36763 2547
rect 37139 2513 37229 2547
rect 31024 2400 31544 2406
rect 8360 2368 8528 2384
rect 8360 2312 8376 2368
rect 8510 2312 8528 2368
rect 8360 2294 8528 2312
rect 14914 2373 15082 2389
rect 14914 2317 14930 2373
rect 15064 2317 15082 2373
rect 14914 2299 15082 2317
rect 21563 2361 21731 2377
rect 21563 2305 21579 2361
rect 21713 2305 21731 2361
rect 31024 2330 31458 2400
rect 31025 2329 31458 2330
rect 31531 2329 31544 2400
rect 33130 2380 33164 2396
rect 36671 2395 36763 2429
rect 37139 2395 37155 2429
rect 33904 2348 33920 2382
rect 33954 2348 33970 2382
rect 33130 2330 33164 2346
rect 31025 2322 31544 2329
rect 21563 2287 21731 2305
rect 33508 2298 33542 2314
rect 31724 2261 31780 2278
rect 8127 2207 8143 2241
rect 8177 2207 8193 2241
rect 8245 2207 8261 2241
rect 8295 2207 8311 2241
rect 14681 2212 14697 2246
rect 14731 2212 14747 2246
rect 14799 2212 14815 2246
rect 14849 2212 14865 2246
rect 21330 2200 21346 2234
rect 21380 2200 21396 2234
rect 21448 2200 21464 2234
rect 21498 2200 21514 2234
rect 31724 2227 31730 2261
rect 31764 2227 31780 2261
rect 31724 2210 31780 2227
rect 31905 2245 31939 2261
rect 8084 2157 8118 2173
rect 8084 1765 8118 1781
rect 8202 2157 8236 2173
rect 8202 1765 8236 1781
rect 8320 2157 8354 2173
rect 14638 2162 14672 2178
rect 8320 1765 8354 1781
rect 8437 1957 8471 1973
rect 8437 1765 8471 1781
rect 8555 1957 8589 1973
rect 8555 1765 8589 1781
rect 14638 1770 14672 1786
rect 14756 2162 14790 2178
rect 14756 1770 14790 1786
rect 14874 2162 14908 2178
rect 21287 2150 21321 2166
rect 14874 1770 14908 1786
rect 14991 1962 15025 1978
rect 14991 1770 15025 1786
rect 15109 1962 15143 1978
rect 15109 1770 15143 1786
rect 21287 1758 21321 1774
rect 21405 2150 21439 2166
rect 21405 1758 21439 1774
rect 21523 2150 21557 2166
rect 21523 1758 21557 1774
rect 21640 1950 21674 1966
rect 21640 1758 21674 1774
rect 21758 1950 21792 1966
rect 30027 1878 30195 1894
rect 30027 1808 30043 1878
rect 30179 1808 30195 1878
rect 32023 2245 32057 2261
rect 31905 1853 31939 1869
rect 32022 1869 32023 1916
rect 32141 2245 32175 2261
rect 32057 1869 32058 1916
rect 30027 1792 30195 1808
rect 32022 1811 32058 1869
rect 32259 2245 32293 2261
rect 32141 1853 32175 1869
rect 32257 1869 32259 1916
rect 32257 1811 32293 1869
rect 32377 2245 32411 2261
rect 32377 1853 32411 1869
rect 32495 2245 32529 2261
rect 32613 2245 32647 2261
rect 32529 1869 32531 1915
rect 32495 1811 32531 1869
rect 32775 2040 32845 2044
rect 32775 1949 32779 2040
rect 32841 1949 32845 2040
rect 32775 1944 32845 1949
rect 32613 1853 32647 1869
rect 32790 1811 32831 1944
rect 33508 1906 33542 1922
rect 33626 2298 33660 2314
rect 33626 1906 33660 1922
rect 33744 2298 33778 2314
rect 33861 2298 33895 2314
rect 33861 2106 33895 2122
rect 33979 2298 34013 2314
rect 37190 2311 37229 2513
rect 36747 2277 36763 2311
rect 37139 2277 37229 2311
rect 33979 2106 34013 2122
rect 36672 2164 36763 2198
rect 37139 2164 37155 2198
rect 36672 1962 36711 2164
rect 37190 2080 37229 2277
rect 38080 2238 38096 2272
rect 38272 2238 38288 2272
rect 38080 2120 38096 2154
rect 38272 2120 38288 2154
rect 38084 2080 38284 2120
rect 36747 2046 36763 2080
rect 37139 2046 37229 2080
rect 33744 1906 33778 1922
rect 36475 1920 36585 1936
rect 36672 1928 36763 1962
rect 37139 1928 37155 1962
rect 33551 1838 33567 1872
rect 33601 1838 33617 1872
rect 33669 1838 33685 1872
rect 33719 1838 33735 1872
rect 21758 1758 21792 1774
rect 32022 1771 32831 1811
rect 32041 1770 32831 1771
rect 8480 1697 8496 1731
rect 8530 1697 8546 1731
rect 15034 1702 15050 1736
rect 15084 1702 15100 1736
rect 21683 1690 21699 1724
rect 21733 1690 21749 1724
rect 30564 1688 30834 1722
rect 29738 1638 29772 1654
rect 8598 1580 8614 1614
rect 8648 1580 8664 1614
rect 15152 1585 15168 1619
rect 15202 1585 15218 1619
rect 21801 1573 21817 1607
rect 21851 1573 21867 1607
rect 7847 1520 7881 1536
rect 7847 1328 7881 1344
rect 7965 1520 7999 1536
rect 7965 1328 7999 1344
rect 8083 1520 8117 1536
rect 8083 1328 8117 1344
rect 8201 1520 8235 1536
rect 8201 1328 8235 1344
rect 8319 1520 8353 1536
rect 8319 1328 8353 1344
rect 8437 1520 8471 1536
rect 8437 1328 8471 1344
rect 8555 1520 8589 1536
rect 8555 1328 8589 1344
rect 8673 1520 8707 1536
rect 8673 1294 8707 1344
rect 8791 1520 8825 1536
rect 8791 1328 8825 1344
rect 8909 1520 8943 1536
rect 8909 1294 8943 1344
rect 14401 1525 14435 1541
rect 14401 1333 14435 1349
rect 14519 1525 14553 1541
rect 14519 1333 14553 1349
rect 14637 1525 14671 1541
rect 14637 1333 14671 1349
rect 14755 1525 14789 1541
rect 14755 1333 14789 1349
rect 14873 1525 14907 1541
rect 14873 1333 14907 1349
rect 14991 1525 15025 1541
rect 14991 1333 15025 1349
rect 15109 1525 15143 1541
rect 15109 1333 15143 1349
rect 15227 1525 15261 1541
rect 8673 1260 8943 1294
rect 15227 1299 15261 1349
rect 15345 1525 15379 1541
rect 15345 1333 15379 1349
rect 15463 1525 15497 1541
rect 15463 1299 15497 1349
rect 21050 1513 21084 1529
rect 21050 1321 21084 1337
rect 21168 1513 21202 1529
rect 21168 1321 21202 1337
rect 21286 1513 21320 1529
rect 21286 1321 21320 1337
rect 21404 1513 21438 1529
rect 21404 1321 21438 1337
rect 21522 1513 21556 1529
rect 21522 1321 21556 1337
rect 21640 1513 21674 1529
rect 21640 1321 21674 1337
rect 21758 1513 21792 1529
rect 21758 1321 21792 1337
rect 21876 1513 21910 1529
rect 15227 1265 15497 1299
rect 21876 1287 21910 1337
rect 21994 1513 22028 1529
rect 21994 1321 22028 1337
rect 22112 1513 22146 1529
rect 29738 1446 29772 1462
rect 29856 1638 29890 1654
rect 29856 1446 29890 1462
rect 29974 1638 30008 1654
rect 29974 1446 30008 1462
rect 30092 1638 30126 1654
rect 30092 1446 30126 1462
rect 30210 1638 30244 1654
rect 30210 1446 30244 1462
rect 30328 1638 30362 1654
rect 30328 1446 30362 1462
rect 30446 1638 30480 1654
rect 30446 1446 30480 1462
rect 30564 1638 30598 1688
rect 30564 1446 30598 1462
rect 30682 1638 30716 1654
rect 30682 1446 30716 1462
rect 30800 1638 30834 1688
rect 31919 1681 31986 1697
rect 31919 1647 31935 1681
rect 31969 1647 31986 1681
rect 31919 1631 31986 1647
rect 31750 1614 31784 1630
rect 31750 1564 31784 1580
rect 32096 1529 32130 1770
rect 33784 1767 33952 1785
rect 33784 1711 33800 1767
rect 33934 1711 33952 1767
rect 32566 1681 32633 1697
rect 33784 1695 33952 1711
rect 36475 1724 36493 1920
rect 36569 1724 36585 1920
rect 37190 1844 37229 2046
rect 37725 2034 37810 2050
rect 38080 2046 38096 2080
rect 38472 2046 38488 2080
rect 37338 1986 37354 2020
rect 37388 1986 37404 2020
rect 37725 1974 37738 2034
rect 37793 1974 37810 2034
rect 37725 1958 37810 1974
rect 36747 1810 36763 1844
rect 37139 1810 37229 1844
rect 37440 1916 37525 1932
rect 38080 1928 38096 1962
rect 38472 1928 38488 1962
rect 37440 1856 37453 1916
rect 37508 1856 37525 1916
rect 38721 1862 38807 1878
rect 37440 1840 37525 1856
rect 38080 1810 38096 1844
rect 38472 1810 38488 1844
rect 38573 1843 38607 1859
rect 36475 1708 36585 1724
rect 32566 1647 32583 1681
rect 32617 1647 32633 1681
rect 32566 1631 32633 1647
rect 36672 1692 36763 1726
rect 37139 1692 37155 1726
rect 32873 1613 32907 1629
rect 32185 1563 32201 1597
rect 32235 1563 32251 1597
rect 32303 1564 32319 1598
rect 32353 1564 32369 1598
rect 32873 1563 32907 1579
rect 30800 1446 30834 1462
rect 31603 1513 31637 1529
rect 30489 1368 30505 1402
rect 30539 1368 30555 1402
rect 22112 1287 22146 1337
rect 31603 1321 31637 1337
rect 31721 1513 31755 1529
rect 31721 1321 31755 1337
rect 32023 1513 32057 1529
rect 21876 1253 22146 1287
rect 30371 1251 30387 1285
rect 30421 1251 30437 1285
rect 29975 1201 30009 1217
rect 8136 1174 8304 1190
rect 8136 1104 8152 1174
rect 8288 1104 8304 1174
rect 8136 1088 8304 1104
rect 14690 1179 14858 1195
rect 14690 1109 14706 1179
rect 14842 1109 14858 1179
rect 14690 1093 14858 1109
rect 21339 1167 21507 1183
rect 21339 1097 21355 1167
rect 21491 1097 21507 1167
rect 21339 1081 21507 1097
rect 29975 809 30009 825
rect 30093 1201 30127 1217
rect 30093 809 30127 825
rect 30211 1201 30245 1217
rect 30328 1201 30362 1217
rect 30328 1009 30362 1025
rect 30446 1201 30480 1217
rect 32096 1513 32175 1529
rect 32096 1483 32141 1513
rect 32023 1070 32058 1137
rect 32141 1121 32175 1137
rect 32259 1513 32293 1529
rect 32259 1121 32293 1137
rect 32377 1513 32411 1529
rect 32495 1513 32529 1529
rect 32901 1513 32935 1529
rect 32901 1321 32935 1337
rect 33019 1513 33053 1529
rect 36672 1490 36711 1692
rect 37190 1608 37229 1810
rect 38573 1793 38607 1809
rect 38721 1840 38739 1862
rect 37958 1751 37974 1785
rect 38008 1751 38024 1785
rect 38721 1782 38725 1840
rect 38721 1758 38739 1782
rect 38785 1758 38807 1862
rect 38721 1742 38807 1758
rect 38080 1692 38096 1726
rect 38472 1692 38488 1726
rect 37568 1632 37584 1666
rect 37618 1632 37634 1666
rect 36747 1574 36763 1608
rect 37139 1574 37229 1608
rect 38080 1574 38096 1608
rect 38472 1574 38488 1608
rect 36672 1456 36763 1490
rect 37139 1456 37155 1490
rect 37190 1371 37229 1574
rect 38084 1530 38284 1574
rect 38080 1496 38096 1530
rect 38272 1496 38288 1530
rect 38080 1378 38096 1412
rect 38272 1378 38288 1412
rect 36747 1337 36763 1371
rect 37139 1337 37229 1371
rect 33019 1321 33053 1337
rect 32377 1121 32411 1137
rect 32494 1070 32529 1137
rect 32023 1035 32529 1070
rect 36672 1219 36763 1253
rect 37139 1219 37155 1253
rect 30446 1009 30480 1025
rect 36672 1017 36711 1219
rect 37190 1135 37229 1337
rect 36747 1101 36763 1135
rect 37139 1101 37229 1135
rect 36672 983 36763 1017
rect 37139 983 37155 1017
rect 32170 966 32412 978
rect 32170 864 32217 966
rect 32352 864 32412 966
rect 36947 864 36963 898
rect 37139 864 37232 898
rect 32170 847 32412 864
rect 30211 809 30245 825
rect 30018 741 30034 775
rect 30068 741 30084 775
rect 30136 741 30152 775
rect 30186 741 30202 775
rect 36876 746 36963 780
rect 37139 746 37155 780
rect 30251 670 30419 688
rect 30251 614 30267 670
rect 30401 614 30419 670
rect 30251 598 30419 614
rect 36876 544 36913 746
rect 37193 662 37232 864
rect 36947 628 36963 662
rect 37139 628 37232 662
rect 37313 710 37347 726
rect 37313 660 37347 676
rect 36876 510 36963 544
rect 37139 510 37155 544
rect -2387 319 -2371 353
rect -2195 319 -2179 353
rect -1230 278 15 361
rect 122 278 136 361
rect -1230 265 136 278
rect 2723 355 2914 370
rect 2723 289 2748 355
rect 2892 289 2914 355
rect 2723 268 2914 289
rect -2387 201 -2371 235
rect -2195 201 -2179 235
rect -3612 67 -3596 101
rect -3420 67 -3404 101
<< viali >>
rect 8052 27822 8086 27856
rect 9182 27828 9216 27862
rect 14565 27819 14599 27853
rect 15695 27825 15729 27859
rect 21099 27814 21133 27848
rect 22229 27820 22263 27854
rect 27657 27818 27691 27852
rect 28787 27824 28821 27858
rect 8052 27704 8086 27738
rect 9182 27708 9216 27742
rect 5842 27432 5876 27608
rect 5960 27432 5994 27608
rect 6078 27432 6112 27608
rect 6196 27432 6230 27608
rect 6314 27432 6348 27608
rect 6432 27432 6466 27608
rect 6550 27432 6584 27608
rect 6668 27432 6702 27608
rect 6786 27432 6820 27608
rect 6904 27432 6938 27608
rect 6609 27338 6643 27372
rect 8167 27304 8201 27680
rect 8285 27304 8319 27680
rect 8403 27304 8437 27680
rect 8521 27304 8555 27680
rect 8639 27304 8673 27680
rect 8757 27304 8791 27680
rect 14565 27701 14599 27735
rect 8875 27304 8909 27680
rect 9309 27308 9343 27684
rect 9427 27308 9461 27684
rect 9545 27308 9579 27684
rect 9663 27308 9697 27684
rect 9781 27308 9815 27684
rect 9899 27308 9933 27684
rect 10017 27308 10051 27684
rect 15695 27705 15729 27739
rect 12355 27429 12389 27605
rect 12473 27429 12507 27605
rect 12591 27429 12625 27605
rect 12709 27429 12743 27605
rect 12827 27429 12861 27605
rect 12945 27429 12979 27605
rect 13063 27429 13097 27605
rect 13181 27429 13215 27605
rect 13299 27429 13333 27605
rect 13417 27429 13451 27605
rect 13122 27335 13156 27369
rect 14680 27301 14714 27677
rect 14798 27301 14832 27677
rect 14916 27301 14950 27677
rect 15034 27301 15068 27677
rect 15152 27301 15186 27677
rect 15270 27301 15304 27677
rect 15388 27301 15422 27677
rect 15822 27305 15856 27681
rect 15940 27305 15974 27681
rect 16058 27305 16092 27681
rect 16176 27305 16210 27681
rect 16294 27305 16328 27681
rect 16412 27305 16446 27681
rect 21099 27696 21133 27730
rect 16530 27305 16564 27681
rect 22229 27700 22263 27734
rect 18889 27424 18923 27600
rect 19007 27424 19041 27600
rect 19125 27424 19159 27600
rect 19243 27424 19277 27600
rect 19361 27424 19395 27600
rect 19479 27424 19513 27600
rect 19597 27424 19631 27600
rect 19715 27424 19749 27600
rect 19833 27424 19867 27600
rect 19951 27424 19985 27600
rect 19656 27330 19690 27364
rect 21214 27296 21248 27672
rect 21332 27296 21366 27672
rect 21450 27296 21484 27672
rect 21568 27296 21602 27672
rect 21686 27296 21720 27672
rect 21804 27296 21838 27672
rect 27657 27700 27691 27734
rect 21922 27296 21956 27672
rect 22356 27300 22390 27676
rect 22474 27300 22508 27676
rect 22592 27300 22626 27676
rect 22710 27300 22744 27676
rect 22828 27300 22862 27676
rect 22946 27300 22980 27676
rect 23064 27300 23098 27676
rect 28787 27704 28821 27738
rect 25447 27428 25481 27604
rect 25565 27428 25599 27604
rect 25683 27428 25717 27604
rect 25801 27428 25835 27604
rect 25919 27428 25953 27604
rect 26037 27428 26071 27604
rect 26155 27428 26189 27604
rect 26273 27428 26307 27604
rect 26391 27428 26425 27604
rect 26509 27428 26543 27604
rect 26214 27334 26248 27368
rect 27772 27300 27806 27676
rect 27890 27300 27924 27676
rect 28008 27300 28042 27676
rect 28126 27300 28160 27676
rect 28244 27300 28278 27676
rect 28362 27300 28396 27676
rect 28480 27300 28514 27676
rect 28914 27304 28948 27680
rect 29032 27304 29066 27680
rect 29150 27304 29184 27680
rect 29268 27304 29302 27680
rect 29386 27304 29420 27680
rect 29504 27304 29538 27680
rect 29622 27304 29656 27680
rect 6491 27221 6525 27255
rect 13004 27218 13038 27252
rect 19538 27213 19572 27247
rect 26096 27217 26130 27251
rect 6079 26795 6113 27171
rect 6197 26795 6231 27171
rect 6315 26795 6349 27171
rect 6432 26995 6466 27171
rect 6550 26995 6584 27171
rect 8372 26948 8406 26982
rect 9514 26952 9548 26986
rect 6138 26711 6172 26745
rect 6256 26711 6290 26745
rect 8077 26721 8111 26897
rect 8195 26721 8229 26897
rect 8313 26721 8347 26897
rect 8431 26721 8465 26897
rect 8596 26721 8630 26897
rect 8714 26721 8748 26897
rect 8832 26721 8866 26897
rect 8950 26721 8984 26897
rect 9219 26725 9253 26901
rect 9337 26725 9371 26901
rect 9455 26725 9489 26901
rect 9573 26725 9607 26901
rect 9738 26725 9772 26901
rect 9856 26725 9890 26901
rect 9974 26725 10008 26901
rect 10092 26725 10126 26901
rect 12592 26792 12626 27168
rect 12710 26792 12744 27168
rect 12828 26792 12862 27168
rect 12945 26992 12979 27168
rect 13063 26992 13097 27168
rect 14885 26945 14919 26979
rect 16027 26949 16061 26983
rect 12651 26708 12685 26742
rect 12769 26708 12803 26742
rect 14590 26718 14624 26894
rect 14708 26718 14742 26894
rect 14826 26718 14860 26894
rect 14944 26718 14978 26894
rect 15109 26718 15143 26894
rect 15227 26718 15261 26894
rect 15345 26718 15379 26894
rect 15463 26718 15497 26894
rect 15732 26722 15766 26898
rect 15850 26722 15884 26898
rect 15968 26722 16002 26898
rect 16086 26722 16120 26898
rect 16251 26722 16285 26898
rect 16369 26722 16403 26898
rect 16487 26722 16521 26898
rect 16605 26722 16639 26898
rect 19126 26787 19160 27163
rect 19244 26787 19278 27163
rect 19362 26787 19396 27163
rect 19479 26987 19513 27163
rect 19597 26987 19631 27163
rect 21419 26940 21453 26974
rect 22561 26944 22595 26978
rect 19185 26703 19219 26737
rect 19303 26703 19337 26737
rect 21124 26713 21158 26889
rect 21242 26713 21276 26889
rect 21360 26713 21394 26889
rect 21478 26713 21512 26889
rect 21643 26713 21677 26889
rect 21761 26713 21795 26889
rect 21879 26713 21913 26889
rect 21997 26713 22031 26889
rect 22266 26717 22300 26893
rect 22384 26717 22418 26893
rect 22502 26717 22536 26893
rect 22620 26717 22654 26893
rect 22785 26717 22819 26893
rect 22903 26717 22937 26893
rect 23021 26717 23055 26893
rect 23139 26717 23173 26893
rect 25684 26791 25718 27167
rect 25802 26791 25836 27167
rect 25920 26791 25954 27167
rect 26037 26991 26071 27167
rect 26155 26991 26189 27167
rect 27977 26944 28011 26978
rect 29119 26948 29153 26982
rect 25743 26707 25777 26741
rect 25861 26707 25895 26741
rect 27682 26717 27716 26893
rect 27800 26717 27834 26893
rect 27918 26717 27952 26893
rect 28036 26717 28070 26893
rect 28201 26717 28235 26893
rect 28319 26717 28353 26893
rect 28437 26717 28471 26893
rect 28555 26717 28589 26893
rect 28824 26721 28858 26897
rect 28942 26721 28976 26897
rect 29060 26721 29094 26897
rect 29178 26721 29212 26897
rect 29343 26721 29377 26897
rect 29461 26721 29495 26897
rect 29579 26721 29613 26897
rect 29697 26721 29731 26897
rect 64 25890 118 25939
rect -92 25447 -23 25518
rect -239 25023 -168 25094
rect -382 24573 -311 24634
rect -3592 16221 -3416 16255
rect -3057 16232 -2997 16248
rect -3057 16198 -3043 16232
rect -3043 16198 -3009 16232
rect -3009 16198 -2997 16232
rect -3057 16182 -2997 16198
rect -3592 16103 -3416 16137
rect -2367 16096 -2191 16130
rect -3592 15985 -3416 16019
rect -2468 15949 -2434 15983
rect -2367 15978 -2191 16012
rect -3592 15867 -3416 15901
rect -3099 15794 -2723 15828
rect -3792 15737 -3416 15771
rect -2535 15764 -2501 15798
rect -3099 15676 -2723 15710
rect -2367 15676 -1991 15710
rect -3792 15619 -3416 15653
rect -3099 15558 -2723 15592
rect -3792 15501 -3416 15535
rect -2367 15558 -1991 15592
rect -2451 15498 -2417 15532
rect -3099 15440 -2723 15474
rect -2367 15440 -1991 15474
rect -4047 15380 -4019 15418
rect -4019 15380 -4009 15418
rect -3792 15383 -3416 15417
rect -3099 15322 -2723 15356
rect -3792 15265 -3416 15299
rect -2452 15380 -2418 15414
rect -2367 15322 -1991 15356
rect -1825 15430 -1803 15480
rect -1803 15430 -1783 15480
rect -3099 15204 -2723 15238
rect -2367 15204 -1991 15238
rect -3792 15147 -3416 15181
rect -3099 15086 -2723 15120
rect -3792 15029 -3416 15063
rect -3592 14900 -3416 14934
rect -3247 14838 -3193 14848
rect -3592 14782 -3416 14816
rect -3247 14804 -3237 14838
rect -3237 14804 -3203 14838
rect -3203 14804 -3193 14838
rect -3247 14794 -3193 14804
rect -3592 14664 -3416 14698
rect -2535 15116 -2501 15150
rect -2467 14826 -2433 14860
rect -2367 14798 -2191 14832
rect -2367 14680 -2191 14714
rect -3592 14546 -3416 14580
rect -2695 14514 -2593 14616
rect -3594 14153 -3418 14187
rect -3059 14164 -2999 14180
rect -3059 14130 -3045 14164
rect -3045 14130 -3011 14164
rect -3011 14130 -2999 14164
rect -3059 14114 -2999 14130
rect -3594 14035 -3418 14069
rect -2369 14028 -2193 14062
rect -3594 13917 -3418 13951
rect -2470 13881 -2436 13915
rect -2369 13910 -2193 13944
rect -3594 13799 -3418 13833
rect -3101 13726 -2725 13760
rect -3794 13669 -3418 13703
rect -2537 13696 -2503 13730
rect -3101 13608 -2725 13642
rect -2369 13608 -1993 13642
rect -3794 13551 -3418 13585
rect -3101 13490 -2725 13524
rect -3794 13433 -3418 13467
rect -2369 13490 -1993 13524
rect -2453 13430 -2419 13464
rect -3101 13372 -2725 13406
rect -2369 13372 -1993 13406
rect -4049 13312 -4021 13350
rect -4021 13312 -4011 13350
rect -3794 13315 -3418 13349
rect -3101 13254 -2725 13288
rect -3794 13197 -3418 13231
rect -2454 13312 -2420 13346
rect -2369 13254 -1993 13288
rect -1827 13362 -1805 13412
rect -1805 13362 -1785 13412
rect -3101 13136 -2725 13170
rect -2369 13136 -1993 13170
rect -3794 13079 -3418 13113
rect -3101 13018 -2725 13052
rect -3794 12961 -3418 12995
rect -3594 12832 -3418 12866
rect -3249 12770 -3195 12780
rect -3594 12714 -3418 12748
rect -3249 12736 -3239 12770
rect -3239 12736 -3205 12770
rect -3205 12736 -3195 12770
rect -3249 12726 -3195 12736
rect -3594 12596 -3418 12630
rect -2537 13048 -2503 13082
rect -2469 12758 -2435 12792
rect -2369 12730 -2193 12764
rect -2369 12612 -2193 12646
rect -3594 12478 -3418 12512
rect -2697 12446 -2595 12548
rect -3592 12084 -3416 12118
rect -3057 12095 -2997 12111
rect -3057 12061 -3043 12095
rect -3043 12061 -3009 12095
rect -3009 12061 -2997 12095
rect -3057 12045 -2997 12061
rect -3592 11966 -3416 12000
rect -2367 11959 -2191 11993
rect -3592 11848 -3416 11882
rect -2468 11812 -2434 11846
rect -2367 11841 -2191 11875
rect -3592 11730 -3416 11764
rect -3099 11657 -2723 11691
rect -3792 11600 -3416 11634
rect -2535 11627 -2501 11661
rect -3099 11539 -2723 11573
rect -2367 11539 -1991 11573
rect -3792 11482 -3416 11516
rect -3099 11421 -2723 11455
rect -3792 11364 -3416 11398
rect -2367 11421 -1991 11455
rect -2451 11361 -2417 11395
rect -3099 11303 -2723 11337
rect -2367 11303 -1991 11337
rect -4047 11243 -4019 11281
rect -4019 11243 -4009 11281
rect -3792 11246 -3416 11280
rect -3099 11185 -2723 11219
rect -3792 11128 -3416 11162
rect -2452 11243 -2418 11277
rect -2367 11185 -1991 11219
rect -1825 11293 -1803 11343
rect -1803 11293 -1783 11343
rect -3099 11067 -2723 11101
rect -2367 11067 -1991 11101
rect -3792 11010 -3416 11044
rect -3099 10949 -2723 10983
rect -3792 10892 -3416 10926
rect -3592 10763 -3416 10797
rect -3247 10701 -3193 10711
rect -3592 10645 -3416 10679
rect -3247 10667 -3237 10701
rect -3237 10667 -3203 10701
rect -3203 10667 -3193 10701
rect -3247 10657 -3193 10667
rect -3592 10527 -3416 10561
rect -2535 10979 -2501 11013
rect -2467 10689 -2433 10723
rect -2367 10661 -2191 10695
rect -2367 10543 -2191 10577
rect -3592 10409 -3416 10443
rect -2695 10377 -2593 10479
rect -3594 10016 -3418 10050
rect -3059 10027 -2999 10043
rect -3059 9993 -3045 10027
rect -3045 9993 -3011 10027
rect -3011 9993 -2999 10027
rect -3059 9977 -2999 9993
rect -3594 9898 -3418 9932
rect -2369 9891 -2193 9925
rect -3594 9780 -3418 9814
rect -2470 9744 -2436 9778
rect -2369 9773 -2193 9807
rect -3594 9662 -3418 9696
rect -3101 9589 -2725 9623
rect -3794 9532 -3418 9566
rect -2537 9559 -2503 9593
rect -3101 9471 -2725 9505
rect -2369 9471 -1993 9505
rect -3794 9414 -3418 9448
rect -3101 9353 -2725 9387
rect -3794 9296 -3418 9330
rect -2369 9353 -1993 9387
rect -2453 9293 -2419 9327
rect -3101 9235 -2725 9269
rect -2369 9235 -1993 9269
rect -4049 9175 -4021 9213
rect -4021 9175 -4011 9213
rect -3794 9178 -3418 9212
rect -3101 9117 -2725 9151
rect -3794 9060 -3418 9094
rect -2454 9175 -2420 9209
rect -2369 9117 -1993 9151
rect -1827 9225 -1805 9275
rect -1805 9225 -1785 9275
rect -3101 8999 -2725 9033
rect -2369 8999 -1993 9033
rect -3794 8942 -3418 8976
rect -3101 8881 -2725 8915
rect -3794 8824 -3418 8858
rect -3594 8695 -3418 8729
rect -3249 8633 -3195 8643
rect -3594 8577 -3418 8611
rect -3249 8599 -3239 8633
rect -3239 8599 -3205 8633
rect -3205 8599 -3195 8633
rect -3249 8589 -3195 8599
rect -3594 8459 -3418 8493
rect -2537 8911 -2503 8945
rect -2469 8621 -2435 8655
rect -2369 8593 -2193 8627
rect -2369 8475 -2193 8509
rect -3594 8341 -3418 8375
rect -2697 8309 -2595 8411
rect -3594 7947 -3418 7981
rect -3059 7958 -2999 7974
rect -3059 7924 -3045 7958
rect -3045 7924 -3011 7958
rect -3011 7924 -2999 7958
rect -3059 7908 -2999 7924
rect -3594 7829 -3418 7863
rect -2369 7822 -2193 7856
rect -3594 7711 -3418 7745
rect -2470 7675 -2436 7709
rect -2369 7704 -2193 7738
rect -3594 7593 -3418 7627
rect -3101 7520 -2725 7554
rect -3794 7463 -3418 7497
rect -2537 7490 -2503 7524
rect -3101 7402 -2725 7436
rect -2369 7402 -1993 7436
rect -3794 7345 -3418 7379
rect -3101 7284 -2725 7318
rect -3794 7227 -3418 7261
rect -2369 7284 -1993 7318
rect -2453 7224 -2419 7258
rect -3101 7166 -2725 7200
rect -2369 7166 -1993 7200
rect -4049 7106 -4021 7144
rect -4021 7106 -4011 7144
rect -3794 7109 -3418 7143
rect -3101 7048 -2725 7082
rect -3794 6991 -3418 7025
rect -2454 7106 -2420 7140
rect -2369 7048 -1993 7082
rect -1827 7156 -1805 7206
rect -1805 7156 -1785 7206
rect -3101 6930 -2725 6964
rect -2369 6930 -1993 6964
rect -3794 6873 -3418 6907
rect -3101 6812 -2725 6846
rect -3794 6755 -3418 6789
rect -3594 6626 -3418 6660
rect -3249 6564 -3195 6574
rect -3594 6508 -3418 6542
rect -3249 6530 -3239 6564
rect -3239 6530 -3205 6564
rect -3205 6530 -3195 6564
rect -3249 6520 -3195 6530
rect -3594 6390 -3418 6424
rect -2537 6842 -2503 6876
rect -2469 6552 -2435 6586
rect -2369 6524 -2193 6558
rect -2369 6406 -2193 6440
rect -3594 6272 -3418 6306
rect -2697 6240 -2595 6342
rect -1077 6025 -1011 6087
rect -3596 5879 -3420 5913
rect -3061 5890 -3001 5906
rect -3061 5856 -3047 5890
rect -3047 5856 -3013 5890
rect -3013 5856 -3001 5890
rect -3061 5840 -3001 5856
rect -3596 5761 -3420 5795
rect -2371 5754 -2195 5788
rect -3596 5643 -3420 5677
rect -2472 5607 -2438 5641
rect -2371 5636 -2195 5670
rect -3596 5525 -3420 5559
rect -3103 5452 -2727 5486
rect -3796 5395 -3420 5429
rect -2539 5422 -2505 5456
rect -3103 5334 -2727 5368
rect -2371 5334 -1995 5368
rect -3796 5277 -3420 5311
rect -3103 5216 -2727 5250
rect -3796 5159 -3420 5193
rect -2371 5216 -1995 5250
rect -2455 5156 -2421 5190
rect -3103 5098 -2727 5132
rect -2371 5098 -1995 5132
rect -4051 5038 -4023 5076
rect -4023 5038 -4013 5076
rect -3796 5041 -3420 5075
rect -3103 4980 -2727 5014
rect -3796 4923 -3420 4957
rect -2456 5038 -2422 5072
rect -2371 4980 -1995 5014
rect -1829 5088 -1807 5138
rect -1807 5088 -1787 5138
rect -3103 4862 -2727 4896
rect -2371 4862 -1995 4896
rect -3796 4805 -3420 4839
rect -3103 4744 -2727 4778
rect -3796 4687 -3420 4721
rect -3596 4558 -3420 4592
rect -3251 4496 -3197 4506
rect -3596 4440 -3420 4474
rect -3251 4462 -3241 4496
rect -3241 4462 -3207 4496
rect -3207 4462 -3197 4496
rect -3251 4452 -3197 4462
rect -3596 4322 -3420 4356
rect -2539 4774 -2505 4808
rect -2471 4484 -2437 4518
rect -2371 4456 -2195 4490
rect -2371 4338 -2195 4372
rect -3596 4204 -3420 4238
rect -2699 4172 -2597 4274
rect -1224 3953 -1154 4008
rect -3594 3810 -3418 3844
rect -3059 3821 -2999 3837
rect -3059 3787 -3045 3821
rect -3045 3787 -3011 3821
rect -3011 3787 -2999 3821
rect -3059 3771 -2999 3787
rect -3594 3692 -3418 3726
rect -2369 3685 -2193 3719
rect -3594 3574 -3418 3608
rect -2470 3538 -2436 3572
rect -2369 3567 -2193 3601
rect -3594 3456 -3418 3490
rect -3101 3383 -2725 3417
rect -3794 3326 -3418 3360
rect -2537 3353 -2503 3387
rect -3101 3265 -2725 3299
rect -2369 3265 -1993 3299
rect -3794 3208 -3418 3242
rect -3101 3147 -2725 3181
rect -3794 3090 -3418 3124
rect -2369 3147 -1993 3181
rect -2453 3087 -2419 3121
rect -3101 3029 -2725 3063
rect -2369 3029 -1993 3063
rect -4049 2969 -4021 3007
rect -4021 2969 -4011 3007
rect -3794 2972 -3418 3006
rect -3101 2911 -2725 2945
rect -3794 2854 -3418 2888
rect -2454 2969 -2420 3003
rect -2369 2911 -1993 2945
rect -1827 3019 -1805 3069
rect -1805 3019 -1785 3069
rect -3101 2793 -2725 2827
rect -2369 2793 -1993 2827
rect -3794 2736 -3418 2770
rect -3101 2675 -2725 2709
rect -3794 2618 -3418 2652
rect -3594 2489 -3418 2523
rect -3249 2427 -3195 2437
rect -3594 2371 -3418 2405
rect -3249 2393 -3239 2427
rect -3239 2393 -3205 2427
rect -3205 2393 -3195 2427
rect -3249 2383 -3195 2393
rect -3594 2253 -3418 2287
rect -2537 2705 -2503 2739
rect -2469 2415 -2435 2449
rect -2369 2387 -2193 2421
rect -2369 2269 -2193 2303
rect -3594 2135 -3418 2169
rect -2697 2103 -2595 2205
rect -3596 1742 -3420 1776
rect -3061 1753 -3001 1769
rect -3061 1719 -3047 1753
rect -3047 1719 -3013 1753
rect -3013 1719 -3001 1753
rect -3061 1703 -3001 1719
rect -3596 1624 -3420 1658
rect -2371 1617 -2195 1651
rect -3596 1506 -3420 1540
rect -2472 1470 -2438 1504
rect -2371 1499 -2195 1533
rect -3596 1388 -3420 1422
rect -3103 1315 -2727 1349
rect -3796 1258 -3420 1292
rect -2539 1285 -2505 1319
rect -3103 1197 -2727 1231
rect -2371 1197 -1995 1231
rect -3796 1140 -3420 1174
rect -3103 1079 -2727 1113
rect -3796 1022 -3420 1056
rect -2371 1079 -1995 1113
rect -2455 1019 -2421 1053
rect -3103 961 -2727 995
rect -2371 961 -1995 995
rect -4051 901 -4023 939
rect -4023 901 -4013 939
rect -3796 904 -3420 938
rect -3103 843 -2727 877
rect -3796 786 -3420 820
rect -2456 901 -2422 935
rect -2371 843 -1995 877
rect -1829 951 -1807 1001
rect -1807 951 -1787 1001
rect -3103 725 -2727 759
rect -2371 725 -1995 759
rect -3796 668 -3420 702
rect -3103 607 -2727 641
rect -3796 550 -3420 584
rect -3596 421 -3420 455
rect -3251 359 -3197 369
rect -3596 303 -3420 337
rect -3251 325 -3241 359
rect -3241 325 -3207 359
rect -3207 325 -3197 359
rect -3251 315 -3197 325
rect -3596 185 -3420 219
rect -2539 637 -2505 671
rect -2471 347 -2437 381
rect 5856 25782 5890 25958
rect 5974 25782 6008 25958
rect 6092 25782 6126 25958
rect 6210 25782 6244 25958
rect 6328 25782 6362 25958
rect 6446 25782 6480 25958
rect 6564 25782 6598 25958
rect 6682 25782 6716 25958
rect 6800 25782 6834 25958
rect 6918 25782 6952 25958
rect 12369 25779 12403 25955
rect 12487 25779 12521 25955
rect 12605 25779 12639 25955
rect 12723 25779 12757 25955
rect 12841 25779 12875 25955
rect 12959 25779 12993 25955
rect 13077 25779 13111 25955
rect 13195 25779 13229 25955
rect 13313 25779 13347 25955
rect 13431 25779 13465 25955
rect 18903 25774 18937 25950
rect 19021 25774 19055 25950
rect 19139 25774 19173 25950
rect 19257 25774 19291 25950
rect 19375 25774 19409 25950
rect 19493 25774 19527 25950
rect 19611 25774 19645 25950
rect 19729 25774 19763 25950
rect 19847 25774 19881 25950
rect 19965 25774 19999 25950
rect 25461 25778 25495 25954
rect 25579 25778 25613 25954
rect 25697 25778 25731 25954
rect 25815 25778 25849 25954
rect 25933 25778 25967 25954
rect 26051 25778 26085 25954
rect 26169 25778 26203 25954
rect 26287 25778 26321 25954
rect 26405 25778 26439 25954
rect 26523 25778 26557 25954
rect 6623 25688 6657 25722
rect 13136 25685 13170 25719
rect 19670 25680 19704 25714
rect 26228 25684 26262 25718
rect 6505 25571 6539 25605
rect 6093 25145 6127 25521
rect 6211 25145 6245 25521
rect 6329 25145 6363 25521
rect 6446 25345 6480 25521
rect 6564 25345 6598 25521
rect 7320 25165 7354 25341
rect 7438 25165 7472 25341
rect 7556 25165 7590 25341
rect 7674 25165 7708 25341
rect 7804 25165 7838 25541
rect 7922 25165 7956 25541
rect 8040 25165 8074 25541
rect 8158 25165 8192 25541
rect 8276 25165 8310 25541
rect 8394 25165 8428 25541
rect 8512 25165 8546 25541
rect 8641 25165 8675 25341
rect 8759 25165 8793 25341
rect 8877 25165 8911 25341
rect 8995 25165 9029 25341
rect 9218 25165 9252 25341
rect 9336 25165 9370 25341
rect 9454 25165 9488 25341
rect 9572 25165 9606 25341
rect 9702 25165 9736 25541
rect 9820 25165 9854 25541
rect 9938 25165 9972 25541
rect 10056 25165 10090 25541
rect 10174 25165 10208 25541
rect 13018 25568 13052 25602
rect 10292 25165 10326 25541
rect 10410 25165 10444 25541
rect 10539 25165 10573 25341
rect 10657 25165 10691 25341
rect 10775 25165 10809 25341
rect 10893 25165 10927 25341
rect 12606 25142 12640 25518
rect 12724 25142 12758 25518
rect 12842 25142 12876 25518
rect 12959 25342 12993 25518
rect 13077 25342 13111 25518
rect 6152 25061 6186 25095
rect 6270 25061 6304 25095
rect 13833 25162 13867 25338
rect 13951 25162 13985 25338
rect 14069 25162 14103 25338
rect 14187 25162 14221 25338
rect 14317 25162 14351 25538
rect 14435 25162 14469 25538
rect 14553 25162 14587 25538
rect 14671 25162 14705 25538
rect 14789 25162 14823 25538
rect 14907 25162 14941 25538
rect 15025 25162 15059 25538
rect 15154 25162 15188 25338
rect 15272 25162 15306 25338
rect 15390 25162 15424 25338
rect 15508 25162 15542 25338
rect 15731 25162 15765 25338
rect 15849 25162 15883 25338
rect 15967 25162 16001 25338
rect 16085 25162 16119 25338
rect 16215 25162 16249 25538
rect 16333 25162 16367 25538
rect 16451 25162 16485 25538
rect 16569 25162 16603 25538
rect 16687 25162 16721 25538
rect 19552 25563 19586 25597
rect 16805 25162 16839 25538
rect 16923 25162 16957 25538
rect 17052 25162 17086 25338
rect 17170 25162 17204 25338
rect 17288 25162 17322 25338
rect 17406 25162 17440 25338
rect 19140 25137 19174 25513
rect 19258 25137 19292 25513
rect 19376 25137 19410 25513
rect 19493 25337 19527 25513
rect 19611 25337 19645 25513
rect 12665 25058 12699 25092
rect 12783 25058 12817 25092
rect 20367 25157 20401 25333
rect 20485 25157 20519 25333
rect 20603 25157 20637 25333
rect 20721 25157 20755 25333
rect 20851 25157 20885 25533
rect 20969 25157 21003 25533
rect 21087 25157 21121 25533
rect 21205 25157 21239 25533
rect 21323 25157 21357 25533
rect 21441 25157 21475 25533
rect 21559 25157 21593 25533
rect 21688 25157 21722 25333
rect 21806 25157 21840 25333
rect 21924 25157 21958 25333
rect 22042 25157 22076 25333
rect 22265 25157 22299 25333
rect 22383 25157 22417 25333
rect 22501 25157 22535 25333
rect 22619 25157 22653 25333
rect 22749 25157 22783 25533
rect 22867 25157 22901 25533
rect 22985 25157 23019 25533
rect 23103 25157 23137 25533
rect 23221 25157 23255 25533
rect 26110 25567 26144 25601
rect 23339 25157 23373 25533
rect 23457 25157 23491 25533
rect 23586 25157 23620 25333
rect 23704 25157 23738 25333
rect 23822 25157 23856 25333
rect 23940 25157 23974 25333
rect 25698 25141 25732 25517
rect 25816 25141 25850 25517
rect 25934 25141 25968 25517
rect 26051 25341 26085 25517
rect 26169 25341 26203 25517
rect 19199 25053 19233 25087
rect 19317 25053 19351 25087
rect 26925 25161 26959 25337
rect 27043 25161 27077 25337
rect 27161 25161 27195 25337
rect 27279 25161 27313 25337
rect 27409 25161 27443 25537
rect 27527 25161 27561 25537
rect 27645 25161 27679 25537
rect 27763 25161 27797 25537
rect 27881 25161 27915 25537
rect 27999 25161 28033 25537
rect 28117 25161 28151 25537
rect 28246 25161 28280 25337
rect 28364 25161 28398 25337
rect 28482 25161 28516 25337
rect 28600 25161 28634 25337
rect 28823 25161 28857 25337
rect 28941 25161 28975 25337
rect 29059 25161 29093 25337
rect 29177 25161 29211 25337
rect 29307 25161 29341 25537
rect 29425 25161 29459 25537
rect 29543 25161 29577 25537
rect 29661 25161 29695 25537
rect 29779 25161 29813 25537
rect 29897 25161 29931 25537
rect 30015 25161 30049 25537
rect 30144 25161 30178 25337
rect 30262 25161 30296 25337
rect 30380 25161 30414 25337
rect 30498 25161 30532 25337
rect 34860 25322 34943 25387
rect 25757 25057 25791 25091
rect 25875 25057 25909 25091
rect 8784 24893 8818 24927
rect 10891 24872 10925 24906
rect 15297 24890 15331 24924
rect 7747 24472 7781 24848
rect 7865 24472 7899 24848
rect 5851 24178 5885 24354
rect 5969 24178 6003 24354
rect 6087 24178 6121 24354
rect 6205 24178 6239 24354
rect 6323 24178 6357 24354
rect 6441 24178 6475 24354
rect 6559 24178 6593 24354
rect 6677 24178 6711 24354
rect 6795 24178 6829 24354
rect 7983 24472 8017 24848
rect 8101 24472 8135 24848
rect 8219 24472 8253 24848
rect 8337 24472 8371 24848
rect 8455 24472 8489 24848
rect 9645 24472 9679 24848
rect 9763 24472 9797 24848
rect 9881 24472 9915 24848
rect 9999 24472 10033 24848
rect 10117 24472 10151 24848
rect 10235 24472 10269 24848
rect 17404 24869 17438 24903
rect 21831 24885 21865 24919
rect 10353 24472 10387 24848
rect 14260 24469 14294 24845
rect 14378 24469 14412 24845
rect 6913 24178 6947 24354
rect 7777 24250 7811 24284
rect 7592 24183 7626 24217
rect 8425 24250 8459 24284
rect 9675 24250 9709 24284
rect 8043 24166 8077 24200
rect 8161 24167 8195 24201
rect 8715 24182 8749 24216
rect 9490 24183 9524 24217
rect 10321 24251 10355 24285
rect 9941 24166 9975 24200
rect 10059 24167 10093 24201
rect 10613 24182 10647 24216
rect 6618 24084 6652 24118
rect 6500 23967 6534 24001
rect 7445 23940 7479 24116
rect 6088 23541 6122 23917
rect 6206 23541 6240 23917
rect 6324 23541 6358 23917
rect 6441 23741 6475 23917
rect 7563 23940 7597 24116
rect 6559 23741 6593 23917
rect 7865 23740 7899 24116
rect 7983 23740 8017 24116
rect 8101 23740 8135 24116
rect 8219 23740 8253 24116
rect 8337 23740 8371 24116
rect 8743 23940 8777 24116
rect 8861 23940 8895 24116
rect 9343 23940 9377 24116
rect 9461 23940 9495 24116
rect 9763 23740 9797 24116
rect 9881 23740 9915 24116
rect 9999 23740 10033 24116
rect 10117 23740 10151 24116
rect 10235 23740 10269 24116
rect 10641 23940 10675 24116
rect 10759 23940 10793 24116
rect 6147 23457 6181 23491
rect 6265 23457 6299 23491
rect 12364 24175 12398 24351
rect 12482 24175 12516 24351
rect 12600 24175 12634 24351
rect 12718 24175 12752 24351
rect 12836 24175 12870 24351
rect 12954 24175 12988 24351
rect 13072 24175 13106 24351
rect 13190 24175 13224 24351
rect 13308 24175 13342 24351
rect 14496 24469 14530 24845
rect 14614 24469 14648 24845
rect 14732 24469 14766 24845
rect 14850 24469 14884 24845
rect 14968 24469 15002 24845
rect 16158 24469 16192 24845
rect 16276 24469 16310 24845
rect 16394 24469 16428 24845
rect 16512 24469 16546 24845
rect 16630 24469 16664 24845
rect 16748 24469 16782 24845
rect 23938 24864 23972 24898
rect 28389 24889 28423 24923
rect 16866 24469 16900 24845
rect 20794 24464 20828 24840
rect 20912 24464 20946 24840
rect 13426 24175 13460 24351
rect 14290 24247 14324 24281
rect 14105 24180 14139 24214
rect 14938 24247 14972 24281
rect 16188 24247 16222 24281
rect 14556 24163 14590 24197
rect 14674 24164 14708 24198
rect 15228 24179 15262 24213
rect 16003 24180 16037 24214
rect 16834 24248 16868 24282
rect 16454 24163 16488 24197
rect 16572 24164 16606 24198
rect 17126 24179 17160 24213
rect 13131 24081 13165 24115
rect 13013 23964 13047 23998
rect 13958 23937 13992 24113
rect 12601 23538 12635 23914
rect 12719 23538 12753 23914
rect 12837 23538 12871 23914
rect 12954 23738 12988 23914
rect 14076 23937 14110 24113
rect 13072 23738 13106 23914
rect 14378 23737 14412 24113
rect 14496 23737 14530 24113
rect 14614 23737 14648 24113
rect 14732 23737 14766 24113
rect 14850 23737 14884 24113
rect 15256 23937 15290 24113
rect 15374 23937 15408 24113
rect 15856 23937 15890 24113
rect 15974 23937 16008 24113
rect 16276 23737 16310 24113
rect 16394 23737 16428 24113
rect 16512 23737 16546 24113
rect 16630 23737 16664 24113
rect 16748 23737 16782 24113
rect 17154 23937 17188 24113
rect 17272 23937 17306 24113
rect 12660 23454 12694 23488
rect 12778 23454 12812 23488
rect 18898 24170 18932 24346
rect 19016 24170 19050 24346
rect 19134 24170 19168 24346
rect 19252 24170 19286 24346
rect 19370 24170 19404 24346
rect 19488 24170 19522 24346
rect 19606 24170 19640 24346
rect 19724 24170 19758 24346
rect 19842 24170 19876 24346
rect 21030 24464 21064 24840
rect 21148 24464 21182 24840
rect 21266 24464 21300 24840
rect 21384 24464 21418 24840
rect 21502 24464 21536 24840
rect 22692 24464 22726 24840
rect 22810 24464 22844 24840
rect 22928 24464 22962 24840
rect 23046 24464 23080 24840
rect 23164 24464 23198 24840
rect 23282 24464 23316 24840
rect 30496 24868 30530 24902
rect 23400 24464 23434 24840
rect 27352 24468 27386 24844
rect 27470 24468 27504 24844
rect 19960 24170 19994 24346
rect 20824 24242 20858 24276
rect 20639 24175 20673 24209
rect 21472 24242 21506 24276
rect 22722 24242 22756 24276
rect 21090 24158 21124 24192
rect 21208 24159 21242 24193
rect 21762 24174 21796 24208
rect 22537 24175 22571 24209
rect 23368 24243 23402 24277
rect 22988 24158 23022 24192
rect 23106 24159 23140 24193
rect 23660 24174 23694 24208
rect 19665 24076 19699 24110
rect 19547 23959 19581 23993
rect 20492 23932 20526 24108
rect 19135 23533 19169 23909
rect 19253 23533 19287 23909
rect 19371 23533 19405 23909
rect 19488 23733 19522 23909
rect 20610 23932 20644 24108
rect 19606 23733 19640 23909
rect 20912 23732 20946 24108
rect 21030 23732 21064 24108
rect 21148 23732 21182 24108
rect 21266 23732 21300 24108
rect 21384 23732 21418 24108
rect 21790 23932 21824 24108
rect 21908 23932 21942 24108
rect 22390 23932 22424 24108
rect 22508 23932 22542 24108
rect 22810 23732 22844 24108
rect 22928 23732 22962 24108
rect 23046 23732 23080 24108
rect 23164 23732 23198 24108
rect 23282 23732 23316 24108
rect 23688 23932 23722 24108
rect 23806 23932 23840 24108
rect 19194 23449 19228 23483
rect 19312 23449 19346 23483
rect 25456 24174 25490 24350
rect 25574 24174 25608 24350
rect 25692 24174 25726 24350
rect 25810 24174 25844 24350
rect 25928 24174 25962 24350
rect 26046 24174 26080 24350
rect 26164 24174 26198 24350
rect 26282 24174 26316 24350
rect 26400 24174 26434 24350
rect 27588 24468 27622 24844
rect 27706 24468 27740 24844
rect 27824 24468 27858 24844
rect 27942 24468 27976 24844
rect 28060 24468 28094 24844
rect 29250 24468 29284 24844
rect 29368 24468 29402 24844
rect 29486 24468 29520 24844
rect 29604 24468 29638 24844
rect 29722 24468 29756 24844
rect 29840 24468 29874 24844
rect 29958 24468 29992 24844
rect 26518 24174 26552 24350
rect 27382 24246 27416 24280
rect 27197 24179 27231 24213
rect 28030 24246 28064 24280
rect 29280 24246 29314 24280
rect 27648 24162 27682 24196
rect 27766 24163 27800 24197
rect 28320 24178 28354 24212
rect 29095 24179 29129 24213
rect 32159 24351 32304 24429
rect 29926 24247 29960 24281
rect 29546 24162 29580 24196
rect 29664 24163 29698 24197
rect 30218 24178 30252 24212
rect 26223 24080 26257 24114
rect 26105 23963 26139 23997
rect 27050 23936 27084 24112
rect 25693 23537 25727 23913
rect 25811 23537 25845 23913
rect 25929 23537 25963 23913
rect 26046 23737 26080 23913
rect 27168 23936 27202 24112
rect 26164 23737 26198 23913
rect 27470 23736 27504 24112
rect 27588 23736 27622 24112
rect 27706 23736 27740 24112
rect 27824 23736 27858 24112
rect 27942 23736 27976 24112
rect 28348 23936 28382 24112
rect 28466 23936 28500 24112
rect 28948 23936 28982 24112
rect 29066 23936 29100 24112
rect 29368 23736 29402 24112
rect 29486 23736 29520 24112
rect 29604 23736 29638 24112
rect 29722 23736 29756 24112
rect 29840 23736 29874 24112
rect 30246 23936 30280 24112
rect 30364 23936 30398 24112
rect 25752 23453 25786 23487
rect 25870 23453 25904 23487
rect 32676 22977 32811 23049
rect 33244 22809 33374 22899
rect 37741 25238 37801 25287
rect 36967 25114 37143 25148
rect 36967 24996 37143 25030
rect 36967 24878 37143 24912
rect 37458 24985 37513 25043
rect 37458 24983 37513 24985
rect 36967 24760 37143 24794
rect 36767 24673 37143 24707
rect 36767 24555 37143 24589
rect 36767 24437 37143 24471
rect 36767 24319 37143 24353
rect 36767 24206 37143 24240
rect 38100 24280 38276 24314
rect 38100 24162 38276 24196
rect 36767 24088 37143 24122
rect 36767 23970 37143 24004
rect 36517 23824 36571 23896
rect 38100 24088 38476 24122
rect 37358 24028 37392 24062
rect 37742 24074 37797 24076
rect 37742 24016 37797 24074
rect 36767 23852 37143 23886
rect 38100 23970 38476 24004
rect 37457 23956 37512 23958
rect 37457 23898 37512 23956
rect 38100 23852 38476 23886
rect 36767 23734 37143 23768
rect 38577 23851 38611 23885
rect 37978 23793 38012 23827
rect 38729 23824 38743 23882
rect 38743 23824 38775 23882
rect 38100 23734 38476 23768
rect 37588 23674 37622 23708
rect 36767 23616 37143 23650
rect 38100 23616 38476 23650
rect 36767 23498 37143 23532
rect 38100 23538 38276 23572
rect 38100 23420 38276 23454
rect 36767 23379 37143 23413
rect 36767 23261 37143 23295
rect 36767 23143 37143 23177
rect 36767 23025 37143 23059
rect 36967 22906 37143 22940
rect 6688 22220 6722 22254
rect 7818 22214 7852 22248
rect 13246 22216 13280 22250
rect 14376 22210 14410 22244
rect 19780 22221 19814 22255
rect 20910 22215 20944 22249
rect 36967 22788 37143 22822
rect 36967 22670 37143 22704
rect 37317 22718 37351 22752
rect 36967 22552 37143 22586
rect 26293 22224 26327 22258
rect 27423 22218 27457 22252
rect 6688 22100 6722 22134
rect 5853 21700 5887 22076
rect 5971 21700 6005 22076
rect 6089 21700 6123 22076
rect 6207 21700 6241 22076
rect 6325 21700 6359 22076
rect 6443 21700 6477 22076
rect 7818 22096 7852 22130
rect 6561 21700 6595 22076
rect 6995 21696 7029 22072
rect 7113 21696 7147 22072
rect 7231 21696 7265 22072
rect 7349 21696 7383 22072
rect 7467 21696 7501 22072
rect 7585 21696 7619 22072
rect 13246 22096 13280 22130
rect 7703 21696 7737 22072
rect 8966 21824 9000 22000
rect 9084 21824 9118 22000
rect 9202 21824 9236 22000
rect 9320 21824 9354 22000
rect 9438 21824 9472 22000
rect 9556 21824 9590 22000
rect 9674 21824 9708 22000
rect 9792 21824 9826 22000
rect 9910 21824 9944 22000
rect 10028 21824 10062 22000
rect 9261 21730 9295 21764
rect 12411 21696 12445 22072
rect 12529 21696 12563 22072
rect 12647 21696 12681 22072
rect 12765 21696 12799 22072
rect 12883 21696 12917 22072
rect 13001 21696 13035 22072
rect 14376 22092 14410 22126
rect 19780 22101 19814 22135
rect 13119 21696 13153 22072
rect 13553 21692 13587 22068
rect 13671 21692 13705 22068
rect 13789 21692 13823 22068
rect 13907 21692 13941 22068
rect 14025 21692 14059 22068
rect 14143 21692 14177 22068
rect 14261 21692 14295 22068
rect 15524 21820 15558 21996
rect 15642 21820 15676 21996
rect 15760 21820 15794 21996
rect 15878 21820 15912 21996
rect 15996 21820 16030 21996
rect 16114 21820 16148 21996
rect 16232 21820 16266 21996
rect 16350 21820 16384 21996
rect 16468 21820 16502 21996
rect 16586 21820 16620 21996
rect 15819 21726 15853 21760
rect 18945 21701 18979 22077
rect 19063 21701 19097 22077
rect 19181 21701 19215 22077
rect 19299 21701 19333 22077
rect 19417 21701 19451 22077
rect 19535 21701 19569 22077
rect 20910 22097 20944 22131
rect 19653 21701 19687 22077
rect 20087 21697 20121 22073
rect 20205 21697 20239 22073
rect 20323 21697 20357 22073
rect 20441 21697 20475 22073
rect 20559 21697 20593 22073
rect 20677 21697 20711 22073
rect 26293 22104 26327 22138
rect 20795 21697 20829 22073
rect 22058 21825 22092 22001
rect 22176 21825 22210 22001
rect 22294 21825 22328 22001
rect 22412 21825 22446 22001
rect 22530 21825 22564 22001
rect 22648 21825 22682 22001
rect 22766 21825 22800 22001
rect 22884 21825 22918 22001
rect 23002 21825 23036 22001
rect 23120 21825 23154 22001
rect 22353 21731 22387 21765
rect 25458 21704 25492 22080
rect 25576 21704 25610 22080
rect 25694 21704 25728 22080
rect 25812 21704 25846 22080
rect 25930 21704 25964 22080
rect 26048 21704 26082 22080
rect 27423 22100 27457 22134
rect 26166 21704 26200 22080
rect 26600 21700 26634 22076
rect 26718 21700 26752 22076
rect 26836 21700 26870 22076
rect 26954 21700 26988 22076
rect 27072 21700 27106 22076
rect 27190 21700 27224 22076
rect 27308 21700 27342 22076
rect 28571 21828 28605 22004
rect 28689 21828 28723 22004
rect 28807 21828 28841 22004
rect 28925 21828 28959 22004
rect 29043 21828 29077 22004
rect 29161 21828 29195 22004
rect 29279 21828 29313 22004
rect 29397 21828 29431 22004
rect 29515 21828 29549 22004
rect 29633 21828 29667 22004
rect 28866 21734 28900 21768
rect 9379 21613 9413 21647
rect 15937 21609 15971 21643
rect 22471 21614 22505 21648
rect 28984 21617 29018 21651
rect 9320 21387 9354 21563
rect 6356 21344 6390 21378
rect 7498 21340 7532 21374
rect 9438 21387 9472 21563
rect 5778 21117 5812 21293
rect 5896 21117 5930 21293
rect 6014 21117 6048 21293
rect 6132 21117 6166 21293
rect 6297 21117 6331 21293
rect 6415 21117 6449 21293
rect 6533 21117 6567 21293
rect 6651 21117 6685 21293
rect 6920 21113 6954 21289
rect 7038 21113 7072 21289
rect 7156 21113 7190 21289
rect 7274 21113 7308 21289
rect 7439 21113 7473 21289
rect 7557 21113 7591 21289
rect 7675 21113 7709 21289
rect 7793 21113 7827 21289
rect 9555 21187 9589 21563
rect 9673 21187 9707 21563
rect 9791 21187 9825 21563
rect 15878 21383 15912 21559
rect 12914 21340 12948 21374
rect 14056 21336 14090 21370
rect 15996 21383 16030 21559
rect 9614 21103 9648 21137
rect 9732 21103 9766 21137
rect 12336 21113 12370 21289
rect 12454 21113 12488 21289
rect 12572 21113 12606 21289
rect 12690 21113 12724 21289
rect 12855 21113 12889 21289
rect 12973 21113 13007 21289
rect 13091 21113 13125 21289
rect 13209 21113 13243 21289
rect 13478 21109 13512 21285
rect 13596 21109 13630 21285
rect 13714 21109 13748 21285
rect 13832 21109 13866 21285
rect 13997 21109 14031 21285
rect 14115 21109 14149 21285
rect 14233 21109 14267 21285
rect 14351 21109 14385 21285
rect 16113 21183 16147 21559
rect 16231 21183 16265 21559
rect 16349 21183 16383 21559
rect 22412 21388 22446 21564
rect 19448 21345 19482 21379
rect 20590 21341 20624 21375
rect 22530 21388 22564 21564
rect 16172 21099 16206 21133
rect 16290 21099 16324 21133
rect 18870 21118 18904 21294
rect 18988 21118 19022 21294
rect 19106 21118 19140 21294
rect 19224 21118 19258 21294
rect 19389 21118 19423 21294
rect 19507 21118 19541 21294
rect 19625 21118 19659 21294
rect 19743 21118 19777 21294
rect 20012 21114 20046 21290
rect 20130 21114 20164 21290
rect 20248 21114 20282 21290
rect 20366 21114 20400 21290
rect 20531 21114 20565 21290
rect 20649 21114 20683 21290
rect 20767 21114 20801 21290
rect 20885 21114 20919 21290
rect 22647 21188 22681 21564
rect 22765 21188 22799 21564
rect 22883 21188 22917 21564
rect 28925 21391 28959 21567
rect 25961 21348 25995 21382
rect 27103 21344 27137 21378
rect 29043 21391 29077 21567
rect 22706 21104 22740 21138
rect 22824 21104 22858 21138
rect 25383 21121 25417 21297
rect 25501 21121 25535 21297
rect 25619 21121 25653 21297
rect 25737 21121 25771 21297
rect 25902 21121 25936 21297
rect 26020 21121 26054 21297
rect 26138 21121 26172 21297
rect 26256 21121 26290 21297
rect 26525 21117 26559 21293
rect 26643 21117 26677 21293
rect 26761 21117 26795 21293
rect 26879 21117 26913 21293
rect 27044 21117 27078 21293
rect 27162 21117 27196 21293
rect 27280 21117 27314 21293
rect 27398 21117 27432 21293
rect 29160 21191 29194 21567
rect 29278 21191 29312 21567
rect 29396 21191 29430 21567
rect 29219 21107 29253 21141
rect 29337 21107 29371 21141
rect 10738 20549 10849 20658
rect 8952 20174 8986 20350
rect 9070 20174 9104 20350
rect 9188 20174 9222 20350
rect 9306 20174 9340 20350
rect 9424 20174 9458 20350
rect 9542 20174 9576 20350
rect 9660 20174 9694 20350
rect 9778 20174 9812 20350
rect 9896 20174 9930 20350
rect 10014 20174 10048 20350
rect 9247 20080 9281 20114
rect 4977 19557 5011 19733
rect 5095 19557 5129 19733
rect 5213 19557 5247 19733
rect 5331 19557 5365 19733
rect 5460 19557 5494 19933
rect 5578 19557 5612 19933
rect 5696 19557 5730 19933
rect 5814 19557 5848 19933
rect 5932 19557 5966 19933
rect 6050 19557 6084 19933
rect 6168 19557 6202 19933
rect 6298 19557 6332 19733
rect 6416 19557 6450 19733
rect 6534 19557 6568 19733
rect 6652 19557 6686 19733
rect 6875 19557 6909 19733
rect 6993 19557 7027 19733
rect 7111 19557 7145 19733
rect 7229 19557 7263 19733
rect 7358 19557 7392 19933
rect 7476 19557 7510 19933
rect 7594 19557 7628 19933
rect 9365 19963 9399 19997
rect 7712 19557 7746 19933
rect 7830 19557 7864 19933
rect 7948 19557 7982 19933
rect 8066 19557 8100 19933
rect 8196 19557 8230 19733
rect 8314 19557 8348 19733
rect 8432 19557 8466 19733
rect 8550 19557 8584 19733
rect 9306 19737 9340 19913
rect 9424 19737 9458 19913
rect 9541 19537 9575 19913
rect 9659 19537 9693 19913
rect 9777 19537 9811 19913
rect 9600 19453 9634 19487
rect 9718 19453 9752 19487
rect 4979 19264 5013 19298
rect 7086 19285 7120 19319
rect 5517 18864 5551 19240
rect 5635 18864 5669 19240
rect 4758 18737 4890 18835
rect 5753 18864 5787 19240
rect 5871 18864 5905 19240
rect 5989 18864 6023 19240
rect 6107 18864 6141 19240
rect 6225 18864 6259 19240
rect 7415 18864 7449 19240
rect 7533 18864 7567 19240
rect 7651 18864 7685 19240
rect 7769 18864 7803 19240
rect 7887 18864 7921 19240
rect 8005 18864 8039 19240
rect 8123 18864 8157 19240
rect 5549 18643 5583 18677
rect 5257 18574 5291 18608
rect 5811 18559 5845 18593
rect 5929 18558 5963 18592
rect 6195 18642 6229 18676
rect 7445 18642 7479 18676
rect 6380 18575 6414 18609
rect 7155 18574 7189 18608
rect 7709 18559 7743 18593
rect 7827 18558 7861 18592
rect 8093 18642 8127 18676
rect 8278 18575 8312 18609
rect 8957 18570 8991 18746
rect 9075 18570 9109 18746
rect 9193 18570 9227 18746
rect 9311 18570 9345 18746
rect 9429 18570 9463 18746
rect 9547 18570 9581 18746
rect 9665 18570 9699 18746
rect 9783 18570 9817 18746
rect 9901 18570 9935 18746
rect 10019 18570 10053 18746
rect 5111 18332 5145 18508
rect 5229 18332 5263 18508
rect 5635 18132 5669 18508
rect 5753 18132 5787 18508
rect 5871 18132 5905 18508
rect 5989 18132 6023 18508
rect 6107 18132 6141 18508
rect 6409 18332 6443 18508
rect 6527 18332 6561 18508
rect 7009 18332 7043 18508
rect 7127 18332 7161 18508
rect 7533 18132 7567 18508
rect 7651 18132 7685 18508
rect 7769 18132 7803 18508
rect 7887 18132 7921 18508
rect 8005 18132 8039 18508
rect 8307 18332 8341 18508
rect 8425 18332 8459 18508
rect 9252 18476 9286 18510
rect 9370 18359 9404 18393
rect 9311 18133 9345 18309
rect 9429 18133 9463 18309
rect 9546 17933 9580 18309
rect 9664 17933 9698 18309
rect 9782 17933 9816 18309
rect 9605 17849 9639 17883
rect 9723 17849 9757 17883
rect 17301 20549 17404 20646
rect 15510 20170 15544 20346
rect 15628 20170 15662 20346
rect 15746 20170 15780 20346
rect 15864 20170 15898 20346
rect 15982 20170 16016 20346
rect 16100 20170 16134 20346
rect 16218 20170 16252 20346
rect 16336 20170 16370 20346
rect 16454 20170 16488 20346
rect 16572 20170 16606 20346
rect 15805 20076 15839 20110
rect 11535 19553 11569 19729
rect 11653 19553 11687 19729
rect 11771 19553 11805 19729
rect 11889 19553 11923 19729
rect 12018 19553 12052 19929
rect 12136 19553 12170 19929
rect 12254 19553 12288 19929
rect 12372 19553 12406 19929
rect 12490 19553 12524 19929
rect 12608 19553 12642 19929
rect 12726 19553 12760 19929
rect 12856 19553 12890 19729
rect 12974 19553 13008 19729
rect 13092 19553 13126 19729
rect 13210 19553 13244 19729
rect 13433 19553 13467 19729
rect 13551 19553 13585 19729
rect 13669 19553 13703 19729
rect 13787 19553 13821 19729
rect 13916 19553 13950 19929
rect 14034 19553 14068 19929
rect 14152 19553 14186 19929
rect 15923 19959 15957 19993
rect 14270 19553 14304 19929
rect 14388 19553 14422 19929
rect 14506 19553 14540 19929
rect 14624 19553 14658 19929
rect 14754 19553 14788 19729
rect 14872 19553 14906 19729
rect 14990 19553 15024 19729
rect 15108 19553 15142 19729
rect 15864 19733 15898 19909
rect 15982 19733 16016 19909
rect 16099 19533 16133 19909
rect 16217 19533 16251 19909
rect 16335 19533 16369 19909
rect 16158 19449 16192 19483
rect 16276 19449 16310 19483
rect 11537 19260 11571 19294
rect 13644 19281 13678 19315
rect 12075 18860 12109 19236
rect 12193 18860 12227 19236
rect 11316 18733 11448 18831
rect 12311 18860 12345 19236
rect 12429 18860 12463 19236
rect 12547 18860 12581 19236
rect 12665 18860 12699 19236
rect 12783 18860 12817 19236
rect 13973 18860 14007 19236
rect 14091 18860 14125 19236
rect 14209 18860 14243 19236
rect 14327 18860 14361 19236
rect 14445 18860 14479 19236
rect 14563 18860 14597 19236
rect 14681 18860 14715 19236
rect 12107 18639 12141 18673
rect 11815 18570 11849 18604
rect 12369 18555 12403 18589
rect 12487 18554 12521 18588
rect 12753 18638 12787 18672
rect 14003 18638 14037 18672
rect 12938 18571 12972 18605
rect 13713 18570 13747 18604
rect 14267 18555 14301 18589
rect 14385 18554 14419 18588
rect 14651 18638 14685 18672
rect 14836 18571 14870 18605
rect 15515 18566 15549 18742
rect 15633 18566 15667 18742
rect 15751 18566 15785 18742
rect 15869 18566 15903 18742
rect 15987 18566 16021 18742
rect 16105 18566 16139 18742
rect 16223 18566 16257 18742
rect 16341 18566 16375 18742
rect 16459 18566 16493 18742
rect 16577 18566 16611 18742
rect 11669 18328 11703 18504
rect 11787 18328 11821 18504
rect 12193 18128 12227 18504
rect 12311 18128 12345 18504
rect 12429 18128 12463 18504
rect 12547 18128 12581 18504
rect 12665 18128 12699 18504
rect 12967 18328 13001 18504
rect 13085 18328 13119 18504
rect 13567 18328 13601 18504
rect 13685 18328 13719 18504
rect 14091 18128 14125 18504
rect 14209 18128 14243 18504
rect 14327 18128 14361 18504
rect 14445 18128 14479 18504
rect 14563 18128 14597 18504
rect 14865 18328 14899 18504
rect 14983 18328 15017 18504
rect 15810 18472 15844 18506
rect 15928 18355 15962 18389
rect 15869 18129 15903 18305
rect 15987 18129 16021 18305
rect 16104 17929 16138 18305
rect 16222 17929 16256 18305
rect 16340 17929 16374 18305
rect 16163 17845 16197 17879
rect 16281 17845 16315 17879
rect 23837 20558 23935 20650
rect 22044 20175 22078 20351
rect 22162 20175 22196 20351
rect 22280 20175 22314 20351
rect 22398 20175 22432 20351
rect 22516 20175 22550 20351
rect 22634 20175 22668 20351
rect 22752 20175 22786 20351
rect 22870 20175 22904 20351
rect 22988 20175 23022 20351
rect 23106 20175 23140 20351
rect 22339 20081 22373 20115
rect 18069 19558 18103 19734
rect 18187 19558 18221 19734
rect 18305 19558 18339 19734
rect 18423 19558 18457 19734
rect 18552 19558 18586 19934
rect 18670 19558 18704 19934
rect 18788 19558 18822 19934
rect 18906 19558 18940 19934
rect 19024 19558 19058 19934
rect 19142 19558 19176 19934
rect 19260 19558 19294 19934
rect 19390 19558 19424 19734
rect 19508 19558 19542 19734
rect 19626 19558 19660 19734
rect 19744 19558 19778 19734
rect 19967 19558 20001 19734
rect 20085 19558 20119 19734
rect 20203 19558 20237 19734
rect 20321 19558 20355 19734
rect 20450 19558 20484 19934
rect 20568 19558 20602 19934
rect 20686 19558 20720 19934
rect 22457 19964 22491 19998
rect 20804 19558 20838 19934
rect 20922 19558 20956 19934
rect 21040 19558 21074 19934
rect 21158 19558 21192 19934
rect 21288 19558 21322 19734
rect 21406 19558 21440 19734
rect 21524 19558 21558 19734
rect 21642 19558 21676 19734
rect 22398 19738 22432 19914
rect 22516 19738 22550 19914
rect 22633 19538 22667 19914
rect 22751 19538 22785 19914
rect 22869 19538 22903 19914
rect 22692 19454 22726 19488
rect 22810 19454 22844 19488
rect 18071 19265 18105 19299
rect 20178 19286 20212 19320
rect 18609 18865 18643 19241
rect 18727 18865 18761 19241
rect 17850 18738 17982 18836
rect 18845 18865 18879 19241
rect 18963 18865 18997 19241
rect 19081 18865 19115 19241
rect 19199 18865 19233 19241
rect 19317 18865 19351 19241
rect 20507 18865 20541 19241
rect 20625 18865 20659 19241
rect 20743 18865 20777 19241
rect 20861 18865 20895 19241
rect 20979 18865 21013 19241
rect 21097 18865 21131 19241
rect 21215 18865 21249 19241
rect 18641 18644 18675 18678
rect 18349 18575 18383 18609
rect 18903 18560 18937 18594
rect 19021 18559 19055 18593
rect 19287 18643 19321 18677
rect 20537 18643 20571 18677
rect 19472 18576 19506 18610
rect 20247 18575 20281 18609
rect 20801 18560 20835 18594
rect 20919 18559 20953 18593
rect 21185 18643 21219 18677
rect 21370 18576 21404 18610
rect 22049 18571 22083 18747
rect 22167 18571 22201 18747
rect 22285 18571 22319 18747
rect 22403 18571 22437 18747
rect 22521 18571 22555 18747
rect 22639 18571 22673 18747
rect 22757 18571 22791 18747
rect 22875 18571 22909 18747
rect 22993 18571 23027 18747
rect 23111 18571 23145 18747
rect 18203 18333 18237 18509
rect 18321 18333 18355 18509
rect 18727 18133 18761 18509
rect 18845 18133 18879 18509
rect 18963 18133 18997 18509
rect 19081 18133 19115 18509
rect 19199 18133 19233 18509
rect 19501 18333 19535 18509
rect 19619 18333 19653 18509
rect 20101 18333 20135 18509
rect 20219 18333 20253 18509
rect 20625 18133 20659 18509
rect 20743 18133 20777 18509
rect 20861 18133 20895 18509
rect 20979 18133 21013 18509
rect 21097 18133 21131 18509
rect 21399 18333 21433 18509
rect 21517 18333 21551 18509
rect 22344 18477 22378 18511
rect 22462 18360 22496 18394
rect 22403 18134 22437 18310
rect 22521 18134 22555 18310
rect 22638 17934 22672 18310
rect 22756 17934 22790 18310
rect 22874 17934 22908 18310
rect 22697 17850 22731 17884
rect 22815 17850 22849 17884
rect 28557 20178 28591 20354
rect 28675 20178 28709 20354
rect 28793 20178 28827 20354
rect 28911 20178 28945 20354
rect 29029 20178 29063 20354
rect 29147 20178 29181 20354
rect 29265 20178 29299 20354
rect 29383 20178 29417 20354
rect 29501 20178 29535 20354
rect 29619 20178 29653 20354
rect 28852 20084 28886 20118
rect 24582 19561 24616 19737
rect 24700 19561 24734 19737
rect 24818 19561 24852 19737
rect 24936 19561 24970 19737
rect 25065 19561 25099 19937
rect 25183 19561 25217 19937
rect 25301 19561 25335 19937
rect 25419 19561 25453 19937
rect 25537 19561 25571 19937
rect 25655 19561 25689 19937
rect 25773 19561 25807 19937
rect 25903 19561 25937 19737
rect 26021 19561 26055 19737
rect 26139 19561 26173 19737
rect 26257 19561 26291 19737
rect 26480 19561 26514 19737
rect 26598 19561 26632 19737
rect 26716 19561 26750 19737
rect 26834 19561 26868 19737
rect 26963 19561 26997 19937
rect 27081 19561 27115 19937
rect 27199 19561 27233 19937
rect 28970 19967 29004 20001
rect 27317 19561 27351 19937
rect 27435 19561 27469 19937
rect 27553 19561 27587 19937
rect 27671 19561 27705 19937
rect 27801 19561 27835 19737
rect 27919 19561 27953 19737
rect 28037 19561 28071 19737
rect 28155 19561 28189 19737
rect 28911 19741 28945 19917
rect 29029 19741 29063 19917
rect 29146 19541 29180 19917
rect 29264 19541 29298 19917
rect 29382 19541 29416 19917
rect 29205 19457 29239 19491
rect 29323 19457 29357 19491
rect 24584 19268 24618 19302
rect 26691 19289 26725 19323
rect 25122 18868 25156 19244
rect 25240 18868 25274 19244
rect 24363 18741 24495 18839
rect 25358 18868 25392 19244
rect 25476 18868 25510 19244
rect 25594 18868 25628 19244
rect 25712 18868 25746 19244
rect 25830 18868 25864 19244
rect 27020 18868 27054 19244
rect 27138 18868 27172 19244
rect 27256 18868 27290 19244
rect 27374 18868 27408 19244
rect 27492 18868 27526 19244
rect 27610 18868 27644 19244
rect 27728 18868 27762 19244
rect 25154 18647 25188 18681
rect 24862 18578 24896 18612
rect 25416 18563 25450 18597
rect 25534 18562 25568 18596
rect 25800 18646 25834 18680
rect 27050 18646 27084 18680
rect 25985 18579 26019 18613
rect 26760 18578 26794 18612
rect 27314 18563 27348 18597
rect 27432 18562 27466 18596
rect 27698 18646 27732 18680
rect 27883 18579 27917 18613
rect 28562 18574 28596 18750
rect 28680 18574 28714 18750
rect 28798 18574 28832 18750
rect 28916 18574 28950 18750
rect 29034 18574 29068 18750
rect 29152 18574 29186 18750
rect 29270 18574 29304 18750
rect 29388 18574 29422 18750
rect 29506 18574 29540 18750
rect 29624 18574 29658 18750
rect 24716 18336 24750 18512
rect 24834 18336 24868 18512
rect 25240 18136 25274 18512
rect 25358 18136 25392 18512
rect 25476 18136 25510 18512
rect 25594 18136 25628 18512
rect 25712 18136 25746 18512
rect 26014 18336 26048 18512
rect 26132 18336 26166 18512
rect 26614 18336 26648 18512
rect 26732 18336 26766 18512
rect 27138 18136 27172 18512
rect 27256 18136 27290 18512
rect 27374 18136 27408 18512
rect 27492 18136 27526 18512
rect 27610 18136 27644 18512
rect 27912 18336 27946 18512
rect 28030 18336 28064 18512
rect 28857 18480 28891 18514
rect 28975 18363 29009 18397
rect 28916 18137 28950 18313
rect 29034 18137 29068 18313
rect 29151 17937 29185 18313
rect 29269 17937 29303 18313
rect 29387 17937 29421 18313
rect 29210 17853 29244 17887
rect 29328 17853 29362 17887
rect 23984 16184 24052 16242
rect 17459 16067 17530 16123
rect 34502 22173 34551 22236
rect 37741 22094 37801 22143
rect 36967 21970 37143 22004
rect 36967 21852 37143 21886
rect 36967 21734 37143 21768
rect 37458 21841 37513 21899
rect 37458 21839 37513 21841
rect 36967 21616 37143 21650
rect 36767 21529 37143 21563
rect 36767 21411 37143 21445
rect 36767 21293 37143 21327
rect 36767 21175 37143 21209
rect 36767 21062 37143 21096
rect 38100 21136 38276 21170
rect 38100 21018 38276 21052
rect 36767 20944 37143 20978
rect 36767 20826 37143 20860
rect 36517 20680 36571 20752
rect 38100 20944 38476 20978
rect 37358 20884 37392 20918
rect 37742 20930 37797 20932
rect 37742 20872 37797 20930
rect 36767 20708 37143 20742
rect 38100 20826 38476 20860
rect 37457 20812 37512 20814
rect 37457 20754 37512 20812
rect 38100 20708 38476 20742
rect 36767 20590 37143 20624
rect 38577 20707 38611 20741
rect 37978 20649 38012 20683
rect 38729 20680 38743 20738
rect 38743 20680 38775 20738
rect 38100 20590 38476 20624
rect 37588 20530 37622 20564
rect 36767 20472 37143 20506
rect 38100 20472 38476 20506
rect 36767 20354 37143 20388
rect 38100 20394 38276 20428
rect 38100 20276 38276 20310
rect 36767 20235 37143 20269
rect 36767 20117 37143 20151
rect 36767 19999 37143 20033
rect 36767 19881 37143 19915
rect 36967 19762 37143 19796
rect 36967 19644 37143 19678
rect 36967 19526 37143 19560
rect 37317 19574 37351 19608
rect 36967 19408 37143 19442
rect 10883 15745 10962 15790
rect 8153 15400 8213 15462
rect 14702 15399 14762 15461
rect 21356 15420 21416 15482
rect 30852 15380 30930 15452
rect 7812 15048 7846 15224
rect 7930 15048 7964 15224
rect 8048 15048 8082 15224
rect 8166 15048 8200 15224
rect 8284 15048 8318 15224
rect 8402 15048 8436 15224
rect 8520 15048 8554 15224
rect 8638 15048 8672 15224
rect 8756 15048 8790 15224
rect 8874 15048 8908 15224
rect 14361 15047 14395 15223
rect 14479 15047 14513 15223
rect 14597 15047 14631 15223
rect 14715 15047 14749 15223
rect 14833 15047 14867 15223
rect 14951 15047 14985 15223
rect 15069 15047 15103 15223
rect 15187 15047 15221 15223
rect 15305 15047 15339 15223
rect 15423 15047 15457 15223
rect 21015 15068 21049 15244
rect 21133 15068 21167 15244
rect 21251 15068 21285 15244
rect 21369 15068 21403 15244
rect 21487 15068 21521 15244
rect 21605 15068 21639 15244
rect 21723 15068 21757 15244
rect 21841 15068 21875 15244
rect 21959 15068 21993 15244
rect 22077 15068 22111 15244
rect 30009 15253 30069 15315
rect 32110 15376 32531 15410
rect 32110 15231 32173 15376
rect 32173 15231 32482 15376
rect 32482 15231 32531 15376
rect 32110 15210 32531 15231
rect 8579 14954 8613 14988
rect 15128 14953 15162 14987
rect 21782 14974 21816 15008
rect 29668 14901 29702 15077
rect 8461 14837 8495 14871
rect 15010 14836 15044 14870
rect 21664 14857 21698 14891
rect 29786 14901 29820 15077
rect 29904 14901 29938 15077
rect 30022 14901 30056 15077
rect 30140 14901 30174 15077
rect 30258 14901 30292 15077
rect 30376 14901 30410 15077
rect 30494 14901 30528 15077
rect 30612 14901 30646 15077
rect 30730 14901 30764 15077
rect 8049 14411 8083 14787
rect 8167 14411 8201 14787
rect 8285 14411 8319 14787
rect 8402 14611 8436 14787
rect 8520 14611 8554 14787
rect 14598 14410 14632 14786
rect 14716 14410 14750 14786
rect 14834 14410 14868 14786
rect 14951 14610 14985 14786
rect 15069 14610 15103 14786
rect 21252 14431 21286 14807
rect 21370 14431 21404 14807
rect 21488 14431 21522 14807
rect 21605 14631 21639 14807
rect 30435 14807 30469 14841
rect 21723 14631 21757 14807
rect 30317 14690 30351 14724
rect 8108 14327 8142 14361
rect 8226 14327 8260 14361
rect 14511 14315 14560 14361
rect 14657 14326 14691 14360
rect 14775 14326 14809 14360
rect 21118 14335 21179 14383
rect 21311 14347 21345 14381
rect 21429 14347 21463 14381
rect 8381 14204 8433 14250
rect 66 13871 125 13927
rect 227 14059 288 14109
rect 23 12512 97 12582
rect 14930 14203 14982 14249
rect 7930 13882 7979 13936
rect 21220 14255 21265 14293
rect 21584 14224 21636 14270
rect 29905 14264 29939 14640
rect 30023 14264 30057 14640
rect 30141 14264 30175 14640
rect 30258 14464 30292 14640
rect 30376 14464 30410 14640
rect 31476 14496 31510 14672
rect 31594 14496 31628 14672
rect 31712 14496 31746 14672
rect 31830 14496 31864 14672
rect 31960 14496 31994 14872
rect 32078 14496 32112 14872
rect 32196 14496 32230 14872
rect 32314 14496 32348 14872
rect 32432 14496 32466 14872
rect 32550 14496 32584 14872
rect 32668 14496 32702 14872
rect 33610 14845 33670 14907
rect 32797 14496 32831 14672
rect 32915 14496 32949 14672
rect 33033 14496 33067 14672
rect 33151 14496 33185 14672
rect 33269 14493 33303 14669
rect 33387 14493 33421 14669
rect 33505 14493 33539 14669
rect 33623 14493 33657 14669
rect 33741 14493 33775 14669
rect 33859 14493 33893 14669
rect 33977 14493 34011 14669
rect 34095 14493 34129 14669
rect 34213 14493 34247 14669
rect 34331 14493 34365 14669
rect 34036 14399 34070 14433
rect 33128 14280 33162 14314
rect 33918 14282 33952 14316
rect 29964 14180 29998 14214
rect 30082 14180 30116 14214
rect 31455 14140 31535 14208
rect 31728 14161 31762 14195
rect 30237 14057 30289 14103
rect 380 13491 437 13536
rect 207 12318 320 12402
rect 20 9694 114 9775
rect 21 3919 103 4001
rect 15 821 109 897
rect 1489 13500 1549 13562
rect 1148 13148 1182 13324
rect 1266 13148 1300 13324
rect 1384 13148 1418 13324
rect 1502 13148 1536 13324
rect 1620 13148 1654 13324
rect 1738 13148 1772 13324
rect 1856 13148 1890 13324
rect 1974 13148 2008 13324
rect 2092 13148 2126 13324
rect 2210 13148 2244 13324
rect 1915 13054 1949 13088
rect 1797 12937 1831 12971
rect 499 3919 601 4000
rect 645 12504 734 12580
rect 1385 12511 1419 12887
rect 1503 12511 1537 12887
rect 1621 12511 1655 12887
rect 1738 12711 1772 12887
rect 1856 12711 1890 12887
rect 1444 12427 1478 12461
rect 1562 12427 1596 12461
rect 1139 12342 1195 12386
rect 1717 12304 1769 12350
rect 1481 10915 1541 10977
rect 1140 10563 1174 10739
rect 1258 10563 1292 10739
rect 1376 10563 1410 10739
rect 1494 10563 1528 10739
rect 1612 10563 1646 10739
rect 1730 10563 1764 10739
rect 1848 10563 1882 10739
rect 1966 10563 2000 10739
rect 2084 10563 2118 10739
rect 2202 10563 2236 10739
rect 1907 10469 1941 10503
rect 1789 10352 1823 10386
rect 1377 9926 1411 10302
rect 1495 9926 1529 10302
rect 1613 9926 1647 10302
rect 1730 10126 1764 10302
rect 1848 10126 1882 10302
rect 1436 9842 1470 9876
rect 1554 9842 1588 9876
rect 1709 9719 1761 9765
rect 1462 7637 1522 7699
rect 1121 7285 1155 7461
rect 1239 7285 1273 7461
rect 1357 7285 1391 7461
rect 1475 7285 1509 7461
rect 1593 7285 1627 7461
rect 1711 7285 1745 7461
rect 1829 7285 1863 7461
rect 1947 7285 1981 7461
rect 2065 7285 2099 7461
rect 2183 7285 2217 7461
rect 1888 7191 1922 7225
rect 1770 7074 1804 7108
rect 1358 6648 1392 7024
rect 1476 6648 1510 7024
rect 1594 6648 1628 7024
rect 1711 6848 1745 7024
rect 1829 6848 1863 7024
rect 1417 6564 1451 6598
rect 1535 6564 1569 6598
rect 1083 6474 1143 6527
rect 1690 6441 1742 6487
rect 1478 4877 1538 4939
rect 1137 4525 1171 4701
rect 1255 4525 1289 4701
rect 1373 4525 1407 4701
rect 1491 4525 1525 4701
rect 1609 4525 1643 4701
rect 1727 4525 1761 4701
rect 1845 4525 1879 4701
rect 1963 4525 1997 4701
rect 2081 4525 2115 4701
rect 2199 4525 2233 4701
rect 1904 4431 1938 4465
rect 1786 4314 1820 4348
rect 1374 3888 1408 4264
rect 1492 3888 1526 4264
rect 1610 3888 1644 4264
rect 1727 4088 1761 4264
rect 1845 4088 1879 4264
rect 1433 3804 1467 3838
rect 1551 3804 1585 3838
rect 1706 3681 1758 3727
rect 619 567 763 633
rect 204 422 318 493
rect 4513 13471 4580 13472
rect 4513 13323 4579 13471
rect 4579 13323 4580 13471
rect 6995 13376 7061 13522
rect 7061 13376 7062 13522
rect 6995 13373 7062 13376
rect 6248 13271 6282 13305
rect 8137 13376 8141 13524
rect 8141 13376 8204 13524
rect 8137 13375 8204 13376
rect 7378 13277 7412 13311
rect 11062 13559 11129 13560
rect 11062 13411 11128 13559
rect 11128 13411 11129 13559
rect 13545 13464 13610 13611
rect 13610 13464 13612 13611
rect 13545 13462 13612 13464
rect 12797 13359 12831 13393
rect 14689 13464 14690 13613
rect 14690 13464 14756 13613
rect 13927 13365 13961 13399
rect 17715 13342 17782 13490
rect 17715 13341 17782 13342
rect 20196 13545 20263 13546
rect 20196 13397 20197 13545
rect 20197 13397 20263 13545
rect 12797 13241 12831 13275
rect 6248 13153 6282 13187
rect 7378 13157 7412 13191
rect 13927 13245 13961 13279
rect 4038 12881 4072 13057
rect 4156 12881 4190 13057
rect 4274 12881 4308 13057
rect 4392 12881 4426 13057
rect 4510 12881 4544 13057
rect 4628 12881 4662 13057
rect 4746 12881 4780 13057
rect 4864 12881 4898 13057
rect 4982 12881 5016 13057
rect 5100 12881 5134 13057
rect 4805 12787 4839 12821
rect 6363 12753 6397 13129
rect 6481 12753 6515 13129
rect 6599 12753 6633 13129
rect 6717 12753 6751 13129
rect 6835 12753 6869 13129
rect 6953 12753 6987 13129
rect 7071 12753 7105 13129
rect 7505 12757 7539 13133
rect 7623 12757 7657 13133
rect 7741 12757 7775 13133
rect 7859 12757 7893 13133
rect 7977 12757 8011 13133
rect 8095 12757 8129 13133
rect 8213 12757 8247 13133
rect 10587 12969 10621 13145
rect 10705 12969 10739 13145
rect 10823 12969 10857 13145
rect 10941 12969 10975 13145
rect 11059 12969 11093 13145
rect 11177 12969 11211 13145
rect 11295 12969 11329 13145
rect 11413 12969 11447 13145
rect 11531 12969 11565 13145
rect 11649 12969 11683 13145
rect 11354 12875 11388 12909
rect 12912 12841 12946 13217
rect 13030 12841 13064 13217
rect 13148 12841 13182 13217
rect 13266 12841 13300 13217
rect 13384 12841 13418 13217
rect 13502 12841 13536 13217
rect 13620 12841 13654 13217
rect 14054 12845 14088 13221
rect 14172 12845 14206 13221
rect 14290 12845 14324 13221
rect 14408 12845 14442 13221
rect 14526 12845 14560 13221
rect 14644 12845 14678 13221
rect 19451 13291 19485 13325
rect 21343 13396 21344 13545
rect 21344 13396 21410 13545
rect 20581 13297 20615 13331
rect 24335 13410 24340 13559
rect 24340 13410 24402 13559
rect 26819 13464 26822 13611
rect 26822 13464 26886 13611
rect 26819 13462 26886 13464
rect 26076 13359 26110 13393
rect 27968 13613 28035 13617
rect 27968 13468 27969 13613
rect 27969 13468 28035 13613
rect 27206 13365 27240 13399
rect 26076 13241 26110 13275
rect 14762 12845 14796 13221
rect 19451 13173 19485 13207
rect 20581 13177 20615 13211
rect 17241 12901 17275 13077
rect 17359 12901 17393 13077
rect 17477 12901 17511 13077
rect 17595 12901 17629 13077
rect 17713 12901 17747 13077
rect 17831 12901 17865 13077
rect 17949 12901 17983 13077
rect 18067 12901 18101 13077
rect 18185 12901 18219 13077
rect 18303 12901 18337 13077
rect 18008 12807 18042 12841
rect 11236 12758 11270 12792
rect 19566 12773 19600 13149
rect 19684 12773 19718 13149
rect 19802 12773 19836 13149
rect 19920 12773 19954 13149
rect 20038 12773 20072 13149
rect 20156 12773 20190 13149
rect 27206 13245 27240 13279
rect 20274 12773 20308 13149
rect 20708 12777 20742 13153
rect 20826 12777 20860 13153
rect 20944 12777 20978 13153
rect 21062 12777 21096 13153
rect 21180 12777 21214 13153
rect 21298 12777 21332 13153
rect 21416 12777 21450 13153
rect 23866 12969 23900 13145
rect 23984 12969 24018 13145
rect 24102 12969 24136 13145
rect 24220 12969 24254 13145
rect 24338 12969 24372 13145
rect 24456 12969 24490 13145
rect 24574 12969 24608 13145
rect 24692 12969 24726 13145
rect 24810 12969 24844 13145
rect 24928 12969 24962 13145
rect 24633 12875 24667 12909
rect 26191 12841 26225 13217
rect 26309 12841 26343 13217
rect 26427 12841 26461 13217
rect 26545 12841 26579 13217
rect 26663 12841 26697 13217
rect 26781 12841 26815 13217
rect 26899 12841 26933 13217
rect 27333 12845 27367 13221
rect 27451 12845 27485 13221
rect 27569 12845 27603 13221
rect 27687 12845 27721 13221
rect 27805 12845 27839 13221
rect 27923 12845 27957 13221
rect 28041 12845 28075 13221
rect 24515 12758 24549 12792
rect 4687 12670 4721 12704
rect 4275 12244 4309 12620
rect 4393 12244 4427 12620
rect 4511 12244 4545 12620
rect 4628 12444 4662 12620
rect 4746 12444 4780 12620
rect 6568 12397 6602 12431
rect 7710 12401 7744 12435
rect 4854 12216 5003 12283
rect 4334 12160 4368 12194
rect 4452 12160 4486 12194
rect 6273 12170 6307 12346
rect 6391 12170 6425 12346
rect 6509 12170 6543 12346
rect 6627 12170 6661 12346
rect 6792 12170 6826 12346
rect 6910 12170 6944 12346
rect 7028 12170 7062 12346
rect 7146 12170 7180 12346
rect 7415 12174 7449 12350
rect 7533 12174 7567 12350
rect 7651 12174 7685 12350
rect 7769 12174 7803 12350
rect 7934 12174 7968 12350
rect 8052 12174 8086 12350
rect 8170 12174 8204 12350
rect 8288 12174 8322 12350
rect 10824 12332 10858 12708
rect 10942 12332 10976 12708
rect 11060 12332 11094 12708
rect 11177 12532 11211 12708
rect 11295 12532 11329 12708
rect 17890 12690 17924 12724
rect 13117 12485 13151 12519
rect 14259 12489 14293 12523
rect 11400 12298 11549 12365
rect 10883 12248 10917 12282
rect 11001 12248 11035 12282
rect 12822 12258 12856 12434
rect 12940 12258 12974 12434
rect 13058 12258 13092 12434
rect 13176 12258 13210 12434
rect 13341 12258 13375 12434
rect 13459 12258 13493 12434
rect 13577 12258 13611 12434
rect 13695 12258 13729 12434
rect 13964 12262 13998 12438
rect 14082 12262 14116 12438
rect 14200 12262 14234 12438
rect 14318 12262 14352 12438
rect 14483 12262 14517 12438
rect 14601 12262 14635 12438
rect 14719 12262 14753 12438
rect 14837 12262 14871 12438
rect 17478 12264 17512 12640
rect 17596 12264 17630 12640
rect 17714 12264 17748 12640
rect 17831 12464 17865 12640
rect 17949 12464 17983 12640
rect 19771 12417 19805 12451
rect 20913 12421 20947 12455
rect 18050 12232 18199 12299
rect 17537 12180 17571 12214
rect 17655 12180 17689 12214
rect 19476 12190 19510 12366
rect 19594 12190 19628 12366
rect 19712 12190 19746 12366
rect 19830 12190 19864 12366
rect 19995 12190 20029 12366
rect 20113 12190 20147 12366
rect 20231 12190 20265 12366
rect 20349 12190 20383 12366
rect 20618 12194 20652 12370
rect 20736 12194 20770 12370
rect 20854 12194 20888 12370
rect 20972 12194 21006 12370
rect 21137 12194 21171 12370
rect 21255 12194 21289 12370
rect 21373 12194 21407 12370
rect 21491 12194 21525 12370
rect 24103 12332 24137 12708
rect 24221 12332 24255 12708
rect 24339 12332 24373 12708
rect 24456 12532 24490 12708
rect 24574 12532 24608 12708
rect 30004 12682 30064 12744
rect 26396 12485 26430 12519
rect 27538 12489 27572 12523
rect 24682 12308 24831 12375
rect 24162 12248 24196 12282
rect 24280 12248 24314 12282
rect 26101 12258 26135 12434
rect 26219 12258 26253 12434
rect 26337 12258 26371 12434
rect 26455 12258 26489 12434
rect 26620 12258 26654 12434
rect 26738 12258 26772 12434
rect 26856 12258 26890 12434
rect 26974 12258 27008 12434
rect 27243 12262 27277 12438
rect 27361 12262 27395 12438
rect 27479 12262 27513 12438
rect 27597 12262 27631 12438
rect 27762 12262 27796 12438
rect 27880 12262 27914 12438
rect 27998 12262 28032 12438
rect 28116 12262 28150 12438
rect 29663 12330 29697 12506
rect 29781 12330 29815 12506
rect 29899 12330 29933 12506
rect 30017 12330 30051 12506
rect 30135 12330 30169 12506
rect 30253 12330 30287 12506
rect 30371 12330 30405 12506
rect 30489 12330 30523 12506
rect 30607 12330 30641 12506
rect 30725 12330 30759 12506
rect 30430 12236 30464 12270
rect 30312 12119 30346 12153
rect 4525 11672 4526 11821
rect 4526 11672 4592 11821
rect 6340 11763 6407 11912
rect 7478 11765 7545 11914
rect 11076 11760 11142 11908
rect 11142 11760 11143 11908
rect 11076 11759 11143 11760
rect 12885 11859 12952 12008
rect 14024 11851 14091 12000
rect 17730 11841 17797 11842
rect 17730 11693 17796 11841
rect 17796 11693 17797 11841
rect 19538 11787 19605 11936
rect 20684 11790 20751 11939
rect 24358 11760 24421 11908
rect 24421 11760 24425 11908
rect 24358 11759 24425 11760
rect 26159 11848 26226 11995
rect 26159 11846 26226 11848
rect 27302 11848 27369 11997
rect 4052 11231 4086 11407
rect 4170 11231 4204 11407
rect 4288 11231 4322 11407
rect 4406 11231 4440 11407
rect 4524 11231 4558 11407
rect 4642 11231 4676 11407
rect 4760 11231 4794 11407
rect 4878 11231 4912 11407
rect 4996 11231 5030 11407
rect 5114 11231 5148 11407
rect 8237 11478 8304 11479
rect 8237 11330 8304 11478
rect 10601 11319 10635 11495
rect 10719 11319 10753 11495
rect 10837 11319 10871 11495
rect 10955 11319 10989 11495
rect 11073 11319 11107 11495
rect 11191 11319 11225 11495
rect 11309 11319 11343 11495
rect 11427 11319 11461 11495
rect 11545 11319 11579 11495
rect 11663 11319 11697 11495
rect 29900 11693 29934 12069
rect 30018 11693 30052 12069
rect 30136 11693 30170 12069
rect 30253 11893 30287 12069
rect 30371 11893 30405 12069
rect 14791 11417 14853 11566
rect 14853 11417 14858 11566
rect 11368 11225 11402 11259
rect 17255 11251 17289 11427
rect 17373 11251 17407 11427
rect 17491 11251 17525 11427
rect 17609 11251 17643 11427
rect 17727 11251 17761 11427
rect 17845 11251 17879 11427
rect 17963 11251 17997 11427
rect 18081 11251 18115 11427
rect 18199 11251 18233 11427
rect 18317 11251 18351 11427
rect 21437 11349 21440 11494
rect 21440 11349 21504 11494
rect 21437 11345 21504 11349
rect 23880 11319 23914 11495
rect 23998 11319 24032 11495
rect 24116 11319 24150 11495
rect 24234 11319 24268 11495
rect 24352 11319 24386 11495
rect 24470 11319 24504 11495
rect 24588 11319 24622 11495
rect 24706 11319 24740 11495
rect 24824 11319 24858 11495
rect 24942 11319 24976 11495
rect 29959 11609 29993 11643
rect 30077 11609 30111 11643
rect 28065 11417 28132 11563
rect 28065 11414 28132 11417
rect 30232 11486 30284 11532
rect 24647 11225 24681 11259
rect 4819 11137 4853 11171
rect 11250 11108 11284 11142
rect 4701 11020 4735 11054
rect 3250 10491 3368 10601
rect 4289 10594 4323 10970
rect 4407 10594 4441 10970
rect 4525 10594 4559 10970
rect 4642 10794 4676 10970
rect 4760 10794 4794 10970
rect 4869 10566 5018 10633
rect 5516 10614 5550 10790
rect 5634 10614 5668 10790
rect 5752 10614 5786 10790
rect 5870 10614 5904 10790
rect 6000 10614 6034 10990
rect 6118 10614 6152 10990
rect 6236 10614 6270 10990
rect 6354 10614 6388 10990
rect 6472 10614 6506 10990
rect 6590 10614 6624 10990
rect 6708 10614 6742 10990
rect 6837 10614 6871 10790
rect 6955 10614 6989 10790
rect 7073 10614 7107 10790
rect 7191 10614 7225 10790
rect 7414 10614 7448 10790
rect 7532 10614 7566 10790
rect 7650 10614 7684 10790
rect 7768 10614 7802 10790
rect 7898 10614 7932 10990
rect 8016 10614 8050 10990
rect 8134 10614 8168 10990
rect 8252 10614 8286 10990
rect 8370 10614 8404 10990
rect 8488 10614 8522 10990
rect 8606 10614 8640 10990
rect 8735 10614 8769 10790
rect 8853 10614 8887 10790
rect 8971 10614 9005 10790
rect 9089 10614 9123 10790
rect 10838 10682 10872 11058
rect 10956 10682 10990 11058
rect 11074 10682 11108 11058
rect 11191 10882 11225 11058
rect 11309 10882 11343 11058
rect 11418 10648 11567 10715
rect 12065 10702 12099 10878
rect 12183 10702 12217 10878
rect 12301 10702 12335 10878
rect 12419 10702 12453 10878
rect 12549 10702 12583 11078
rect 12667 10702 12701 11078
rect 12785 10702 12819 11078
rect 12903 10702 12937 11078
rect 13021 10702 13055 11078
rect 18022 11157 18056 11191
rect 13139 10702 13173 11078
rect 13257 10702 13291 11078
rect 13386 10702 13420 10878
rect 13504 10702 13538 10878
rect 13622 10702 13656 10878
rect 13740 10702 13774 10878
rect 13963 10702 13997 10878
rect 14081 10702 14115 10878
rect 14199 10702 14233 10878
rect 14317 10702 14351 10878
rect 14447 10702 14481 11078
rect 14565 10702 14599 11078
rect 14683 10702 14717 11078
rect 14801 10702 14835 11078
rect 14919 10702 14953 11078
rect 24529 11108 24563 11142
rect 15037 10702 15071 11078
rect 15155 10702 15189 11078
rect 17904 11040 17938 11074
rect 15284 10702 15318 10878
rect 15402 10702 15436 10878
rect 15520 10702 15554 10878
rect 15638 10702 15672 10878
rect 10897 10598 10931 10632
rect 11015 10598 11049 10632
rect 4348 10510 4382 10544
rect 4466 10510 4500 10544
rect 16452 10513 16591 10630
rect 17492 10614 17526 10990
rect 17610 10614 17644 10990
rect 17728 10614 17762 10990
rect 17845 10814 17879 10990
rect 17963 10814 17997 10990
rect 18067 10581 18216 10648
rect 18719 10634 18753 10810
rect 18837 10634 18871 10810
rect 18955 10634 18989 10810
rect 19073 10634 19107 10810
rect 19203 10634 19237 11010
rect 19321 10634 19355 11010
rect 19439 10634 19473 11010
rect 19557 10634 19591 11010
rect 19675 10634 19709 11010
rect 19793 10634 19827 11010
rect 19911 10634 19945 11010
rect 20040 10634 20074 10810
rect 20158 10634 20192 10810
rect 20276 10634 20310 10810
rect 20394 10634 20428 10810
rect 20617 10634 20651 10810
rect 20735 10634 20769 10810
rect 20853 10634 20887 10810
rect 20971 10634 21005 10810
rect 21101 10634 21135 11010
rect 21219 10634 21253 11010
rect 21337 10634 21371 11010
rect 21455 10634 21489 11010
rect 21573 10634 21607 11010
rect 21691 10634 21725 11010
rect 21809 10634 21843 11010
rect 21938 10634 21972 10810
rect 22056 10634 22090 10810
rect 22174 10634 22208 10810
rect 22292 10634 22326 10810
rect 24117 10682 24151 11058
rect 24235 10682 24269 11058
rect 24353 10682 24387 11058
rect 24470 10882 24504 11058
rect 24588 10882 24622 11058
rect 24687 10647 24836 10714
rect 25344 10702 25378 10878
rect 25462 10702 25496 10878
rect 25580 10702 25614 10878
rect 25698 10702 25732 10878
rect 25828 10702 25862 11078
rect 25946 10702 25980 11078
rect 26064 10702 26098 11078
rect 26182 10702 26216 11078
rect 26300 10702 26334 11078
rect 26418 10702 26452 11078
rect 26536 10702 26570 11078
rect 26665 10702 26699 10878
rect 26783 10702 26817 10878
rect 26901 10702 26935 10878
rect 27019 10702 27053 10878
rect 27242 10702 27276 10878
rect 27360 10702 27394 10878
rect 27478 10702 27512 10878
rect 27596 10702 27630 10878
rect 27726 10702 27760 11078
rect 27844 10702 27878 11078
rect 27962 10702 27996 11078
rect 28080 10702 28114 11078
rect 28198 10702 28232 11078
rect 28316 10702 28350 11078
rect 28434 10702 28468 11078
rect 28563 10702 28597 10878
rect 28681 10702 28715 10878
rect 28799 10702 28833 10878
rect 28917 10702 28951 10878
rect 24176 10598 24210 10632
rect 24294 10598 24328 10632
rect 17551 10530 17585 10564
rect 17669 10530 17703 10564
rect 13529 10430 13563 10464
rect 15636 10409 15670 10443
rect 6980 10342 7014 10376
rect 9087 10321 9121 10355
rect 4523 10068 4588 10215
rect 4588 10068 4590 10215
rect 4523 10066 4590 10068
rect 5943 9921 5977 10297
rect 6061 9921 6095 10297
rect 4047 9627 4081 9803
rect 4165 9627 4199 9803
rect 4283 9627 4317 9803
rect 4401 9627 4435 9803
rect 4519 9627 4553 9803
rect 4637 9627 4671 9803
rect 4755 9627 4789 9803
rect 4873 9627 4907 9803
rect 4991 9627 5025 9803
rect 6179 9921 6213 10297
rect 6297 9921 6331 10297
rect 6415 9921 6449 10297
rect 6533 9921 6567 10297
rect 6651 9921 6685 10297
rect 7841 9921 7875 10297
rect 7959 9921 7993 10297
rect 8077 9921 8111 10297
rect 8195 9921 8229 10297
rect 8313 9921 8347 10297
rect 8431 9921 8465 10297
rect 8549 9921 8583 10297
rect 11068 10305 11135 10308
rect 11068 10159 11070 10305
rect 11070 10159 11135 10305
rect 12492 10009 12526 10385
rect 12610 10009 12644 10385
rect 5109 9627 5143 9803
rect 5973 9699 6007 9733
rect 5788 9632 5822 9666
rect 6621 9699 6655 9733
rect 7871 9699 7905 9733
rect 6239 9615 6273 9649
rect 6357 9616 6391 9650
rect 6911 9631 6945 9665
rect 7686 9632 7720 9666
rect 8517 9700 8551 9734
rect 8137 9615 8171 9649
rect 8255 9616 8289 9650
rect 8809 9631 8843 9665
rect 4814 9533 4848 9567
rect 4696 9416 4730 9450
rect 5641 9389 5675 9565
rect 4284 8990 4318 9366
rect 4402 8990 4436 9366
rect 4520 8990 4554 9366
rect 4637 9190 4671 9366
rect 5759 9389 5793 9565
rect 4755 9190 4789 9366
rect 6061 9189 6095 9565
rect 6179 9189 6213 9565
rect 6297 9189 6331 9565
rect 6415 9189 6449 9565
rect 6533 9189 6567 9565
rect 6939 9389 6973 9565
rect 7057 9389 7091 9565
rect 7539 9389 7573 9565
rect 7657 9389 7691 9565
rect 7959 9189 7993 9565
rect 8077 9189 8111 9565
rect 8195 9189 8229 9565
rect 8313 9189 8347 9565
rect 8431 9189 8465 9565
rect 8837 9389 8871 9565
rect 8955 9389 8989 9565
rect 4867 8958 5016 9025
rect 4343 8906 4377 8940
rect 4461 8906 4495 8940
rect 6280 8723 6347 8872
rect 10596 9715 10630 9891
rect 10714 9715 10748 9891
rect 10832 9715 10866 9891
rect 10950 9715 10984 9891
rect 11068 9715 11102 9891
rect 11186 9715 11220 9891
rect 11304 9715 11338 9891
rect 11422 9715 11456 9891
rect 11540 9715 11574 9891
rect 12728 10009 12762 10385
rect 12846 10009 12880 10385
rect 12964 10009 12998 10385
rect 13082 10009 13116 10385
rect 13200 10009 13234 10385
rect 14390 10009 14424 10385
rect 14508 10009 14542 10385
rect 14626 10009 14660 10385
rect 14744 10009 14778 10385
rect 14862 10009 14896 10385
rect 14980 10009 15014 10385
rect 15098 10009 15132 10385
rect 11658 9715 11692 9891
rect 12522 9787 12556 9821
rect 12337 9720 12371 9754
rect 13170 9787 13204 9821
rect 14420 9787 14454 9821
rect 12788 9703 12822 9737
rect 12906 9704 12940 9738
rect 13460 9719 13494 9753
rect 14235 9720 14269 9754
rect 15759 9882 15891 9980
rect 15066 9788 15100 9822
rect 14686 9703 14720 9737
rect 14804 9704 14838 9738
rect 15358 9719 15392 9753
rect 11363 9621 11397 9655
rect 11245 9504 11279 9538
rect 12190 9477 12224 9653
rect 10833 9078 10867 9454
rect 10951 9078 10985 9454
rect 11069 9078 11103 9454
rect 11186 9278 11220 9454
rect 12308 9477 12342 9653
rect 11304 9278 11338 9454
rect 12610 9277 12644 9653
rect 12728 9277 12762 9653
rect 12846 9277 12880 9653
rect 12964 9277 12998 9653
rect 13082 9277 13116 9653
rect 13488 9477 13522 9653
rect 13606 9477 13640 9653
rect 14088 9477 14122 9653
rect 14206 9477 14240 9653
rect 14508 9277 14542 9653
rect 14626 9277 14660 9653
rect 14744 9277 14778 9653
rect 14862 9277 14896 9653
rect 14980 9277 15014 9653
rect 15386 9477 15420 9653
rect 15504 9477 15538 9653
rect 11415 9047 11564 9114
rect 10892 8994 10926 9028
rect 11010 8994 11044 9028
rect 12829 8808 12896 8957
rect 26808 10430 26842 10464
rect 28915 10409 28949 10443
rect 20183 10362 20217 10396
rect 22290 10341 22324 10375
rect 17725 10237 17792 10239
rect 17725 10090 17791 10237
rect 17791 10090 17792 10237
rect 19146 9941 19180 10317
rect 19264 9941 19298 10317
rect 17250 9647 17284 9823
rect 17368 9647 17402 9823
rect 17486 9647 17520 9823
rect 17604 9647 17638 9823
rect 17722 9647 17756 9823
rect 17840 9647 17874 9823
rect 17958 9647 17992 9823
rect 18076 9647 18110 9823
rect 18194 9647 18228 9823
rect 19382 9941 19416 10317
rect 19500 9941 19534 10317
rect 19618 9941 19652 10317
rect 19736 9941 19770 10317
rect 19854 9941 19888 10317
rect 21044 9941 21078 10317
rect 21162 9941 21196 10317
rect 21280 9941 21314 10317
rect 21398 9941 21432 10317
rect 21516 9941 21550 10317
rect 21634 9941 21668 10317
rect 21752 9941 21786 10317
rect 24350 10156 24416 10300
rect 24416 10156 24417 10300
rect 24350 10151 24417 10156
rect 25771 10009 25805 10385
rect 25889 10009 25923 10385
rect 18312 9647 18346 9823
rect 19176 9719 19210 9753
rect 18991 9652 19025 9686
rect 19824 9719 19858 9753
rect 21074 9719 21108 9753
rect 19442 9635 19476 9669
rect 19560 9636 19594 9670
rect 20114 9651 20148 9685
rect 20889 9652 20923 9686
rect 22874 9811 22970 9911
rect 21720 9720 21754 9754
rect 23875 9715 23909 9891
rect 23993 9715 24027 9891
rect 24111 9715 24145 9891
rect 24229 9715 24263 9891
rect 24347 9715 24381 9891
rect 24465 9715 24499 9891
rect 24583 9715 24617 9891
rect 24701 9715 24735 9891
rect 24819 9715 24853 9891
rect 26007 10009 26041 10385
rect 26125 10009 26159 10385
rect 26243 10009 26277 10385
rect 26361 10009 26395 10385
rect 26479 10009 26513 10385
rect 27669 10009 27703 10385
rect 27787 10009 27821 10385
rect 27905 10009 27939 10385
rect 28023 10009 28057 10385
rect 28141 10009 28175 10385
rect 28259 10009 28293 10385
rect 28377 10009 28411 10385
rect 24937 9715 24971 9891
rect 25801 9787 25835 9821
rect 25616 9720 25650 9754
rect 21340 9635 21374 9669
rect 21458 9636 21492 9670
rect 22012 9651 22046 9685
rect 26449 9787 26483 9821
rect 27699 9787 27733 9821
rect 26067 9703 26101 9737
rect 26185 9704 26219 9738
rect 26739 9719 26773 9753
rect 27514 9720 27548 9754
rect 29038 9882 29170 9980
rect 28345 9788 28379 9822
rect 27965 9703 27999 9737
rect 28083 9704 28117 9738
rect 28637 9719 28671 9753
rect 24642 9621 24676 9655
rect 18017 9553 18051 9587
rect 17899 9436 17933 9470
rect 18844 9409 18878 9585
rect 17487 9010 17521 9386
rect 17605 9010 17639 9386
rect 17723 9010 17757 9386
rect 17840 9210 17874 9386
rect 18962 9409 18996 9585
rect 17958 9210 17992 9386
rect 19264 9209 19298 9585
rect 19382 9209 19416 9585
rect 19500 9209 19534 9585
rect 19618 9209 19652 9585
rect 19736 9209 19770 9585
rect 20142 9409 20176 9585
rect 20260 9409 20294 9585
rect 20742 9409 20776 9585
rect 20860 9409 20894 9585
rect 21162 9209 21196 9585
rect 21280 9209 21314 9585
rect 21398 9209 21432 9585
rect 21516 9209 21550 9585
rect 21634 9209 21668 9585
rect 22040 9409 22074 9585
rect 22158 9409 22192 9585
rect 24524 9504 24558 9538
rect 25469 9477 25503 9653
rect 24112 9078 24146 9454
rect 24230 9078 24264 9454
rect 24348 9078 24382 9454
rect 24465 9278 24499 9454
rect 25587 9477 25621 9653
rect 24583 9278 24617 9454
rect 25889 9277 25923 9653
rect 26007 9277 26041 9653
rect 26125 9277 26159 9653
rect 26243 9277 26277 9653
rect 26361 9277 26395 9653
rect 26767 9477 26801 9653
rect 26885 9477 26919 9653
rect 27367 9477 27401 9653
rect 27485 9477 27519 9653
rect 27787 9277 27821 9653
rect 27905 9277 27939 9653
rect 28023 9277 28057 9653
rect 28141 9277 28175 9653
rect 28259 9277 28293 9653
rect 28665 9477 28699 9653
rect 28783 9477 28817 9653
rect 30004 9649 30064 9711
rect 29663 9297 29697 9473
rect 29781 9297 29815 9473
rect 29899 9297 29933 9473
rect 30017 9297 30051 9473
rect 30135 9297 30169 9473
rect 30253 9297 30287 9473
rect 30371 9297 30405 9473
rect 30489 9297 30523 9473
rect 30607 9297 30641 9473
rect 30725 9297 30759 9473
rect 30430 9203 30464 9237
rect 18069 8976 18218 9043
rect 24693 9042 24842 9109
rect 30312 9086 30346 9120
rect 24171 8994 24205 9028
rect 24289 8994 24323 9028
rect 17546 8926 17580 8960
rect 17664 8926 17698 8960
rect 19478 8742 19545 8891
rect 26109 8808 26176 8957
rect 29900 8660 29934 9036
rect 30018 8660 30052 9036
rect 30136 8660 30170 9036
rect 30253 8860 30287 9036
rect 30371 8860 30405 9036
rect 16431 8497 16501 8565
rect 22414 8491 22520 8590
rect 23523 8491 23629 8590
rect 29959 8576 29993 8610
rect 30077 8576 30111 8610
rect 30232 8453 30284 8499
rect 31903 13803 31937 14179
rect 32021 13803 32055 14179
rect 32139 13803 32173 14179
rect 32257 13803 32291 14179
rect 32375 13803 32409 14179
rect 32493 13803 32527 14179
rect 32611 13803 32645 14179
rect 32777 13883 32839 13974
rect 33506 13856 33540 14232
rect 33624 13856 33658 14232
rect 33742 13856 33776 14232
rect 33859 14056 33893 14232
rect 33977 14056 34011 14232
rect 37737 18962 37797 19011
rect 36963 18838 37139 18872
rect 36963 18720 37139 18754
rect 36963 18602 37139 18636
rect 37454 18709 37509 18767
rect 37454 18707 37509 18709
rect 36963 18484 37139 18518
rect 36763 18397 37139 18431
rect 36763 18279 37139 18313
rect 36763 18161 37139 18195
rect 36763 18043 37139 18077
rect 36763 17930 37139 17964
rect 38096 18004 38272 18038
rect 38096 17886 38272 17920
rect 36763 17812 37139 17846
rect 36763 17694 37139 17728
rect 36513 17548 36567 17620
rect 38096 17812 38472 17846
rect 37354 17752 37388 17786
rect 37738 17798 37793 17800
rect 37738 17740 37793 17798
rect 36763 17576 37139 17610
rect 38096 17694 38472 17728
rect 37453 17680 37508 17682
rect 37453 17622 37508 17680
rect 38096 17576 38472 17610
rect 36763 17458 37139 17492
rect 38573 17575 38607 17609
rect 37974 17517 38008 17551
rect 38725 17548 38739 17606
rect 38739 17548 38771 17606
rect 38096 17458 38472 17492
rect 37584 17398 37618 17432
rect 36763 17340 37139 17374
rect 38096 17340 38472 17374
rect 36763 17222 37139 17256
rect 38096 17262 38272 17296
rect 38096 17144 38272 17178
rect 36763 17103 37139 17137
rect 36763 16985 37139 17019
rect 36763 16867 37139 16901
rect 36763 16749 37139 16783
rect 36963 16630 37139 16664
rect 36963 16512 37139 16546
rect 36963 16394 37139 16428
rect 37313 16442 37347 16476
rect 36963 16276 37139 16310
rect 36963 15694 37139 15728
rect 36963 15576 37139 15610
rect 36963 15458 37139 15492
rect 37454 15565 37509 15623
rect 37454 15563 37509 15565
rect 36963 15340 37139 15374
rect 36763 15253 37139 15287
rect 36763 15135 37139 15169
rect 36763 15017 37139 15051
rect 36763 14899 37139 14933
rect 36763 14786 37139 14820
rect 38096 14860 38272 14894
rect 38096 14742 38272 14776
rect 36763 14668 37139 14702
rect 36763 14550 37139 14584
rect 36513 14404 36567 14476
rect 38096 14668 38472 14702
rect 37354 14608 37388 14642
rect 37738 14654 37793 14656
rect 37738 14596 37793 14654
rect 36763 14432 37139 14466
rect 38096 14550 38472 14584
rect 37453 14536 37508 14538
rect 37453 14478 37508 14536
rect 38096 14432 38472 14466
rect 36763 14314 37139 14348
rect 38573 14431 38607 14465
rect 37974 14373 38008 14407
rect 38725 14404 38739 14462
rect 38739 14404 38771 14462
rect 38096 14314 38472 14348
rect 37584 14254 37618 14288
rect 36763 14196 37139 14230
rect 38096 14196 38472 14230
rect 36763 14078 37139 14112
rect 38096 14118 38272 14152
rect 38096 14000 38272 14034
rect 34254 13883 34377 13977
rect 36763 13959 37139 13993
rect 36763 13841 37139 13875
rect 33565 13772 33599 13806
rect 33683 13772 33717 13806
rect 31933 13581 31967 13615
rect 31748 13514 31782 13548
rect 33838 13649 33890 13695
rect 36763 13723 37139 13757
rect 32581 13581 32615 13615
rect 36763 13605 37139 13639
rect 32199 13497 32233 13531
rect 32317 13498 32351 13532
rect 32871 13513 32905 13547
rect 36963 13486 37139 13520
rect 31601 13271 31635 13447
rect 31719 13271 31753 13447
rect 32021 13071 32055 13447
rect 32139 13071 32173 13447
rect 32257 13071 32291 13447
rect 32375 13071 32409 13447
rect 32493 13071 32527 13447
rect 32899 13271 32933 13447
rect 33017 13271 33051 13447
rect 36963 13368 37139 13402
rect 36963 13250 37139 13284
rect 37313 13298 37347 13332
rect 36963 13132 37139 13166
rect 32215 12798 32350 12900
rect 37741 12616 37801 12665
rect 32112 11285 32533 11319
rect 32112 11140 32175 11285
rect 32175 11140 32484 11285
rect 32484 11140 32533 11285
rect 32112 11119 32533 11140
rect 31478 10405 31512 10581
rect 31596 10405 31630 10581
rect 31714 10405 31748 10581
rect 31832 10405 31866 10581
rect 31962 10405 31996 10781
rect 32080 10405 32114 10781
rect 32198 10405 32232 10781
rect 32316 10405 32350 10781
rect 32434 10405 32468 10781
rect 32552 10405 32586 10781
rect 32670 10405 32704 10781
rect 33612 10754 33672 10816
rect 32799 10405 32833 10581
rect 32917 10405 32951 10581
rect 33035 10405 33069 10581
rect 33153 10405 33187 10581
rect 33271 10402 33305 10578
rect 33389 10402 33423 10578
rect 33507 10402 33541 10578
rect 33625 10402 33659 10578
rect 33743 10402 33777 10578
rect 33861 10402 33895 10578
rect 33979 10402 34013 10578
rect 34097 10402 34131 10578
rect 34215 10402 34249 10578
rect 34333 10402 34367 10578
rect 34038 10308 34072 10342
rect 33130 10189 33164 10223
rect 33920 10191 33954 10225
rect 31730 10070 31764 10104
rect 31905 9712 31939 10088
rect 32023 9712 32057 10088
rect 32141 9712 32175 10088
rect 32259 9712 32293 10088
rect 32377 9712 32411 10088
rect 32495 9712 32529 10088
rect 32613 9712 32647 10088
rect 32779 9792 32841 9883
rect 33508 9765 33542 10141
rect 33626 9765 33660 10141
rect 33744 9765 33778 10141
rect 33861 9965 33895 10141
rect 33979 9965 34013 10141
rect 34226 10060 34353 10131
rect 33567 9681 33601 9715
rect 33685 9681 33719 9715
rect 31935 9490 31969 9524
rect 31750 9423 31784 9457
rect 33840 9558 33892 9604
rect 32583 9490 32617 9524
rect 32201 9406 32235 9440
rect 32319 9407 32353 9441
rect 32873 9422 32907 9456
rect 31603 9180 31637 9356
rect 31721 9180 31755 9356
rect 32023 8980 32057 9356
rect 32141 8980 32175 9356
rect 32259 8980 32293 9356
rect 32377 8980 32411 9356
rect 32495 8980 32529 9356
rect 32901 9180 32935 9356
rect 33019 9180 33053 9356
rect 32217 8707 32352 8809
rect 4501 7691 4568 7692
rect 4501 7543 4504 7691
rect 4504 7543 4568 7691
rect 6981 7745 7048 7747
rect 6981 7598 6986 7745
rect 6986 7598 7048 7745
rect 6240 7491 6274 7525
rect 8137 7596 8200 7744
rect 8200 7596 8204 7744
rect 8137 7595 8204 7596
rect 7370 7497 7404 7531
rect 11056 7689 11123 7690
rect 11056 7541 11122 7689
rect 11122 7541 11123 7689
rect 13537 7594 13604 7743
rect 12791 7489 12825 7523
rect 14685 7594 14751 7743
rect 14751 7594 14752 7743
rect 13921 7495 13955 7529
rect 16430 7680 16500 7748
rect 6240 7373 6274 7407
rect 7370 7377 7404 7411
rect 4030 7101 4064 7277
rect 4148 7101 4182 7277
rect 4266 7101 4300 7277
rect 4384 7101 4418 7277
rect 4502 7101 4536 7277
rect 4620 7101 4654 7277
rect 4738 7101 4772 7277
rect 4856 7101 4890 7277
rect 4974 7101 5008 7277
rect 5092 7101 5126 7277
rect 4797 7007 4831 7041
rect 6355 6973 6389 7349
rect 6473 6973 6507 7349
rect 6591 6973 6625 7349
rect 6709 6973 6743 7349
rect 6827 6973 6861 7349
rect 6945 6973 6979 7349
rect 12791 7371 12825 7405
rect 7063 6973 7097 7349
rect 7497 6977 7531 7353
rect 7615 6977 7649 7353
rect 7733 6977 7767 7353
rect 7851 6977 7885 7353
rect 7969 6977 8003 7353
rect 8087 6977 8121 7353
rect 8205 6977 8239 7353
rect 13921 7375 13955 7409
rect 10581 7099 10615 7275
rect 10699 7099 10733 7275
rect 10817 7099 10851 7275
rect 10935 7099 10969 7275
rect 11053 7099 11087 7275
rect 11171 7099 11205 7275
rect 11289 7099 11323 7275
rect 11407 7099 11441 7275
rect 11525 7099 11559 7275
rect 11643 7099 11677 7275
rect 11348 7005 11382 7039
rect 12906 6971 12940 7347
rect 13024 6971 13058 7347
rect 13142 6971 13176 7347
rect 13260 6971 13294 7347
rect 13378 6971 13412 7347
rect 13496 6971 13530 7347
rect 13614 6971 13648 7347
rect 14048 6975 14082 7351
rect 14166 6975 14200 7351
rect 14284 6975 14318 7351
rect 14402 6975 14436 7351
rect 14520 6975 14554 7351
rect 14638 6975 14672 7351
rect 14756 6975 14790 7351
rect 17707 7541 17710 7687
rect 17710 7541 17774 7687
rect 17707 7538 17774 7541
rect 20192 7744 20259 7747
rect 20192 7598 20259 7744
rect 19446 7490 19480 7524
rect 21341 7595 21406 7744
rect 21406 7595 21408 7744
rect 20576 7496 20610 7530
rect 24331 7691 24398 7692
rect 24331 7543 24332 7691
rect 24332 7543 24398 7691
rect 26810 7596 26814 7740
rect 26814 7596 26877 7740
rect 26810 7591 26877 7596
rect 26068 7491 26102 7525
rect 27958 7745 28025 7746
rect 27958 7597 27961 7745
rect 27961 7597 28025 7745
rect 30075 7729 30135 7791
rect 27198 7497 27232 7531
rect 32112 7790 32533 7824
rect 32112 7645 32175 7790
rect 32175 7645 32484 7790
rect 32484 7645 32533 7790
rect 32112 7624 32533 7645
rect 19446 7372 19480 7406
rect 20576 7376 20610 7410
rect 4679 6890 4713 6924
rect 11230 6888 11264 6922
rect 4267 6464 4301 6840
rect 4385 6464 4419 6840
rect 4503 6464 4537 6840
rect 4620 6664 4654 6840
rect 4738 6664 4772 6840
rect 6560 6617 6594 6651
rect 7702 6621 7736 6655
rect 4844 6429 4993 6496
rect 4326 6380 4360 6414
rect 4444 6380 4478 6414
rect 6265 6390 6299 6566
rect 6383 6390 6417 6566
rect 6501 6390 6535 6566
rect 6619 6390 6653 6566
rect 6784 6390 6818 6566
rect 6902 6390 6936 6566
rect 7020 6390 7054 6566
rect 7138 6390 7172 6566
rect 7407 6394 7441 6570
rect 7525 6394 7559 6570
rect 7643 6394 7677 6570
rect 7761 6394 7795 6570
rect 7926 6394 7960 6570
rect 8044 6394 8078 6570
rect 8162 6394 8196 6570
rect 8280 6394 8314 6570
rect 10818 6462 10852 6838
rect 10936 6462 10970 6838
rect 11054 6462 11088 6838
rect 11171 6662 11205 6838
rect 11289 6662 11323 6838
rect 13111 6615 13145 6649
rect 14253 6619 14287 6653
rect 11394 6423 11543 6490
rect 10877 6378 10911 6412
rect 10995 6378 11029 6412
rect 12816 6388 12850 6564
rect 12934 6388 12968 6564
rect 13052 6388 13086 6564
rect 13170 6388 13204 6564
rect 13335 6388 13369 6564
rect 13453 6388 13487 6564
rect 13571 6388 13605 6564
rect 13689 6388 13723 6564
rect 13958 6392 13992 6568
rect 14076 6392 14110 6568
rect 14194 6392 14228 6568
rect 14312 6392 14346 6568
rect 14477 6392 14511 6568
rect 14595 6392 14629 6568
rect 14713 6392 14747 6568
rect 14831 6392 14865 6568
rect 4522 5892 4585 6039
rect 4585 5892 4589 6039
rect 4522 5890 4589 5892
rect 6321 5986 6388 6135
rect 7474 5981 7541 6130
rect 11067 6039 11134 6046
rect 11067 5897 11069 6039
rect 11069 5897 11134 6039
rect 12879 5983 12946 6132
rect 14020 5976 14087 6121
rect 14020 5972 14087 5976
rect 4044 5451 4078 5627
rect 4162 5451 4196 5627
rect 4280 5451 4314 5627
rect 4398 5451 4432 5627
rect 4516 5451 4550 5627
rect 4634 5451 4668 5627
rect 4752 5451 4786 5627
rect 4870 5451 4904 5627
rect 4988 5451 5022 5627
rect 5106 5451 5140 5627
rect 8228 5549 8229 5698
rect 8229 5549 8295 5698
rect 10595 5449 10629 5625
rect 10713 5449 10747 5625
rect 10831 5449 10865 5625
rect 10949 5449 10983 5625
rect 11067 5449 11101 5625
rect 11185 5449 11219 5625
rect 11303 5449 11337 5625
rect 11421 5449 11455 5625
rect 11539 5449 11573 5625
rect 11657 5449 11691 5625
rect 14784 5696 14851 5697
rect 14784 5548 14847 5696
rect 14847 5548 14851 5696
rect 4811 5357 4845 5391
rect 11362 5355 11396 5389
rect 4693 5240 4727 5274
rect 4281 4814 4315 5190
rect 4399 4814 4433 5190
rect 4517 4814 4551 5190
rect 4634 5014 4668 5190
rect 4752 5014 4786 5190
rect 4852 4779 5001 4846
rect 5508 4834 5542 5010
rect 5626 4834 5660 5010
rect 5744 4834 5778 5010
rect 5862 4834 5896 5010
rect 5992 4834 6026 5210
rect 6110 4834 6144 5210
rect 6228 4834 6262 5210
rect 6346 4834 6380 5210
rect 6464 4834 6498 5210
rect 6582 4834 6616 5210
rect 6700 4834 6734 5210
rect 6829 4834 6863 5010
rect 6947 4834 6981 5010
rect 7065 4834 7099 5010
rect 7183 4834 7217 5010
rect 7406 4834 7440 5010
rect 7524 4834 7558 5010
rect 7642 4834 7676 5010
rect 7760 4834 7794 5010
rect 7890 4834 7924 5210
rect 8008 4834 8042 5210
rect 8126 4834 8160 5210
rect 8244 4834 8278 5210
rect 8362 4834 8396 5210
rect 11244 5238 11278 5272
rect 8480 4834 8514 5210
rect 8598 4834 8632 5210
rect 8727 4834 8761 5010
rect 8845 4834 8879 5010
rect 8963 4834 8997 5010
rect 9081 4834 9115 5010
rect 10832 4812 10866 5188
rect 10950 4812 10984 5188
rect 11068 4812 11102 5188
rect 11185 5012 11219 5188
rect 11303 5012 11337 5188
rect 4340 4730 4374 4764
rect 4458 4730 4492 4764
rect 11410 4778 11559 4845
rect 12059 4832 12093 5008
rect 12177 4832 12211 5008
rect 12295 4832 12329 5008
rect 12413 4832 12447 5008
rect 12543 4832 12577 5208
rect 12661 4832 12695 5208
rect 12779 4832 12813 5208
rect 12897 4832 12931 5208
rect 13015 4832 13049 5208
rect 13133 4832 13167 5208
rect 13251 4832 13285 5208
rect 13380 4832 13414 5008
rect 13498 4832 13532 5008
rect 13616 4832 13650 5008
rect 13734 4832 13768 5008
rect 13957 4832 13991 5008
rect 14075 4832 14109 5008
rect 14193 4832 14227 5008
rect 14311 4832 14345 5008
rect 14441 4832 14475 5208
rect 14559 4832 14593 5208
rect 14677 4832 14711 5208
rect 14795 4832 14829 5208
rect 14913 4832 14947 5208
rect 15031 4832 15065 5208
rect 15149 4832 15183 5208
rect 15278 4832 15312 5008
rect 15396 4832 15430 5008
rect 15514 4832 15548 5008
rect 15632 4832 15666 5008
rect 10891 4728 10925 4762
rect 11009 4728 11043 4762
rect 6972 4562 7006 4596
rect 9079 4541 9113 4575
rect 13523 4560 13557 4594
rect 4511 4437 4578 4440
rect 4511 4291 4513 4437
rect 4513 4291 4578 4437
rect 5935 4141 5969 4517
rect 6053 4141 6087 4517
rect 4039 3847 4073 4023
rect 4157 3847 4191 4023
rect 4275 3847 4309 4023
rect 4393 3847 4427 4023
rect 4511 3847 4545 4023
rect 4629 3847 4663 4023
rect 4747 3847 4781 4023
rect 4865 3847 4899 4023
rect 4983 3847 5017 4023
rect 6171 4141 6205 4517
rect 6289 4141 6323 4517
rect 6407 4141 6441 4517
rect 6525 4141 6559 4517
rect 6643 4141 6677 4517
rect 7833 4141 7867 4517
rect 7951 4141 7985 4517
rect 8069 4141 8103 4517
rect 8187 4141 8221 4517
rect 8305 4141 8339 4517
rect 8423 4141 8457 4517
rect 15630 4539 15664 4573
rect 8541 4141 8575 4517
rect 11067 4286 11131 4435
rect 11131 4286 11134 4435
rect 12486 4139 12520 4515
rect 12604 4139 12638 4515
rect 5101 3847 5135 4023
rect 5965 3919 5999 3953
rect 5780 3852 5814 3886
rect 6613 3919 6647 3953
rect 7863 3919 7897 3953
rect 6231 3835 6265 3869
rect 6349 3836 6383 3870
rect 6903 3851 6937 3885
rect 7678 3852 7712 3886
rect 9202 4014 9334 4112
rect 8509 3920 8543 3954
rect 8129 3835 8163 3869
rect 8247 3836 8281 3870
rect 8801 3851 8835 3885
rect 10590 3845 10624 4021
rect 10708 3845 10742 4021
rect 10826 3845 10860 4021
rect 10944 3845 10978 4021
rect 11062 3845 11096 4021
rect 11180 3845 11214 4021
rect 11298 3845 11332 4021
rect 11416 3845 11450 4021
rect 11534 3845 11568 4021
rect 12722 4139 12756 4515
rect 12840 4139 12874 4515
rect 12958 4139 12992 4515
rect 13076 4139 13110 4515
rect 13194 4139 13228 4515
rect 14384 4139 14418 4515
rect 14502 4139 14536 4515
rect 14620 4139 14654 4515
rect 14738 4139 14772 4515
rect 14856 4139 14890 4515
rect 14974 4139 15008 4515
rect 15092 4139 15126 4515
rect 11652 3845 11686 4021
rect 12516 3917 12550 3951
rect 12331 3850 12365 3884
rect 4806 3753 4840 3787
rect 4688 3636 4722 3670
rect 5633 3609 5667 3785
rect 4276 3210 4310 3586
rect 4394 3210 4428 3586
rect 4512 3210 4546 3586
rect 4629 3410 4663 3586
rect 5751 3609 5785 3785
rect 4747 3410 4781 3586
rect 6053 3409 6087 3785
rect 6171 3409 6205 3785
rect 6289 3409 6323 3785
rect 6407 3409 6441 3785
rect 6525 3409 6559 3785
rect 6931 3609 6965 3785
rect 7049 3609 7083 3785
rect 7531 3609 7565 3785
rect 7649 3609 7683 3785
rect 7951 3409 7985 3785
rect 8069 3409 8103 3785
rect 8187 3409 8221 3785
rect 8305 3409 8339 3785
rect 8423 3409 8457 3785
rect 8829 3609 8863 3785
rect 13164 3917 13198 3951
rect 14414 3917 14448 3951
rect 12782 3833 12816 3867
rect 12900 3834 12934 3868
rect 13454 3849 13488 3883
rect 14229 3850 14263 3884
rect 15060 3918 15094 3952
rect 14680 3833 14714 3867
rect 14798 3834 14832 3868
rect 15352 3849 15386 3883
rect 8947 3609 8981 3785
rect 11357 3751 11391 3785
rect 11239 3634 11273 3668
rect 12184 3607 12218 3783
rect 4852 3187 5001 3254
rect 10827 3208 10861 3584
rect 10945 3208 10979 3584
rect 11063 3208 11097 3584
rect 11180 3408 11214 3584
rect 12302 3607 12336 3783
rect 11298 3408 11332 3584
rect 12604 3407 12638 3783
rect 12722 3407 12756 3783
rect 12840 3407 12874 3783
rect 12958 3407 12992 3783
rect 13076 3407 13110 3783
rect 13482 3607 13516 3783
rect 13600 3607 13634 3783
rect 14082 3607 14116 3783
rect 14200 3607 14234 3783
rect 14502 3407 14536 3783
rect 14620 3407 14654 3783
rect 14738 3407 14772 3783
rect 14856 3407 14890 3783
rect 14974 3407 15008 3783
rect 15380 3607 15414 3783
rect 15498 3607 15532 3783
rect 4335 3126 4369 3160
rect 4453 3126 4487 3160
rect 11399 3178 11548 3245
rect 10886 3124 10920 3158
rect 11004 3124 11038 3158
rect 6273 2937 6340 3086
rect 12821 2936 12888 3085
rect 17236 7100 17270 7276
rect 17354 7100 17388 7276
rect 17472 7100 17506 7276
rect 17590 7100 17624 7276
rect 17708 7100 17742 7276
rect 17826 7100 17860 7276
rect 17944 7100 17978 7276
rect 18062 7100 18096 7276
rect 18180 7100 18214 7276
rect 18298 7100 18332 7276
rect 18003 7006 18037 7040
rect 19561 6972 19595 7348
rect 19679 6972 19713 7348
rect 19797 6972 19831 7348
rect 19915 6972 19949 7348
rect 20033 6972 20067 7348
rect 20151 6972 20185 7348
rect 26068 7373 26102 7407
rect 20269 6972 20303 7348
rect 20703 6976 20737 7352
rect 20821 6976 20855 7352
rect 20939 6976 20973 7352
rect 21057 6976 21091 7352
rect 21175 6976 21209 7352
rect 21293 6976 21327 7352
rect 21411 6976 21445 7352
rect 27198 7377 27232 7411
rect 23858 7101 23892 7277
rect 23976 7101 24010 7277
rect 24094 7101 24128 7277
rect 24212 7101 24246 7277
rect 24330 7101 24364 7277
rect 24448 7101 24482 7277
rect 24566 7101 24600 7277
rect 24684 7101 24718 7277
rect 24802 7101 24836 7277
rect 24920 7101 24954 7277
rect 24625 7007 24659 7041
rect 26183 6973 26217 7349
rect 26301 6973 26335 7349
rect 26419 6973 26453 7349
rect 26537 6973 26571 7349
rect 26655 6973 26689 7349
rect 26773 6973 26807 7349
rect 29734 7377 29768 7553
rect 26891 6973 26925 7349
rect 27325 6977 27359 7353
rect 27443 6977 27477 7353
rect 27561 6977 27595 7353
rect 27679 6977 27713 7353
rect 27797 6977 27831 7353
rect 27915 6977 27949 7353
rect 29852 7377 29886 7553
rect 29970 7377 30004 7553
rect 30088 7377 30122 7553
rect 30206 7377 30240 7553
rect 30324 7377 30358 7553
rect 30442 7377 30476 7553
rect 30560 7377 30594 7553
rect 30678 7377 30712 7553
rect 30796 7377 30830 7553
rect 28033 6977 28067 7353
rect 30501 7283 30535 7317
rect 30383 7166 30417 7200
rect 17885 6889 17919 6923
rect 24507 6890 24541 6924
rect 17473 6463 17507 6839
rect 17591 6463 17625 6839
rect 17709 6463 17743 6839
rect 17826 6663 17860 6839
rect 17944 6663 17978 6839
rect 19766 6616 19800 6650
rect 20908 6620 20942 6654
rect 18055 6432 18204 6499
rect 17532 6379 17566 6413
rect 17650 6379 17684 6413
rect 19471 6389 19505 6565
rect 19589 6389 19623 6565
rect 19707 6389 19741 6565
rect 19825 6389 19859 6565
rect 19990 6389 20024 6565
rect 20108 6389 20142 6565
rect 20226 6389 20260 6565
rect 20344 6389 20378 6565
rect 20613 6393 20647 6569
rect 20731 6393 20765 6569
rect 20849 6393 20883 6569
rect 20967 6393 21001 6569
rect 21132 6393 21166 6569
rect 21250 6393 21284 6569
rect 21368 6393 21402 6569
rect 21486 6393 21520 6569
rect 24095 6464 24129 6840
rect 24213 6464 24247 6840
rect 24331 6464 24365 6840
rect 24448 6664 24482 6840
rect 24566 6664 24600 6840
rect 29971 6740 30005 7116
rect 30089 6740 30123 7116
rect 30207 6740 30241 7116
rect 30324 6940 30358 7116
rect 30442 6940 30476 7116
rect 31478 6910 31512 7086
rect 31596 6910 31630 7086
rect 31714 6910 31748 7086
rect 31832 6910 31866 7086
rect 31962 6910 31996 7286
rect 32080 6910 32114 7286
rect 32198 6910 32232 7286
rect 32316 6910 32350 7286
rect 32434 6910 32468 7286
rect 32552 6910 32586 7286
rect 32670 6910 32704 7286
rect 33612 7259 33672 7321
rect 32799 6910 32833 7086
rect 32917 6910 32951 7086
rect 33035 6910 33069 7086
rect 33153 6910 33187 7086
rect 33271 6907 33305 7083
rect 33389 6907 33423 7083
rect 33507 6907 33541 7083
rect 33625 6907 33659 7083
rect 33743 6907 33777 7083
rect 33861 6907 33895 7083
rect 33979 6907 34013 7083
rect 34097 6907 34131 7083
rect 34215 6907 34249 7083
rect 34333 6907 34367 7083
rect 34038 6813 34072 6847
rect 33130 6694 33164 6728
rect 33920 6696 33954 6730
rect 30030 6656 30064 6690
rect 30148 6656 30182 6690
rect 26388 6617 26422 6651
rect 27530 6621 27564 6655
rect 24671 6437 24820 6504
rect 24154 6380 24188 6414
rect 24272 6380 24306 6414
rect 26093 6390 26127 6566
rect 26211 6390 26245 6566
rect 26329 6390 26363 6566
rect 26447 6390 26481 6566
rect 26612 6390 26646 6566
rect 26730 6390 26764 6566
rect 26848 6390 26882 6566
rect 26966 6390 27000 6566
rect 27235 6394 27269 6570
rect 27353 6394 27387 6570
rect 27471 6394 27505 6570
rect 27589 6394 27623 6570
rect 27754 6394 27788 6570
rect 27872 6394 27906 6570
rect 27990 6394 28024 6570
rect 28108 6394 28142 6570
rect 30303 6533 30355 6579
rect 31730 6575 31764 6609
rect 31905 6217 31939 6593
rect 32023 6217 32057 6593
rect 17727 6040 17794 6041
rect 17727 5892 17791 6040
rect 17791 5892 17794 6040
rect 19531 5987 19598 6136
rect 20677 5990 20744 6139
rect 24346 6041 24413 6042
rect 24346 5893 24413 6041
rect 26162 5991 26229 6140
rect 27296 5982 27363 6131
rect 32141 6217 32175 6593
rect 32259 6217 32293 6593
rect 32377 6217 32411 6593
rect 32495 6217 32529 6593
rect 32613 6217 32647 6593
rect 32779 6297 32841 6388
rect 33508 6270 33542 6646
rect 33626 6270 33660 6646
rect 33744 6270 33778 6646
rect 33861 6470 33895 6646
rect 33979 6470 34013 6646
rect 36967 12492 37143 12526
rect 36967 12374 37143 12408
rect 36967 12256 37143 12290
rect 37458 12363 37513 12421
rect 37458 12361 37513 12363
rect 36967 12138 37143 12172
rect 36767 12051 37143 12085
rect 36767 11933 37143 11967
rect 36767 11815 37143 11849
rect 36767 11697 37143 11731
rect 36767 11584 37143 11618
rect 38100 11658 38276 11692
rect 38100 11540 38276 11574
rect 36767 11466 37143 11500
rect 36767 11348 37143 11382
rect 36517 11202 36571 11274
rect 38100 11466 38476 11500
rect 37358 11406 37392 11440
rect 37742 11452 37797 11454
rect 37742 11394 37797 11452
rect 36767 11230 37143 11264
rect 38100 11348 38476 11382
rect 37457 11334 37512 11336
rect 37457 11276 37512 11334
rect 38100 11230 38476 11264
rect 36767 11112 37143 11146
rect 38577 11229 38611 11263
rect 37978 11171 38012 11205
rect 38729 11202 38743 11260
rect 38743 11202 38775 11260
rect 38100 11112 38476 11146
rect 37588 11052 37622 11086
rect 36767 10994 37143 11028
rect 38100 10994 38476 11028
rect 36767 10876 37143 10910
rect 38100 10916 38276 10950
rect 38100 10798 38276 10832
rect 36767 10757 37143 10791
rect 36767 10639 37143 10673
rect 36767 10521 37143 10555
rect 36767 10403 37143 10437
rect 36967 10284 37143 10318
rect 36967 10166 37143 10200
rect 36967 10048 37143 10082
rect 37317 10096 37351 10130
rect 36967 9930 37143 9964
rect 36967 9348 37143 9382
rect 36967 9230 37143 9264
rect 36967 9112 37143 9146
rect 37458 9219 37513 9277
rect 37458 9217 37513 9219
rect 36967 8994 37143 9028
rect 36767 8907 37143 8941
rect 36767 8789 37143 8823
rect 36767 8671 37143 8705
rect 36767 8553 37143 8587
rect 36767 8440 37143 8474
rect 38100 8514 38276 8548
rect 38100 8396 38276 8430
rect 36767 8322 37143 8356
rect 36767 8204 37143 8238
rect 36517 8058 36571 8130
rect 38100 8322 38476 8356
rect 37358 8262 37392 8296
rect 37742 8308 37797 8310
rect 37742 8250 37797 8308
rect 36767 8086 37143 8120
rect 38100 8204 38476 8238
rect 37457 8190 37512 8192
rect 37457 8132 37512 8190
rect 38100 8086 38476 8120
rect 36767 7968 37143 8002
rect 38577 8085 38611 8119
rect 37978 8027 38012 8061
rect 38729 8058 38743 8116
rect 38743 8058 38775 8116
rect 38100 7968 38476 8002
rect 37588 7908 37622 7942
rect 36767 7850 37143 7884
rect 38100 7850 38476 7884
rect 36767 7732 37143 7766
rect 38100 7772 38276 7806
rect 38100 7654 38276 7688
rect 36767 7613 37143 7647
rect 36767 7495 37143 7529
rect 36767 7377 37143 7411
rect 36767 7259 37143 7293
rect 36967 7140 37143 7174
rect 36967 7022 37143 7056
rect 36967 6904 37143 6938
rect 37317 6952 37351 6986
rect 36967 6786 37143 6820
rect 34662 6418 34728 6486
rect 34434 6303 34529 6375
rect 37737 6340 37797 6389
rect 33567 6186 33601 6220
rect 33685 6186 33719 6220
rect 36963 6216 37139 6250
rect 31935 5995 31969 6029
rect 31750 5928 31784 5962
rect 33840 6063 33892 6109
rect 32583 5995 32617 6029
rect 36963 6098 37139 6132
rect 36963 5980 37139 6014
rect 32201 5911 32235 5945
rect 32319 5912 32353 5946
rect 32873 5927 32907 5961
rect 37454 6087 37509 6145
rect 37454 6085 37509 6087
rect 17250 5450 17284 5626
rect 17368 5450 17402 5626
rect 17486 5450 17520 5626
rect 17604 5450 17638 5626
rect 17722 5450 17756 5626
rect 17840 5450 17874 5626
rect 17958 5450 17992 5626
rect 18076 5450 18110 5626
rect 18194 5450 18228 5626
rect 18312 5450 18346 5626
rect 21438 5697 21505 5699
rect 21438 5550 21502 5697
rect 21502 5550 21505 5697
rect 23872 5451 23906 5627
rect 23990 5451 24024 5627
rect 24108 5451 24142 5627
rect 24226 5451 24260 5627
rect 24344 5451 24378 5627
rect 24462 5451 24496 5627
rect 24580 5451 24614 5627
rect 24698 5451 24732 5627
rect 24816 5451 24850 5627
rect 24934 5451 24968 5627
rect 28059 5549 28124 5697
rect 28124 5549 28126 5697
rect 28059 5548 28126 5549
rect 31603 5685 31637 5861
rect 31721 5685 31755 5861
rect 32023 5485 32057 5861
rect 32141 5485 32175 5861
rect 32259 5485 32293 5861
rect 32377 5485 32411 5861
rect 32495 5485 32529 5861
rect 32901 5685 32935 5861
rect 36963 5862 37139 5896
rect 33019 5685 33053 5861
rect 36763 5775 37139 5809
rect 36763 5657 37139 5691
rect 36763 5539 37139 5573
rect 36763 5421 37139 5455
rect 18017 5356 18051 5390
rect 24639 5357 24673 5391
rect 17899 5239 17933 5273
rect 17487 4813 17521 5189
rect 17605 4813 17639 5189
rect 17723 4813 17757 5189
rect 17840 5013 17874 5189
rect 17958 5013 17992 5189
rect 18066 4781 18215 4848
rect 18714 4833 18748 5009
rect 18832 4833 18866 5009
rect 18950 4833 18984 5009
rect 19068 4833 19102 5009
rect 19198 4833 19232 5209
rect 19316 4833 19350 5209
rect 19434 4833 19468 5209
rect 19552 4833 19586 5209
rect 19670 4833 19704 5209
rect 19788 4833 19822 5209
rect 19906 4833 19940 5209
rect 20035 4833 20069 5009
rect 20153 4833 20187 5009
rect 20271 4833 20305 5009
rect 20389 4833 20423 5009
rect 20612 4833 20646 5009
rect 20730 4833 20764 5009
rect 20848 4833 20882 5009
rect 20966 4833 21000 5009
rect 21096 4833 21130 5209
rect 21214 4833 21248 5209
rect 21332 4833 21366 5209
rect 21450 4833 21484 5209
rect 21568 4833 21602 5209
rect 24521 5240 24555 5274
rect 21686 4833 21720 5209
rect 21804 4833 21838 5209
rect 21933 4833 21967 5009
rect 22051 4833 22085 5009
rect 22169 4833 22203 5009
rect 22287 4833 22321 5009
rect 24109 4814 24143 5190
rect 24227 4814 24261 5190
rect 24345 4814 24379 5190
rect 24462 5014 24496 5190
rect 24580 5014 24614 5190
rect 17546 4729 17580 4763
rect 17664 4729 17698 4763
rect 24689 4788 24838 4855
rect 25336 4834 25370 5010
rect 25454 4834 25488 5010
rect 25572 4834 25606 5010
rect 25690 4834 25724 5010
rect 25820 4834 25854 5210
rect 25938 4834 25972 5210
rect 26056 4834 26090 5210
rect 26174 4834 26208 5210
rect 26292 4834 26326 5210
rect 26410 4834 26444 5210
rect 26528 4834 26562 5210
rect 26657 4834 26691 5010
rect 26775 4834 26809 5010
rect 26893 4834 26927 5010
rect 27011 4834 27045 5010
rect 27234 4834 27268 5010
rect 27352 4834 27386 5010
rect 27470 4834 27504 5010
rect 27588 4834 27622 5010
rect 27718 4834 27752 5210
rect 27836 4834 27870 5210
rect 27954 4834 27988 5210
rect 28072 4834 28106 5210
rect 28190 4834 28224 5210
rect 28308 4834 28342 5210
rect 28426 4834 28460 5210
rect 32217 5212 32352 5314
rect 36763 5308 37139 5342
rect 38096 5382 38272 5416
rect 38096 5264 38272 5298
rect 36763 5190 37139 5224
rect 36763 5072 37139 5106
rect 28555 4834 28589 5010
rect 28673 4834 28707 5010
rect 28791 4834 28825 5010
rect 28909 4834 28943 5010
rect 36513 4926 36567 4998
rect 38096 5190 38472 5224
rect 37354 5130 37388 5164
rect 37738 5176 37793 5178
rect 37738 5118 37793 5176
rect 36763 4954 37139 4988
rect 38096 5072 38472 5106
rect 37453 5058 37508 5060
rect 37453 5000 37508 5058
rect 38096 4954 38472 4988
rect 36763 4836 37139 4870
rect 24168 4730 24202 4764
rect 24286 4730 24320 4764
rect 30072 4659 30132 4721
rect 38573 4953 38607 4987
rect 37974 4895 38008 4929
rect 38725 4926 38739 4984
rect 38739 4926 38771 4984
rect 38096 4836 38472 4870
rect 37584 4776 37618 4810
rect 36763 4718 37139 4752
rect 38096 4718 38472 4752
rect 20178 4561 20212 4595
rect 36763 4600 37139 4634
rect 22285 4540 22319 4574
rect 26800 4562 26834 4596
rect 17722 4287 17786 4433
rect 17786 4287 17789 4433
rect 17722 4284 17789 4287
rect 19141 4140 19175 4516
rect 19259 4140 19293 4516
rect 17245 3846 17279 4022
rect 17363 3846 17397 4022
rect 17481 3846 17515 4022
rect 17599 3846 17633 4022
rect 17717 3846 17751 4022
rect 17835 3846 17869 4022
rect 17953 3846 17987 4022
rect 18071 3846 18105 4022
rect 18189 3846 18223 4022
rect 19377 4140 19411 4516
rect 19495 4140 19529 4516
rect 19613 4140 19647 4516
rect 19731 4140 19765 4516
rect 19849 4140 19883 4516
rect 21039 4140 21073 4516
rect 21157 4140 21191 4516
rect 21275 4140 21309 4516
rect 21393 4140 21427 4516
rect 21511 4140 21545 4516
rect 21629 4140 21663 4516
rect 28907 4541 28941 4575
rect 21747 4140 21781 4516
rect 24343 4288 24408 4433
rect 24408 4288 24410 4433
rect 24343 4284 24410 4288
rect 25763 4141 25797 4517
rect 25881 4141 25915 4517
rect 18307 3846 18341 4022
rect 19171 3918 19205 3952
rect 18986 3851 19020 3885
rect 19819 3918 19853 3952
rect 21069 3918 21103 3952
rect 19437 3834 19471 3868
rect 19555 3835 19589 3869
rect 20109 3850 20143 3884
rect 20884 3851 20918 3885
rect 22408 4013 22540 4111
rect 21715 3919 21749 3953
rect 21335 3834 21369 3868
rect 21453 3835 21487 3869
rect 22007 3850 22041 3884
rect 23867 3847 23901 4023
rect 23985 3847 24019 4023
rect 24103 3847 24137 4023
rect 24221 3847 24255 4023
rect 24339 3847 24373 4023
rect 24457 3847 24491 4023
rect 24575 3847 24609 4023
rect 24693 3847 24727 4023
rect 24811 3847 24845 4023
rect 25999 4141 26033 4517
rect 26117 4141 26151 4517
rect 26235 4141 26269 4517
rect 26353 4141 26387 4517
rect 26471 4141 26505 4517
rect 27661 4141 27695 4517
rect 27779 4141 27813 4517
rect 27897 4141 27931 4517
rect 28015 4141 28049 4517
rect 28133 4141 28167 4517
rect 28251 4141 28285 4517
rect 28369 4141 28403 4517
rect 29731 4307 29765 4483
rect 29849 4307 29883 4483
rect 29967 4307 30001 4483
rect 30085 4307 30119 4483
rect 30203 4307 30237 4483
rect 30321 4307 30355 4483
rect 30439 4307 30473 4483
rect 30557 4307 30591 4483
rect 30675 4307 30709 4483
rect 38096 4640 38272 4674
rect 38096 4522 38272 4556
rect 30793 4307 30827 4483
rect 36763 4481 37139 4515
rect 36763 4363 37139 4397
rect 30498 4213 30532 4247
rect 36763 4245 37139 4279
rect 24929 3847 24963 4023
rect 25793 3919 25827 3953
rect 25608 3852 25642 3886
rect 26441 3919 26475 3953
rect 27691 3919 27725 3953
rect 26059 3835 26093 3869
rect 26177 3836 26211 3870
rect 26731 3851 26765 3885
rect 27506 3852 27540 3886
rect 29030 4014 29162 4112
rect 30380 4096 30414 4130
rect 36763 4127 37139 4161
rect 28337 3920 28371 3954
rect 27957 3835 27991 3869
rect 28075 3836 28109 3870
rect 28629 3851 28663 3885
rect 18012 3752 18046 3786
rect 17894 3635 17928 3669
rect 18839 3608 18873 3784
rect 17482 3209 17516 3585
rect 17600 3209 17634 3585
rect 17718 3209 17752 3585
rect 17835 3409 17869 3585
rect 18957 3608 18991 3784
rect 17953 3409 17987 3585
rect 19259 3408 19293 3784
rect 19377 3408 19411 3784
rect 19495 3408 19529 3784
rect 19613 3408 19647 3784
rect 19731 3408 19765 3784
rect 20137 3608 20171 3784
rect 20255 3608 20289 3784
rect 20737 3608 20771 3784
rect 20855 3608 20889 3784
rect 21157 3408 21191 3784
rect 21275 3408 21309 3784
rect 21393 3408 21427 3784
rect 21511 3408 21545 3784
rect 21629 3408 21663 3784
rect 22035 3608 22069 3784
rect 22153 3608 22187 3784
rect 24634 3753 24668 3787
rect 24516 3636 24550 3670
rect 25461 3609 25495 3785
rect 18069 3172 18215 3239
rect 18215 3172 18218 3239
rect 24104 3210 24138 3586
rect 24222 3210 24256 3586
rect 24340 3210 24374 3586
rect 24457 3410 24491 3586
rect 25579 3609 25613 3785
rect 24575 3410 24609 3586
rect 25881 3409 25915 3785
rect 25999 3409 26033 3785
rect 26117 3409 26151 3785
rect 26235 3409 26269 3785
rect 26353 3409 26387 3785
rect 26759 3609 26793 3785
rect 26877 3609 26911 3785
rect 27359 3609 27393 3785
rect 27477 3609 27511 3785
rect 27779 3409 27813 3785
rect 27897 3409 27931 3785
rect 28015 3409 28049 3785
rect 28133 3409 28167 3785
rect 28251 3409 28285 3785
rect 28657 3609 28691 3785
rect 28775 3609 28809 3785
rect 29968 3670 30002 4046
rect 30086 3670 30120 4046
rect 30204 3670 30238 4046
rect 30321 3870 30355 4046
rect 30439 3870 30473 4046
rect 36963 4008 37139 4042
rect 36963 3890 37139 3924
rect 36963 3772 37139 3806
rect 37313 3820 37347 3854
rect 36963 3654 37139 3688
rect 30027 3586 30061 3620
rect 30145 3586 30179 3620
rect 30300 3463 30352 3509
rect 32112 3442 32533 3476
rect 32112 3297 32175 3442
rect 32175 3297 32484 3442
rect 32484 3297 32533 3442
rect 32112 3276 32533 3297
rect 34797 3275 34890 3341
rect 17541 3125 17575 3159
rect 17659 3125 17693 3159
rect 24680 3171 24829 3238
rect 16430 2922 16500 2990
rect 24163 3126 24197 3160
rect 24281 3126 24315 3160
rect 37737 3196 37797 3245
rect 19471 2937 19538 3086
rect 26099 2943 26166 3092
rect 36963 3072 37139 3106
rect 31478 2562 31512 2738
rect 31596 2562 31630 2738
rect 31714 2562 31748 2738
rect 31832 2562 31866 2738
rect 31962 2562 31996 2938
rect 32080 2562 32114 2938
rect 32198 2562 32232 2938
rect 32316 2562 32350 2938
rect 32434 2562 32468 2938
rect 32552 2562 32586 2938
rect 32670 2562 32704 2938
rect 33612 2911 33672 2973
rect 36963 2954 37139 2988
rect 36963 2836 37139 2870
rect 32799 2562 32833 2738
rect 32917 2562 32951 2738
rect 33035 2562 33069 2738
rect 33153 2562 33187 2738
rect 33271 2559 33305 2735
rect 33389 2559 33423 2735
rect 33507 2559 33541 2735
rect 33625 2559 33659 2735
rect 33743 2559 33777 2735
rect 33861 2559 33895 2735
rect 33979 2559 34013 2735
rect 34097 2559 34131 2735
rect 34215 2559 34249 2735
rect 37454 2943 37509 3001
rect 37454 2941 37509 2943
rect 34333 2559 34367 2735
rect 36963 2718 37139 2752
rect 36763 2631 37139 2665
rect 34038 2465 34072 2499
rect 36763 2513 37139 2547
rect 8416 2318 8468 2364
rect 14970 2323 15022 2369
rect 21619 2311 21671 2357
rect 31458 2329 31531 2400
rect 36763 2395 37139 2429
rect 33130 2346 33164 2380
rect 33920 2348 33954 2382
rect 8143 2207 8177 2241
rect 8261 2207 8295 2241
rect 14697 2212 14731 2246
rect 14815 2212 14849 2246
rect 21346 2200 21380 2234
rect 21464 2200 21498 2234
rect 31730 2227 31764 2261
rect 8084 1781 8118 2157
rect 8202 1781 8236 2157
rect 8320 1781 8354 2157
rect 8437 1781 8471 1957
rect 8555 1781 8589 1957
rect 14638 1786 14672 2162
rect 14756 1786 14790 2162
rect 14874 1786 14908 2162
rect 14991 1786 15025 1962
rect 15109 1786 15143 1962
rect 21287 1774 21321 2150
rect 21405 1774 21439 2150
rect 21523 1774 21557 2150
rect 21640 1774 21674 1950
rect 21758 1774 21792 1950
rect 30079 1814 30139 1876
rect 31905 1869 31939 2245
rect 32023 1869 32057 2245
rect 32141 1869 32175 2245
rect 32259 1869 32293 2245
rect 32377 1869 32411 2245
rect 32495 1869 32529 2245
rect 32613 1869 32647 2245
rect 32779 1949 32841 2040
rect 33508 1922 33542 2298
rect 33626 1922 33660 2298
rect 33744 1922 33778 2298
rect 33861 2122 33895 2298
rect 33979 2122 34013 2298
rect 36763 2277 37139 2311
rect 36763 2164 37139 2198
rect 38096 2238 38272 2272
rect 38096 2120 38272 2154
rect 36763 2046 37139 2080
rect 36763 1928 37139 1962
rect 33567 1838 33601 1872
rect 33685 1838 33719 1872
rect 8496 1697 8530 1731
rect 15050 1702 15084 1736
rect 21699 1690 21733 1724
rect 8614 1580 8648 1614
rect 15168 1585 15202 1619
rect 21817 1573 21851 1607
rect 7847 1344 7881 1520
rect 7965 1344 7999 1520
rect 8083 1344 8117 1520
rect 8201 1344 8235 1520
rect 8319 1344 8353 1520
rect 8437 1344 8471 1520
rect 8555 1344 8589 1520
rect 8673 1344 8707 1520
rect 8791 1344 8825 1520
rect 8909 1344 8943 1520
rect 14401 1349 14435 1525
rect 14519 1349 14553 1525
rect 14637 1349 14671 1525
rect 14755 1349 14789 1525
rect 14873 1349 14907 1525
rect 14991 1349 15025 1525
rect 15109 1349 15143 1525
rect 15227 1349 15261 1525
rect 15345 1349 15379 1525
rect 15463 1349 15497 1525
rect 21050 1337 21084 1513
rect 21168 1337 21202 1513
rect 21286 1337 21320 1513
rect 21404 1337 21438 1513
rect 21522 1337 21556 1513
rect 21640 1337 21674 1513
rect 21758 1337 21792 1513
rect 21876 1337 21910 1513
rect 21994 1337 22028 1513
rect 22112 1337 22146 1513
rect 29738 1462 29772 1638
rect 29856 1462 29890 1638
rect 29974 1462 30008 1638
rect 30092 1462 30126 1638
rect 30210 1462 30244 1638
rect 30328 1462 30362 1638
rect 30446 1462 30480 1638
rect 30564 1462 30598 1638
rect 30682 1462 30716 1638
rect 30800 1462 30834 1638
rect 31935 1647 31969 1681
rect 31750 1580 31784 1614
rect 33840 1715 33892 1761
rect 36513 1782 36567 1854
rect 38096 2046 38472 2080
rect 37354 1986 37388 2020
rect 37738 2032 37793 2034
rect 37738 1974 37793 2032
rect 36763 1810 37139 1844
rect 38096 1928 38472 1962
rect 37453 1914 37508 1916
rect 37453 1856 37508 1914
rect 38096 1810 38472 1844
rect 32583 1647 32617 1681
rect 36763 1692 37139 1726
rect 32201 1563 32235 1597
rect 32319 1564 32353 1598
rect 32873 1579 32907 1613
rect 30505 1368 30539 1402
rect 31603 1337 31637 1513
rect 31721 1337 31755 1513
rect 30387 1251 30421 1285
rect 8188 1106 8248 1168
rect 14742 1111 14802 1173
rect 21391 1099 21451 1161
rect 29975 825 30009 1201
rect 30093 825 30127 1201
rect 30211 825 30245 1201
rect 30328 1025 30362 1201
rect 30446 1025 30480 1201
rect 32023 1137 32057 1513
rect 32141 1137 32175 1513
rect 32259 1137 32293 1513
rect 32377 1137 32411 1513
rect 32495 1137 32529 1513
rect 32901 1337 32935 1513
rect 33019 1337 33053 1513
rect 38573 1809 38607 1843
rect 37974 1751 38008 1785
rect 38725 1782 38739 1840
rect 38739 1782 38771 1840
rect 38096 1692 38472 1726
rect 37584 1632 37618 1666
rect 36763 1574 37139 1608
rect 38096 1574 38472 1608
rect 36763 1456 37139 1490
rect 38096 1496 38272 1530
rect 38096 1378 38272 1412
rect 36763 1337 37139 1371
rect 36763 1219 37139 1253
rect 36763 1101 37139 1135
rect 36763 983 37139 1017
rect 32217 864 32352 966
rect 36963 864 37139 898
rect 30034 741 30068 775
rect 30152 741 30186 775
rect 36963 746 37139 780
rect 30307 618 30359 664
rect 36963 628 37139 662
rect 37313 676 37347 710
rect 36963 510 37139 544
rect -2371 319 -2195 353
rect 15 278 122 361
rect 2748 289 2892 355
rect -2371 201 -2195 235
rect -3596 67 -3420 101
rect -2699 35 -2597 137
<< metal1 >>
rect 4376 28316 4538 28575
rect 4375 28302 4538 28316
rect 4375 28180 4391 28302
rect 4522 28180 4538 28302
rect 4375 28130 4538 28180
rect 6239 27906 6459 27926
rect 6239 27798 6283 27906
rect 6415 27798 6459 27906
rect 8036 27864 8092 27872
rect 6239 27756 6459 27798
rect 7110 27856 8092 27864
rect 7110 27822 8052 27856
rect 8086 27822 8092 27856
rect 8755 27852 8765 27960
rect 8897 27897 8907 27960
rect 8897 27886 8909 27897
rect 8897 27852 8910 27886
rect 9166 27876 9222 27878
rect 7110 27806 8092 27822
rect 8765 27814 8910 27852
rect 7110 27805 8089 27806
rect 5843 27726 6820 27756
rect 5843 27620 5875 27726
rect 6079 27620 6111 27726
rect 6315 27620 6347 27726
rect 6551 27620 6583 27726
rect 6786 27620 6820 27726
rect 5836 27608 5882 27620
rect 5836 27432 5842 27608
rect 5876 27432 5882 27608
rect 5836 27420 5882 27432
rect 5954 27608 6000 27620
rect 5954 27432 5960 27608
rect 5994 27432 6000 27608
rect 5954 27420 6000 27432
rect 6072 27608 6118 27620
rect 6072 27432 6078 27608
rect 6112 27432 6118 27608
rect 6072 27420 6118 27432
rect 6190 27608 6236 27620
rect 6190 27432 6196 27608
rect 6230 27432 6236 27608
rect 6190 27420 6236 27432
rect 6308 27608 6354 27620
rect 6308 27432 6314 27608
rect 6348 27432 6354 27608
rect 6308 27420 6354 27432
rect 6426 27608 6472 27620
rect 6426 27432 6432 27608
rect 6466 27432 6472 27608
rect 6426 27420 6472 27432
rect 6544 27608 6590 27620
rect 6544 27432 6550 27608
rect 6584 27432 6590 27608
rect 6544 27420 6590 27432
rect 6662 27608 6708 27620
rect 6662 27432 6668 27608
rect 6702 27432 6708 27608
rect 6662 27420 6708 27432
rect 6780 27608 6826 27620
rect 6780 27432 6786 27608
rect 6820 27432 6826 27608
rect 6780 27420 6826 27432
rect 6898 27608 6944 27620
rect 6898 27432 6904 27608
rect 6938 27432 6944 27608
rect 6898 27420 6944 27432
rect 5959 27326 5995 27420
rect 6195 27326 6231 27420
rect 6431 27327 6467 27420
rect 6593 27372 6659 27379
rect 6593 27338 6609 27372
rect 6643 27338 6659 27372
rect 6593 27327 6659 27338
rect 6431 27326 6659 27327
rect 5959 27297 6659 27326
rect 5959 27296 6541 27297
rect 341 27256 740 27257
rect -4186 27078 740 27256
rect 6079 27183 6113 27296
rect 6475 27255 6541 27296
rect 6475 27221 6491 27255
rect 6525 27221 6541 27255
rect 6475 27214 6541 27221
rect 6903 27215 6938 27420
rect 7110 27215 7177 27805
rect 8869 27782 8910 27814
rect 9156 27810 9166 27876
rect 9222 27810 9232 27876
rect 9902 27852 9912 27960
rect 10044 27897 10054 27960
rect 12752 27903 12972 27923
rect 10044 27886 10056 27897
rect 10044 27852 10057 27886
rect 9912 27814 10057 27852
rect 10016 27786 10057 27814
rect 8285 27754 8555 27782
rect 8026 27688 8036 27754
rect 8102 27688 8112 27754
rect 8285 27692 8319 27754
rect 8521 27692 8555 27754
rect 8639 27754 8910 27782
rect 9427 27758 9697 27786
rect 8639 27692 8673 27754
rect 8875 27692 8910 27754
rect 9051 27742 9222 27758
rect 9051 27708 9182 27742
rect 9216 27708 9222 27742
rect 9051 27692 9222 27708
rect 9427 27696 9461 27758
rect 9663 27696 9697 27758
rect 9781 27758 10057 27786
rect 9781 27696 9815 27758
rect 10017 27696 10057 27758
rect 12752 27795 12796 27903
rect 12928 27795 12972 27903
rect 14549 27861 14605 27869
rect 12752 27753 12972 27795
rect 13623 27853 14605 27861
rect 13623 27819 14565 27853
rect 14599 27819 14605 27853
rect 15268 27849 15278 27957
rect 15410 27894 15420 27957
rect 15410 27883 15422 27894
rect 15410 27849 15423 27883
rect 15679 27873 15735 27875
rect 13623 27803 14605 27819
rect 15278 27811 15423 27849
rect 13623 27802 14602 27803
rect 8161 27680 8207 27692
rect 8161 27304 8167 27680
rect 8201 27304 8207 27680
rect 8161 27292 8207 27304
rect 8279 27680 8325 27692
rect 8279 27304 8285 27680
rect 8319 27304 8325 27680
rect 8279 27292 8325 27304
rect 8397 27680 8443 27692
rect 8397 27304 8403 27680
rect 8437 27304 8443 27680
rect 8397 27292 8443 27304
rect 8515 27680 8561 27692
rect 8515 27304 8521 27680
rect 8555 27304 8561 27680
rect 8515 27292 8561 27304
rect 8633 27680 8679 27692
rect 8633 27304 8639 27680
rect 8673 27304 8679 27680
rect 8633 27292 8679 27304
rect 8751 27680 8797 27692
rect 8751 27304 8757 27680
rect 8791 27304 8797 27680
rect 8751 27292 8797 27304
rect 8869 27680 8915 27692
rect 8869 27304 8875 27680
rect 8909 27304 8915 27680
rect 8869 27292 8915 27304
rect 6903 27187 7177 27215
rect 6549 27183 7177 27187
rect -4189 26648 572 26831
rect 646 26816 740 27078
rect 6073 27171 6119 27183
rect 646 26778 5190 26816
rect 6073 26795 6079 27171
rect 6113 26795 6119 27171
rect 6073 26783 6119 26795
rect 6191 27171 6237 27183
rect 6191 26795 6197 27171
rect 6231 26795 6237 27171
rect 6191 26783 6237 26795
rect 6309 27171 6355 27183
rect 6309 26795 6315 27171
rect 6349 26819 6355 27171
rect 6426 27171 6472 27183
rect 6426 26995 6432 27171
rect 6466 26995 6472 27171
rect 6426 26983 6472 26995
rect 6544 27171 7177 27183
rect 6544 26995 6550 27171
rect 6584 27158 7177 27171
rect 8167 27250 8201 27292
rect 8403 27250 8437 27292
rect 8167 27222 8437 27250
rect 8521 27251 8555 27292
rect 8757 27251 8791 27292
rect 8521 27222 8791 27251
rect 8167 27174 8201 27222
rect 6584 26995 6590 27158
rect 8167 27144 8230 27174
rect 6544 26983 6590 26995
rect 8195 27052 8230 27144
rect 8195 27016 8422 27052
rect 8692 27041 8702 27138
rect 8801 27041 8811 27138
rect 8875 27109 8909 27292
rect 8875 27055 8984 27109
rect 6432 26867 6467 26983
rect 8195 26909 8230 27016
rect 8356 26982 8422 27016
rect 8356 26948 8372 26982
rect 8406 26948 8422 26982
rect 8703 27040 8800 27041
rect 8703 26973 8760 27040
rect 8356 26942 8422 26948
rect 8597 26937 8866 26973
rect 8597 26909 8630 26937
rect 8833 26909 8866 26937
rect 8950 26909 8984 27055
rect 8071 26897 8117 26909
rect 6563 26867 6671 26877
rect 6432 26819 6563 26867
rect 6349 26795 6563 26819
rect 6309 26783 6563 26795
rect 6315 26779 6563 26783
rect 646 26751 5951 26778
rect 646 26745 6188 26751
rect 646 26711 6138 26745
rect 6172 26711 6188 26745
rect 646 26695 6188 26711
rect 6240 26745 6306 26751
rect 6240 26711 6256 26745
rect 6290 26711 6306 26745
rect 6489 26735 6563 26779
rect 6563 26725 6671 26735
rect 646 26679 5951 26695
rect 646 26678 5888 26679
rect 646 26674 5423 26678
rect 4901 26673 5190 26674
rect -4192 26227 432 26418
rect -195 25994 288 25995
rect -4186 25939 288 25994
rect -4186 25890 64 25939
rect 118 25890 288 25939
rect -4186 25808 288 25890
rect -4186 25806 -131 25808
rect -4189 25518 125 25562
rect -4189 25447 -92 25518
rect -23 25447 125 25518
rect -4189 25376 125 25447
rect -4192 25094 -14 25137
rect -4192 25023 -239 25094
rect -168 25023 -14 25094
rect -4192 24955 -14 25023
rect -4186 24634 -143 24689
rect -4186 24573 -382 24634
rect -311 24573 -143 24634
rect -4186 24503 -143 24573
rect -217 24303 -143 24503
rect -1161 24264 -276 24265
rect -4189 24073 -276 24264
rect -1183 23828 -429 23829
rect -4192 23652 -429 23828
rect -1183 23650 -429 23652
rect -1168 23415 -588 23418
rect -4190 23393 -588 23415
rect -4190 23256 -832 23393
rect -674 23256 -588 23393
rect -4190 23232 -588 23256
rect -4193 22994 -1108 22995
rect -4193 22802 -723 22994
rect -4196 22381 -858 22555
rect -4190 21941 -998 22130
rect -4193 21511 -1135 21690
rect -4196 21090 -1273 21265
rect -4193 20661 -1415 20846
rect -4196 20231 -1568 20415
rect -3222 20009 -3134 20011
rect -4199 19810 -3134 20009
rect -3255 16262 -3134 19810
rect -3604 16255 -3404 16261
rect -3604 16221 -3592 16255
rect -3416 16221 -3335 16255
rect -3604 16215 -3404 16221
rect -3604 16137 -3404 16143
rect -3950 16103 -3592 16137
rect -3416 16103 -3404 16137
rect -3950 15771 -3907 16103
rect -3604 16097 -3404 16103
rect -3370 16130 -3335 16221
rect -3253 16236 -3134 16262
rect -3063 16248 -2991 16261
rect -3187 16215 -3134 16236
rect -3067 16184 -3057 16248
rect -2996 16184 -2986 16248
rect -3063 16182 -3057 16184
rect -2997 16182 -2991 16184
rect -3063 16170 -2991 16182
rect -3253 16160 -3187 16170
rect -2379 16130 -2179 16136
rect -3370 16096 -2367 16130
rect -2191 16096 -2179 16130
rect -3604 16019 -3404 16025
rect -3604 15985 -3592 16019
rect -3416 15985 -3404 16019
rect -3604 15979 -3404 15985
rect -3604 15901 -3404 15907
rect -3604 15867 -3592 15901
rect -3416 15867 -3404 15901
rect -3604 15861 -3404 15867
rect -3592 15777 -3416 15861
rect -3111 15828 -2711 15834
rect -3273 15794 -3099 15828
rect -2723 15794 -2711 15828
rect -2551 15814 -2508 16096
rect -2379 16090 -2179 16096
rect -2379 16013 -2179 16018
rect -2379 16012 -1853 16013
rect -2480 15983 -2418 15989
rect -2480 15949 -2468 15983
rect -2434 15949 -2418 15983
rect -2379 15978 -2367 16012
rect -2191 15979 -1853 16012
rect -2191 15978 -2179 15979
rect -2379 15972 -2179 15978
rect -2480 15933 -2418 15949
rect -3804 15771 -3404 15777
rect -3950 15737 -3792 15771
rect -3416 15737 -3404 15771
rect -3950 15535 -3907 15737
rect -3804 15731 -3404 15737
rect -3804 15653 -3404 15659
rect -3804 15619 -3792 15653
rect -3416 15619 -3335 15653
rect -3804 15613 -3404 15619
rect -3804 15535 -3404 15541
rect -3950 15501 -3792 15535
rect -3416 15501 -3404 15535
rect -3950 15466 -3907 15501
rect -3804 15495 -3404 15501
rect -4033 15438 -3907 15466
rect -4055 15428 -3907 15438
rect -4001 15374 -3907 15428
rect -3804 15417 -3404 15423
rect -3370 15417 -3335 15619
rect -3273 15592 -3235 15794
rect -3111 15788 -2711 15794
rect -2546 15798 -2495 15814
rect -2546 15764 -2535 15798
rect -2501 15764 -2495 15798
rect -2546 15747 -2495 15764
rect -3111 15710 -2711 15716
rect -3111 15676 -3099 15710
rect -2723 15676 -2711 15710
rect -3111 15670 -2711 15676
rect -3111 15592 -2711 15598
rect -3273 15558 -3099 15592
rect -2723 15558 -2711 15592
rect -3273 15417 -3235 15558
rect -3111 15552 -2711 15558
rect -2467 15548 -2418 15933
rect -2379 15710 -1979 15716
rect -2379 15676 -2367 15710
rect -1991 15676 -1979 15710
rect -2379 15670 -1979 15676
rect -2379 15592 -1979 15598
rect -2379 15558 -2367 15592
rect -1991 15558 -1979 15592
rect -2379 15552 -1979 15558
rect -2467 15532 -2410 15548
rect -2467 15498 -2451 15532
rect -2417 15498 -2410 15532
rect -2467 15482 -2410 15498
rect -1885 15520 -1853 15979
rect -1885 15486 -1768 15520
rect -3111 15474 -2711 15480
rect -3111 15440 -3099 15474
rect -2723 15440 -2711 15474
rect -3111 15434 -2711 15440
rect -2379 15474 -1979 15480
rect -2379 15440 -2367 15474
rect -1991 15440 -1979 15474
rect -2379 15434 -1979 15440
rect -3804 15383 -3792 15417
rect -3416 15383 -3235 15417
rect -3804 15377 -3404 15383
rect -4055 15364 -3907 15374
rect -4033 15332 -3907 15364
rect -3950 15299 -3907 15332
rect -3273 15356 -3235 15383
rect -2467 15414 -2408 15430
rect -2467 15380 -2452 15414
rect -2418 15380 -2408 15414
rect -2467 15363 -2408 15380
rect -1885 15424 -1831 15486
rect -1773 15424 -1768 15486
rect -1885 15388 -1768 15424
rect -3111 15356 -2711 15362
rect -3273 15322 -3099 15356
rect -2723 15322 -2711 15356
rect -3804 15299 -3404 15305
rect -3950 15265 -3792 15299
rect -3416 15265 -3404 15299
rect -3950 15063 -3907 15265
rect -3804 15259 -3404 15265
rect -3804 15181 -3404 15187
rect -3804 15147 -3792 15181
rect -3416 15147 -3404 15181
rect -3804 15141 -3404 15147
rect -3273 15120 -3235 15322
rect -3111 15316 -2711 15322
rect -3111 15238 -2711 15244
rect -3111 15204 -3099 15238
rect -2723 15204 -2711 15238
rect -3111 15198 -2711 15204
rect -2546 15150 -2495 15167
rect -3111 15120 -2711 15126
rect -3273 15086 -3099 15120
rect -2723 15086 -2711 15120
rect -2546 15116 -2535 15150
rect -2501 15116 -2495 15150
rect -2546 15100 -2495 15116
rect -3111 15080 -2711 15086
rect -3804 15063 -3404 15069
rect -3950 15029 -3792 15063
rect -3416 15029 -3404 15063
rect -3950 14698 -3907 15029
rect -3804 15023 -3404 15029
rect -3592 14940 -3416 15023
rect -2551 14987 -2508 15100
rect -3604 14934 -3404 14940
rect -3604 14900 -3592 14934
rect -3416 14900 -3404 14934
rect -3604 14894 -3404 14900
rect -3253 14848 -3187 14860
rect -3604 14816 -3404 14822
rect -3604 14782 -3592 14816
rect -3416 14782 -3335 14816
rect -3253 14794 -3247 14848
rect -3193 14794 -3187 14848
rect -3253 14782 -3187 14794
rect -3604 14776 -3404 14782
rect -3370 14714 -3335 14782
rect -2552 14714 -2507 14987
rect -2467 14876 -2418 15363
rect -2379 15356 -1979 15362
rect -1885 15356 -1853 15388
rect -2379 15322 -2367 15356
rect -1991 15322 -1853 15356
rect -2379 15316 -1979 15322
rect -2379 15238 -1979 15244
rect -2379 15204 -2367 15238
rect -1991 15204 -1979 15238
rect -2379 15198 -1979 15204
rect -2479 14860 -2417 14876
rect -2479 14826 -2467 14860
rect -2433 14826 -2417 14860
rect -2479 14820 -2417 14826
rect -2379 14832 -2179 14838
rect -1885 14832 -1853 15322
rect -2379 14798 -2367 14832
rect -2191 14799 -1853 14832
rect -2191 14798 -2179 14799
rect -2379 14792 -2179 14798
rect -2379 14714 -2179 14720
rect -3604 14698 -3404 14704
rect -3950 14664 -3592 14698
rect -3416 14664 -3404 14698
rect -3604 14658 -3404 14664
rect -3370 14680 -2367 14714
rect -2191 14680 -2179 14714
rect -3604 14580 -3404 14586
rect -3370 14580 -3335 14680
rect -2379 14674 -2179 14680
rect -3604 14546 -3592 14580
rect -3416 14546 -3335 14580
rect -2701 14616 -2587 14628
rect -3604 14540 -3404 14546
rect -2701 14514 -2695 14616
rect -2593 14514 -2587 14616
rect -2701 14502 -2587 14514
rect -1657 14351 -1568 20231
rect -3255 14265 -1568 14351
rect -3255 14195 -3188 14265
rect -3606 14187 -3406 14193
rect -3606 14153 -3594 14187
rect -3418 14153 -3337 14187
rect -3606 14147 -3406 14153
rect -3606 14069 -3406 14075
rect -3952 14035 -3594 14069
rect -3418 14035 -3406 14069
rect -3952 13703 -3909 14035
rect -3606 14029 -3406 14035
rect -3372 14062 -3337 14153
rect -3255 14168 -3189 14195
rect -3066 14180 -2993 14193
rect -3066 14115 -3059 14180
rect -3065 14114 -3059 14115
rect -2999 14114 -2993 14180
rect -3065 14102 -2993 14114
rect -3255 14092 -3189 14102
rect -2381 14062 -2181 14068
rect -3372 14028 -2369 14062
rect -2193 14028 -2181 14062
rect -3606 13951 -3406 13957
rect -3606 13917 -3594 13951
rect -3418 13917 -3406 13951
rect -3606 13911 -3406 13917
rect -3606 13833 -3406 13839
rect -3606 13799 -3594 13833
rect -3418 13799 -3406 13833
rect -3606 13793 -3406 13799
rect -3594 13709 -3418 13793
rect -3113 13760 -2713 13766
rect -3275 13726 -3101 13760
rect -2725 13726 -2713 13760
rect -2553 13746 -2510 14028
rect -2381 14022 -2181 14028
rect -2381 13945 -2181 13950
rect -2381 13944 -1855 13945
rect -2482 13915 -2420 13921
rect -2482 13881 -2470 13915
rect -2436 13881 -2420 13915
rect -2381 13910 -2369 13944
rect -2193 13911 -1855 13944
rect -2193 13910 -2181 13911
rect -2381 13904 -2181 13910
rect -2482 13865 -2420 13881
rect -3806 13703 -3406 13709
rect -3952 13669 -3794 13703
rect -3418 13669 -3406 13703
rect -3952 13467 -3909 13669
rect -3806 13663 -3406 13669
rect -3806 13585 -3406 13591
rect -3806 13551 -3794 13585
rect -3418 13551 -3337 13585
rect -3806 13545 -3406 13551
rect -3806 13467 -3406 13473
rect -3952 13433 -3794 13467
rect -3418 13433 -3406 13467
rect -3952 13398 -3909 13433
rect -3806 13427 -3406 13433
rect -4035 13370 -3909 13398
rect -4057 13360 -3909 13370
rect -4003 13306 -3909 13360
rect -3806 13349 -3406 13355
rect -3372 13349 -3337 13551
rect -3275 13524 -3237 13726
rect -3113 13720 -2713 13726
rect -2548 13730 -2497 13746
rect -2548 13696 -2537 13730
rect -2503 13696 -2497 13730
rect -2548 13679 -2497 13696
rect -3113 13642 -2713 13648
rect -3113 13608 -3101 13642
rect -2725 13608 -2713 13642
rect -3113 13602 -2713 13608
rect -3113 13524 -2713 13530
rect -3275 13490 -3101 13524
rect -2725 13490 -2713 13524
rect -3275 13349 -3237 13490
rect -3113 13484 -2713 13490
rect -2469 13480 -2420 13865
rect -2381 13642 -1981 13648
rect -2381 13608 -2369 13642
rect -1993 13608 -1981 13642
rect -2381 13602 -1981 13608
rect -2381 13524 -1981 13530
rect -2381 13490 -2369 13524
rect -1993 13490 -1981 13524
rect -2381 13484 -1981 13490
rect -2469 13464 -2412 13480
rect -2469 13430 -2453 13464
rect -2419 13430 -2412 13464
rect -2469 13414 -2412 13430
rect -1887 13452 -1855 13911
rect -1887 13418 -1770 13452
rect -3113 13406 -2713 13412
rect -3113 13372 -3101 13406
rect -2725 13372 -2713 13406
rect -3113 13366 -2713 13372
rect -2381 13406 -1981 13412
rect -2381 13372 -2369 13406
rect -1993 13372 -1981 13406
rect -2381 13366 -1981 13372
rect -3806 13315 -3794 13349
rect -3418 13315 -3237 13349
rect -3806 13309 -3406 13315
rect -4057 13296 -3909 13306
rect -4035 13264 -3909 13296
rect -3952 13231 -3909 13264
rect -3275 13288 -3237 13315
rect -2469 13346 -2410 13362
rect -2469 13312 -2454 13346
rect -2420 13312 -2410 13346
rect -2469 13295 -2410 13312
rect -1887 13356 -1833 13418
rect -1775 13356 -1770 13418
rect -1887 13320 -1770 13356
rect -3113 13288 -2713 13294
rect -3275 13254 -3101 13288
rect -2725 13254 -2713 13288
rect -3806 13231 -3406 13237
rect -3952 13197 -3794 13231
rect -3418 13197 -3406 13231
rect -3952 12995 -3909 13197
rect -3806 13191 -3406 13197
rect -3806 13113 -3406 13119
rect -3806 13079 -3794 13113
rect -3418 13079 -3406 13113
rect -3806 13073 -3406 13079
rect -3275 13052 -3237 13254
rect -3113 13248 -2713 13254
rect -3113 13170 -2713 13176
rect -3113 13136 -3101 13170
rect -2725 13136 -2713 13170
rect -3113 13130 -2713 13136
rect -2548 13082 -2497 13099
rect -3113 13052 -2713 13058
rect -3275 13018 -3101 13052
rect -2725 13018 -2713 13052
rect -2548 13048 -2537 13082
rect -2503 13048 -2497 13082
rect -2548 13032 -2497 13048
rect -3113 13012 -2713 13018
rect -3806 12995 -3406 13001
rect -3952 12961 -3794 12995
rect -3418 12961 -3406 12995
rect -3952 12630 -3909 12961
rect -3806 12955 -3406 12961
rect -3594 12872 -3418 12955
rect -2553 12919 -2510 13032
rect -3606 12866 -3406 12872
rect -3606 12832 -3594 12866
rect -3418 12832 -3406 12866
rect -3606 12826 -3406 12832
rect -3255 12780 -3189 12792
rect -3606 12748 -3406 12754
rect -3606 12714 -3594 12748
rect -3418 12714 -3337 12748
rect -3255 12726 -3249 12780
rect -3195 12726 -3189 12780
rect -3255 12714 -3189 12726
rect -3606 12708 -3406 12714
rect -3372 12646 -3337 12714
rect -2554 12646 -2509 12919
rect -2469 12808 -2420 13295
rect -2381 13288 -1981 13294
rect -1887 13288 -1855 13320
rect -2381 13254 -2369 13288
rect -1993 13254 -1855 13288
rect -2381 13248 -1981 13254
rect -2381 13170 -1981 13176
rect -2381 13136 -2369 13170
rect -1993 13136 -1981 13170
rect -2381 13130 -1981 13136
rect -2481 12792 -2419 12808
rect -2481 12758 -2469 12792
rect -2435 12758 -2419 12792
rect -2481 12752 -2419 12758
rect -2381 12764 -2181 12770
rect -1887 12764 -1855 13254
rect -2381 12730 -2369 12764
rect -2193 12731 -1855 12764
rect -2193 12730 -2181 12731
rect -2381 12724 -2181 12730
rect -2381 12646 -2181 12652
rect -3606 12630 -3406 12636
rect -3952 12596 -3594 12630
rect -3418 12596 -3406 12630
rect -3606 12590 -3406 12596
rect -3372 12612 -2369 12646
rect -2193 12612 -2181 12646
rect -3606 12512 -3406 12518
rect -3372 12512 -3337 12612
rect -2381 12606 -2181 12612
rect -3606 12478 -3594 12512
rect -3418 12478 -3337 12512
rect -2703 12548 -2589 12560
rect -3606 12472 -3406 12478
rect -2703 12446 -2697 12548
rect -2595 12446 -2589 12548
rect -2703 12434 -2589 12446
rect -1494 12481 -1415 20661
rect -1494 12296 -1414 12481
rect -3254 12210 -1414 12296
rect -3604 12118 -3404 12124
rect -3604 12084 -3592 12118
rect -3416 12084 -3335 12118
rect -3254 12114 -3187 12210
rect -3604 12078 -3404 12084
rect -3604 12000 -3404 12006
rect -3950 11966 -3592 12000
rect -3416 11966 -3404 12000
rect -3950 11634 -3907 11966
rect -3604 11960 -3404 11966
rect -3370 11993 -3335 12084
rect -3253 12099 -3187 12114
rect -3063 12111 -2991 12125
rect -3063 12045 -3057 12111
rect -2997 12108 -2991 12111
rect -2996 12048 -2991 12108
rect -2997 12045 -2991 12048
rect -3063 12033 -2991 12045
rect -3253 12023 -3187 12033
rect -2379 11993 -2179 11999
rect -3370 11959 -2367 11993
rect -2191 11959 -2179 11993
rect -3604 11882 -3404 11888
rect -3604 11848 -3592 11882
rect -3416 11848 -3404 11882
rect -3604 11842 -3404 11848
rect -3604 11764 -3404 11770
rect -3604 11730 -3592 11764
rect -3416 11730 -3404 11764
rect -3604 11724 -3404 11730
rect -3592 11640 -3416 11724
rect -3111 11691 -2711 11697
rect -3273 11657 -3099 11691
rect -2723 11657 -2711 11691
rect -2551 11677 -2508 11959
rect -2379 11953 -2179 11959
rect -2379 11876 -2179 11881
rect -2379 11875 -1853 11876
rect -2480 11846 -2418 11852
rect -2480 11812 -2468 11846
rect -2434 11812 -2418 11846
rect -2379 11841 -2367 11875
rect -2191 11842 -1853 11875
rect -2191 11841 -2179 11842
rect -2379 11835 -2179 11841
rect -2480 11796 -2418 11812
rect -3804 11634 -3404 11640
rect -3950 11600 -3792 11634
rect -3416 11600 -3404 11634
rect -3950 11398 -3907 11600
rect -3804 11594 -3404 11600
rect -3804 11516 -3404 11522
rect -3804 11482 -3792 11516
rect -3416 11482 -3335 11516
rect -3804 11476 -3404 11482
rect -3804 11398 -3404 11404
rect -3950 11364 -3792 11398
rect -3416 11364 -3404 11398
rect -3950 11329 -3907 11364
rect -3804 11358 -3404 11364
rect -4033 11301 -3907 11329
rect -4055 11291 -3907 11301
rect -4001 11237 -3907 11291
rect -3804 11280 -3404 11286
rect -3370 11280 -3335 11482
rect -3273 11455 -3235 11657
rect -3111 11651 -2711 11657
rect -2546 11661 -2495 11677
rect -2546 11627 -2535 11661
rect -2501 11627 -2495 11661
rect -2546 11610 -2495 11627
rect -3111 11573 -2711 11579
rect -3111 11539 -3099 11573
rect -2723 11539 -2711 11573
rect -3111 11533 -2711 11539
rect -3111 11455 -2711 11461
rect -3273 11421 -3099 11455
rect -2723 11421 -2711 11455
rect -3273 11280 -3235 11421
rect -3111 11415 -2711 11421
rect -2467 11411 -2418 11796
rect -2379 11573 -1979 11579
rect -2379 11539 -2367 11573
rect -1991 11539 -1979 11573
rect -2379 11533 -1979 11539
rect -2379 11455 -1979 11461
rect -2379 11421 -2367 11455
rect -1991 11421 -1979 11455
rect -2379 11415 -1979 11421
rect -2467 11395 -2410 11411
rect -2467 11361 -2451 11395
rect -2417 11361 -2410 11395
rect -2467 11345 -2410 11361
rect -1885 11383 -1853 11842
rect -1885 11349 -1768 11383
rect -3111 11337 -2711 11343
rect -3111 11303 -3099 11337
rect -2723 11303 -2711 11337
rect -3111 11297 -2711 11303
rect -2379 11337 -1979 11343
rect -2379 11303 -2367 11337
rect -1991 11303 -1979 11337
rect -2379 11297 -1979 11303
rect -3804 11246 -3792 11280
rect -3416 11246 -3235 11280
rect -3804 11240 -3404 11246
rect -4055 11227 -3907 11237
rect -4033 11195 -3907 11227
rect -3950 11162 -3907 11195
rect -3273 11219 -3235 11246
rect -2467 11277 -2408 11293
rect -2467 11243 -2452 11277
rect -2418 11243 -2408 11277
rect -2467 11226 -2408 11243
rect -1885 11287 -1831 11349
rect -1773 11287 -1768 11349
rect -1885 11251 -1768 11287
rect -3111 11219 -2711 11225
rect -3273 11185 -3099 11219
rect -2723 11185 -2711 11219
rect -3804 11162 -3404 11168
rect -3950 11128 -3792 11162
rect -3416 11128 -3404 11162
rect -3950 10926 -3907 11128
rect -3804 11122 -3404 11128
rect -3804 11044 -3404 11050
rect -3804 11010 -3792 11044
rect -3416 11010 -3404 11044
rect -3804 11004 -3404 11010
rect -3273 10983 -3235 11185
rect -3111 11179 -2711 11185
rect -3111 11101 -2711 11107
rect -3111 11067 -3099 11101
rect -2723 11067 -2711 11101
rect -3111 11061 -2711 11067
rect -2546 11013 -2495 11030
rect -3111 10983 -2711 10989
rect -3273 10949 -3099 10983
rect -2723 10949 -2711 10983
rect -2546 10979 -2535 11013
rect -2501 10979 -2495 11013
rect -2546 10963 -2495 10979
rect -3111 10943 -2711 10949
rect -3804 10926 -3404 10932
rect -3950 10892 -3792 10926
rect -3416 10892 -3404 10926
rect -3950 10561 -3907 10892
rect -3804 10886 -3404 10892
rect -3592 10803 -3416 10886
rect -2551 10850 -2508 10963
rect -3604 10797 -3404 10803
rect -3604 10763 -3592 10797
rect -3416 10763 -3404 10797
rect -3604 10757 -3404 10763
rect -3253 10711 -3187 10723
rect -3604 10679 -3404 10685
rect -3604 10645 -3592 10679
rect -3416 10645 -3335 10679
rect -3253 10657 -3247 10711
rect -3193 10657 -3187 10711
rect -3253 10645 -3187 10657
rect -3604 10639 -3404 10645
rect -3370 10577 -3335 10645
rect -2552 10577 -2507 10850
rect -2467 10739 -2418 11226
rect -2379 11219 -1979 11225
rect -1885 11219 -1853 11251
rect -2379 11185 -2367 11219
rect -1991 11185 -1853 11219
rect -2379 11179 -1979 11185
rect -2379 11101 -1979 11107
rect -2379 11067 -2367 11101
rect -1991 11067 -1979 11101
rect -2379 11061 -1979 11067
rect -2479 10723 -2417 10739
rect -2479 10689 -2467 10723
rect -2433 10689 -2417 10723
rect -2479 10683 -2417 10689
rect -2379 10695 -2179 10701
rect -1885 10695 -1853 11185
rect -2379 10661 -2367 10695
rect -2191 10662 -1853 10695
rect -2191 10661 -2179 10662
rect -2379 10655 -2179 10661
rect -2379 10577 -2179 10583
rect -3604 10561 -3404 10567
rect -3950 10527 -3592 10561
rect -3416 10527 -3404 10561
rect -3604 10521 -3404 10527
rect -3370 10543 -2367 10577
rect -2191 10543 -2179 10577
rect -3604 10443 -3404 10449
rect -3370 10443 -3335 10543
rect -2379 10537 -2179 10543
rect -3604 10409 -3592 10443
rect -3416 10409 -3335 10443
rect -2701 10479 -2587 10491
rect -3604 10403 -3404 10409
rect -2701 10377 -2695 10479
rect -2593 10377 -2587 10479
rect -2701 10365 -2587 10377
rect -1350 10294 -1273 21090
rect -1216 12389 -1135 21511
rect -1219 12315 -1209 12389
rect -1143 12315 -1133 12389
rect -1350 10230 -1342 10294
rect -1280 10230 -1272 10294
rect -1350 10222 -1273 10230
rect -3255 10143 -1273 10222
rect -3606 10050 -3406 10056
rect -3606 10016 -3594 10050
rect -3418 10016 -3337 10050
rect -3606 10010 -3406 10016
rect -3606 9932 -3406 9938
rect -3952 9898 -3594 9932
rect -3418 9898 -3406 9932
rect -3952 9566 -3909 9898
rect -3606 9892 -3406 9898
rect -3372 9925 -3337 10016
rect -3255 10031 -3189 10143
rect -3065 10043 -2993 10056
rect -3065 9977 -3059 10043
rect -2999 9977 -2993 10043
rect -3065 9965 -2993 9977
rect -3255 9955 -3189 9965
rect -2381 9925 -2181 9931
rect -3372 9891 -2369 9925
rect -2193 9891 -2181 9925
rect -3606 9814 -3406 9820
rect -3606 9780 -3594 9814
rect -3418 9780 -3406 9814
rect -3606 9774 -3406 9780
rect -3606 9696 -3406 9702
rect -3606 9662 -3594 9696
rect -3418 9662 -3406 9696
rect -3606 9656 -3406 9662
rect -3594 9572 -3418 9656
rect -3113 9623 -2713 9629
rect -3275 9589 -3101 9623
rect -2725 9589 -2713 9623
rect -2553 9609 -2510 9891
rect -2381 9885 -2181 9891
rect -2381 9808 -2181 9813
rect -2381 9807 -1855 9808
rect -2482 9778 -2420 9784
rect -2482 9744 -2470 9778
rect -2436 9744 -2420 9778
rect -2381 9773 -2369 9807
rect -2193 9774 -1855 9807
rect -2193 9773 -2181 9774
rect -2381 9767 -2181 9773
rect -2482 9728 -2420 9744
rect -3806 9566 -3406 9572
rect -3952 9532 -3794 9566
rect -3418 9532 -3406 9566
rect -3952 9330 -3909 9532
rect -3806 9526 -3406 9532
rect -3806 9448 -3406 9454
rect -3806 9414 -3794 9448
rect -3418 9414 -3337 9448
rect -3806 9408 -3406 9414
rect -3806 9330 -3406 9336
rect -3952 9296 -3794 9330
rect -3418 9296 -3406 9330
rect -3952 9261 -3909 9296
rect -3806 9290 -3406 9296
rect -4035 9233 -3909 9261
rect -4057 9223 -3909 9233
rect -4003 9169 -3909 9223
rect -3806 9212 -3406 9218
rect -3372 9212 -3337 9414
rect -3275 9387 -3237 9589
rect -3113 9583 -2713 9589
rect -2548 9593 -2497 9609
rect -2548 9559 -2537 9593
rect -2503 9559 -2497 9593
rect -2548 9542 -2497 9559
rect -3113 9505 -2713 9511
rect -3113 9471 -3101 9505
rect -2725 9471 -2713 9505
rect -3113 9465 -2713 9471
rect -3113 9387 -2713 9393
rect -3275 9353 -3101 9387
rect -2725 9353 -2713 9387
rect -3275 9212 -3237 9353
rect -3113 9347 -2713 9353
rect -2469 9343 -2420 9728
rect -2381 9505 -1981 9511
rect -2381 9471 -2369 9505
rect -1993 9471 -1981 9505
rect -2381 9465 -1981 9471
rect -2381 9387 -1981 9393
rect -2381 9353 -2369 9387
rect -1993 9353 -1981 9387
rect -2381 9347 -1981 9353
rect -2469 9327 -2412 9343
rect -2469 9293 -2453 9327
rect -2419 9293 -2412 9327
rect -2469 9277 -2412 9293
rect -1887 9315 -1855 9774
rect -1887 9281 -1770 9315
rect -3113 9269 -2713 9275
rect -3113 9235 -3101 9269
rect -2725 9235 -2713 9269
rect -3113 9229 -2713 9235
rect -2381 9269 -1981 9275
rect -2381 9235 -2369 9269
rect -1993 9235 -1981 9269
rect -2381 9229 -1981 9235
rect -3806 9178 -3794 9212
rect -3418 9178 -3237 9212
rect -3806 9172 -3406 9178
rect -4057 9159 -3909 9169
rect -4035 9127 -3909 9159
rect -3952 9094 -3909 9127
rect -3275 9151 -3237 9178
rect -2469 9209 -2410 9225
rect -2469 9175 -2454 9209
rect -2420 9175 -2410 9209
rect -2469 9158 -2410 9175
rect -1887 9219 -1833 9281
rect -1775 9219 -1770 9281
rect -1887 9183 -1770 9219
rect -3113 9151 -2713 9157
rect -3275 9117 -3101 9151
rect -2725 9117 -2713 9151
rect -3806 9094 -3406 9100
rect -3952 9060 -3794 9094
rect -3418 9060 -3406 9094
rect -3952 8858 -3909 9060
rect -3806 9054 -3406 9060
rect -3806 8976 -3406 8982
rect -3806 8942 -3794 8976
rect -3418 8942 -3406 8976
rect -3806 8936 -3406 8942
rect -3275 8915 -3237 9117
rect -3113 9111 -2713 9117
rect -3113 9033 -2713 9039
rect -3113 8999 -3101 9033
rect -2725 8999 -2713 9033
rect -3113 8993 -2713 8999
rect -2548 8945 -2497 8962
rect -3113 8915 -2713 8921
rect -3275 8881 -3101 8915
rect -2725 8881 -2713 8915
rect -2548 8911 -2537 8945
rect -2503 8911 -2497 8945
rect -2548 8895 -2497 8911
rect -3113 8875 -2713 8881
rect -3806 8858 -3406 8864
rect -3952 8824 -3794 8858
rect -3418 8824 -3406 8858
rect -3952 8493 -3909 8824
rect -3806 8818 -3406 8824
rect -3594 8735 -3418 8818
rect -2553 8782 -2510 8895
rect -3606 8729 -3406 8735
rect -3606 8695 -3594 8729
rect -3418 8695 -3406 8729
rect -3606 8689 -3406 8695
rect -3255 8643 -3189 8655
rect -3606 8611 -3406 8617
rect -3606 8577 -3594 8611
rect -3418 8577 -3337 8611
rect -3255 8589 -3249 8643
rect -3195 8589 -3189 8643
rect -3255 8577 -3189 8589
rect -3606 8571 -3406 8577
rect -3372 8509 -3337 8577
rect -2554 8509 -2509 8782
rect -2469 8671 -2420 9158
rect -2381 9151 -1981 9157
rect -1887 9151 -1855 9183
rect -2381 9117 -2369 9151
rect -1993 9117 -1855 9151
rect -2381 9111 -1981 9117
rect -2381 9033 -1981 9039
rect -2381 8999 -2369 9033
rect -1993 8999 -1981 9033
rect -2381 8993 -1981 8999
rect -2481 8655 -2419 8671
rect -2481 8621 -2469 8655
rect -2435 8621 -2419 8655
rect -2481 8615 -2419 8621
rect -2381 8627 -2181 8633
rect -1887 8627 -1855 9117
rect -2381 8593 -2369 8627
rect -2193 8594 -1855 8627
rect -2193 8593 -2181 8594
rect -2381 8587 -2181 8593
rect -2381 8509 -2181 8515
rect -3606 8493 -3406 8499
rect -3952 8459 -3594 8493
rect -3418 8459 -3406 8493
rect -3606 8453 -3406 8459
rect -3372 8475 -2369 8509
rect -2193 8475 -2181 8509
rect -3606 8375 -3406 8381
rect -3372 8375 -3337 8475
rect -2381 8469 -2181 8475
rect -3606 8341 -3594 8375
rect -3418 8341 -3337 8375
rect -2703 8411 -2589 8423
rect -3606 8335 -3406 8341
rect -2703 8309 -2697 8411
rect -2595 8309 -2589 8411
rect -2703 8297 -2589 8309
rect -1216 8153 -1135 12315
rect -3255 8074 -1135 8153
rect -3606 7981 -3406 7987
rect -3606 7947 -3594 7981
rect -3418 7947 -3337 7981
rect -3606 7941 -3406 7947
rect -3606 7863 -3406 7869
rect -3952 7829 -3594 7863
rect -3418 7829 -3406 7863
rect -3952 7497 -3909 7829
rect -3606 7823 -3406 7829
rect -3372 7856 -3337 7947
rect -3255 7973 -3188 8074
rect -3065 7974 -2993 7989
rect -3255 7962 -3189 7973
rect -3065 7971 -3059 7974
rect -2999 7971 -2993 7974
rect -3068 7910 -3059 7971
rect -2999 7910 -2992 7971
rect -3065 7908 -3059 7910
rect -2999 7908 -2993 7910
rect -3065 7896 -2993 7908
rect -3255 7886 -3189 7896
rect -2381 7856 -2181 7862
rect -3372 7822 -2369 7856
rect -2193 7822 -2181 7856
rect -3606 7745 -3406 7751
rect -3606 7711 -3594 7745
rect -3418 7711 -3406 7745
rect -3606 7705 -3406 7711
rect -3606 7627 -3406 7633
rect -3606 7593 -3594 7627
rect -3418 7593 -3406 7627
rect -3606 7587 -3406 7593
rect -3594 7503 -3418 7587
rect -3113 7554 -2713 7560
rect -3275 7520 -3101 7554
rect -2725 7520 -2713 7554
rect -2553 7540 -2510 7822
rect -2381 7816 -2181 7822
rect -2381 7739 -2181 7744
rect -2381 7738 -1855 7739
rect -2482 7709 -2420 7715
rect -2482 7675 -2470 7709
rect -2436 7675 -2420 7709
rect -2381 7704 -2369 7738
rect -2193 7705 -1855 7738
rect -2193 7704 -2181 7705
rect -2381 7698 -2181 7704
rect -2482 7659 -2420 7675
rect -3806 7497 -3406 7503
rect -3952 7463 -3794 7497
rect -3418 7463 -3406 7497
rect -3952 7261 -3909 7463
rect -3806 7457 -3406 7463
rect -3806 7379 -3406 7385
rect -3806 7345 -3794 7379
rect -3418 7345 -3337 7379
rect -3806 7339 -3406 7345
rect -3806 7261 -3406 7267
rect -3952 7227 -3794 7261
rect -3418 7227 -3406 7261
rect -3952 7192 -3909 7227
rect -3806 7221 -3406 7227
rect -4035 7164 -3909 7192
rect -4057 7154 -3909 7164
rect -4003 7100 -3909 7154
rect -3806 7143 -3406 7149
rect -3372 7143 -3337 7345
rect -3275 7318 -3237 7520
rect -3113 7514 -2713 7520
rect -2548 7524 -2497 7540
rect -2548 7490 -2537 7524
rect -2503 7490 -2497 7524
rect -2548 7473 -2497 7490
rect -3113 7436 -2713 7442
rect -3113 7402 -3101 7436
rect -2725 7402 -2713 7436
rect -3113 7396 -2713 7402
rect -3113 7318 -2713 7324
rect -3275 7284 -3101 7318
rect -2725 7284 -2713 7318
rect -3275 7143 -3237 7284
rect -3113 7278 -2713 7284
rect -2469 7274 -2420 7659
rect -2381 7436 -1981 7442
rect -2381 7402 -2369 7436
rect -1993 7402 -1981 7436
rect -2381 7396 -1981 7402
rect -2381 7318 -1981 7324
rect -2381 7284 -2369 7318
rect -1993 7284 -1981 7318
rect -2381 7278 -1981 7284
rect -2469 7258 -2412 7274
rect -2469 7224 -2453 7258
rect -2419 7224 -2412 7258
rect -2469 7208 -2412 7224
rect -1887 7246 -1855 7705
rect -1887 7212 -1770 7246
rect -3113 7200 -2713 7206
rect -3113 7166 -3101 7200
rect -2725 7166 -2713 7200
rect -3113 7160 -2713 7166
rect -2381 7200 -1981 7206
rect -2381 7166 -2369 7200
rect -1993 7166 -1981 7200
rect -2381 7160 -1981 7166
rect -3806 7109 -3794 7143
rect -3418 7109 -3237 7143
rect -3806 7103 -3406 7109
rect -4057 7090 -3909 7100
rect -4035 7058 -3909 7090
rect -3952 7025 -3909 7058
rect -3275 7082 -3237 7109
rect -2469 7140 -2410 7156
rect -2469 7106 -2454 7140
rect -2420 7106 -2410 7140
rect -2469 7089 -2410 7106
rect -1887 7150 -1833 7212
rect -1775 7150 -1770 7212
rect -1887 7114 -1770 7150
rect -3113 7082 -2713 7088
rect -3275 7048 -3101 7082
rect -2725 7048 -2713 7082
rect -3806 7025 -3406 7031
rect -3952 6991 -3794 7025
rect -3418 6991 -3406 7025
rect -3952 6789 -3909 6991
rect -3806 6985 -3406 6991
rect -3806 6907 -3406 6913
rect -3806 6873 -3794 6907
rect -3418 6873 -3406 6907
rect -3806 6867 -3406 6873
rect -3275 6846 -3237 7048
rect -3113 7042 -2713 7048
rect -3113 6964 -2713 6970
rect -3113 6930 -3101 6964
rect -2725 6930 -2713 6964
rect -3113 6924 -2713 6930
rect -2548 6876 -2497 6893
rect -3113 6846 -2713 6852
rect -3275 6812 -3101 6846
rect -2725 6812 -2713 6846
rect -2548 6842 -2537 6876
rect -2503 6842 -2497 6876
rect -2548 6826 -2497 6842
rect -3113 6806 -2713 6812
rect -3806 6789 -3406 6795
rect -3952 6755 -3794 6789
rect -3418 6755 -3406 6789
rect -3952 6424 -3909 6755
rect -3806 6749 -3406 6755
rect -3594 6666 -3418 6749
rect -2553 6713 -2510 6826
rect -3606 6660 -3406 6666
rect -3606 6626 -3594 6660
rect -3418 6626 -3406 6660
rect -3606 6620 -3406 6626
rect -3255 6574 -3189 6586
rect -3606 6542 -3406 6548
rect -3606 6508 -3594 6542
rect -3418 6508 -3337 6542
rect -3255 6520 -3249 6574
rect -3195 6520 -3189 6574
rect -3255 6508 -3189 6520
rect -3606 6502 -3406 6508
rect -3372 6440 -3337 6508
rect -2554 6440 -2509 6713
rect -2469 6602 -2420 7089
rect -2381 7082 -1981 7088
rect -1887 7082 -1855 7114
rect -2381 7048 -2369 7082
rect -1993 7048 -1855 7082
rect -2381 7042 -1981 7048
rect -2381 6964 -1981 6970
rect -2381 6930 -2369 6964
rect -1993 6930 -1981 6964
rect -2381 6924 -1981 6930
rect -2481 6586 -2419 6602
rect -2481 6552 -2469 6586
rect -2435 6552 -2419 6586
rect -2481 6546 -2419 6552
rect -2381 6558 -2181 6564
rect -1887 6558 -1855 7048
rect -2381 6524 -2369 6558
rect -2193 6525 -1855 6558
rect -2193 6524 -2181 6525
rect -2381 6518 -2181 6524
rect -2381 6440 -2181 6446
rect -3606 6424 -3406 6430
rect -3952 6390 -3594 6424
rect -3418 6390 -3406 6424
rect -3606 6384 -3406 6390
rect -3372 6406 -2369 6440
rect -2193 6406 -2181 6440
rect -3606 6306 -3406 6312
rect -3372 6306 -3337 6406
rect -2381 6400 -2181 6406
rect -3606 6272 -3594 6306
rect -3418 6272 -3337 6306
rect -2703 6342 -2589 6354
rect -3606 6266 -3406 6272
rect -2703 6240 -2697 6342
rect -2595 6240 -2589 6342
rect -2703 6228 -2589 6240
rect -1077 6099 -998 21941
rect -3257 6087 -998 6099
rect -3257 6025 -1077 6087
rect -1011 6025 -998 6087
rect -3257 6011 -998 6025
rect -3608 5913 -3408 5919
rect -3608 5879 -3596 5913
rect -3420 5879 -3339 5913
rect -3608 5873 -3408 5879
rect -3608 5795 -3408 5801
rect -3954 5761 -3596 5795
rect -3420 5761 -3408 5795
rect -3954 5429 -3911 5761
rect -3608 5755 -3408 5761
rect -3374 5788 -3339 5879
rect -3257 5894 -3191 6011
rect -3067 5906 -2995 5924
rect -3067 5904 -3061 5906
rect -3001 5904 -2995 5906
rect -3069 5842 -3061 5904
rect -3001 5842 -2993 5904
rect -3067 5840 -3061 5842
rect -3001 5840 -2995 5842
rect -3067 5828 -2995 5840
rect -3257 5818 -3191 5828
rect -2383 5788 -2183 5794
rect -3374 5754 -2371 5788
rect -2195 5754 -2183 5788
rect -3608 5677 -3408 5683
rect -3608 5643 -3596 5677
rect -3420 5643 -3408 5677
rect -3608 5637 -3408 5643
rect -3608 5559 -3408 5565
rect -3608 5525 -3596 5559
rect -3420 5525 -3408 5559
rect -3608 5519 -3408 5525
rect -3596 5435 -3420 5519
rect -3115 5486 -2715 5492
rect -3277 5452 -3103 5486
rect -2727 5452 -2715 5486
rect -2555 5472 -2512 5754
rect -2383 5748 -2183 5754
rect -2383 5671 -2183 5676
rect -2383 5670 -1857 5671
rect -2484 5641 -2422 5647
rect -2484 5607 -2472 5641
rect -2438 5607 -2422 5641
rect -2383 5636 -2371 5670
rect -2195 5637 -1857 5670
rect -2195 5636 -2183 5637
rect -2383 5630 -2183 5636
rect -2484 5591 -2422 5607
rect -3808 5429 -3408 5435
rect -3954 5395 -3796 5429
rect -3420 5395 -3408 5429
rect -3954 5193 -3911 5395
rect -3808 5389 -3408 5395
rect -3808 5311 -3408 5317
rect -3808 5277 -3796 5311
rect -3420 5277 -3339 5311
rect -3808 5271 -3408 5277
rect -3808 5193 -3408 5199
rect -3954 5159 -3796 5193
rect -3420 5159 -3408 5193
rect -3954 5124 -3911 5159
rect -3808 5153 -3408 5159
rect -4037 5096 -3911 5124
rect -4059 5086 -3911 5096
rect -4005 5032 -3911 5086
rect -3808 5075 -3408 5081
rect -3374 5075 -3339 5277
rect -3277 5250 -3239 5452
rect -3115 5446 -2715 5452
rect -2550 5456 -2499 5472
rect -2550 5422 -2539 5456
rect -2505 5422 -2499 5456
rect -2550 5405 -2499 5422
rect -3115 5368 -2715 5374
rect -3115 5334 -3103 5368
rect -2727 5334 -2715 5368
rect -3115 5328 -2715 5334
rect -3115 5250 -2715 5256
rect -3277 5216 -3103 5250
rect -2727 5216 -2715 5250
rect -3277 5075 -3239 5216
rect -3115 5210 -2715 5216
rect -2471 5206 -2422 5591
rect -2383 5368 -1983 5374
rect -2383 5334 -2371 5368
rect -1995 5334 -1983 5368
rect -2383 5328 -1983 5334
rect -2383 5250 -1983 5256
rect -2383 5216 -2371 5250
rect -1995 5216 -1983 5250
rect -2383 5210 -1983 5216
rect -2471 5190 -2414 5206
rect -2471 5156 -2455 5190
rect -2421 5156 -2414 5190
rect -2471 5140 -2414 5156
rect -1889 5178 -1857 5637
rect -1889 5144 -1772 5178
rect -3115 5132 -2715 5138
rect -3115 5098 -3103 5132
rect -2727 5098 -2715 5132
rect -3115 5092 -2715 5098
rect -2383 5132 -1983 5138
rect -2383 5098 -2371 5132
rect -1995 5098 -1983 5132
rect -2383 5092 -1983 5098
rect -3808 5041 -3796 5075
rect -3420 5041 -3239 5075
rect -3808 5035 -3408 5041
rect -4059 5022 -3911 5032
rect -4037 4990 -3911 5022
rect -3954 4957 -3911 4990
rect -3277 5014 -3239 5041
rect -2471 5072 -2412 5088
rect -2471 5038 -2456 5072
rect -2422 5038 -2412 5072
rect -2471 5021 -2412 5038
rect -1889 5082 -1835 5144
rect -1777 5082 -1772 5144
rect -1889 5046 -1772 5082
rect -3115 5014 -2715 5020
rect -3277 4980 -3103 5014
rect -2727 4980 -2715 5014
rect -3808 4957 -3408 4963
rect -3954 4923 -3796 4957
rect -3420 4923 -3408 4957
rect -3954 4721 -3911 4923
rect -3808 4917 -3408 4923
rect -3808 4839 -3408 4845
rect -3808 4805 -3796 4839
rect -3420 4805 -3408 4839
rect -3808 4799 -3408 4805
rect -3277 4778 -3239 4980
rect -3115 4974 -2715 4980
rect -3115 4896 -2715 4902
rect -3115 4862 -3103 4896
rect -2727 4862 -2715 4896
rect -3115 4856 -2715 4862
rect -2550 4808 -2499 4825
rect -3115 4778 -2715 4784
rect -3277 4744 -3103 4778
rect -2727 4744 -2715 4778
rect -2550 4774 -2539 4808
rect -2505 4774 -2499 4808
rect -2550 4758 -2499 4774
rect -3115 4738 -2715 4744
rect -3808 4721 -3408 4727
rect -3954 4687 -3796 4721
rect -3420 4687 -3408 4721
rect -3954 4356 -3911 4687
rect -3808 4681 -3408 4687
rect -3596 4598 -3420 4681
rect -2555 4645 -2512 4758
rect -3608 4592 -3408 4598
rect -3608 4558 -3596 4592
rect -3420 4558 -3408 4592
rect -3608 4552 -3408 4558
rect -3257 4506 -3191 4518
rect -3608 4474 -3408 4480
rect -3608 4440 -3596 4474
rect -3420 4440 -3339 4474
rect -3257 4452 -3251 4506
rect -3197 4452 -3191 4506
rect -3257 4440 -3191 4452
rect -3608 4434 -3408 4440
rect -3374 4372 -3339 4440
rect -2556 4372 -2511 4645
rect -2471 4534 -2422 5021
rect -2383 5014 -1983 5020
rect -1889 5014 -1857 5046
rect -2383 4980 -2371 5014
rect -1995 4980 -1857 5014
rect -2383 4974 -1983 4980
rect -2383 4896 -1983 4902
rect -2383 4862 -2371 4896
rect -1995 4862 -1983 4896
rect -2383 4856 -1983 4862
rect -2483 4518 -2421 4534
rect -2483 4484 -2471 4518
rect -2437 4484 -2421 4518
rect -2483 4478 -2421 4484
rect -2383 4490 -2183 4496
rect -1889 4490 -1857 4980
rect -2383 4456 -2371 4490
rect -2195 4457 -1857 4490
rect -2195 4456 -2183 4457
rect -2383 4450 -2183 4456
rect -2383 4372 -2183 4378
rect -3608 4356 -3408 4362
rect -3954 4322 -3596 4356
rect -3420 4322 -3408 4356
rect -3608 4316 -3408 4322
rect -3374 4338 -2371 4372
rect -2195 4338 -2183 4372
rect -3608 4238 -3408 4244
rect -3374 4238 -3339 4338
rect -2383 4332 -2183 4338
rect -3608 4204 -3596 4238
rect -3420 4204 -3339 4238
rect -2705 4274 -2591 4286
rect -3608 4198 -3408 4204
rect -2705 4172 -2699 4274
rect -2597 4172 -2591 4274
rect -2705 4160 -2591 4172
rect -933 4019 -858 22381
rect -3255 4008 -858 4019
rect -3255 3953 -1224 4008
rect -1154 3953 -858 4008
rect -3255 3941 -858 3953
rect -3606 3844 -3406 3850
rect -3606 3810 -3594 3844
rect -3418 3810 -3337 3844
rect -3606 3804 -3406 3810
rect -3606 3726 -3406 3732
rect -3952 3692 -3594 3726
rect -3418 3692 -3406 3726
rect -3952 3360 -3909 3692
rect -3606 3686 -3406 3692
rect -3372 3719 -3337 3810
rect -3255 3825 -3189 3941
rect -3065 3837 -2993 3858
rect -3065 3771 -3059 3837
rect -2999 3771 -2993 3837
rect -3065 3759 -2993 3771
rect -3255 3749 -3189 3759
rect -2381 3719 -2181 3725
rect -3372 3685 -2369 3719
rect -2193 3685 -2181 3719
rect -3606 3608 -3406 3614
rect -3606 3574 -3594 3608
rect -3418 3574 -3406 3608
rect -3606 3568 -3406 3574
rect -3606 3490 -3406 3496
rect -3606 3456 -3594 3490
rect -3418 3456 -3406 3490
rect -3606 3450 -3406 3456
rect -3594 3366 -3418 3450
rect -3113 3417 -2713 3423
rect -3275 3383 -3101 3417
rect -2725 3383 -2713 3417
rect -2553 3403 -2510 3685
rect -2381 3679 -2181 3685
rect -2381 3602 -2181 3607
rect -2381 3601 -1855 3602
rect -2482 3572 -2420 3578
rect -2482 3538 -2470 3572
rect -2436 3538 -2420 3572
rect -2381 3567 -2369 3601
rect -2193 3568 -1855 3601
rect -2193 3567 -2181 3568
rect -2381 3561 -2181 3567
rect -2482 3522 -2420 3538
rect -3806 3360 -3406 3366
rect -3952 3326 -3794 3360
rect -3418 3326 -3406 3360
rect -3952 3124 -3909 3326
rect -3806 3320 -3406 3326
rect -3806 3242 -3406 3248
rect -3806 3208 -3794 3242
rect -3418 3208 -3337 3242
rect -3806 3202 -3406 3208
rect -3806 3124 -3406 3130
rect -3952 3090 -3794 3124
rect -3418 3090 -3406 3124
rect -3952 3055 -3909 3090
rect -3806 3084 -3406 3090
rect -4035 3027 -3909 3055
rect -4057 3017 -3909 3027
rect -4003 2963 -3909 3017
rect -3806 3006 -3406 3012
rect -3372 3006 -3337 3208
rect -3275 3181 -3237 3383
rect -3113 3377 -2713 3383
rect -2548 3387 -2497 3403
rect -2548 3353 -2537 3387
rect -2503 3353 -2497 3387
rect -2548 3336 -2497 3353
rect -3113 3299 -2713 3305
rect -3113 3265 -3101 3299
rect -2725 3265 -2713 3299
rect -3113 3259 -2713 3265
rect -3113 3181 -2713 3187
rect -3275 3147 -3101 3181
rect -2725 3147 -2713 3181
rect -3275 3006 -3237 3147
rect -3113 3141 -2713 3147
rect -2469 3137 -2420 3522
rect -2381 3299 -1981 3305
rect -2381 3265 -2369 3299
rect -1993 3265 -1981 3299
rect -2381 3259 -1981 3265
rect -2381 3181 -1981 3187
rect -2381 3147 -2369 3181
rect -1993 3147 -1981 3181
rect -2381 3141 -1981 3147
rect -2469 3121 -2412 3137
rect -2469 3087 -2453 3121
rect -2419 3087 -2412 3121
rect -2469 3071 -2412 3087
rect -1887 3109 -1855 3568
rect -1887 3075 -1770 3109
rect -3113 3063 -2713 3069
rect -3113 3029 -3101 3063
rect -2725 3029 -2713 3063
rect -3113 3023 -2713 3029
rect -2381 3063 -1981 3069
rect -2381 3029 -2369 3063
rect -1993 3029 -1981 3063
rect -2381 3023 -1981 3029
rect -3806 2972 -3794 3006
rect -3418 2972 -3237 3006
rect -3806 2966 -3406 2972
rect -4057 2953 -3909 2963
rect -4035 2921 -3909 2953
rect -3952 2888 -3909 2921
rect -3275 2945 -3237 2972
rect -2469 3003 -2410 3019
rect -2469 2969 -2454 3003
rect -2420 2969 -2410 3003
rect -2469 2952 -2410 2969
rect -1887 3013 -1833 3075
rect -1775 3013 -1770 3075
rect -1887 2977 -1770 3013
rect -3113 2945 -2713 2951
rect -3275 2911 -3101 2945
rect -2725 2911 -2713 2945
rect -3806 2888 -3406 2894
rect -3952 2854 -3794 2888
rect -3418 2854 -3406 2888
rect -3952 2652 -3909 2854
rect -3806 2848 -3406 2854
rect -3806 2770 -3406 2776
rect -3806 2736 -3794 2770
rect -3418 2736 -3406 2770
rect -3806 2730 -3406 2736
rect -3275 2709 -3237 2911
rect -3113 2905 -2713 2911
rect -3113 2827 -2713 2833
rect -3113 2793 -3101 2827
rect -2725 2793 -2713 2827
rect -3113 2787 -2713 2793
rect -2548 2739 -2497 2756
rect -3113 2709 -2713 2715
rect -3275 2675 -3101 2709
rect -2725 2675 -2713 2709
rect -2548 2705 -2537 2739
rect -2503 2705 -2497 2739
rect -2548 2689 -2497 2705
rect -3113 2669 -2713 2675
rect -3806 2652 -3406 2658
rect -3952 2618 -3794 2652
rect -3418 2618 -3406 2652
rect -3952 2287 -3909 2618
rect -3806 2612 -3406 2618
rect -3594 2529 -3418 2612
rect -2553 2576 -2510 2689
rect -3606 2523 -3406 2529
rect -3606 2489 -3594 2523
rect -3418 2489 -3406 2523
rect -3606 2483 -3406 2489
rect -3255 2437 -3189 2449
rect -3606 2405 -3406 2411
rect -3606 2371 -3594 2405
rect -3418 2371 -3337 2405
rect -3255 2383 -3249 2437
rect -3195 2383 -3189 2437
rect -3255 2371 -3189 2383
rect -3606 2365 -3406 2371
rect -3372 2303 -3337 2371
rect -2554 2303 -2509 2576
rect -2469 2465 -2420 2952
rect -2381 2945 -1981 2951
rect -1887 2945 -1855 2977
rect -2381 2911 -2369 2945
rect -1993 2911 -1855 2945
rect -2381 2905 -1981 2911
rect -2381 2827 -1981 2833
rect -2381 2793 -2369 2827
rect -1993 2793 -1981 2827
rect -2381 2787 -1981 2793
rect -2481 2449 -2419 2465
rect -2481 2415 -2469 2449
rect -2435 2415 -2419 2449
rect -2481 2409 -2419 2415
rect -2381 2421 -2181 2427
rect -1887 2421 -1855 2911
rect -2381 2387 -2369 2421
rect -2193 2388 -1855 2421
rect -2193 2387 -2181 2388
rect -2381 2381 -2181 2387
rect -2381 2303 -2181 2309
rect -3606 2287 -3406 2293
rect -3952 2253 -3594 2287
rect -3418 2253 -3406 2287
rect -3606 2247 -3406 2253
rect -3372 2269 -2369 2303
rect -2193 2269 -2181 2303
rect -3606 2169 -3406 2175
rect -3372 2169 -3337 2269
rect -2381 2263 -2181 2269
rect -3606 2135 -3594 2169
rect -3418 2135 -3337 2169
rect -2703 2205 -2589 2217
rect -3606 2129 -3406 2135
rect -2703 2103 -2697 2205
rect -2595 2103 -2589 2205
rect -2703 2091 -2589 2103
rect -798 1940 -723 22802
rect -661 22993 -588 23232
rect -661 16334 -586 22993
rect -661 16282 -651 16334
rect -590 16282 -580 16334
rect -661 14246 -586 16282
rect -514 15963 -429 23650
rect -349 16140 -276 24073
rect -216 16296 -143 24303
rect -86 24616 -14 24955
rect -86 16447 -13 24616
rect 52 16599 125 25376
rect 194 22750 288 25808
rect 354 22940 432 26227
rect 491 23084 572 26648
rect 5330 24780 5423 26674
rect 5486 26615 5952 26637
rect 6240 26615 6306 26711
rect 8071 26721 8077 26897
rect 8111 26721 8117 26897
rect 8071 26709 8117 26721
rect 8189 26897 8235 26909
rect 8189 26721 8195 26897
rect 8229 26721 8235 26897
rect 8189 26709 8235 26721
rect 8307 26897 8353 26909
rect 8307 26721 8313 26897
rect 8347 26721 8353 26897
rect 8307 26709 8353 26721
rect 8425 26897 8471 26909
rect 8425 26721 8431 26897
rect 8465 26842 8471 26897
rect 8590 26897 8636 26909
rect 8590 26842 8596 26897
rect 8465 26754 8596 26842
rect 8465 26721 8471 26754
rect 8425 26709 8471 26721
rect 8590 26721 8596 26754
rect 8630 26721 8636 26897
rect 8590 26709 8636 26721
rect 8708 26897 8754 26909
rect 8708 26721 8714 26897
rect 8748 26721 8754 26897
rect 8708 26709 8754 26721
rect 8826 26897 8872 26909
rect 8826 26721 8832 26897
rect 8866 26721 8872 26897
rect 8826 26709 8872 26721
rect 8944 26897 8990 26909
rect 8944 26721 8950 26897
rect 8984 26721 8990 26897
rect 8944 26709 8990 26721
rect 8077 26670 8111 26709
rect 8313 26670 8347 26709
rect 8077 26635 8347 26670
rect 8714 26671 8747 26709
rect 8950 26671 8983 26709
rect 8714 26635 8983 26671
rect 5486 26567 6306 26615
rect 8111 26634 8347 26635
rect 5486 26536 5952 26567
rect 8111 26560 8243 26634
rect 5486 26280 5591 26536
rect 8101 26452 8111 26560
rect 8243 26452 8253 26560
rect 5486 26174 5549 26280
rect 5661 26174 5671 26280
rect 6253 26256 6473 26276
rect 5486 26163 5635 26174
rect 5486 24986 5591 26163
rect 6253 26148 6297 26256
rect 6429 26148 6473 26256
rect 6253 26106 6473 26148
rect 9051 26121 9113 27692
rect 9303 27684 9349 27696
rect 9303 27308 9309 27684
rect 9343 27308 9349 27684
rect 9303 27296 9349 27308
rect 9421 27684 9467 27696
rect 9421 27308 9427 27684
rect 9461 27308 9467 27684
rect 9421 27296 9467 27308
rect 9539 27684 9585 27696
rect 9539 27308 9545 27684
rect 9579 27308 9585 27684
rect 9539 27296 9585 27308
rect 9657 27684 9703 27696
rect 9657 27308 9663 27684
rect 9697 27308 9703 27684
rect 9657 27296 9703 27308
rect 9775 27684 9821 27696
rect 9775 27308 9781 27684
rect 9815 27308 9821 27684
rect 9775 27296 9821 27308
rect 9893 27684 9939 27696
rect 9893 27308 9899 27684
rect 9933 27308 9939 27684
rect 9893 27296 9939 27308
rect 10011 27684 10057 27696
rect 10011 27308 10017 27684
rect 10051 27308 10057 27684
rect 12356 27723 13333 27753
rect 12356 27617 12388 27723
rect 12592 27617 12624 27723
rect 12828 27617 12860 27723
rect 13064 27617 13096 27723
rect 13299 27617 13333 27723
rect 12349 27605 12395 27617
rect 12349 27429 12355 27605
rect 12389 27429 12395 27605
rect 12349 27417 12395 27429
rect 12467 27605 12513 27617
rect 12467 27429 12473 27605
rect 12507 27429 12513 27605
rect 12467 27417 12513 27429
rect 12585 27605 12631 27617
rect 12585 27429 12591 27605
rect 12625 27429 12631 27605
rect 12585 27417 12631 27429
rect 12703 27605 12749 27617
rect 12703 27429 12709 27605
rect 12743 27429 12749 27605
rect 12703 27417 12749 27429
rect 12821 27605 12867 27617
rect 12821 27429 12827 27605
rect 12861 27429 12867 27605
rect 12821 27417 12867 27429
rect 12939 27605 12985 27617
rect 12939 27429 12945 27605
rect 12979 27429 12985 27605
rect 12939 27417 12985 27429
rect 13057 27605 13103 27617
rect 13057 27429 13063 27605
rect 13097 27429 13103 27605
rect 13057 27417 13103 27429
rect 13175 27605 13221 27617
rect 13175 27429 13181 27605
rect 13215 27429 13221 27605
rect 13175 27417 13221 27429
rect 13293 27605 13339 27617
rect 13293 27429 13299 27605
rect 13333 27429 13339 27605
rect 13293 27417 13339 27429
rect 13411 27605 13457 27617
rect 13411 27429 13417 27605
rect 13451 27429 13457 27605
rect 13411 27417 13457 27429
rect 10011 27296 10057 27308
rect 12472 27323 12508 27417
rect 12708 27323 12744 27417
rect 12944 27324 12980 27417
rect 13106 27369 13172 27376
rect 13106 27335 13122 27369
rect 13156 27335 13172 27369
rect 13106 27324 13172 27335
rect 12944 27323 13172 27324
rect 9309 27254 9343 27296
rect 9545 27254 9579 27296
rect 9309 27226 9579 27254
rect 9663 27255 9697 27296
rect 9899 27255 9933 27296
rect 9663 27226 9933 27255
rect 9309 27178 9343 27226
rect 9309 27148 9372 27178
rect 9337 27056 9372 27148
rect 9844 27118 9944 27139
rect 9844 27064 9858 27118
rect 9923 27064 9944 27118
rect 9844 27059 9944 27064
rect 10017 27113 10051 27296
rect 12472 27294 13172 27323
rect 12472 27293 13054 27294
rect 12592 27180 12626 27293
rect 12988 27252 13054 27293
rect 12988 27218 13004 27252
rect 13038 27218 13054 27252
rect 12988 27211 13054 27218
rect 13416 27212 13451 27417
rect 13623 27212 13690 27802
rect 15382 27779 15423 27811
rect 15669 27807 15679 27873
rect 15735 27807 15745 27873
rect 16415 27849 16425 27957
rect 16557 27894 16567 27957
rect 19286 27898 19506 27918
rect 16557 27883 16569 27894
rect 16557 27849 16570 27883
rect 16425 27811 16570 27849
rect 16529 27783 16570 27811
rect 14798 27751 15068 27779
rect 14539 27685 14549 27751
rect 14615 27685 14625 27751
rect 14798 27689 14832 27751
rect 15034 27689 15068 27751
rect 15152 27751 15423 27779
rect 15940 27755 16210 27783
rect 15152 27689 15186 27751
rect 15388 27689 15423 27751
rect 15564 27739 15735 27755
rect 15564 27705 15695 27739
rect 15729 27705 15735 27739
rect 15564 27689 15735 27705
rect 15940 27693 15974 27755
rect 16176 27693 16210 27755
rect 16294 27755 16570 27783
rect 16294 27693 16328 27755
rect 16530 27693 16570 27755
rect 19286 27790 19330 27898
rect 19462 27790 19506 27898
rect 21083 27856 21139 27864
rect 19286 27748 19506 27790
rect 20157 27848 21139 27856
rect 20157 27814 21099 27848
rect 21133 27814 21139 27848
rect 21802 27844 21812 27952
rect 21944 27889 21954 27952
rect 21944 27878 21956 27889
rect 21944 27844 21957 27878
rect 22213 27868 22269 27870
rect 20157 27798 21139 27814
rect 21812 27806 21957 27844
rect 20157 27797 21136 27798
rect 14674 27677 14720 27689
rect 14674 27301 14680 27677
rect 14714 27301 14720 27677
rect 14674 27289 14720 27301
rect 14792 27677 14838 27689
rect 14792 27301 14798 27677
rect 14832 27301 14838 27677
rect 14792 27289 14838 27301
rect 14910 27677 14956 27689
rect 14910 27301 14916 27677
rect 14950 27301 14956 27677
rect 14910 27289 14956 27301
rect 15028 27677 15074 27689
rect 15028 27301 15034 27677
rect 15068 27301 15074 27677
rect 15028 27289 15074 27301
rect 15146 27677 15192 27689
rect 15146 27301 15152 27677
rect 15186 27301 15192 27677
rect 15146 27289 15192 27301
rect 15264 27677 15310 27689
rect 15264 27301 15270 27677
rect 15304 27301 15310 27677
rect 15264 27289 15310 27301
rect 15382 27677 15428 27689
rect 15382 27301 15388 27677
rect 15422 27301 15428 27677
rect 15382 27289 15428 27301
rect 13416 27184 13690 27212
rect 13062 27180 13690 27184
rect 12586 27168 12632 27180
rect 11019 27127 11126 27129
rect 10017 27059 10126 27113
rect 9337 27020 9564 27056
rect 9337 26913 9372 27020
rect 9498 26986 9564 27020
rect 9498 26952 9514 26986
rect 9548 26952 9564 26986
rect 9845 27044 9942 27059
rect 9845 26977 9902 27044
rect 9498 26946 9564 26952
rect 9739 26941 10008 26977
rect 9739 26913 9772 26941
rect 9975 26913 10008 26941
rect 10092 26913 10126 27059
rect 10943 27052 10953 27127
rect 11021 27052 11126 27127
rect 10970 27051 11126 27052
rect 9213 26901 9259 26913
rect 9213 26725 9219 26901
rect 9253 26725 9259 26901
rect 9213 26713 9259 26725
rect 9331 26901 9377 26913
rect 9331 26725 9337 26901
rect 9371 26725 9377 26901
rect 9331 26713 9377 26725
rect 9449 26901 9495 26913
rect 9449 26725 9455 26901
rect 9489 26725 9495 26901
rect 9449 26713 9495 26725
rect 9567 26901 9613 26913
rect 9567 26725 9573 26901
rect 9607 26846 9613 26901
rect 9732 26901 9778 26913
rect 9732 26846 9738 26901
rect 9607 26758 9738 26846
rect 9607 26725 9613 26758
rect 9567 26713 9613 26725
rect 9732 26725 9738 26758
rect 9772 26725 9778 26901
rect 9732 26713 9778 26725
rect 9850 26901 9896 26913
rect 9850 26725 9856 26901
rect 9890 26725 9896 26901
rect 9850 26713 9896 26725
rect 9968 26901 10014 26913
rect 9968 26725 9974 26901
rect 10008 26725 10014 26901
rect 9968 26713 10014 26725
rect 10086 26901 10132 26913
rect 10086 26725 10092 26901
rect 10126 26725 10132 26901
rect 10086 26713 10132 26725
rect 9219 26674 9253 26713
rect 9455 26674 9489 26713
rect 9219 26638 9489 26674
rect 9856 26675 9889 26713
rect 10092 26675 10125 26713
rect 9856 26639 10125 26675
rect 9219 26637 9385 26638
rect 9253 26558 9385 26637
rect 9243 26450 9253 26558
rect 9385 26450 9395 26558
rect 5857 26076 6834 26106
rect 9051 26104 9114 26121
rect 8976 26100 9114 26104
rect 5857 25970 5889 26076
rect 6093 25970 6125 26076
rect 6329 25970 6361 26076
rect 6565 25970 6597 26076
rect 6800 25970 6834 26076
rect 7144 26066 9114 26100
rect 7142 26037 9114 26066
rect 7142 26021 7188 26037
rect 8976 26035 9114 26037
rect 5850 25958 5896 25970
rect 5850 25782 5856 25958
rect 5890 25782 5896 25958
rect 5850 25770 5896 25782
rect 5968 25958 6014 25970
rect 5968 25782 5974 25958
rect 6008 25782 6014 25958
rect 5968 25770 6014 25782
rect 6086 25958 6132 25970
rect 6086 25782 6092 25958
rect 6126 25782 6132 25958
rect 6086 25770 6132 25782
rect 6204 25958 6250 25970
rect 6204 25782 6210 25958
rect 6244 25782 6250 25958
rect 6204 25770 6250 25782
rect 6322 25958 6368 25970
rect 6322 25782 6328 25958
rect 6362 25782 6368 25958
rect 6322 25770 6368 25782
rect 6440 25958 6486 25970
rect 6440 25782 6446 25958
rect 6480 25782 6486 25958
rect 6440 25770 6486 25782
rect 6558 25958 6604 25970
rect 6558 25782 6564 25958
rect 6598 25782 6604 25958
rect 6558 25770 6604 25782
rect 6676 25958 6722 25970
rect 6676 25782 6682 25958
rect 6716 25782 6722 25958
rect 6676 25770 6722 25782
rect 6794 25958 6840 25970
rect 6794 25782 6800 25958
rect 6834 25782 6840 25958
rect 6794 25770 6840 25782
rect 6912 25958 6958 25970
rect 6912 25782 6918 25958
rect 6952 25782 6958 25958
rect 6912 25770 6958 25782
rect 5973 25676 6009 25770
rect 6209 25676 6245 25770
rect 6445 25677 6481 25770
rect 6607 25722 6673 25729
rect 6607 25688 6623 25722
rect 6657 25688 6673 25722
rect 6607 25677 6673 25688
rect 6445 25676 6673 25677
rect 5973 25647 6673 25676
rect 5973 25646 6555 25647
rect 6093 25533 6127 25646
rect 6489 25605 6555 25646
rect 6489 25571 6505 25605
rect 6539 25571 6555 25605
rect 6489 25564 6555 25571
rect 6917 25552 6952 25770
rect 7141 25569 7188 26021
rect 8100 25805 8110 25913
rect 8242 25805 8252 25913
rect 9998 25805 10008 25913
rect 10140 25805 10150 25913
rect 8110 25765 8242 25805
rect 10008 25765 10140 25805
rect 8109 25699 8242 25765
rect 10007 25699 10140 25765
rect 7438 25656 8911 25699
rect 7141 25553 7187 25569
rect 7106 25552 7187 25553
rect 6917 25537 7187 25552
rect 6563 25533 7187 25537
rect 6087 25521 6133 25533
rect 5822 25043 5832 25161
rect 5950 25129 5960 25161
rect 6087 25145 6093 25521
rect 6127 25145 6133 25521
rect 6087 25133 6133 25145
rect 6205 25521 6251 25533
rect 6205 25145 6211 25521
rect 6245 25145 6251 25521
rect 6205 25133 6251 25145
rect 6323 25521 6369 25533
rect 6323 25145 6329 25521
rect 6363 25169 6369 25521
rect 6440 25521 6486 25533
rect 6440 25345 6446 25521
rect 6480 25345 6486 25521
rect 6440 25333 6486 25345
rect 6558 25521 7187 25533
rect 6558 25345 6564 25521
rect 6598 25509 7187 25521
rect 6598 25508 6840 25509
rect 6598 25345 6604 25508
rect 7106 25507 7187 25509
rect 7438 25353 7472 25656
rect 7804 25553 7838 25656
rect 8040 25553 8074 25656
rect 8276 25553 8310 25656
rect 8512 25553 8546 25656
rect 7798 25541 7844 25553
rect 6558 25333 6604 25345
rect 7314 25341 7360 25353
rect 6446 25217 6481 25333
rect 6577 25217 6685 25227
rect 6446 25169 6577 25217
rect 6363 25145 6577 25169
rect 6323 25133 6577 25145
rect 6329 25129 6577 25133
rect 5950 25101 5965 25129
rect 5950 25095 6202 25101
rect 5950 25061 6152 25095
rect 6186 25061 6202 25095
rect 5950 25045 6202 25061
rect 6254 25095 6320 25101
rect 6254 25061 6270 25095
rect 6304 25061 6320 25095
rect 6503 25085 6577 25129
rect 7314 25165 7320 25341
rect 7354 25165 7360 25341
rect 7314 25153 7360 25165
rect 7432 25341 7478 25353
rect 7432 25165 7438 25341
rect 7472 25165 7478 25341
rect 7432 25153 7478 25165
rect 7550 25341 7596 25353
rect 7550 25165 7556 25341
rect 7590 25165 7596 25341
rect 7550 25153 7596 25165
rect 7668 25341 7714 25353
rect 7798 25341 7804 25541
rect 7668 25165 7674 25341
rect 7708 25165 7804 25341
rect 7838 25165 7844 25541
rect 7668 25153 7714 25165
rect 7798 25153 7844 25165
rect 7916 25541 7962 25553
rect 7916 25165 7922 25541
rect 7956 25165 7962 25541
rect 7916 25153 7962 25165
rect 8034 25541 8080 25553
rect 8034 25165 8040 25541
rect 8074 25165 8080 25541
rect 8034 25153 8080 25165
rect 8152 25541 8198 25553
rect 8152 25165 8158 25541
rect 8192 25165 8198 25541
rect 8152 25153 8198 25165
rect 8270 25541 8316 25553
rect 8270 25165 8276 25541
rect 8310 25165 8316 25541
rect 8270 25153 8316 25165
rect 8388 25541 8434 25553
rect 8388 25165 8394 25541
rect 8428 25165 8434 25541
rect 8388 25153 8434 25165
rect 8506 25541 8552 25553
rect 8506 25165 8512 25541
rect 8546 25341 8552 25541
rect 8877 25353 8911 25656
rect 9336 25656 10809 25699
rect 9336 25353 9370 25656
rect 9702 25553 9736 25656
rect 9938 25553 9972 25656
rect 10174 25553 10208 25656
rect 10410 25553 10444 25656
rect 9696 25541 9742 25553
rect 8635 25341 8681 25353
rect 8546 25165 8641 25341
rect 8675 25165 8681 25341
rect 8506 25153 8552 25165
rect 8635 25153 8681 25165
rect 8753 25341 8799 25353
rect 8753 25165 8759 25341
rect 8793 25165 8799 25341
rect 8753 25153 8799 25165
rect 8871 25341 8917 25353
rect 8871 25165 8877 25341
rect 8911 25165 8917 25341
rect 8871 25153 8917 25165
rect 8989 25341 9035 25353
rect 8989 25165 8995 25341
rect 9029 25165 9035 25341
rect 8989 25153 9035 25165
rect 9212 25341 9258 25353
rect 9212 25165 9218 25341
rect 9252 25165 9258 25341
rect 9212 25153 9258 25165
rect 9330 25341 9376 25353
rect 9330 25165 9336 25341
rect 9370 25165 9376 25341
rect 9330 25153 9376 25165
rect 9448 25341 9494 25353
rect 9448 25165 9454 25341
rect 9488 25165 9494 25341
rect 9448 25153 9494 25165
rect 9566 25341 9612 25353
rect 9696 25341 9702 25541
rect 9566 25165 9572 25341
rect 9606 25165 9702 25341
rect 9736 25165 9742 25541
rect 9566 25153 9612 25165
rect 9696 25153 9742 25165
rect 9814 25541 9860 25553
rect 9814 25165 9820 25541
rect 9854 25165 9860 25541
rect 9814 25153 9860 25165
rect 9932 25541 9978 25553
rect 9932 25165 9938 25541
rect 9972 25165 9978 25541
rect 9932 25153 9978 25165
rect 10050 25541 10096 25553
rect 10050 25165 10056 25541
rect 10090 25165 10096 25541
rect 10050 25153 10096 25165
rect 10168 25541 10214 25553
rect 10168 25165 10174 25541
rect 10208 25165 10214 25541
rect 10168 25153 10214 25165
rect 10286 25541 10332 25553
rect 10286 25165 10292 25541
rect 10326 25165 10332 25541
rect 10286 25153 10332 25165
rect 10404 25541 10450 25553
rect 10404 25165 10410 25541
rect 10444 25341 10450 25541
rect 10775 25353 10809 25656
rect 10533 25341 10579 25353
rect 10444 25165 10539 25341
rect 10573 25165 10579 25341
rect 10404 25153 10450 25165
rect 10533 25153 10579 25165
rect 10651 25341 10697 25353
rect 10651 25165 10657 25341
rect 10691 25165 10697 25341
rect 10651 25153 10697 25165
rect 10769 25341 10815 25353
rect 10769 25165 10775 25341
rect 10809 25165 10815 25341
rect 10769 25153 10815 25165
rect 10887 25341 10933 25353
rect 10887 25165 10893 25341
rect 10927 25165 10933 25341
rect 11019 25307 11126 27051
rect 11414 26838 11703 26864
rect 11414 26694 11432 26838
rect 11668 26775 11703 26838
rect 12586 26792 12592 27168
rect 12626 26792 12632 27168
rect 12586 26780 12632 26792
rect 12704 27168 12750 27180
rect 12704 26792 12710 27168
rect 12744 26792 12750 27168
rect 12704 26780 12750 26792
rect 12822 27168 12868 27180
rect 12822 26792 12828 27168
rect 12862 26816 12868 27168
rect 12939 27168 12985 27180
rect 12939 26992 12945 27168
rect 12979 26992 12985 27168
rect 12939 26980 12985 26992
rect 13057 27168 13690 27180
rect 13057 26992 13063 27168
rect 13097 27155 13690 27168
rect 14680 27247 14714 27289
rect 14916 27247 14950 27289
rect 14680 27219 14950 27247
rect 15034 27248 15068 27289
rect 15270 27248 15304 27289
rect 15034 27219 15304 27248
rect 14680 27171 14714 27219
rect 13097 26992 13103 27155
rect 14680 27141 14743 27171
rect 13057 26980 13103 26992
rect 14708 27049 14743 27141
rect 14708 27013 14935 27049
rect 15205 27038 15215 27135
rect 15314 27038 15324 27135
rect 15388 27106 15422 27289
rect 15388 27052 15497 27106
rect 12945 26864 12980 26980
rect 14708 26906 14743 27013
rect 14869 26979 14935 27013
rect 14869 26945 14885 26979
rect 14919 26945 14935 26979
rect 15216 27037 15313 27038
rect 15216 26970 15273 27037
rect 14869 26939 14935 26945
rect 15110 26934 15379 26970
rect 15110 26906 15143 26934
rect 15346 26906 15379 26934
rect 15463 26906 15497 27052
rect 14584 26894 14630 26906
rect 13076 26864 13184 26874
rect 12945 26816 13076 26864
rect 12862 26792 13076 26816
rect 12822 26780 13076 26792
rect 12828 26776 13076 26780
rect 11668 26748 12464 26775
rect 11668 26742 12701 26748
rect 11668 26708 12651 26742
rect 12685 26708 12701 26742
rect 11668 26694 12701 26708
rect 11414 26692 12701 26694
rect 12753 26742 12819 26748
rect 12753 26708 12769 26742
rect 12803 26708 12819 26742
rect 13002 26732 13076 26776
rect 13076 26722 13184 26732
rect 11414 26676 12464 26692
rect 11414 26675 12401 26676
rect 11414 26671 11936 26675
rect 11414 26670 11703 26671
rect 11431 25307 11719 25310
rect 11019 25191 11719 25307
rect 11019 25188 11126 25191
rect 10887 25153 10933 25165
rect 6577 25075 6685 25085
rect 7320 25119 7354 25153
rect 7922 25119 7956 25153
rect 8158 25119 8192 25153
rect 7320 25084 7479 25119
rect 7922 25084 8192 25119
rect 8759 25119 8793 25153
rect 8995 25119 9029 25153
rect 8759 25084 9029 25119
rect 9218 25119 9252 25153
rect 9820 25119 9854 25153
rect 10056 25119 10090 25153
rect 9218 25084 9377 25119
rect 9820 25084 10090 25119
rect 10657 25119 10691 25153
rect 10893 25119 10927 25153
rect 10657 25084 10927 25119
rect 11431 25148 11719 25191
rect 5950 25043 5965 25045
rect 5865 25029 5965 25043
rect 5865 24986 5965 24987
rect 5486 24965 5965 24986
rect 6254 24965 6320 25061
rect 5486 24917 6320 24965
rect 5486 24888 5965 24917
rect 5486 24886 5591 24888
rect 5865 24887 5965 24888
rect 5319 24701 5329 24780
rect 5422 24701 5432 24780
rect 5330 23527 5423 24701
rect 6248 24652 6468 24672
rect 6248 24544 6292 24652
rect 6424 24544 6468 24652
rect 6248 24502 6468 24544
rect 5852 24472 6829 24502
rect 5852 24366 5884 24472
rect 6088 24366 6120 24472
rect 6324 24366 6356 24472
rect 6560 24366 6592 24472
rect 6795 24366 6829 24472
rect 5845 24354 5891 24366
rect 5845 24178 5851 24354
rect 5885 24178 5891 24354
rect 5845 24166 5891 24178
rect 5963 24354 6009 24366
rect 5963 24178 5969 24354
rect 6003 24178 6009 24354
rect 5963 24166 6009 24178
rect 6081 24354 6127 24366
rect 6081 24178 6087 24354
rect 6121 24178 6127 24354
rect 6081 24166 6127 24178
rect 6199 24354 6245 24366
rect 6199 24178 6205 24354
rect 6239 24178 6245 24354
rect 6199 24166 6245 24178
rect 6317 24354 6363 24366
rect 6317 24178 6323 24354
rect 6357 24178 6363 24354
rect 6317 24166 6363 24178
rect 6435 24354 6481 24366
rect 6435 24178 6441 24354
rect 6475 24178 6481 24354
rect 6435 24166 6481 24178
rect 6553 24354 6599 24366
rect 6553 24178 6559 24354
rect 6593 24178 6599 24354
rect 6553 24166 6599 24178
rect 6671 24354 6717 24366
rect 6671 24178 6677 24354
rect 6711 24178 6717 24354
rect 6671 24166 6717 24178
rect 6789 24354 6835 24366
rect 6789 24178 6795 24354
rect 6829 24178 6835 24354
rect 6789 24166 6835 24178
rect 6907 24354 6953 24366
rect 6907 24178 6913 24354
rect 6947 24178 6953 24354
rect 6907 24166 6953 24178
rect 7445 24300 7479 25084
rect 8158 25022 8192 25084
rect 7747 24984 8489 25022
rect 7747 24860 7781 24984
rect 7983 24860 8017 24984
rect 8219 24860 8253 24984
rect 8455 24860 8489 24984
rect 8745 24877 8755 24943
rect 8818 24877 8828 24943
rect 7741 24848 7787 24860
rect 7741 24472 7747 24848
rect 7781 24472 7787 24848
rect 7741 24460 7787 24472
rect 7859 24848 7905 24860
rect 7859 24472 7865 24848
rect 7899 24472 7905 24848
rect 7859 24460 7905 24472
rect 7977 24848 8023 24860
rect 7977 24472 7983 24848
rect 8017 24472 8023 24848
rect 7977 24460 8023 24472
rect 8095 24848 8141 24860
rect 8095 24472 8101 24848
rect 8135 24472 8141 24848
rect 8095 24460 8141 24472
rect 8213 24848 8259 24860
rect 8213 24472 8219 24848
rect 8253 24472 8259 24848
rect 8213 24460 8259 24472
rect 8331 24848 8377 24860
rect 8331 24472 8337 24848
rect 8371 24472 8377 24848
rect 8331 24460 8377 24472
rect 8449 24848 8495 24860
rect 8449 24472 8455 24848
rect 8489 24472 8495 24848
rect 8449 24460 8495 24472
rect 8861 24301 8895 25084
rect 8588 24300 8895 24301
rect 7445 24295 7761 24300
rect 8475 24295 8895 24300
rect 7445 24284 7828 24295
rect 7445 24257 7777 24284
rect 5968 24072 6004 24166
rect 6204 24072 6240 24166
rect 6440 24073 6476 24166
rect 6602 24118 6668 24125
rect 6602 24084 6618 24118
rect 6652 24084 6668 24118
rect 6602 24073 6668 24084
rect 6440 24072 6668 24073
rect 5968 24043 6668 24072
rect 5968 24042 6550 24043
rect 6088 23929 6122 24042
rect 6484 24001 6550 24042
rect 6484 23967 6500 24001
rect 6534 23967 6550 24001
rect 6484 23960 6550 23967
rect 6912 23933 6947 24166
rect 7445 24128 7479 24257
rect 7761 24250 7777 24257
rect 7811 24250 7828 24284
rect 7761 24244 7828 24250
rect 8408 24284 8895 24295
rect 8408 24250 8425 24284
rect 8459 24257 8895 24284
rect 8459 24250 8475 24257
rect 8588 24256 8895 24257
rect 8408 24244 8475 24250
rect 7586 24217 7642 24229
rect 7586 24183 7592 24217
rect 7626 24216 7642 24217
rect 8699 24216 8755 24228
rect 7626 24200 8093 24216
rect 7626 24183 8043 24200
rect 7586 24167 8043 24183
rect 8027 24166 8043 24167
rect 8077 24166 8093 24200
rect 8027 24159 8093 24166
rect 8145 24201 8715 24216
rect 8145 24167 8161 24201
rect 8195 24182 8715 24201
rect 8749 24182 8755 24216
rect 8195 24167 8755 24182
rect 8145 24157 8212 24167
rect 8699 24166 8755 24167
rect 8861 24128 8895 24256
rect 9343 24300 9377 25084
rect 10056 25022 10090 25084
rect 9645 24984 10387 25022
rect 9645 24860 9679 24984
rect 9881 24860 9915 24984
rect 10117 24860 10151 24984
rect 10353 24860 10387 24984
rect 9639 24848 9685 24860
rect 9639 24472 9645 24848
rect 9679 24472 9685 24848
rect 9639 24460 9685 24472
rect 9757 24848 9803 24860
rect 9757 24472 9763 24848
rect 9797 24472 9803 24848
rect 9757 24460 9803 24472
rect 9875 24848 9921 24860
rect 9875 24472 9881 24848
rect 9915 24472 9921 24848
rect 9875 24460 9921 24472
rect 9993 24848 10039 24860
rect 9993 24472 9999 24848
rect 10033 24472 10039 24848
rect 9993 24460 10039 24472
rect 10111 24848 10157 24860
rect 10111 24472 10117 24848
rect 10151 24472 10157 24848
rect 10111 24460 10157 24472
rect 10229 24848 10275 24860
rect 10229 24472 10235 24848
rect 10269 24472 10275 24848
rect 10229 24460 10275 24472
rect 10347 24848 10393 24860
rect 10347 24472 10353 24848
rect 10387 24472 10393 24848
rect 10347 24460 10393 24472
rect 10759 24301 10793 25084
rect 11431 25042 11567 25148
rect 11679 25146 11719 25148
rect 11685 25135 11719 25146
rect 11431 25040 11573 25042
rect 11685 25040 11720 25135
rect 11431 25031 11720 25040
rect 11431 25030 11719 25031
rect 11431 25029 11687 25030
rect 10371 24300 10440 24301
rect 10486 24300 10793 24301
rect 9343 24295 9659 24300
rect 10371 24296 10793 24300
rect 9343 24284 9726 24295
rect 9343 24257 9675 24284
rect 9343 24128 9377 24257
rect 9659 24250 9675 24257
rect 9709 24250 9726 24284
rect 9659 24244 9726 24250
rect 10304 24285 10793 24296
rect 10304 24251 10321 24285
rect 10355 24257 10793 24285
rect 10355 24251 10371 24257
rect 10486 24256 10793 24257
rect 10304 24245 10371 24251
rect 9484 24217 9540 24229
rect 9484 24183 9490 24217
rect 9524 24216 9540 24217
rect 10597 24216 10653 24228
rect 9524 24200 9991 24216
rect 9524 24183 9941 24200
rect 9484 24167 9941 24183
rect 9925 24166 9941 24167
rect 9975 24166 9991 24200
rect 9925 24159 9991 24166
rect 10043 24201 10613 24216
rect 10043 24167 10059 24201
rect 10093 24182 10613 24201
rect 10647 24182 10653 24216
rect 10093 24167 10653 24182
rect 10043 24157 10110 24167
rect 10597 24166 10653 24167
rect 10759 24128 10793 24256
rect 10874 24906 10941 24930
rect 10874 24872 10891 24906
rect 10925 24872 10941 24906
rect 6558 23929 6947 23933
rect 6082 23917 6128 23929
rect 6082 23541 6088 23917
rect 6122 23541 6128 23917
rect 6082 23529 6128 23541
rect 6200 23917 6246 23929
rect 6200 23541 6206 23917
rect 6240 23541 6246 23917
rect 6200 23529 6246 23541
rect 6318 23917 6364 23929
rect 6318 23541 6324 23917
rect 6358 23565 6364 23917
rect 6435 23917 6481 23929
rect 6435 23741 6441 23917
rect 6475 23741 6481 23917
rect 6435 23729 6481 23741
rect 6553 23917 6947 23929
rect 7439 24116 7485 24128
rect 7439 23940 7445 24116
rect 7479 23940 7485 24116
rect 7439 23928 7485 23940
rect 7557 24116 7603 24128
rect 7557 23940 7563 24116
rect 7597 23940 7603 24116
rect 7557 23928 7603 23940
rect 7859 24116 7905 24128
rect 6553 23741 6559 23917
rect 6593 23904 6947 23917
rect 6593 23741 6599 23904
rect 6869 23901 6947 23904
rect 6869 23849 6879 23901
rect 6942 23849 6952 23901
rect 6874 23843 6947 23849
rect 6553 23729 6599 23741
rect 6441 23613 6476 23729
rect 7562 23634 7596 23928
rect 7859 23740 7865 24116
rect 7899 23740 7905 24116
rect 7859 23728 7905 23740
rect 7977 24116 8023 24128
rect 7977 23740 7983 24116
rect 8017 23740 8023 24116
rect 7977 23728 8023 23740
rect 8095 24116 8141 24128
rect 8095 23740 8101 24116
rect 8135 23740 8141 24116
rect 8095 23728 8141 23740
rect 8213 24116 8259 24128
rect 8213 23740 8219 24116
rect 8253 23740 8259 24116
rect 8213 23728 8259 23740
rect 8331 24116 8377 24128
rect 8331 23740 8337 24116
rect 8371 23740 8377 24116
rect 8737 24116 8783 24128
rect 8737 23940 8743 24116
rect 8777 23940 8783 24116
rect 8737 23928 8783 23940
rect 8855 24116 8901 24128
rect 8855 23940 8861 24116
rect 8895 23940 8901 24116
rect 8855 23928 8901 23940
rect 9337 24116 9383 24128
rect 9337 23940 9343 24116
rect 9377 23940 9383 24116
rect 9337 23928 9383 23940
rect 9455 24116 9501 24128
rect 9455 23940 9461 24116
rect 9495 23940 9501 24116
rect 9455 23928 9501 23940
rect 9757 24116 9803 24128
rect 8331 23728 8377 23740
rect 8219 23634 8253 23728
rect 8743 23634 8776 23928
rect 6572 23613 6680 23623
rect 6441 23565 6572 23613
rect 6358 23541 6572 23565
rect 6318 23529 6572 23541
rect 5330 23525 5915 23527
rect 6324 23525 6572 23529
rect 5330 23497 5960 23525
rect 5330 23491 6197 23497
rect 5330 23457 6147 23491
rect 6181 23457 6197 23491
rect 5330 23441 6197 23457
rect 6249 23491 6315 23497
rect 6249 23457 6265 23491
rect 6299 23457 6315 23491
rect 6498 23481 6572 23525
rect 7562 23602 8776 23634
rect 9460 23634 9494 23928
rect 9757 23740 9763 24116
rect 9797 23740 9803 24116
rect 9757 23728 9803 23740
rect 9875 24116 9921 24128
rect 9875 23740 9881 24116
rect 9915 23740 9921 24116
rect 9875 23728 9921 23740
rect 9993 24116 10039 24128
rect 9993 23740 9999 24116
rect 10033 23740 10039 24116
rect 9993 23728 10039 23740
rect 10111 24116 10157 24128
rect 10111 23740 10117 24116
rect 10151 23740 10157 24116
rect 10111 23728 10157 23740
rect 10229 24116 10275 24128
rect 10229 23740 10235 24116
rect 10269 23740 10275 24116
rect 10635 24116 10681 24128
rect 10635 23940 10641 24116
rect 10675 23940 10681 24116
rect 10635 23928 10681 23940
rect 10753 24116 10799 24128
rect 10753 23940 10759 24116
rect 10793 23940 10799 24116
rect 10753 23928 10799 23940
rect 10229 23728 10275 23740
rect 10117 23634 10151 23728
rect 10641 23634 10674 23928
rect 9460 23602 10674 23634
rect 8055 23517 8187 23602
rect 9953 23517 10085 23602
rect 6572 23471 6680 23481
rect 5330 23425 5960 23441
rect 5330 23421 5915 23425
rect 5330 23420 5431 23421
rect 5860 23372 5960 23383
rect 5824 23266 5834 23372
rect 5946 23361 5960 23372
rect 6249 23361 6315 23457
rect 8045 23409 8055 23517
rect 8187 23409 8197 23517
rect 9943 23409 9953 23517
rect 10085 23409 10095 23517
rect 10874 23489 10941 24872
rect 11843 24777 11936 26671
rect 11999 26612 12465 26634
rect 12753 26612 12819 26708
rect 14584 26718 14590 26894
rect 14624 26718 14630 26894
rect 14584 26706 14630 26718
rect 14702 26894 14748 26906
rect 14702 26718 14708 26894
rect 14742 26718 14748 26894
rect 14702 26706 14748 26718
rect 14820 26894 14866 26906
rect 14820 26718 14826 26894
rect 14860 26718 14866 26894
rect 14820 26706 14866 26718
rect 14938 26894 14984 26906
rect 14938 26718 14944 26894
rect 14978 26839 14984 26894
rect 15103 26894 15149 26906
rect 15103 26839 15109 26894
rect 14978 26751 15109 26839
rect 14978 26718 14984 26751
rect 14938 26706 14984 26718
rect 15103 26718 15109 26751
rect 15143 26718 15149 26894
rect 15103 26706 15149 26718
rect 15221 26894 15267 26906
rect 15221 26718 15227 26894
rect 15261 26718 15267 26894
rect 15221 26706 15267 26718
rect 15339 26894 15385 26906
rect 15339 26718 15345 26894
rect 15379 26718 15385 26894
rect 15339 26706 15385 26718
rect 15457 26894 15503 26906
rect 15457 26718 15463 26894
rect 15497 26718 15503 26894
rect 15457 26706 15503 26718
rect 14590 26667 14624 26706
rect 14826 26667 14860 26706
rect 14590 26632 14860 26667
rect 15227 26668 15260 26706
rect 15463 26668 15496 26706
rect 15227 26632 15496 26668
rect 11999 26564 12819 26612
rect 14624 26631 14860 26632
rect 11999 26533 12465 26564
rect 14624 26557 14756 26631
rect 11999 26277 12104 26533
rect 14614 26449 14624 26557
rect 14756 26449 14766 26557
rect 11999 26171 12062 26277
rect 12174 26171 12184 26277
rect 12766 26253 12986 26273
rect 11999 26160 12148 26171
rect 11999 24983 12104 26160
rect 12766 26145 12810 26253
rect 12942 26145 12986 26253
rect 12766 26103 12986 26145
rect 15564 26118 15626 27689
rect 15816 27681 15862 27693
rect 15816 27305 15822 27681
rect 15856 27305 15862 27681
rect 15816 27293 15862 27305
rect 15934 27681 15980 27693
rect 15934 27305 15940 27681
rect 15974 27305 15980 27681
rect 15934 27293 15980 27305
rect 16052 27681 16098 27693
rect 16052 27305 16058 27681
rect 16092 27305 16098 27681
rect 16052 27293 16098 27305
rect 16170 27681 16216 27693
rect 16170 27305 16176 27681
rect 16210 27305 16216 27681
rect 16170 27293 16216 27305
rect 16288 27681 16334 27693
rect 16288 27305 16294 27681
rect 16328 27305 16334 27681
rect 16288 27293 16334 27305
rect 16406 27681 16452 27693
rect 16406 27305 16412 27681
rect 16446 27305 16452 27681
rect 16406 27293 16452 27305
rect 16524 27681 16570 27693
rect 16524 27305 16530 27681
rect 16564 27305 16570 27681
rect 18890 27718 19867 27748
rect 18890 27612 18922 27718
rect 19126 27612 19158 27718
rect 19362 27612 19394 27718
rect 19598 27612 19630 27718
rect 19833 27612 19867 27718
rect 18883 27600 18929 27612
rect 18883 27424 18889 27600
rect 18923 27424 18929 27600
rect 18883 27412 18929 27424
rect 19001 27600 19047 27612
rect 19001 27424 19007 27600
rect 19041 27424 19047 27600
rect 19001 27412 19047 27424
rect 19119 27600 19165 27612
rect 19119 27424 19125 27600
rect 19159 27424 19165 27600
rect 19119 27412 19165 27424
rect 19237 27600 19283 27612
rect 19237 27424 19243 27600
rect 19277 27424 19283 27600
rect 19237 27412 19283 27424
rect 19355 27600 19401 27612
rect 19355 27424 19361 27600
rect 19395 27424 19401 27600
rect 19355 27412 19401 27424
rect 19473 27600 19519 27612
rect 19473 27424 19479 27600
rect 19513 27424 19519 27600
rect 19473 27412 19519 27424
rect 19591 27600 19637 27612
rect 19591 27424 19597 27600
rect 19631 27424 19637 27600
rect 19591 27412 19637 27424
rect 19709 27600 19755 27612
rect 19709 27424 19715 27600
rect 19749 27424 19755 27600
rect 19709 27412 19755 27424
rect 19827 27600 19873 27612
rect 19827 27424 19833 27600
rect 19867 27424 19873 27600
rect 19827 27412 19873 27424
rect 19945 27600 19991 27612
rect 19945 27424 19951 27600
rect 19985 27424 19991 27600
rect 19945 27412 19991 27424
rect 16524 27293 16570 27305
rect 19006 27318 19042 27412
rect 19242 27318 19278 27412
rect 19478 27319 19514 27412
rect 19640 27364 19706 27371
rect 19640 27330 19656 27364
rect 19690 27330 19706 27364
rect 19640 27319 19706 27330
rect 19478 27318 19706 27319
rect 15822 27251 15856 27293
rect 16058 27251 16092 27293
rect 15822 27223 16092 27251
rect 16176 27252 16210 27293
rect 16412 27252 16446 27293
rect 16176 27223 16446 27252
rect 15822 27175 15856 27223
rect 15822 27145 15885 27175
rect 15850 27053 15885 27145
rect 16357 27115 16457 27136
rect 16357 27061 16371 27115
rect 16436 27061 16457 27115
rect 16357 27056 16457 27061
rect 16530 27110 16564 27293
rect 19006 27289 19706 27318
rect 19006 27288 19588 27289
rect 19126 27175 19160 27288
rect 19522 27247 19588 27288
rect 19522 27213 19538 27247
rect 19572 27213 19588 27247
rect 19522 27206 19588 27213
rect 19950 27207 19985 27412
rect 20157 27207 20224 27797
rect 21916 27774 21957 27806
rect 22203 27802 22213 27868
rect 22269 27802 22279 27868
rect 22949 27844 22959 27952
rect 23091 27889 23101 27952
rect 25844 27902 26064 27922
rect 23091 27878 23103 27889
rect 23091 27844 23104 27878
rect 22959 27806 23104 27844
rect 23063 27778 23104 27806
rect 21332 27746 21602 27774
rect 21073 27680 21083 27746
rect 21149 27680 21159 27746
rect 21332 27684 21366 27746
rect 21568 27684 21602 27746
rect 21686 27746 21957 27774
rect 22474 27750 22744 27778
rect 21686 27684 21720 27746
rect 21922 27684 21957 27746
rect 22098 27734 22269 27750
rect 22098 27700 22229 27734
rect 22263 27700 22269 27734
rect 22098 27684 22269 27700
rect 22474 27688 22508 27750
rect 22710 27688 22744 27750
rect 22828 27750 23104 27778
rect 25844 27794 25888 27902
rect 26020 27794 26064 27902
rect 27641 27860 27697 27868
rect 25844 27752 26064 27794
rect 26715 27852 27697 27860
rect 26715 27818 27657 27852
rect 27691 27818 27697 27852
rect 28360 27848 28370 27956
rect 28502 27893 28512 27956
rect 28502 27882 28514 27893
rect 28502 27848 28515 27882
rect 28771 27872 28827 27874
rect 26715 27802 27697 27818
rect 28370 27810 28515 27848
rect 26715 27801 27694 27802
rect 22828 27688 22862 27750
rect 23064 27688 23104 27750
rect 21208 27672 21254 27684
rect 21208 27296 21214 27672
rect 21248 27296 21254 27672
rect 21208 27284 21254 27296
rect 21326 27672 21372 27684
rect 21326 27296 21332 27672
rect 21366 27296 21372 27672
rect 21326 27284 21372 27296
rect 21444 27672 21490 27684
rect 21444 27296 21450 27672
rect 21484 27296 21490 27672
rect 21444 27284 21490 27296
rect 21562 27672 21608 27684
rect 21562 27296 21568 27672
rect 21602 27296 21608 27672
rect 21562 27284 21608 27296
rect 21680 27672 21726 27684
rect 21680 27296 21686 27672
rect 21720 27296 21726 27672
rect 21680 27284 21726 27296
rect 21798 27672 21844 27684
rect 21798 27296 21804 27672
rect 21838 27296 21844 27672
rect 21798 27284 21844 27296
rect 21916 27672 21962 27684
rect 21916 27296 21922 27672
rect 21956 27296 21962 27672
rect 21916 27284 21962 27296
rect 19950 27179 20224 27207
rect 19596 27175 20224 27179
rect 19120 27163 19166 27175
rect 17539 27124 17638 27128
rect 16530 27056 16639 27110
rect 15850 27017 16077 27053
rect 15850 26910 15885 27017
rect 16011 26983 16077 27017
rect 16011 26949 16027 26983
rect 16061 26949 16077 26983
rect 16358 27041 16455 27056
rect 16358 26974 16415 27041
rect 16011 26943 16077 26949
rect 16252 26938 16521 26974
rect 16252 26910 16285 26938
rect 16488 26910 16521 26938
rect 16605 26910 16639 27056
rect 17456 27049 17466 27124
rect 17534 27049 17638 27124
rect 17483 27048 17638 27049
rect 15726 26898 15772 26910
rect 15726 26722 15732 26898
rect 15766 26722 15772 26898
rect 15726 26710 15772 26722
rect 15844 26898 15890 26910
rect 15844 26722 15850 26898
rect 15884 26722 15890 26898
rect 15844 26710 15890 26722
rect 15962 26898 16008 26910
rect 15962 26722 15968 26898
rect 16002 26722 16008 26898
rect 15962 26710 16008 26722
rect 16080 26898 16126 26910
rect 16080 26722 16086 26898
rect 16120 26843 16126 26898
rect 16245 26898 16291 26910
rect 16245 26843 16251 26898
rect 16120 26755 16251 26843
rect 16120 26722 16126 26755
rect 16080 26710 16126 26722
rect 16245 26722 16251 26755
rect 16285 26722 16291 26898
rect 16245 26710 16291 26722
rect 16363 26898 16409 26910
rect 16363 26722 16369 26898
rect 16403 26722 16409 26898
rect 16363 26710 16409 26722
rect 16481 26898 16527 26910
rect 16481 26722 16487 26898
rect 16521 26722 16527 26898
rect 16481 26710 16527 26722
rect 16599 26898 16645 26910
rect 16599 26722 16605 26898
rect 16639 26722 16645 26898
rect 16599 26710 16645 26722
rect 15732 26671 15766 26710
rect 15968 26671 16002 26710
rect 15732 26635 16002 26671
rect 16369 26672 16402 26710
rect 16605 26672 16638 26710
rect 16369 26636 16638 26672
rect 15732 26634 15898 26635
rect 15766 26555 15898 26634
rect 15756 26447 15766 26555
rect 15898 26447 15908 26555
rect 12370 26073 13347 26103
rect 15564 26101 15627 26118
rect 15489 26097 15627 26101
rect 12370 25967 12402 26073
rect 12606 25967 12638 26073
rect 12842 25967 12874 26073
rect 13078 25967 13110 26073
rect 13313 25967 13347 26073
rect 13657 26063 15627 26097
rect 13655 26034 15627 26063
rect 13655 26018 13701 26034
rect 15489 26032 15627 26034
rect 12363 25955 12409 25967
rect 12363 25779 12369 25955
rect 12403 25779 12409 25955
rect 12363 25767 12409 25779
rect 12481 25955 12527 25967
rect 12481 25779 12487 25955
rect 12521 25779 12527 25955
rect 12481 25767 12527 25779
rect 12599 25955 12645 25967
rect 12599 25779 12605 25955
rect 12639 25779 12645 25955
rect 12599 25767 12645 25779
rect 12717 25955 12763 25967
rect 12717 25779 12723 25955
rect 12757 25779 12763 25955
rect 12717 25767 12763 25779
rect 12835 25955 12881 25967
rect 12835 25779 12841 25955
rect 12875 25779 12881 25955
rect 12835 25767 12881 25779
rect 12953 25955 12999 25967
rect 12953 25779 12959 25955
rect 12993 25779 12999 25955
rect 12953 25767 12999 25779
rect 13071 25955 13117 25967
rect 13071 25779 13077 25955
rect 13111 25779 13117 25955
rect 13071 25767 13117 25779
rect 13189 25955 13235 25967
rect 13189 25779 13195 25955
rect 13229 25779 13235 25955
rect 13189 25767 13235 25779
rect 13307 25955 13353 25967
rect 13307 25779 13313 25955
rect 13347 25779 13353 25955
rect 13307 25767 13353 25779
rect 13425 25955 13471 25967
rect 13425 25779 13431 25955
rect 13465 25779 13471 25955
rect 13425 25767 13471 25779
rect 12486 25673 12522 25767
rect 12722 25673 12758 25767
rect 12958 25674 12994 25767
rect 13120 25719 13186 25726
rect 13120 25685 13136 25719
rect 13170 25685 13186 25719
rect 13120 25674 13186 25685
rect 12958 25673 13186 25674
rect 12486 25644 13186 25673
rect 12486 25643 13068 25644
rect 12606 25530 12640 25643
rect 13002 25602 13068 25643
rect 13002 25568 13018 25602
rect 13052 25568 13068 25602
rect 13002 25561 13068 25568
rect 13430 25549 13465 25767
rect 13654 25566 13701 26018
rect 14613 25802 14623 25910
rect 14755 25802 14765 25910
rect 16511 25802 16521 25910
rect 16653 25802 16663 25910
rect 14623 25762 14755 25802
rect 16521 25762 16653 25802
rect 14622 25696 14755 25762
rect 16520 25696 16653 25762
rect 13951 25653 15424 25696
rect 13654 25550 13700 25566
rect 13619 25549 13700 25550
rect 13430 25534 13700 25549
rect 13076 25530 13700 25534
rect 12600 25518 12646 25530
rect 12335 25040 12345 25158
rect 12463 25126 12473 25158
rect 12600 25142 12606 25518
rect 12640 25142 12646 25518
rect 12600 25130 12646 25142
rect 12718 25518 12764 25530
rect 12718 25142 12724 25518
rect 12758 25142 12764 25518
rect 12718 25130 12764 25142
rect 12836 25518 12882 25530
rect 12836 25142 12842 25518
rect 12876 25166 12882 25518
rect 12953 25518 12999 25530
rect 12953 25342 12959 25518
rect 12993 25342 12999 25518
rect 12953 25330 12999 25342
rect 13071 25518 13700 25530
rect 13071 25342 13077 25518
rect 13111 25506 13700 25518
rect 13111 25505 13353 25506
rect 13111 25342 13117 25505
rect 13619 25504 13700 25506
rect 13951 25350 13985 25653
rect 14317 25550 14351 25653
rect 14553 25550 14587 25653
rect 14789 25550 14823 25653
rect 15025 25550 15059 25653
rect 14311 25538 14357 25550
rect 13071 25330 13117 25342
rect 13827 25338 13873 25350
rect 12959 25214 12994 25330
rect 13090 25214 13198 25224
rect 12959 25166 13090 25214
rect 12876 25142 13090 25166
rect 12836 25130 13090 25142
rect 12842 25126 13090 25130
rect 12463 25098 12478 25126
rect 12463 25092 12715 25098
rect 12463 25058 12665 25092
rect 12699 25058 12715 25092
rect 12463 25042 12715 25058
rect 12767 25092 12833 25098
rect 12767 25058 12783 25092
rect 12817 25058 12833 25092
rect 13016 25082 13090 25126
rect 13827 25162 13833 25338
rect 13867 25162 13873 25338
rect 13827 25150 13873 25162
rect 13945 25338 13991 25350
rect 13945 25162 13951 25338
rect 13985 25162 13991 25338
rect 13945 25150 13991 25162
rect 14063 25338 14109 25350
rect 14063 25162 14069 25338
rect 14103 25162 14109 25338
rect 14063 25150 14109 25162
rect 14181 25338 14227 25350
rect 14311 25338 14317 25538
rect 14181 25162 14187 25338
rect 14221 25162 14317 25338
rect 14351 25162 14357 25538
rect 14181 25150 14227 25162
rect 14311 25150 14357 25162
rect 14429 25538 14475 25550
rect 14429 25162 14435 25538
rect 14469 25162 14475 25538
rect 14429 25150 14475 25162
rect 14547 25538 14593 25550
rect 14547 25162 14553 25538
rect 14587 25162 14593 25538
rect 14547 25150 14593 25162
rect 14665 25538 14711 25550
rect 14665 25162 14671 25538
rect 14705 25162 14711 25538
rect 14665 25150 14711 25162
rect 14783 25538 14829 25550
rect 14783 25162 14789 25538
rect 14823 25162 14829 25538
rect 14783 25150 14829 25162
rect 14901 25538 14947 25550
rect 14901 25162 14907 25538
rect 14941 25162 14947 25538
rect 14901 25150 14947 25162
rect 15019 25538 15065 25550
rect 15019 25162 15025 25538
rect 15059 25338 15065 25538
rect 15390 25350 15424 25653
rect 15849 25653 17322 25696
rect 15849 25350 15883 25653
rect 16215 25550 16249 25653
rect 16451 25550 16485 25653
rect 16687 25550 16721 25653
rect 16923 25550 16957 25653
rect 16209 25538 16255 25550
rect 15148 25338 15194 25350
rect 15059 25162 15154 25338
rect 15188 25162 15194 25338
rect 15019 25150 15065 25162
rect 15148 25150 15194 25162
rect 15266 25338 15312 25350
rect 15266 25162 15272 25338
rect 15306 25162 15312 25338
rect 15266 25150 15312 25162
rect 15384 25338 15430 25350
rect 15384 25162 15390 25338
rect 15424 25162 15430 25338
rect 15384 25150 15430 25162
rect 15502 25338 15548 25350
rect 15502 25162 15508 25338
rect 15542 25162 15548 25338
rect 15502 25150 15548 25162
rect 15725 25338 15771 25350
rect 15725 25162 15731 25338
rect 15765 25162 15771 25338
rect 15725 25150 15771 25162
rect 15843 25338 15889 25350
rect 15843 25162 15849 25338
rect 15883 25162 15889 25338
rect 15843 25150 15889 25162
rect 15961 25338 16007 25350
rect 15961 25162 15967 25338
rect 16001 25162 16007 25338
rect 15961 25150 16007 25162
rect 16079 25338 16125 25350
rect 16209 25338 16215 25538
rect 16079 25162 16085 25338
rect 16119 25162 16215 25338
rect 16249 25162 16255 25538
rect 16079 25150 16125 25162
rect 16209 25150 16255 25162
rect 16327 25538 16373 25550
rect 16327 25162 16333 25538
rect 16367 25162 16373 25538
rect 16327 25150 16373 25162
rect 16445 25538 16491 25550
rect 16445 25162 16451 25538
rect 16485 25162 16491 25538
rect 16445 25150 16491 25162
rect 16563 25538 16609 25550
rect 16563 25162 16569 25538
rect 16603 25162 16609 25538
rect 16563 25150 16609 25162
rect 16681 25538 16727 25550
rect 16681 25162 16687 25538
rect 16721 25162 16727 25538
rect 16681 25150 16727 25162
rect 16799 25538 16845 25550
rect 16799 25162 16805 25538
rect 16839 25162 16845 25538
rect 16799 25150 16845 25162
rect 16917 25538 16963 25550
rect 16917 25162 16923 25538
rect 16957 25338 16963 25538
rect 17288 25350 17322 25653
rect 17046 25338 17092 25350
rect 16957 25162 17052 25338
rect 17086 25162 17092 25338
rect 16917 25150 16963 25162
rect 17046 25150 17092 25162
rect 17164 25338 17210 25350
rect 17164 25162 17170 25338
rect 17204 25162 17210 25338
rect 17164 25150 17210 25162
rect 17282 25338 17328 25350
rect 17282 25162 17288 25338
rect 17322 25162 17328 25338
rect 17282 25150 17328 25162
rect 17400 25338 17446 25350
rect 17400 25162 17406 25338
rect 17440 25162 17446 25338
rect 17539 25302 17638 27048
rect 17948 26845 18237 26864
rect 17948 26688 17969 26845
rect 18202 26770 18237 26845
rect 19120 26787 19126 27163
rect 19160 26787 19166 27163
rect 19120 26775 19166 26787
rect 19238 27163 19284 27175
rect 19238 26787 19244 27163
rect 19278 26787 19284 27163
rect 19238 26775 19284 26787
rect 19356 27163 19402 27175
rect 19356 26787 19362 27163
rect 19396 26811 19402 27163
rect 19473 27163 19519 27175
rect 19473 26987 19479 27163
rect 19513 26987 19519 27163
rect 19473 26975 19519 26987
rect 19591 27163 20224 27175
rect 19591 26987 19597 27163
rect 19631 27150 20224 27163
rect 21214 27242 21248 27284
rect 21450 27242 21484 27284
rect 21214 27214 21484 27242
rect 21568 27243 21602 27284
rect 21804 27243 21838 27284
rect 21568 27214 21838 27243
rect 21214 27166 21248 27214
rect 19631 26987 19637 27150
rect 21214 27136 21277 27166
rect 19591 26975 19637 26987
rect 21242 27044 21277 27136
rect 21242 27008 21469 27044
rect 21739 27033 21749 27130
rect 21848 27033 21858 27130
rect 21922 27101 21956 27284
rect 21922 27047 22031 27101
rect 19479 26859 19514 26975
rect 21242 26901 21277 27008
rect 21403 26974 21469 27008
rect 21403 26940 21419 26974
rect 21453 26940 21469 26974
rect 21750 27032 21847 27033
rect 21750 26965 21807 27032
rect 21403 26934 21469 26940
rect 21644 26929 21913 26965
rect 21644 26901 21677 26929
rect 21880 26901 21913 26929
rect 21997 26901 22031 27047
rect 21118 26889 21164 26901
rect 19610 26859 19718 26869
rect 19479 26811 19610 26859
rect 19396 26787 19610 26811
rect 19356 26775 19610 26787
rect 19362 26771 19610 26775
rect 18202 26743 18998 26770
rect 18202 26737 19235 26743
rect 18202 26703 19185 26737
rect 19219 26703 19235 26737
rect 18202 26688 19235 26703
rect 17948 26687 19235 26688
rect 19287 26737 19353 26743
rect 19287 26703 19303 26737
rect 19337 26703 19353 26737
rect 19536 26727 19610 26771
rect 19610 26717 19718 26727
rect 17948 26671 18998 26687
rect 17948 26670 18935 26671
rect 17948 26666 18470 26670
rect 17948 26665 18237 26666
rect 17965 25302 18253 25305
rect 17539 25192 18253 25302
rect 17400 25150 17446 25162
rect 13090 25072 13198 25082
rect 13833 25116 13867 25150
rect 14435 25116 14469 25150
rect 14671 25116 14705 25150
rect 13833 25081 13992 25116
rect 14435 25081 14705 25116
rect 15272 25116 15306 25150
rect 15508 25116 15542 25150
rect 15272 25081 15542 25116
rect 15731 25116 15765 25150
rect 16333 25116 16367 25150
rect 16569 25116 16603 25150
rect 15731 25081 15890 25116
rect 16333 25081 16603 25116
rect 17170 25116 17204 25150
rect 17406 25116 17440 25150
rect 17170 25081 17440 25116
rect 17965 25143 18253 25192
rect 12463 25040 12478 25042
rect 12378 25026 12478 25040
rect 12378 24983 12478 24984
rect 11999 24962 12478 24983
rect 12767 24962 12833 25058
rect 11999 24914 12833 24962
rect 11999 24885 12478 24914
rect 11999 24883 12104 24885
rect 12378 24884 12478 24885
rect 11832 24698 11842 24777
rect 11935 24698 11945 24777
rect 11843 23524 11936 24698
rect 12761 24649 12981 24669
rect 12761 24541 12805 24649
rect 12937 24541 12981 24649
rect 12761 24499 12981 24541
rect 12365 24469 13342 24499
rect 12365 24363 12397 24469
rect 12601 24363 12633 24469
rect 12837 24363 12869 24469
rect 13073 24363 13105 24469
rect 13308 24363 13342 24469
rect 12358 24351 12404 24363
rect 12358 24175 12364 24351
rect 12398 24175 12404 24351
rect 12358 24163 12404 24175
rect 12476 24351 12522 24363
rect 12476 24175 12482 24351
rect 12516 24175 12522 24351
rect 12476 24163 12522 24175
rect 12594 24351 12640 24363
rect 12594 24175 12600 24351
rect 12634 24175 12640 24351
rect 12594 24163 12640 24175
rect 12712 24351 12758 24363
rect 12712 24175 12718 24351
rect 12752 24175 12758 24351
rect 12712 24163 12758 24175
rect 12830 24351 12876 24363
rect 12830 24175 12836 24351
rect 12870 24175 12876 24351
rect 12830 24163 12876 24175
rect 12948 24351 12994 24363
rect 12948 24175 12954 24351
rect 12988 24175 12994 24351
rect 12948 24163 12994 24175
rect 13066 24351 13112 24363
rect 13066 24175 13072 24351
rect 13106 24175 13112 24351
rect 13066 24163 13112 24175
rect 13184 24351 13230 24363
rect 13184 24175 13190 24351
rect 13224 24175 13230 24351
rect 13184 24163 13230 24175
rect 13302 24351 13348 24363
rect 13302 24175 13308 24351
rect 13342 24175 13348 24351
rect 13302 24163 13348 24175
rect 13420 24351 13466 24363
rect 13420 24175 13426 24351
rect 13460 24175 13466 24351
rect 13420 24163 13466 24175
rect 13958 24297 13992 25081
rect 14671 25019 14705 25081
rect 14260 24981 15002 25019
rect 14260 24857 14294 24981
rect 14496 24857 14530 24981
rect 14732 24857 14766 24981
rect 14968 24857 15002 24981
rect 15258 24874 15268 24940
rect 15331 24874 15341 24940
rect 14254 24845 14300 24857
rect 14254 24469 14260 24845
rect 14294 24469 14300 24845
rect 14254 24457 14300 24469
rect 14372 24845 14418 24857
rect 14372 24469 14378 24845
rect 14412 24469 14418 24845
rect 14372 24457 14418 24469
rect 14490 24845 14536 24857
rect 14490 24469 14496 24845
rect 14530 24469 14536 24845
rect 14490 24457 14536 24469
rect 14608 24845 14654 24857
rect 14608 24469 14614 24845
rect 14648 24469 14654 24845
rect 14608 24457 14654 24469
rect 14726 24845 14772 24857
rect 14726 24469 14732 24845
rect 14766 24469 14772 24845
rect 14726 24457 14772 24469
rect 14844 24845 14890 24857
rect 14844 24469 14850 24845
rect 14884 24469 14890 24845
rect 14844 24457 14890 24469
rect 14962 24845 15008 24857
rect 14962 24469 14968 24845
rect 15002 24469 15008 24845
rect 14962 24457 15008 24469
rect 15374 24298 15408 25081
rect 15101 24297 15408 24298
rect 13958 24292 14274 24297
rect 14988 24292 15408 24297
rect 13958 24281 14341 24292
rect 13958 24254 14290 24281
rect 12481 24069 12517 24163
rect 12717 24069 12753 24163
rect 12953 24070 12989 24163
rect 13115 24115 13181 24122
rect 13115 24081 13131 24115
rect 13165 24081 13181 24115
rect 13115 24070 13181 24081
rect 12953 24069 13181 24070
rect 12481 24040 13181 24069
rect 12481 24039 13063 24040
rect 12601 23926 12635 24039
rect 12997 23998 13063 24039
rect 12997 23964 13013 23998
rect 13047 23964 13063 23998
rect 12997 23957 13063 23964
rect 13425 23930 13460 24163
rect 13958 24125 13992 24254
rect 14274 24247 14290 24254
rect 14324 24247 14341 24281
rect 14274 24241 14341 24247
rect 14921 24281 15408 24292
rect 14921 24247 14938 24281
rect 14972 24254 15408 24281
rect 14972 24247 14988 24254
rect 15101 24253 15408 24254
rect 14921 24241 14988 24247
rect 14099 24214 14155 24226
rect 14099 24180 14105 24214
rect 14139 24213 14155 24214
rect 15212 24213 15268 24225
rect 14139 24197 14606 24213
rect 14139 24180 14556 24197
rect 14099 24164 14556 24180
rect 14540 24163 14556 24164
rect 14590 24163 14606 24197
rect 14540 24156 14606 24163
rect 14658 24198 15228 24213
rect 14658 24164 14674 24198
rect 14708 24179 15228 24198
rect 15262 24179 15268 24213
rect 14708 24164 15268 24179
rect 14658 24154 14725 24164
rect 15212 24163 15268 24164
rect 15374 24125 15408 24253
rect 15856 24297 15890 25081
rect 16569 25019 16603 25081
rect 16158 24981 16900 25019
rect 16158 24857 16192 24981
rect 16394 24857 16428 24981
rect 16630 24857 16664 24981
rect 16866 24857 16900 24981
rect 16152 24845 16198 24857
rect 16152 24469 16158 24845
rect 16192 24469 16198 24845
rect 16152 24457 16198 24469
rect 16270 24845 16316 24857
rect 16270 24469 16276 24845
rect 16310 24469 16316 24845
rect 16270 24457 16316 24469
rect 16388 24845 16434 24857
rect 16388 24469 16394 24845
rect 16428 24469 16434 24845
rect 16388 24457 16434 24469
rect 16506 24845 16552 24857
rect 16506 24469 16512 24845
rect 16546 24469 16552 24845
rect 16506 24457 16552 24469
rect 16624 24845 16670 24857
rect 16624 24469 16630 24845
rect 16664 24469 16670 24845
rect 16624 24457 16670 24469
rect 16742 24845 16788 24857
rect 16742 24469 16748 24845
rect 16782 24469 16788 24845
rect 16742 24457 16788 24469
rect 16860 24845 16906 24857
rect 16860 24469 16866 24845
rect 16900 24469 16906 24845
rect 16860 24457 16906 24469
rect 17272 24298 17306 25081
rect 17965 25037 18101 25143
rect 18213 25141 18253 25143
rect 18219 25130 18253 25141
rect 17965 25035 18107 25037
rect 18219 25035 18254 25130
rect 17965 25026 18254 25035
rect 17965 25025 18253 25026
rect 17965 25024 18221 25025
rect 16884 24297 16953 24298
rect 16999 24297 17306 24298
rect 15856 24292 16172 24297
rect 16884 24293 17306 24297
rect 15856 24281 16239 24292
rect 15856 24254 16188 24281
rect 15856 24125 15890 24254
rect 16172 24247 16188 24254
rect 16222 24247 16239 24281
rect 16172 24241 16239 24247
rect 16817 24282 17306 24293
rect 16817 24248 16834 24282
rect 16868 24254 17306 24282
rect 16868 24248 16884 24254
rect 16999 24253 17306 24254
rect 16817 24242 16884 24248
rect 15997 24214 16053 24226
rect 15997 24180 16003 24214
rect 16037 24213 16053 24214
rect 17110 24213 17166 24225
rect 16037 24197 16504 24213
rect 16037 24180 16454 24197
rect 15997 24164 16454 24180
rect 16438 24163 16454 24164
rect 16488 24163 16504 24197
rect 16438 24156 16504 24163
rect 16556 24198 17126 24213
rect 16556 24164 16572 24198
rect 16606 24179 17126 24198
rect 17160 24179 17166 24213
rect 16606 24164 17166 24179
rect 16556 24154 16623 24164
rect 17110 24163 17166 24164
rect 17272 24125 17306 24253
rect 17387 24903 17454 24927
rect 17387 24869 17404 24903
rect 17438 24869 17454 24903
rect 13071 23926 13460 23930
rect 12595 23914 12641 23926
rect 12595 23538 12601 23914
rect 12635 23538 12641 23914
rect 12595 23526 12641 23538
rect 12713 23914 12759 23926
rect 12713 23538 12719 23914
rect 12753 23538 12759 23914
rect 12713 23526 12759 23538
rect 12831 23914 12877 23926
rect 12831 23538 12837 23914
rect 12871 23562 12877 23914
rect 12948 23914 12994 23926
rect 12948 23738 12954 23914
rect 12988 23738 12994 23914
rect 12948 23726 12994 23738
rect 13066 23914 13460 23926
rect 13952 24113 13998 24125
rect 13952 23937 13958 24113
rect 13992 23937 13998 24113
rect 13952 23925 13998 23937
rect 14070 24113 14116 24125
rect 14070 23937 14076 24113
rect 14110 23937 14116 24113
rect 14070 23925 14116 23937
rect 14372 24113 14418 24125
rect 13066 23738 13072 23914
rect 13106 23901 13460 23914
rect 13106 23738 13112 23901
rect 13382 23898 13460 23901
rect 13382 23846 13392 23898
rect 13455 23846 13465 23898
rect 13387 23840 13460 23846
rect 13066 23726 13112 23738
rect 12954 23610 12989 23726
rect 14075 23631 14109 23925
rect 14372 23737 14378 24113
rect 14412 23737 14418 24113
rect 14372 23725 14418 23737
rect 14490 24113 14536 24125
rect 14490 23737 14496 24113
rect 14530 23737 14536 24113
rect 14490 23725 14536 23737
rect 14608 24113 14654 24125
rect 14608 23737 14614 24113
rect 14648 23737 14654 24113
rect 14608 23725 14654 23737
rect 14726 24113 14772 24125
rect 14726 23737 14732 24113
rect 14766 23737 14772 24113
rect 14726 23725 14772 23737
rect 14844 24113 14890 24125
rect 14844 23737 14850 24113
rect 14884 23737 14890 24113
rect 15250 24113 15296 24125
rect 15250 23937 15256 24113
rect 15290 23937 15296 24113
rect 15250 23925 15296 23937
rect 15368 24113 15414 24125
rect 15368 23937 15374 24113
rect 15408 23937 15414 24113
rect 15368 23925 15414 23937
rect 15850 24113 15896 24125
rect 15850 23937 15856 24113
rect 15890 23937 15896 24113
rect 15850 23925 15896 23937
rect 15968 24113 16014 24125
rect 15968 23937 15974 24113
rect 16008 23937 16014 24113
rect 15968 23925 16014 23937
rect 16270 24113 16316 24125
rect 14844 23725 14890 23737
rect 14732 23631 14766 23725
rect 15256 23631 15289 23925
rect 13085 23610 13193 23620
rect 12954 23562 13085 23610
rect 12871 23538 13085 23562
rect 12831 23526 13085 23538
rect 11843 23522 12428 23524
rect 12837 23522 13085 23526
rect 11843 23494 12473 23522
rect 5946 23313 6315 23361
rect 5946 23283 5960 23313
rect 5946 23266 5956 23283
rect 6248 23210 6314 23313
rect 10874 23210 10940 23489
rect 11843 23488 12710 23494
rect 11843 23454 12660 23488
rect 12694 23454 12710 23488
rect 11843 23438 12710 23454
rect 12762 23488 12828 23494
rect 12762 23454 12778 23488
rect 12812 23454 12828 23488
rect 13011 23478 13085 23522
rect 14075 23599 15289 23631
rect 15973 23631 16007 23925
rect 16270 23737 16276 24113
rect 16310 23737 16316 24113
rect 16270 23725 16316 23737
rect 16388 24113 16434 24125
rect 16388 23737 16394 24113
rect 16428 23737 16434 24113
rect 16388 23725 16434 23737
rect 16506 24113 16552 24125
rect 16506 23737 16512 24113
rect 16546 23737 16552 24113
rect 16506 23725 16552 23737
rect 16624 24113 16670 24125
rect 16624 23737 16630 24113
rect 16664 23737 16670 24113
rect 16624 23725 16670 23737
rect 16742 24113 16788 24125
rect 16742 23737 16748 24113
rect 16782 23737 16788 24113
rect 17148 24113 17194 24125
rect 17148 23937 17154 24113
rect 17188 23937 17194 24113
rect 17148 23925 17194 23937
rect 17266 24113 17312 24125
rect 17266 23937 17272 24113
rect 17306 23937 17312 24113
rect 17266 23925 17312 23937
rect 16742 23725 16788 23737
rect 16630 23631 16664 23725
rect 17154 23631 17187 23925
rect 15973 23599 17187 23631
rect 14568 23514 14700 23599
rect 16466 23514 16598 23599
rect 13085 23468 13193 23478
rect 11843 23422 12473 23438
rect 11843 23418 12428 23422
rect 11843 23417 11944 23418
rect 12373 23369 12473 23380
rect 12337 23263 12347 23369
rect 12459 23358 12473 23369
rect 12762 23358 12828 23454
rect 14558 23406 14568 23514
rect 14700 23406 14710 23514
rect 16456 23406 16466 23514
rect 16598 23406 16608 23514
rect 17387 23486 17454 24869
rect 18377 24772 18470 26666
rect 18533 26607 18999 26629
rect 19287 26607 19353 26703
rect 21118 26713 21124 26889
rect 21158 26713 21164 26889
rect 21118 26701 21164 26713
rect 21236 26889 21282 26901
rect 21236 26713 21242 26889
rect 21276 26713 21282 26889
rect 21236 26701 21282 26713
rect 21354 26889 21400 26901
rect 21354 26713 21360 26889
rect 21394 26713 21400 26889
rect 21354 26701 21400 26713
rect 21472 26889 21518 26901
rect 21472 26713 21478 26889
rect 21512 26834 21518 26889
rect 21637 26889 21683 26901
rect 21637 26834 21643 26889
rect 21512 26746 21643 26834
rect 21512 26713 21518 26746
rect 21472 26701 21518 26713
rect 21637 26713 21643 26746
rect 21677 26713 21683 26889
rect 21637 26701 21683 26713
rect 21755 26889 21801 26901
rect 21755 26713 21761 26889
rect 21795 26713 21801 26889
rect 21755 26701 21801 26713
rect 21873 26889 21919 26901
rect 21873 26713 21879 26889
rect 21913 26713 21919 26889
rect 21873 26701 21919 26713
rect 21991 26889 22037 26901
rect 21991 26713 21997 26889
rect 22031 26713 22037 26889
rect 21991 26701 22037 26713
rect 21124 26662 21158 26701
rect 21360 26662 21394 26701
rect 21124 26627 21394 26662
rect 21761 26663 21794 26701
rect 21997 26663 22030 26701
rect 21761 26627 22030 26663
rect 18533 26559 19353 26607
rect 21158 26626 21394 26627
rect 18533 26528 18999 26559
rect 21158 26552 21290 26626
rect 18533 26272 18638 26528
rect 21148 26444 21158 26552
rect 21290 26444 21300 26552
rect 18533 26166 18596 26272
rect 18708 26166 18718 26272
rect 19300 26248 19520 26268
rect 18533 26155 18682 26166
rect 18533 24978 18638 26155
rect 19300 26140 19344 26248
rect 19476 26140 19520 26248
rect 19300 26098 19520 26140
rect 22098 26113 22160 27684
rect 22350 27676 22396 27688
rect 22350 27300 22356 27676
rect 22390 27300 22396 27676
rect 22350 27288 22396 27300
rect 22468 27676 22514 27688
rect 22468 27300 22474 27676
rect 22508 27300 22514 27676
rect 22468 27288 22514 27300
rect 22586 27676 22632 27688
rect 22586 27300 22592 27676
rect 22626 27300 22632 27676
rect 22586 27288 22632 27300
rect 22704 27676 22750 27688
rect 22704 27300 22710 27676
rect 22744 27300 22750 27676
rect 22704 27288 22750 27300
rect 22822 27676 22868 27688
rect 22822 27300 22828 27676
rect 22862 27300 22868 27676
rect 22822 27288 22868 27300
rect 22940 27676 22986 27688
rect 22940 27300 22946 27676
rect 22980 27300 22986 27676
rect 22940 27288 22986 27300
rect 23058 27676 23104 27688
rect 23058 27300 23064 27676
rect 23098 27300 23104 27676
rect 25448 27722 26425 27752
rect 25448 27616 25480 27722
rect 25684 27616 25716 27722
rect 25920 27616 25952 27722
rect 26156 27616 26188 27722
rect 26391 27616 26425 27722
rect 25441 27604 25487 27616
rect 25441 27428 25447 27604
rect 25481 27428 25487 27604
rect 25441 27416 25487 27428
rect 25559 27604 25605 27616
rect 25559 27428 25565 27604
rect 25599 27428 25605 27604
rect 25559 27416 25605 27428
rect 25677 27604 25723 27616
rect 25677 27428 25683 27604
rect 25717 27428 25723 27604
rect 25677 27416 25723 27428
rect 25795 27604 25841 27616
rect 25795 27428 25801 27604
rect 25835 27428 25841 27604
rect 25795 27416 25841 27428
rect 25913 27604 25959 27616
rect 25913 27428 25919 27604
rect 25953 27428 25959 27604
rect 25913 27416 25959 27428
rect 26031 27604 26077 27616
rect 26031 27428 26037 27604
rect 26071 27428 26077 27604
rect 26031 27416 26077 27428
rect 26149 27604 26195 27616
rect 26149 27428 26155 27604
rect 26189 27428 26195 27604
rect 26149 27416 26195 27428
rect 26267 27604 26313 27616
rect 26267 27428 26273 27604
rect 26307 27428 26313 27604
rect 26267 27416 26313 27428
rect 26385 27604 26431 27616
rect 26385 27428 26391 27604
rect 26425 27428 26431 27604
rect 26385 27416 26431 27428
rect 26503 27604 26549 27616
rect 26503 27428 26509 27604
rect 26543 27428 26549 27604
rect 26503 27416 26549 27428
rect 23058 27288 23104 27300
rect 25564 27322 25600 27416
rect 25800 27322 25836 27416
rect 26036 27323 26072 27416
rect 26198 27368 26264 27375
rect 26198 27334 26214 27368
rect 26248 27334 26264 27368
rect 26198 27323 26264 27334
rect 26036 27322 26264 27323
rect 25564 27293 26264 27322
rect 25564 27292 26146 27293
rect 22356 27246 22390 27288
rect 22592 27246 22626 27288
rect 22356 27218 22626 27246
rect 22710 27247 22744 27288
rect 22946 27247 22980 27288
rect 22710 27218 22980 27247
rect 22356 27170 22390 27218
rect 22356 27140 22419 27170
rect 22384 27048 22419 27140
rect 22891 27110 22991 27131
rect 22891 27056 22905 27110
rect 22970 27056 22991 27110
rect 22891 27051 22991 27056
rect 23064 27105 23098 27288
rect 25684 27179 25718 27292
rect 26080 27251 26146 27292
rect 26080 27217 26096 27251
rect 26130 27217 26146 27251
rect 26080 27210 26146 27217
rect 26508 27211 26543 27416
rect 26715 27211 26782 27801
rect 28474 27778 28515 27810
rect 28761 27806 28771 27872
rect 28827 27806 28837 27872
rect 29507 27848 29517 27956
rect 29649 27893 29659 27956
rect 29649 27882 29661 27893
rect 29649 27848 29662 27882
rect 29517 27810 29662 27848
rect 29621 27782 29662 27810
rect 27890 27750 28160 27778
rect 27631 27684 27641 27750
rect 27707 27684 27717 27750
rect 27890 27688 27924 27750
rect 28126 27688 28160 27750
rect 28244 27750 28515 27778
rect 29032 27754 29302 27782
rect 28244 27688 28278 27750
rect 28480 27688 28515 27750
rect 28656 27738 28827 27754
rect 28656 27704 28787 27738
rect 28821 27704 28827 27738
rect 28656 27688 28827 27704
rect 29032 27692 29066 27754
rect 29268 27692 29302 27754
rect 29386 27754 29662 27782
rect 29386 27692 29420 27754
rect 29622 27692 29662 27754
rect 27766 27676 27812 27688
rect 27766 27300 27772 27676
rect 27806 27300 27812 27676
rect 27766 27288 27812 27300
rect 27884 27676 27930 27688
rect 27884 27300 27890 27676
rect 27924 27300 27930 27676
rect 27884 27288 27930 27300
rect 28002 27676 28048 27688
rect 28002 27300 28008 27676
rect 28042 27300 28048 27676
rect 28002 27288 28048 27300
rect 28120 27676 28166 27688
rect 28120 27300 28126 27676
rect 28160 27300 28166 27676
rect 28120 27288 28166 27300
rect 28238 27676 28284 27688
rect 28238 27300 28244 27676
rect 28278 27300 28284 27676
rect 28238 27288 28284 27300
rect 28356 27676 28402 27688
rect 28356 27300 28362 27676
rect 28396 27300 28402 27676
rect 28356 27288 28402 27300
rect 28474 27676 28520 27688
rect 28474 27300 28480 27676
rect 28514 27300 28520 27676
rect 28474 27288 28520 27300
rect 26508 27183 26782 27211
rect 26154 27179 26782 27183
rect 25678 27167 25724 27179
rect 24076 27119 24168 27122
rect 23064 27051 23173 27105
rect 22384 27012 22611 27048
rect 22384 26905 22419 27012
rect 22545 26978 22611 27012
rect 22545 26944 22561 26978
rect 22595 26944 22611 26978
rect 22892 27036 22989 27051
rect 22892 26969 22949 27036
rect 22545 26938 22611 26944
rect 22786 26933 23055 26969
rect 22786 26905 22819 26933
rect 23022 26905 23055 26933
rect 23139 26905 23173 27051
rect 23990 27044 24000 27119
rect 24068 27044 24168 27119
rect 24017 27043 24168 27044
rect 22260 26893 22306 26905
rect 22260 26717 22266 26893
rect 22300 26717 22306 26893
rect 22260 26705 22306 26717
rect 22378 26893 22424 26905
rect 22378 26717 22384 26893
rect 22418 26717 22424 26893
rect 22378 26705 22424 26717
rect 22496 26893 22542 26905
rect 22496 26717 22502 26893
rect 22536 26717 22542 26893
rect 22496 26705 22542 26717
rect 22614 26893 22660 26905
rect 22614 26717 22620 26893
rect 22654 26838 22660 26893
rect 22779 26893 22825 26905
rect 22779 26838 22785 26893
rect 22654 26750 22785 26838
rect 22654 26717 22660 26750
rect 22614 26705 22660 26717
rect 22779 26717 22785 26750
rect 22819 26717 22825 26893
rect 22779 26705 22825 26717
rect 22897 26893 22943 26905
rect 22897 26717 22903 26893
rect 22937 26717 22943 26893
rect 22897 26705 22943 26717
rect 23015 26893 23061 26905
rect 23015 26717 23021 26893
rect 23055 26717 23061 26893
rect 23015 26705 23061 26717
rect 23133 26893 23179 26905
rect 23133 26717 23139 26893
rect 23173 26717 23179 26893
rect 23133 26705 23179 26717
rect 22266 26666 22300 26705
rect 22502 26666 22536 26705
rect 22266 26630 22536 26666
rect 22903 26667 22936 26705
rect 23139 26667 23172 26705
rect 22903 26631 23172 26667
rect 22266 26629 22432 26630
rect 22300 26550 22432 26629
rect 22290 26442 22300 26550
rect 22432 26442 22442 26550
rect 18904 26068 19881 26098
rect 22098 26096 22161 26113
rect 22023 26092 22161 26096
rect 18904 25962 18936 26068
rect 19140 25962 19172 26068
rect 19376 25962 19408 26068
rect 19612 25962 19644 26068
rect 19847 25962 19881 26068
rect 20191 26058 22161 26092
rect 20189 26029 22161 26058
rect 20189 26013 20235 26029
rect 22023 26027 22161 26029
rect 18897 25950 18943 25962
rect 18897 25774 18903 25950
rect 18937 25774 18943 25950
rect 18897 25762 18943 25774
rect 19015 25950 19061 25962
rect 19015 25774 19021 25950
rect 19055 25774 19061 25950
rect 19015 25762 19061 25774
rect 19133 25950 19179 25962
rect 19133 25774 19139 25950
rect 19173 25774 19179 25950
rect 19133 25762 19179 25774
rect 19251 25950 19297 25962
rect 19251 25774 19257 25950
rect 19291 25774 19297 25950
rect 19251 25762 19297 25774
rect 19369 25950 19415 25962
rect 19369 25774 19375 25950
rect 19409 25774 19415 25950
rect 19369 25762 19415 25774
rect 19487 25950 19533 25962
rect 19487 25774 19493 25950
rect 19527 25774 19533 25950
rect 19487 25762 19533 25774
rect 19605 25950 19651 25962
rect 19605 25774 19611 25950
rect 19645 25774 19651 25950
rect 19605 25762 19651 25774
rect 19723 25950 19769 25962
rect 19723 25774 19729 25950
rect 19763 25774 19769 25950
rect 19723 25762 19769 25774
rect 19841 25950 19887 25962
rect 19841 25774 19847 25950
rect 19881 25774 19887 25950
rect 19841 25762 19887 25774
rect 19959 25950 20005 25962
rect 19959 25774 19965 25950
rect 19999 25774 20005 25950
rect 19959 25762 20005 25774
rect 19020 25668 19056 25762
rect 19256 25668 19292 25762
rect 19492 25669 19528 25762
rect 19654 25714 19720 25721
rect 19654 25680 19670 25714
rect 19704 25680 19720 25714
rect 19654 25669 19720 25680
rect 19492 25668 19720 25669
rect 19020 25639 19720 25668
rect 19020 25638 19602 25639
rect 19140 25525 19174 25638
rect 19536 25597 19602 25638
rect 19536 25563 19552 25597
rect 19586 25563 19602 25597
rect 19536 25556 19602 25563
rect 19964 25544 19999 25762
rect 20188 25561 20235 26013
rect 21147 25797 21157 25905
rect 21289 25797 21299 25905
rect 23045 25797 23055 25905
rect 23187 25797 23197 25905
rect 21157 25757 21289 25797
rect 23055 25757 23187 25797
rect 21156 25691 21289 25757
rect 23054 25691 23187 25757
rect 20485 25648 21958 25691
rect 20188 25545 20234 25561
rect 20153 25544 20234 25545
rect 19964 25529 20234 25544
rect 19610 25525 20234 25529
rect 19134 25513 19180 25525
rect 18869 25035 18879 25153
rect 18997 25121 19007 25153
rect 19134 25137 19140 25513
rect 19174 25137 19180 25513
rect 19134 25125 19180 25137
rect 19252 25513 19298 25525
rect 19252 25137 19258 25513
rect 19292 25137 19298 25513
rect 19252 25125 19298 25137
rect 19370 25513 19416 25525
rect 19370 25137 19376 25513
rect 19410 25161 19416 25513
rect 19487 25513 19533 25525
rect 19487 25337 19493 25513
rect 19527 25337 19533 25513
rect 19487 25325 19533 25337
rect 19605 25513 20234 25525
rect 19605 25337 19611 25513
rect 19645 25501 20234 25513
rect 19645 25500 19887 25501
rect 19645 25337 19651 25500
rect 20153 25499 20234 25501
rect 20485 25345 20519 25648
rect 20851 25545 20885 25648
rect 21087 25545 21121 25648
rect 21323 25545 21357 25648
rect 21559 25545 21593 25648
rect 20845 25533 20891 25545
rect 19605 25325 19651 25337
rect 20361 25333 20407 25345
rect 19493 25209 19528 25325
rect 19624 25209 19732 25219
rect 19493 25161 19624 25209
rect 19410 25137 19624 25161
rect 19370 25125 19624 25137
rect 19376 25121 19624 25125
rect 18997 25093 19012 25121
rect 18997 25087 19249 25093
rect 18997 25053 19199 25087
rect 19233 25053 19249 25087
rect 18997 25037 19249 25053
rect 19301 25087 19367 25093
rect 19301 25053 19317 25087
rect 19351 25053 19367 25087
rect 19550 25077 19624 25121
rect 20361 25157 20367 25333
rect 20401 25157 20407 25333
rect 20361 25145 20407 25157
rect 20479 25333 20525 25345
rect 20479 25157 20485 25333
rect 20519 25157 20525 25333
rect 20479 25145 20525 25157
rect 20597 25333 20643 25345
rect 20597 25157 20603 25333
rect 20637 25157 20643 25333
rect 20597 25145 20643 25157
rect 20715 25333 20761 25345
rect 20845 25333 20851 25533
rect 20715 25157 20721 25333
rect 20755 25157 20851 25333
rect 20885 25157 20891 25533
rect 20715 25145 20761 25157
rect 20845 25145 20891 25157
rect 20963 25533 21009 25545
rect 20963 25157 20969 25533
rect 21003 25157 21009 25533
rect 20963 25145 21009 25157
rect 21081 25533 21127 25545
rect 21081 25157 21087 25533
rect 21121 25157 21127 25533
rect 21081 25145 21127 25157
rect 21199 25533 21245 25545
rect 21199 25157 21205 25533
rect 21239 25157 21245 25533
rect 21199 25145 21245 25157
rect 21317 25533 21363 25545
rect 21317 25157 21323 25533
rect 21357 25157 21363 25533
rect 21317 25145 21363 25157
rect 21435 25533 21481 25545
rect 21435 25157 21441 25533
rect 21475 25157 21481 25533
rect 21435 25145 21481 25157
rect 21553 25533 21599 25545
rect 21553 25157 21559 25533
rect 21593 25333 21599 25533
rect 21924 25345 21958 25648
rect 22383 25648 23856 25691
rect 22383 25345 22417 25648
rect 22749 25545 22783 25648
rect 22985 25545 23019 25648
rect 23221 25545 23255 25648
rect 23457 25545 23491 25648
rect 22743 25533 22789 25545
rect 21682 25333 21728 25345
rect 21593 25157 21688 25333
rect 21722 25157 21728 25333
rect 21553 25145 21599 25157
rect 21682 25145 21728 25157
rect 21800 25333 21846 25345
rect 21800 25157 21806 25333
rect 21840 25157 21846 25333
rect 21800 25145 21846 25157
rect 21918 25333 21964 25345
rect 21918 25157 21924 25333
rect 21958 25157 21964 25333
rect 21918 25145 21964 25157
rect 22036 25333 22082 25345
rect 22036 25157 22042 25333
rect 22076 25157 22082 25333
rect 22036 25145 22082 25157
rect 22259 25333 22305 25345
rect 22259 25157 22265 25333
rect 22299 25157 22305 25333
rect 22259 25145 22305 25157
rect 22377 25333 22423 25345
rect 22377 25157 22383 25333
rect 22417 25157 22423 25333
rect 22377 25145 22423 25157
rect 22495 25333 22541 25345
rect 22495 25157 22501 25333
rect 22535 25157 22541 25333
rect 22495 25145 22541 25157
rect 22613 25333 22659 25345
rect 22743 25333 22749 25533
rect 22613 25157 22619 25333
rect 22653 25157 22749 25333
rect 22783 25157 22789 25533
rect 22613 25145 22659 25157
rect 22743 25145 22789 25157
rect 22861 25533 22907 25545
rect 22861 25157 22867 25533
rect 22901 25157 22907 25533
rect 22861 25145 22907 25157
rect 22979 25533 23025 25545
rect 22979 25157 22985 25533
rect 23019 25157 23025 25533
rect 22979 25145 23025 25157
rect 23097 25533 23143 25545
rect 23097 25157 23103 25533
rect 23137 25157 23143 25533
rect 23097 25145 23143 25157
rect 23215 25533 23261 25545
rect 23215 25157 23221 25533
rect 23255 25157 23261 25533
rect 23215 25145 23261 25157
rect 23333 25533 23379 25545
rect 23333 25157 23339 25533
rect 23373 25157 23379 25533
rect 23333 25145 23379 25157
rect 23451 25533 23497 25545
rect 23451 25157 23457 25533
rect 23491 25333 23497 25533
rect 23822 25345 23856 25648
rect 23580 25333 23626 25345
rect 23491 25157 23586 25333
rect 23620 25157 23626 25333
rect 23451 25145 23497 25157
rect 23580 25145 23626 25157
rect 23698 25333 23744 25345
rect 23698 25157 23704 25333
rect 23738 25157 23744 25333
rect 23698 25145 23744 25157
rect 23816 25333 23862 25345
rect 23816 25157 23822 25333
rect 23856 25157 23862 25333
rect 23816 25145 23862 25157
rect 23934 25333 23980 25345
rect 23934 25157 23940 25333
rect 23974 25157 23980 25333
rect 24076 25307 24168 27043
rect 24506 26846 24795 26865
rect 24506 26683 24529 26846
rect 24776 26774 24795 26846
rect 25678 26791 25684 27167
rect 25718 26791 25724 27167
rect 25678 26779 25724 26791
rect 25796 27167 25842 27179
rect 25796 26791 25802 27167
rect 25836 26791 25842 27167
rect 25796 26779 25842 26791
rect 25914 27167 25960 27179
rect 25914 26791 25920 27167
rect 25954 26815 25960 27167
rect 26031 27167 26077 27179
rect 26031 26991 26037 27167
rect 26071 26991 26077 27167
rect 26031 26979 26077 26991
rect 26149 27167 26782 27179
rect 26149 26991 26155 27167
rect 26189 27154 26782 27167
rect 27772 27246 27806 27288
rect 28008 27246 28042 27288
rect 27772 27218 28042 27246
rect 28126 27247 28160 27288
rect 28362 27247 28396 27288
rect 28126 27218 28396 27247
rect 27772 27170 27806 27218
rect 26189 26991 26195 27154
rect 27772 27140 27835 27170
rect 26149 26979 26195 26991
rect 27800 27048 27835 27140
rect 27800 27012 28027 27048
rect 28297 27037 28307 27134
rect 28406 27037 28416 27134
rect 28480 27105 28514 27288
rect 28480 27051 28589 27105
rect 26037 26863 26072 26979
rect 27800 26905 27835 27012
rect 27961 26978 28027 27012
rect 27961 26944 27977 26978
rect 28011 26944 28027 26978
rect 28308 27036 28405 27037
rect 28308 26969 28365 27036
rect 27961 26938 28027 26944
rect 28202 26933 28471 26969
rect 28202 26905 28235 26933
rect 28438 26905 28471 26933
rect 28555 26905 28589 27051
rect 27676 26893 27722 26905
rect 26168 26863 26276 26873
rect 26037 26815 26168 26863
rect 25954 26791 26168 26815
rect 25914 26779 26168 26791
rect 25920 26775 26168 26779
rect 24776 26747 25556 26774
rect 24776 26741 25793 26747
rect 24776 26707 25743 26741
rect 25777 26707 25793 26741
rect 24776 26691 25793 26707
rect 25845 26741 25911 26747
rect 25845 26707 25861 26741
rect 25895 26707 25911 26741
rect 26094 26731 26168 26775
rect 26168 26721 26276 26731
rect 24776 26683 25556 26691
rect 24506 26675 25556 26683
rect 24506 26674 25493 26675
rect 24506 26670 25028 26674
rect 24506 26669 24795 26670
rect 24523 25307 24811 25309
rect 24076 25191 24811 25307
rect 23934 25145 23980 25157
rect 24523 25147 24811 25191
rect 19624 25067 19732 25077
rect 20367 25111 20401 25145
rect 20969 25111 21003 25145
rect 21205 25111 21239 25145
rect 20367 25076 20526 25111
rect 20969 25076 21239 25111
rect 21806 25111 21840 25145
rect 22042 25111 22076 25145
rect 21806 25076 22076 25111
rect 22265 25111 22299 25145
rect 22867 25111 22901 25145
rect 23103 25111 23137 25145
rect 22265 25076 22424 25111
rect 22867 25076 23137 25111
rect 23704 25111 23738 25145
rect 23940 25111 23974 25145
rect 23704 25076 23974 25111
rect 18997 25035 19012 25037
rect 18912 25021 19012 25035
rect 18912 24978 19012 24979
rect 18533 24957 19012 24978
rect 19301 24957 19367 25053
rect 18533 24909 19367 24957
rect 18533 24880 19012 24909
rect 18533 24878 18638 24880
rect 18912 24879 19012 24880
rect 18366 24693 18376 24772
rect 18469 24693 18479 24772
rect 18377 23519 18470 24693
rect 19295 24644 19515 24664
rect 19295 24536 19339 24644
rect 19471 24536 19515 24644
rect 19295 24494 19515 24536
rect 18899 24464 19876 24494
rect 18899 24358 18931 24464
rect 19135 24358 19167 24464
rect 19371 24358 19403 24464
rect 19607 24358 19639 24464
rect 19842 24358 19876 24464
rect 18892 24346 18938 24358
rect 18892 24170 18898 24346
rect 18932 24170 18938 24346
rect 18892 24158 18938 24170
rect 19010 24346 19056 24358
rect 19010 24170 19016 24346
rect 19050 24170 19056 24346
rect 19010 24158 19056 24170
rect 19128 24346 19174 24358
rect 19128 24170 19134 24346
rect 19168 24170 19174 24346
rect 19128 24158 19174 24170
rect 19246 24346 19292 24358
rect 19246 24170 19252 24346
rect 19286 24170 19292 24346
rect 19246 24158 19292 24170
rect 19364 24346 19410 24358
rect 19364 24170 19370 24346
rect 19404 24170 19410 24346
rect 19364 24158 19410 24170
rect 19482 24346 19528 24358
rect 19482 24170 19488 24346
rect 19522 24170 19528 24346
rect 19482 24158 19528 24170
rect 19600 24346 19646 24358
rect 19600 24170 19606 24346
rect 19640 24170 19646 24346
rect 19600 24158 19646 24170
rect 19718 24346 19764 24358
rect 19718 24170 19724 24346
rect 19758 24170 19764 24346
rect 19718 24158 19764 24170
rect 19836 24346 19882 24358
rect 19836 24170 19842 24346
rect 19876 24170 19882 24346
rect 19836 24158 19882 24170
rect 19954 24346 20000 24358
rect 19954 24170 19960 24346
rect 19994 24170 20000 24346
rect 19954 24158 20000 24170
rect 20492 24292 20526 25076
rect 21205 25014 21239 25076
rect 20794 24976 21536 25014
rect 20794 24852 20828 24976
rect 21030 24852 21064 24976
rect 21266 24852 21300 24976
rect 21502 24852 21536 24976
rect 21792 24869 21802 24935
rect 21865 24869 21875 24935
rect 20788 24840 20834 24852
rect 20788 24464 20794 24840
rect 20828 24464 20834 24840
rect 20788 24452 20834 24464
rect 20906 24840 20952 24852
rect 20906 24464 20912 24840
rect 20946 24464 20952 24840
rect 20906 24452 20952 24464
rect 21024 24840 21070 24852
rect 21024 24464 21030 24840
rect 21064 24464 21070 24840
rect 21024 24452 21070 24464
rect 21142 24840 21188 24852
rect 21142 24464 21148 24840
rect 21182 24464 21188 24840
rect 21142 24452 21188 24464
rect 21260 24840 21306 24852
rect 21260 24464 21266 24840
rect 21300 24464 21306 24840
rect 21260 24452 21306 24464
rect 21378 24840 21424 24852
rect 21378 24464 21384 24840
rect 21418 24464 21424 24840
rect 21378 24452 21424 24464
rect 21496 24840 21542 24852
rect 21496 24464 21502 24840
rect 21536 24464 21542 24840
rect 21496 24452 21542 24464
rect 21908 24293 21942 25076
rect 21635 24292 21942 24293
rect 20492 24287 20808 24292
rect 21522 24287 21942 24292
rect 20492 24276 20875 24287
rect 20492 24249 20824 24276
rect 19015 24064 19051 24158
rect 19251 24064 19287 24158
rect 19487 24065 19523 24158
rect 19649 24110 19715 24117
rect 19649 24076 19665 24110
rect 19699 24076 19715 24110
rect 19649 24065 19715 24076
rect 19487 24064 19715 24065
rect 19015 24035 19715 24064
rect 19015 24034 19597 24035
rect 19135 23921 19169 24034
rect 19531 23993 19597 24034
rect 19531 23959 19547 23993
rect 19581 23959 19597 23993
rect 19531 23952 19597 23959
rect 19959 23925 19994 24158
rect 20492 24120 20526 24249
rect 20808 24242 20824 24249
rect 20858 24242 20875 24276
rect 20808 24236 20875 24242
rect 21455 24276 21942 24287
rect 21455 24242 21472 24276
rect 21506 24249 21942 24276
rect 21506 24242 21522 24249
rect 21635 24248 21942 24249
rect 21455 24236 21522 24242
rect 20633 24209 20689 24221
rect 20633 24175 20639 24209
rect 20673 24208 20689 24209
rect 21746 24208 21802 24220
rect 20673 24192 21140 24208
rect 20673 24175 21090 24192
rect 20633 24159 21090 24175
rect 21074 24158 21090 24159
rect 21124 24158 21140 24192
rect 21074 24151 21140 24158
rect 21192 24193 21762 24208
rect 21192 24159 21208 24193
rect 21242 24174 21762 24193
rect 21796 24174 21802 24208
rect 21242 24159 21802 24174
rect 21192 24149 21259 24159
rect 21746 24158 21802 24159
rect 21908 24120 21942 24248
rect 22390 24292 22424 25076
rect 23103 25014 23137 25076
rect 22692 24976 23434 25014
rect 22692 24852 22726 24976
rect 22928 24852 22962 24976
rect 23164 24852 23198 24976
rect 23400 24852 23434 24976
rect 22686 24840 22732 24852
rect 22686 24464 22692 24840
rect 22726 24464 22732 24840
rect 22686 24452 22732 24464
rect 22804 24840 22850 24852
rect 22804 24464 22810 24840
rect 22844 24464 22850 24840
rect 22804 24452 22850 24464
rect 22922 24840 22968 24852
rect 22922 24464 22928 24840
rect 22962 24464 22968 24840
rect 22922 24452 22968 24464
rect 23040 24840 23086 24852
rect 23040 24464 23046 24840
rect 23080 24464 23086 24840
rect 23040 24452 23086 24464
rect 23158 24840 23204 24852
rect 23158 24464 23164 24840
rect 23198 24464 23204 24840
rect 23158 24452 23204 24464
rect 23276 24840 23322 24852
rect 23276 24464 23282 24840
rect 23316 24464 23322 24840
rect 23276 24452 23322 24464
rect 23394 24840 23440 24852
rect 23394 24464 23400 24840
rect 23434 24464 23440 24840
rect 23394 24452 23440 24464
rect 23806 24293 23840 25076
rect 24523 25041 24659 25147
rect 24771 25145 24811 25147
rect 24777 25134 24811 25145
rect 24523 25039 24665 25041
rect 24777 25039 24812 25134
rect 24523 25030 24812 25039
rect 24523 25029 24811 25030
rect 24523 25028 24779 25029
rect 23418 24292 23487 24293
rect 23533 24292 23840 24293
rect 22390 24287 22706 24292
rect 23418 24288 23840 24292
rect 22390 24276 22773 24287
rect 22390 24249 22722 24276
rect 22390 24120 22424 24249
rect 22706 24242 22722 24249
rect 22756 24242 22773 24276
rect 22706 24236 22773 24242
rect 23351 24277 23840 24288
rect 23351 24243 23368 24277
rect 23402 24249 23840 24277
rect 23402 24243 23418 24249
rect 23533 24248 23840 24249
rect 23351 24237 23418 24243
rect 22531 24209 22587 24221
rect 22531 24175 22537 24209
rect 22571 24208 22587 24209
rect 23644 24208 23700 24220
rect 22571 24192 23038 24208
rect 22571 24175 22988 24192
rect 22531 24159 22988 24175
rect 22972 24158 22988 24159
rect 23022 24158 23038 24192
rect 22972 24151 23038 24158
rect 23090 24193 23660 24208
rect 23090 24159 23106 24193
rect 23140 24174 23660 24193
rect 23694 24174 23700 24208
rect 23140 24159 23700 24174
rect 23090 24149 23157 24159
rect 23644 24158 23700 24159
rect 23806 24120 23840 24248
rect 23921 24898 23988 24922
rect 23921 24864 23938 24898
rect 23972 24864 23988 24898
rect 19605 23921 19994 23925
rect 19129 23909 19175 23921
rect 19129 23533 19135 23909
rect 19169 23533 19175 23909
rect 19129 23521 19175 23533
rect 19247 23909 19293 23921
rect 19247 23533 19253 23909
rect 19287 23533 19293 23909
rect 19247 23521 19293 23533
rect 19365 23909 19411 23921
rect 19365 23533 19371 23909
rect 19405 23557 19411 23909
rect 19482 23909 19528 23921
rect 19482 23733 19488 23909
rect 19522 23733 19528 23909
rect 19482 23721 19528 23733
rect 19600 23909 19994 23921
rect 20486 24108 20532 24120
rect 20486 23932 20492 24108
rect 20526 23932 20532 24108
rect 20486 23920 20532 23932
rect 20604 24108 20650 24120
rect 20604 23932 20610 24108
rect 20644 23932 20650 24108
rect 20604 23920 20650 23932
rect 20906 24108 20952 24120
rect 19600 23733 19606 23909
rect 19640 23896 19994 23909
rect 19640 23733 19646 23896
rect 19916 23893 19994 23896
rect 19916 23841 19926 23893
rect 19989 23841 19999 23893
rect 19921 23835 19994 23841
rect 19600 23721 19646 23733
rect 19488 23605 19523 23721
rect 20609 23626 20643 23920
rect 20906 23732 20912 24108
rect 20946 23732 20952 24108
rect 20906 23720 20952 23732
rect 21024 24108 21070 24120
rect 21024 23732 21030 24108
rect 21064 23732 21070 24108
rect 21024 23720 21070 23732
rect 21142 24108 21188 24120
rect 21142 23732 21148 24108
rect 21182 23732 21188 24108
rect 21142 23720 21188 23732
rect 21260 24108 21306 24120
rect 21260 23732 21266 24108
rect 21300 23732 21306 24108
rect 21260 23720 21306 23732
rect 21378 24108 21424 24120
rect 21378 23732 21384 24108
rect 21418 23732 21424 24108
rect 21784 24108 21830 24120
rect 21784 23932 21790 24108
rect 21824 23932 21830 24108
rect 21784 23920 21830 23932
rect 21902 24108 21948 24120
rect 21902 23932 21908 24108
rect 21942 23932 21948 24108
rect 21902 23920 21948 23932
rect 22384 24108 22430 24120
rect 22384 23932 22390 24108
rect 22424 23932 22430 24108
rect 22384 23920 22430 23932
rect 22502 24108 22548 24120
rect 22502 23932 22508 24108
rect 22542 23932 22548 24108
rect 22502 23920 22548 23932
rect 22804 24108 22850 24120
rect 21378 23720 21424 23732
rect 21266 23626 21300 23720
rect 21790 23626 21823 23920
rect 19619 23605 19727 23615
rect 19488 23557 19619 23605
rect 19405 23533 19619 23557
rect 19365 23521 19619 23533
rect 18377 23517 18962 23519
rect 19371 23517 19619 23521
rect 18377 23489 19007 23517
rect 12459 23310 12828 23358
rect 12459 23280 12473 23310
rect 12459 23263 12469 23280
rect 6246 23130 10940 23210
rect 12761 23207 12827 23310
rect 17387 23207 17453 23486
rect 18377 23483 19244 23489
rect 18377 23449 19194 23483
rect 19228 23449 19244 23483
rect 18377 23433 19244 23449
rect 19296 23483 19362 23489
rect 19296 23449 19312 23483
rect 19346 23449 19362 23483
rect 19545 23473 19619 23517
rect 20609 23594 21823 23626
rect 22507 23626 22541 23920
rect 22804 23732 22810 24108
rect 22844 23732 22850 24108
rect 22804 23720 22850 23732
rect 22922 24108 22968 24120
rect 22922 23732 22928 24108
rect 22962 23732 22968 24108
rect 22922 23720 22968 23732
rect 23040 24108 23086 24120
rect 23040 23732 23046 24108
rect 23080 23732 23086 24108
rect 23040 23720 23086 23732
rect 23158 24108 23204 24120
rect 23158 23732 23164 24108
rect 23198 23732 23204 24108
rect 23158 23720 23204 23732
rect 23276 24108 23322 24120
rect 23276 23732 23282 24108
rect 23316 23732 23322 24108
rect 23682 24108 23728 24120
rect 23682 23932 23688 24108
rect 23722 23932 23728 24108
rect 23682 23920 23728 23932
rect 23800 24108 23846 24120
rect 23800 23932 23806 24108
rect 23840 23932 23846 24108
rect 23800 23920 23846 23932
rect 23276 23720 23322 23732
rect 23164 23626 23198 23720
rect 23688 23626 23721 23920
rect 22507 23594 23721 23626
rect 21102 23509 21234 23594
rect 23000 23509 23132 23594
rect 19619 23463 19727 23473
rect 18377 23417 19007 23433
rect 18377 23413 18962 23417
rect 18377 23412 18478 23413
rect 18907 23364 19007 23375
rect 18871 23258 18881 23364
rect 18993 23353 19007 23364
rect 19296 23353 19362 23449
rect 21092 23401 21102 23509
rect 21234 23401 21244 23509
rect 22990 23401 23000 23509
rect 23132 23401 23142 23509
rect 23921 23481 23988 24864
rect 24935 24776 25028 26670
rect 25091 26611 25557 26633
rect 25845 26611 25911 26707
rect 27676 26717 27682 26893
rect 27716 26717 27722 26893
rect 27676 26705 27722 26717
rect 27794 26893 27840 26905
rect 27794 26717 27800 26893
rect 27834 26717 27840 26893
rect 27794 26705 27840 26717
rect 27912 26893 27958 26905
rect 27912 26717 27918 26893
rect 27952 26717 27958 26893
rect 27912 26705 27958 26717
rect 28030 26893 28076 26905
rect 28030 26717 28036 26893
rect 28070 26838 28076 26893
rect 28195 26893 28241 26905
rect 28195 26838 28201 26893
rect 28070 26750 28201 26838
rect 28070 26717 28076 26750
rect 28030 26705 28076 26717
rect 28195 26717 28201 26750
rect 28235 26717 28241 26893
rect 28195 26705 28241 26717
rect 28313 26893 28359 26905
rect 28313 26717 28319 26893
rect 28353 26717 28359 26893
rect 28313 26705 28359 26717
rect 28431 26893 28477 26905
rect 28431 26717 28437 26893
rect 28471 26717 28477 26893
rect 28431 26705 28477 26717
rect 28549 26893 28595 26905
rect 28549 26717 28555 26893
rect 28589 26717 28595 26893
rect 28549 26705 28595 26717
rect 27682 26666 27716 26705
rect 27918 26666 27952 26705
rect 27682 26631 27952 26666
rect 28319 26667 28352 26705
rect 28555 26667 28588 26705
rect 28319 26631 28588 26667
rect 25091 26563 25911 26611
rect 27716 26630 27952 26631
rect 25091 26532 25557 26563
rect 27716 26556 27848 26630
rect 25091 26276 25196 26532
rect 27706 26448 27716 26556
rect 27848 26448 27858 26556
rect 25091 26170 25154 26276
rect 25266 26170 25276 26276
rect 25858 26252 26078 26272
rect 25091 26159 25240 26170
rect 25091 24982 25196 26159
rect 25858 26144 25902 26252
rect 26034 26144 26078 26252
rect 25858 26102 26078 26144
rect 28656 26117 28718 27688
rect 28908 27680 28954 27692
rect 28908 27304 28914 27680
rect 28948 27304 28954 27680
rect 28908 27292 28954 27304
rect 29026 27680 29072 27692
rect 29026 27304 29032 27680
rect 29066 27304 29072 27680
rect 29026 27292 29072 27304
rect 29144 27680 29190 27692
rect 29144 27304 29150 27680
rect 29184 27304 29190 27680
rect 29144 27292 29190 27304
rect 29262 27680 29308 27692
rect 29262 27304 29268 27680
rect 29302 27304 29308 27680
rect 29262 27292 29308 27304
rect 29380 27680 29426 27692
rect 29380 27304 29386 27680
rect 29420 27304 29426 27680
rect 29380 27292 29426 27304
rect 29498 27680 29544 27692
rect 29498 27304 29504 27680
rect 29538 27304 29544 27680
rect 29498 27292 29544 27304
rect 29616 27680 29662 27692
rect 29616 27304 29622 27680
rect 29656 27304 29662 27680
rect 29616 27292 29662 27304
rect 28914 27250 28948 27292
rect 29150 27250 29184 27292
rect 28914 27222 29184 27250
rect 29268 27251 29302 27292
rect 29504 27251 29538 27292
rect 29268 27222 29538 27251
rect 28914 27174 28948 27222
rect 28914 27144 28977 27174
rect 28942 27052 28977 27144
rect 29449 27114 29549 27135
rect 29449 27060 29463 27114
rect 29528 27060 29549 27114
rect 29449 27055 29549 27060
rect 29622 27109 29656 27292
rect 30656 27123 31022 27125
rect 29622 27055 29731 27109
rect 28942 27016 29169 27052
rect 28942 26909 28977 27016
rect 29103 26982 29169 27016
rect 29103 26948 29119 26982
rect 29153 26948 29169 26982
rect 29450 27040 29547 27055
rect 29450 26973 29507 27040
rect 29103 26942 29169 26948
rect 29344 26937 29613 26973
rect 29344 26909 29377 26937
rect 29580 26909 29613 26937
rect 29697 26909 29731 27055
rect 30548 27048 30558 27123
rect 30626 27048 31022 27123
rect 30575 27047 31022 27048
rect 30621 27043 31022 27047
rect 28818 26897 28864 26909
rect 28818 26721 28824 26897
rect 28858 26721 28864 26897
rect 28818 26709 28864 26721
rect 28936 26897 28982 26909
rect 28936 26721 28942 26897
rect 28976 26721 28982 26897
rect 28936 26709 28982 26721
rect 29054 26897 29100 26909
rect 29054 26721 29060 26897
rect 29094 26721 29100 26897
rect 29054 26709 29100 26721
rect 29172 26897 29218 26909
rect 29172 26721 29178 26897
rect 29212 26842 29218 26897
rect 29337 26897 29383 26909
rect 29337 26842 29343 26897
rect 29212 26754 29343 26842
rect 29212 26721 29218 26754
rect 29172 26709 29218 26721
rect 29337 26721 29343 26754
rect 29377 26721 29383 26897
rect 29337 26709 29383 26721
rect 29455 26897 29501 26909
rect 29455 26721 29461 26897
rect 29495 26721 29501 26897
rect 29455 26709 29501 26721
rect 29573 26897 29619 26909
rect 29573 26721 29579 26897
rect 29613 26721 29619 26897
rect 29573 26709 29619 26721
rect 29691 26897 29737 26909
rect 29691 26721 29697 26897
rect 29731 26721 29737 26897
rect 29691 26709 29737 26721
rect 28824 26670 28858 26709
rect 29060 26670 29094 26709
rect 28824 26634 29094 26670
rect 29461 26671 29494 26709
rect 29697 26671 29730 26709
rect 29461 26635 29730 26671
rect 28824 26633 28990 26634
rect 28858 26554 28990 26633
rect 28848 26446 28858 26554
rect 28990 26446 29000 26554
rect 30895 26125 31022 27043
rect 25462 26072 26439 26102
rect 28656 26100 28719 26117
rect 28581 26096 28719 26100
rect 25462 25966 25494 26072
rect 25698 25966 25730 26072
rect 25934 25966 25966 26072
rect 26170 25966 26202 26072
rect 26405 25966 26439 26072
rect 26749 26062 28719 26096
rect 26747 26033 28719 26062
rect 26747 26017 26793 26033
rect 28581 26031 28719 26033
rect 30897 26018 31020 26125
rect 25455 25954 25501 25966
rect 25455 25778 25461 25954
rect 25495 25778 25501 25954
rect 25455 25766 25501 25778
rect 25573 25954 25619 25966
rect 25573 25778 25579 25954
rect 25613 25778 25619 25954
rect 25573 25766 25619 25778
rect 25691 25954 25737 25966
rect 25691 25778 25697 25954
rect 25731 25778 25737 25954
rect 25691 25766 25737 25778
rect 25809 25954 25855 25966
rect 25809 25778 25815 25954
rect 25849 25778 25855 25954
rect 25809 25766 25855 25778
rect 25927 25954 25973 25966
rect 25927 25778 25933 25954
rect 25967 25778 25973 25954
rect 25927 25766 25973 25778
rect 26045 25954 26091 25966
rect 26045 25778 26051 25954
rect 26085 25778 26091 25954
rect 26045 25766 26091 25778
rect 26163 25954 26209 25966
rect 26163 25778 26169 25954
rect 26203 25778 26209 25954
rect 26163 25766 26209 25778
rect 26281 25954 26327 25966
rect 26281 25778 26287 25954
rect 26321 25778 26327 25954
rect 26281 25766 26327 25778
rect 26399 25954 26445 25966
rect 26399 25778 26405 25954
rect 26439 25778 26445 25954
rect 26399 25766 26445 25778
rect 26517 25954 26563 25966
rect 26517 25778 26523 25954
rect 26557 25778 26563 25954
rect 26517 25766 26563 25778
rect 25578 25672 25614 25766
rect 25814 25672 25850 25766
rect 26050 25673 26086 25766
rect 26212 25718 26278 25725
rect 26212 25684 26228 25718
rect 26262 25684 26278 25718
rect 26212 25673 26278 25684
rect 26050 25672 26278 25673
rect 25578 25643 26278 25672
rect 25578 25642 26160 25643
rect 25698 25529 25732 25642
rect 26094 25601 26160 25642
rect 26094 25567 26110 25601
rect 26144 25567 26160 25601
rect 26094 25560 26160 25567
rect 26522 25548 26557 25766
rect 26746 25565 26793 26017
rect 27705 25801 27715 25909
rect 27847 25801 27857 25909
rect 29603 25801 29613 25909
rect 29745 25801 29755 25909
rect 27715 25761 27847 25801
rect 29613 25761 29745 25801
rect 27714 25695 27847 25761
rect 29612 25695 29745 25761
rect 27043 25652 28516 25695
rect 26746 25549 26792 25565
rect 26711 25548 26792 25549
rect 26522 25533 26792 25548
rect 26168 25529 26792 25533
rect 25692 25517 25738 25529
rect 25427 25039 25437 25157
rect 25555 25125 25565 25157
rect 25692 25141 25698 25517
rect 25732 25141 25738 25517
rect 25692 25129 25738 25141
rect 25810 25517 25856 25529
rect 25810 25141 25816 25517
rect 25850 25141 25856 25517
rect 25810 25129 25856 25141
rect 25928 25517 25974 25529
rect 25928 25141 25934 25517
rect 25968 25165 25974 25517
rect 26045 25517 26091 25529
rect 26045 25341 26051 25517
rect 26085 25341 26091 25517
rect 26045 25329 26091 25341
rect 26163 25517 26792 25529
rect 26163 25341 26169 25517
rect 26203 25505 26792 25517
rect 26203 25504 26445 25505
rect 26203 25341 26209 25504
rect 26711 25503 26792 25505
rect 27043 25349 27077 25652
rect 27409 25549 27443 25652
rect 27645 25549 27679 25652
rect 27881 25549 27915 25652
rect 28117 25549 28151 25652
rect 27403 25537 27449 25549
rect 26163 25329 26209 25341
rect 26919 25337 26965 25349
rect 26051 25213 26086 25329
rect 26182 25213 26290 25223
rect 26051 25165 26182 25213
rect 25968 25141 26182 25165
rect 25928 25129 26182 25141
rect 25934 25125 26182 25129
rect 25555 25097 25570 25125
rect 25555 25091 25807 25097
rect 25555 25057 25757 25091
rect 25791 25057 25807 25091
rect 25555 25041 25807 25057
rect 25859 25091 25925 25097
rect 25859 25057 25875 25091
rect 25909 25057 25925 25091
rect 26108 25081 26182 25125
rect 26919 25161 26925 25337
rect 26959 25161 26965 25337
rect 26919 25149 26965 25161
rect 27037 25337 27083 25349
rect 27037 25161 27043 25337
rect 27077 25161 27083 25337
rect 27037 25149 27083 25161
rect 27155 25337 27201 25349
rect 27155 25161 27161 25337
rect 27195 25161 27201 25337
rect 27155 25149 27201 25161
rect 27273 25337 27319 25349
rect 27403 25337 27409 25537
rect 27273 25161 27279 25337
rect 27313 25161 27409 25337
rect 27443 25161 27449 25537
rect 27273 25149 27319 25161
rect 27403 25149 27449 25161
rect 27521 25537 27567 25549
rect 27521 25161 27527 25537
rect 27561 25161 27567 25537
rect 27521 25149 27567 25161
rect 27639 25537 27685 25549
rect 27639 25161 27645 25537
rect 27679 25161 27685 25537
rect 27639 25149 27685 25161
rect 27757 25537 27803 25549
rect 27757 25161 27763 25537
rect 27797 25161 27803 25537
rect 27757 25149 27803 25161
rect 27875 25537 27921 25549
rect 27875 25161 27881 25537
rect 27915 25161 27921 25537
rect 27875 25149 27921 25161
rect 27993 25537 28039 25549
rect 27993 25161 27999 25537
rect 28033 25161 28039 25537
rect 27993 25149 28039 25161
rect 28111 25537 28157 25549
rect 28111 25161 28117 25537
rect 28151 25337 28157 25537
rect 28482 25349 28516 25652
rect 28941 25652 30414 25695
rect 28941 25349 28975 25652
rect 29307 25549 29341 25652
rect 29543 25549 29577 25652
rect 29779 25549 29813 25652
rect 30015 25549 30049 25652
rect 29301 25537 29347 25549
rect 28240 25337 28286 25349
rect 28151 25161 28246 25337
rect 28280 25161 28286 25337
rect 28111 25149 28157 25161
rect 28240 25149 28286 25161
rect 28358 25337 28404 25349
rect 28358 25161 28364 25337
rect 28398 25161 28404 25337
rect 28358 25149 28404 25161
rect 28476 25337 28522 25349
rect 28476 25161 28482 25337
rect 28516 25161 28522 25337
rect 28476 25149 28522 25161
rect 28594 25337 28640 25349
rect 28594 25161 28600 25337
rect 28634 25161 28640 25337
rect 28594 25149 28640 25161
rect 28817 25337 28863 25349
rect 28817 25161 28823 25337
rect 28857 25161 28863 25337
rect 28817 25149 28863 25161
rect 28935 25337 28981 25349
rect 28935 25161 28941 25337
rect 28975 25161 28981 25337
rect 28935 25149 28981 25161
rect 29053 25337 29099 25349
rect 29053 25161 29059 25337
rect 29093 25161 29099 25337
rect 29053 25149 29099 25161
rect 29171 25337 29217 25349
rect 29301 25337 29307 25537
rect 29171 25161 29177 25337
rect 29211 25161 29307 25337
rect 29341 25161 29347 25537
rect 29171 25149 29217 25161
rect 29301 25149 29347 25161
rect 29419 25537 29465 25549
rect 29419 25161 29425 25537
rect 29459 25161 29465 25537
rect 29419 25149 29465 25161
rect 29537 25537 29583 25549
rect 29537 25161 29543 25537
rect 29577 25161 29583 25537
rect 29537 25149 29583 25161
rect 29655 25537 29701 25549
rect 29655 25161 29661 25537
rect 29695 25161 29701 25537
rect 29655 25149 29701 25161
rect 29773 25537 29819 25549
rect 29773 25161 29779 25537
rect 29813 25161 29819 25537
rect 29773 25149 29819 25161
rect 29891 25537 29937 25549
rect 29891 25161 29897 25537
rect 29931 25161 29937 25537
rect 29891 25149 29937 25161
rect 30009 25537 30055 25549
rect 30009 25161 30015 25537
rect 30049 25337 30055 25537
rect 30380 25349 30414 25652
rect 30138 25337 30184 25349
rect 30049 25161 30144 25337
rect 30178 25161 30184 25337
rect 30009 25149 30055 25161
rect 30138 25149 30184 25161
rect 30256 25337 30302 25349
rect 30256 25161 30262 25337
rect 30296 25161 30302 25337
rect 30256 25149 30302 25161
rect 30374 25337 30420 25349
rect 30374 25161 30380 25337
rect 30414 25161 30420 25337
rect 30374 25149 30420 25161
rect 30492 25337 30538 25349
rect 30492 25161 30498 25337
rect 30532 25161 30538 25337
rect 30492 25149 30538 25161
rect 26182 25071 26290 25081
rect 26925 25115 26959 25149
rect 27527 25115 27561 25149
rect 27763 25115 27797 25149
rect 26925 25080 27084 25115
rect 27527 25080 27797 25115
rect 28364 25115 28398 25149
rect 28600 25115 28634 25149
rect 28364 25080 28634 25115
rect 28823 25115 28857 25149
rect 29425 25115 29459 25149
rect 29661 25115 29695 25149
rect 28823 25080 28982 25115
rect 29425 25080 29695 25115
rect 30262 25115 30296 25149
rect 30498 25115 30532 25149
rect 30262 25080 30532 25115
rect 25555 25039 25570 25041
rect 25470 25025 25570 25039
rect 25470 24982 25570 24983
rect 25091 24961 25570 24982
rect 25859 24961 25925 25057
rect 25091 24913 25925 24961
rect 25091 24884 25570 24913
rect 25091 24882 25196 24884
rect 25470 24883 25570 24884
rect 24924 24697 24934 24776
rect 25027 24697 25037 24776
rect 24935 23523 25028 24697
rect 25853 24648 26073 24668
rect 25853 24540 25897 24648
rect 26029 24540 26073 24648
rect 25853 24498 26073 24540
rect 25457 24468 26434 24498
rect 25457 24362 25489 24468
rect 25693 24362 25725 24468
rect 25929 24362 25961 24468
rect 26165 24362 26197 24468
rect 26400 24362 26434 24468
rect 25450 24350 25496 24362
rect 25450 24174 25456 24350
rect 25490 24174 25496 24350
rect 25450 24162 25496 24174
rect 25568 24350 25614 24362
rect 25568 24174 25574 24350
rect 25608 24174 25614 24350
rect 25568 24162 25614 24174
rect 25686 24350 25732 24362
rect 25686 24174 25692 24350
rect 25726 24174 25732 24350
rect 25686 24162 25732 24174
rect 25804 24350 25850 24362
rect 25804 24174 25810 24350
rect 25844 24174 25850 24350
rect 25804 24162 25850 24174
rect 25922 24350 25968 24362
rect 25922 24174 25928 24350
rect 25962 24174 25968 24350
rect 25922 24162 25968 24174
rect 26040 24350 26086 24362
rect 26040 24174 26046 24350
rect 26080 24174 26086 24350
rect 26040 24162 26086 24174
rect 26158 24350 26204 24362
rect 26158 24174 26164 24350
rect 26198 24174 26204 24350
rect 26158 24162 26204 24174
rect 26276 24350 26322 24362
rect 26276 24174 26282 24350
rect 26316 24174 26322 24350
rect 26276 24162 26322 24174
rect 26394 24350 26440 24362
rect 26394 24174 26400 24350
rect 26434 24174 26440 24350
rect 26394 24162 26440 24174
rect 26512 24350 26558 24362
rect 26512 24174 26518 24350
rect 26552 24174 26558 24350
rect 26512 24162 26558 24174
rect 27050 24296 27084 25080
rect 27763 25018 27797 25080
rect 27352 24980 28094 25018
rect 27352 24856 27386 24980
rect 27588 24856 27622 24980
rect 27824 24856 27858 24980
rect 28060 24856 28094 24980
rect 28350 24873 28360 24939
rect 28423 24873 28433 24939
rect 27346 24844 27392 24856
rect 27346 24468 27352 24844
rect 27386 24468 27392 24844
rect 27346 24456 27392 24468
rect 27464 24844 27510 24856
rect 27464 24468 27470 24844
rect 27504 24468 27510 24844
rect 27464 24456 27510 24468
rect 27582 24844 27628 24856
rect 27582 24468 27588 24844
rect 27622 24468 27628 24844
rect 27582 24456 27628 24468
rect 27700 24844 27746 24856
rect 27700 24468 27706 24844
rect 27740 24468 27746 24844
rect 27700 24456 27746 24468
rect 27818 24844 27864 24856
rect 27818 24468 27824 24844
rect 27858 24468 27864 24844
rect 27818 24456 27864 24468
rect 27936 24844 27982 24856
rect 27936 24468 27942 24844
rect 27976 24468 27982 24844
rect 27936 24456 27982 24468
rect 28054 24844 28100 24856
rect 28054 24468 28060 24844
rect 28094 24468 28100 24844
rect 28054 24456 28100 24468
rect 28466 24297 28500 25080
rect 28193 24296 28500 24297
rect 27050 24291 27366 24296
rect 28080 24291 28500 24296
rect 27050 24280 27433 24291
rect 27050 24253 27382 24280
rect 25573 24068 25609 24162
rect 25809 24068 25845 24162
rect 26045 24069 26081 24162
rect 26207 24114 26273 24121
rect 26207 24080 26223 24114
rect 26257 24080 26273 24114
rect 26207 24069 26273 24080
rect 26045 24068 26273 24069
rect 25573 24039 26273 24068
rect 25573 24038 26155 24039
rect 25693 23925 25727 24038
rect 26089 23997 26155 24038
rect 26089 23963 26105 23997
rect 26139 23963 26155 23997
rect 26089 23956 26155 23963
rect 26517 23929 26552 24162
rect 27050 24124 27084 24253
rect 27366 24246 27382 24253
rect 27416 24246 27433 24280
rect 27366 24240 27433 24246
rect 28013 24280 28500 24291
rect 28013 24246 28030 24280
rect 28064 24253 28500 24280
rect 28064 24246 28080 24253
rect 28193 24252 28500 24253
rect 28013 24240 28080 24246
rect 27191 24213 27247 24225
rect 27191 24179 27197 24213
rect 27231 24212 27247 24213
rect 28304 24212 28360 24224
rect 27231 24196 27698 24212
rect 27231 24179 27648 24196
rect 27191 24163 27648 24179
rect 27632 24162 27648 24163
rect 27682 24162 27698 24196
rect 27632 24155 27698 24162
rect 27750 24197 28320 24212
rect 27750 24163 27766 24197
rect 27800 24178 28320 24197
rect 28354 24178 28360 24212
rect 27800 24163 28360 24178
rect 27750 24153 27817 24163
rect 28304 24162 28360 24163
rect 28466 24124 28500 24252
rect 28948 24296 28982 25080
rect 29661 25018 29695 25080
rect 29250 24980 29992 25018
rect 29250 24856 29284 24980
rect 29486 24856 29520 24980
rect 29722 24856 29756 24980
rect 29958 24856 29992 24980
rect 29244 24844 29290 24856
rect 29244 24468 29250 24844
rect 29284 24468 29290 24844
rect 29244 24456 29290 24468
rect 29362 24844 29408 24856
rect 29362 24468 29368 24844
rect 29402 24468 29408 24844
rect 29362 24456 29408 24468
rect 29480 24844 29526 24856
rect 29480 24468 29486 24844
rect 29520 24468 29526 24844
rect 29480 24456 29526 24468
rect 29598 24844 29644 24856
rect 29598 24468 29604 24844
rect 29638 24468 29644 24844
rect 29598 24456 29644 24468
rect 29716 24844 29762 24856
rect 29716 24468 29722 24844
rect 29756 24468 29762 24844
rect 29716 24456 29762 24468
rect 29834 24844 29880 24856
rect 29834 24468 29840 24844
rect 29874 24468 29880 24844
rect 29834 24456 29880 24468
rect 29952 24844 29998 24856
rect 29952 24468 29958 24844
rect 29992 24468 29998 24844
rect 29952 24456 29998 24468
rect 30364 24297 30398 25080
rect 29976 24296 30045 24297
rect 30091 24296 30398 24297
rect 28948 24291 29264 24296
rect 29976 24292 30398 24296
rect 28948 24280 29331 24291
rect 28948 24253 29280 24280
rect 28948 24124 28982 24253
rect 29264 24246 29280 24253
rect 29314 24246 29331 24280
rect 29264 24240 29331 24246
rect 29909 24281 30398 24292
rect 29909 24247 29926 24281
rect 29960 24253 30398 24281
rect 29960 24247 29976 24253
rect 30091 24252 30398 24253
rect 29909 24241 29976 24247
rect 29089 24213 29145 24225
rect 29089 24179 29095 24213
rect 29129 24212 29145 24213
rect 30202 24212 30258 24224
rect 29129 24196 29596 24212
rect 29129 24179 29546 24196
rect 29089 24163 29546 24179
rect 29530 24162 29546 24163
rect 29580 24162 29596 24196
rect 29530 24155 29596 24162
rect 29648 24197 30218 24212
rect 29648 24163 29664 24197
rect 29698 24178 30218 24197
rect 30252 24178 30258 24212
rect 29698 24163 30258 24178
rect 29648 24153 29715 24163
rect 30202 24162 30258 24163
rect 30364 24124 30398 24252
rect 30479 24902 30546 24926
rect 30479 24868 30496 24902
rect 30530 24868 30546 24902
rect 26163 23925 26552 23929
rect 25687 23913 25733 23925
rect 25687 23537 25693 23913
rect 25727 23537 25733 23913
rect 25687 23525 25733 23537
rect 25805 23913 25851 23925
rect 25805 23537 25811 23913
rect 25845 23537 25851 23913
rect 25805 23525 25851 23537
rect 25923 23913 25969 23925
rect 25923 23537 25929 23913
rect 25963 23561 25969 23913
rect 26040 23913 26086 23925
rect 26040 23737 26046 23913
rect 26080 23737 26086 23913
rect 26040 23725 26086 23737
rect 26158 23913 26552 23925
rect 27044 24112 27090 24124
rect 27044 23936 27050 24112
rect 27084 23936 27090 24112
rect 27044 23924 27090 23936
rect 27162 24112 27208 24124
rect 27162 23936 27168 24112
rect 27202 23936 27208 24112
rect 27162 23924 27208 23936
rect 27464 24112 27510 24124
rect 26158 23737 26164 23913
rect 26198 23900 26552 23913
rect 26198 23737 26204 23900
rect 26474 23897 26552 23900
rect 26474 23845 26484 23897
rect 26547 23845 26557 23897
rect 26479 23839 26552 23845
rect 26158 23725 26204 23737
rect 26046 23609 26081 23725
rect 27167 23630 27201 23924
rect 27464 23736 27470 24112
rect 27504 23736 27510 24112
rect 27464 23724 27510 23736
rect 27582 24112 27628 24124
rect 27582 23736 27588 24112
rect 27622 23736 27628 24112
rect 27582 23724 27628 23736
rect 27700 24112 27746 24124
rect 27700 23736 27706 24112
rect 27740 23736 27746 24112
rect 27700 23724 27746 23736
rect 27818 24112 27864 24124
rect 27818 23736 27824 24112
rect 27858 23736 27864 24112
rect 27818 23724 27864 23736
rect 27936 24112 27982 24124
rect 27936 23736 27942 24112
rect 27976 23736 27982 24112
rect 28342 24112 28388 24124
rect 28342 23936 28348 24112
rect 28382 23936 28388 24112
rect 28342 23924 28388 23936
rect 28460 24112 28506 24124
rect 28460 23936 28466 24112
rect 28500 23936 28506 24112
rect 28460 23924 28506 23936
rect 28942 24112 28988 24124
rect 28942 23936 28948 24112
rect 28982 23936 28988 24112
rect 28942 23924 28988 23936
rect 29060 24112 29106 24124
rect 29060 23936 29066 24112
rect 29100 23936 29106 24112
rect 29060 23924 29106 23936
rect 29362 24112 29408 24124
rect 27936 23724 27982 23736
rect 27824 23630 27858 23724
rect 28348 23630 28381 23924
rect 26177 23609 26285 23619
rect 26046 23561 26177 23609
rect 25963 23537 26177 23561
rect 25923 23525 26177 23537
rect 24935 23521 25520 23523
rect 25929 23521 26177 23525
rect 24935 23493 25565 23521
rect 24935 23487 25802 23493
rect 18993 23305 19362 23353
rect 18993 23275 19007 23305
rect 18993 23258 19003 23275
rect 12759 23127 17453 23207
rect 19295 23202 19361 23305
rect 23921 23202 23987 23481
rect 24935 23453 25752 23487
rect 25786 23453 25802 23487
rect 24935 23437 25802 23453
rect 25854 23487 25920 23493
rect 25854 23453 25870 23487
rect 25904 23453 25920 23487
rect 26103 23477 26177 23521
rect 27167 23598 28381 23630
rect 29065 23630 29099 23924
rect 29362 23736 29368 24112
rect 29402 23736 29408 24112
rect 29362 23724 29408 23736
rect 29480 24112 29526 24124
rect 29480 23736 29486 24112
rect 29520 23736 29526 24112
rect 29480 23724 29526 23736
rect 29598 24112 29644 24124
rect 29598 23736 29604 24112
rect 29638 23736 29644 24112
rect 29598 23724 29644 23736
rect 29716 24112 29762 24124
rect 29716 23736 29722 24112
rect 29756 23736 29762 24112
rect 29716 23724 29762 23736
rect 29834 24112 29880 24124
rect 29834 23736 29840 24112
rect 29874 23736 29880 24112
rect 30240 24112 30286 24124
rect 30240 23936 30246 24112
rect 30280 23936 30286 24112
rect 30240 23924 30286 23936
rect 30358 24112 30404 24124
rect 30358 23936 30364 24112
rect 30398 23936 30404 24112
rect 30358 23924 30404 23936
rect 29834 23724 29880 23736
rect 29722 23630 29756 23724
rect 30246 23630 30279 23924
rect 29065 23598 30279 23630
rect 27660 23513 27792 23598
rect 29558 23513 29690 23598
rect 26177 23467 26285 23477
rect 24935 23421 25565 23437
rect 24935 23417 25520 23421
rect 24935 23416 25036 23417
rect 25465 23368 25565 23379
rect 25429 23262 25439 23368
rect 25551 23357 25565 23368
rect 25854 23357 25920 23453
rect 27650 23405 27660 23513
rect 27792 23405 27802 23513
rect 29548 23405 29558 23513
rect 29690 23405 29700 23513
rect 30479 23485 30546 24868
rect 25551 23309 25920 23357
rect 25551 23279 25565 23309
rect 25551 23262 25561 23279
rect 25853 23206 25919 23309
rect 30479 23206 30545 23485
rect 19293 23122 23987 23202
rect 25851 23126 30545 23206
rect 491 23083 890 23084
rect 491 23072 11412 23083
rect 491 22994 11268 23072
rect 11396 22994 11412 23072
rect 491 22980 11412 22994
rect 354 22921 17915 22940
rect 354 22810 17781 22921
rect 17892 22810 17915 22921
rect 354 22797 17915 22810
rect 354 22796 17703 22797
rect 194 22738 24516 22750
rect 194 22620 24369 22738
rect 24503 22620 24516 22738
rect 194 22606 24516 22620
rect 5850 22289 5860 22352
rect 5848 22278 5860 22289
rect 5847 22244 5860 22278
rect 5992 22244 6002 22352
rect 6997 22289 7007 22352
rect 6995 22278 7007 22289
rect 6682 22268 6738 22270
rect 5847 22206 5992 22244
rect 5847 22178 5888 22206
rect 6672 22202 6682 22268
rect 6738 22202 6748 22268
rect 6994 22244 7007 22278
rect 7139 22244 7149 22352
rect 9445 22298 9665 22318
rect 7812 22256 7868 22264
rect 7812 22248 8794 22256
rect 6994 22206 7139 22244
rect 7812 22214 7818 22248
rect 7852 22214 8794 22248
rect 5847 22150 6123 22178
rect 5847 22088 5887 22150
rect 6089 22088 6123 22150
rect 6207 22150 6477 22178
rect 6994 22174 7035 22206
rect 7812 22198 8794 22214
rect 7815 22197 8794 22198
rect 6207 22088 6241 22150
rect 6443 22088 6477 22150
rect 6682 22134 6853 22150
rect 6682 22100 6688 22134
rect 6722 22100 6853 22134
rect 5847 22076 5893 22088
rect 5847 21700 5853 22076
rect 5887 21700 5893 22076
rect 5847 21688 5893 21700
rect 5965 22076 6011 22088
rect 5965 21700 5971 22076
rect 6005 21700 6011 22076
rect 5965 21688 6011 21700
rect 6083 22076 6129 22088
rect 6083 21700 6089 22076
rect 6123 21700 6129 22076
rect 6083 21688 6129 21700
rect 6201 22076 6247 22088
rect 6201 21700 6207 22076
rect 6241 21700 6247 22076
rect 6201 21688 6247 21700
rect 6319 22076 6365 22088
rect 6319 21700 6325 22076
rect 6359 21700 6365 22076
rect 6319 21688 6365 21700
rect 6437 22076 6483 22088
rect 6437 21700 6443 22076
rect 6477 21700 6483 22076
rect 6437 21688 6483 21700
rect 6555 22076 6601 22088
rect 6682 22084 6853 22100
rect 6994 22146 7265 22174
rect 6994 22084 7029 22146
rect 7231 22084 7265 22146
rect 7349 22146 7619 22174
rect 7349 22084 7383 22146
rect 7585 22084 7619 22146
rect 6555 21700 6561 22076
rect 6595 21700 6601 22076
rect 6555 21688 6601 21700
rect 5853 21505 5887 21688
rect 5971 21647 6005 21688
rect 6207 21647 6241 21688
rect 5971 21618 6241 21647
rect 6325 21646 6359 21688
rect 6561 21646 6595 21688
rect 6325 21618 6595 21646
rect 6561 21570 6595 21618
rect 6532 21540 6595 21570
rect 5778 21451 5887 21505
rect 5960 21510 6060 21531
rect 5960 21456 5981 21510
rect 6046 21456 6060 21510
rect 5960 21451 6060 21456
rect 5778 21305 5812 21451
rect 5962 21436 6059 21451
rect 6532 21448 6567 21540
rect 6002 21369 6059 21436
rect 6340 21412 6567 21448
rect 6340 21378 6406 21412
rect 5896 21333 6165 21369
rect 6340 21344 6356 21378
rect 6390 21344 6406 21378
rect 6340 21338 6406 21344
rect 5896 21305 5929 21333
rect 6132 21305 6165 21333
rect 6532 21305 6567 21412
rect 5772 21293 5818 21305
rect 5772 21117 5778 21293
rect 5812 21117 5818 21293
rect 5772 21105 5818 21117
rect 5890 21293 5936 21305
rect 5890 21117 5896 21293
rect 5930 21117 5936 21293
rect 5890 21105 5936 21117
rect 6008 21293 6054 21305
rect 6008 21117 6014 21293
rect 6048 21117 6054 21293
rect 6008 21105 6054 21117
rect 6126 21293 6172 21305
rect 6126 21117 6132 21293
rect 6166 21238 6172 21293
rect 6291 21293 6337 21305
rect 6291 21238 6297 21293
rect 6166 21150 6297 21238
rect 6166 21117 6172 21150
rect 6126 21105 6172 21117
rect 6291 21117 6297 21150
rect 6331 21117 6337 21293
rect 6291 21105 6337 21117
rect 6409 21293 6455 21305
rect 6409 21117 6415 21293
rect 6449 21117 6455 21293
rect 6409 21105 6455 21117
rect 6527 21293 6573 21305
rect 6527 21117 6533 21293
rect 6567 21117 6573 21293
rect 6527 21105 6573 21117
rect 6645 21293 6691 21305
rect 6645 21117 6651 21293
rect 6685 21117 6691 21293
rect 6645 21105 6691 21117
rect 5779 21067 5812 21105
rect 6015 21067 6048 21105
rect 5779 21031 6048 21067
rect 6415 21066 6449 21105
rect 6651 21066 6685 21105
rect 6415 21030 6685 21066
rect 6519 21029 6685 21030
rect 6519 20950 6651 21029
rect 6509 20842 6519 20950
rect 6651 20842 6661 20950
rect 6791 20513 6853 22084
rect 6989 22072 7035 22084
rect 6989 21696 6995 22072
rect 7029 21696 7035 22072
rect 6989 21684 7035 21696
rect 7107 22072 7153 22084
rect 7107 21696 7113 22072
rect 7147 21696 7153 22072
rect 7107 21684 7153 21696
rect 7225 22072 7271 22084
rect 7225 21696 7231 22072
rect 7265 21696 7271 22072
rect 7225 21684 7271 21696
rect 7343 22072 7389 22084
rect 7343 21696 7349 22072
rect 7383 21696 7389 22072
rect 7343 21684 7389 21696
rect 7461 22072 7507 22084
rect 7461 21696 7467 22072
rect 7501 21696 7507 22072
rect 7461 21684 7507 21696
rect 7579 22072 7625 22084
rect 7579 21696 7585 22072
rect 7619 21696 7625 22072
rect 7579 21684 7625 21696
rect 7697 22072 7743 22084
rect 7792 22080 7802 22146
rect 7868 22080 7878 22146
rect 7697 21696 7703 22072
rect 7737 21696 7743 22072
rect 7697 21684 7743 21696
rect 6995 21501 7029 21684
rect 7113 21643 7147 21684
rect 7349 21643 7383 21684
rect 7113 21614 7383 21643
rect 7467 21642 7501 21684
rect 7703 21642 7737 21684
rect 7467 21614 7737 21642
rect 7703 21566 7737 21614
rect 7674 21536 7737 21566
rect 8727 21607 8794 22197
rect 9445 22190 9489 22298
rect 9621 22190 9665 22298
rect 12408 22285 12418 22348
rect 12406 22274 12418 22285
rect 9445 22148 9665 22190
rect 12405 22240 12418 22274
rect 12550 22240 12560 22348
rect 13555 22285 13565 22348
rect 13553 22274 13565 22285
rect 13240 22264 13296 22266
rect 12405 22202 12550 22240
rect 12405 22174 12446 22202
rect 13230 22198 13240 22264
rect 13296 22198 13306 22264
rect 13552 22240 13565 22274
rect 13697 22240 13707 22348
rect 16003 22294 16223 22314
rect 14370 22252 14426 22260
rect 14370 22244 15352 22252
rect 13552 22202 13697 22240
rect 14370 22210 14376 22244
rect 14410 22210 15352 22244
rect 9084 22118 10061 22148
rect 9084 22012 9118 22118
rect 9321 22012 9353 22118
rect 9557 22012 9589 22118
rect 9793 22012 9825 22118
rect 10029 22012 10061 22118
rect 12405 22146 12681 22174
rect 12405 22084 12445 22146
rect 12647 22084 12681 22146
rect 12765 22146 13035 22174
rect 13552 22170 13593 22202
rect 14370 22194 15352 22210
rect 14373 22193 15352 22194
rect 12765 22084 12799 22146
rect 13001 22084 13035 22146
rect 13240 22130 13411 22146
rect 13240 22096 13246 22130
rect 13280 22096 13411 22130
rect 12405 22072 12451 22084
rect 8960 22000 9006 22012
rect 8960 21824 8966 22000
rect 9000 21824 9006 22000
rect 8960 21812 9006 21824
rect 9078 22000 9124 22012
rect 9078 21824 9084 22000
rect 9118 21824 9124 22000
rect 9078 21812 9124 21824
rect 9196 22000 9242 22012
rect 9196 21824 9202 22000
rect 9236 21824 9242 22000
rect 9196 21812 9242 21824
rect 9314 22000 9360 22012
rect 9314 21824 9320 22000
rect 9354 21824 9360 22000
rect 9314 21812 9360 21824
rect 9432 22000 9478 22012
rect 9432 21824 9438 22000
rect 9472 21824 9478 22000
rect 9432 21812 9478 21824
rect 9550 22000 9596 22012
rect 9550 21824 9556 22000
rect 9590 21824 9596 22000
rect 9550 21812 9596 21824
rect 9668 22000 9714 22012
rect 9668 21824 9674 22000
rect 9708 21824 9714 22000
rect 9668 21812 9714 21824
rect 9786 22000 9832 22012
rect 9786 21824 9792 22000
rect 9826 21824 9832 22000
rect 9786 21812 9832 21824
rect 9904 22000 9950 22012
rect 9904 21824 9910 22000
rect 9944 21824 9950 22000
rect 9904 21812 9950 21824
rect 10022 22000 10068 22012
rect 10022 21824 10028 22000
rect 10062 21824 10068 22000
rect 10022 21812 10068 21824
rect 8966 21607 9001 21812
rect 9245 21764 9311 21771
rect 9245 21730 9261 21764
rect 9295 21730 9311 21764
rect 9245 21719 9311 21730
rect 9437 21719 9473 21812
rect 9245 21718 9473 21719
rect 9673 21718 9709 21812
rect 9909 21718 9945 21812
rect 9245 21689 9945 21718
rect 8727 21579 9001 21607
rect 9363 21688 9945 21689
rect 12405 21696 12411 22072
rect 12445 21696 12451 22072
rect 9363 21647 9429 21688
rect 9363 21613 9379 21647
rect 9413 21613 9429 21647
rect 9363 21606 9429 21613
rect 8727 21575 9355 21579
rect 9791 21575 9825 21688
rect 12405 21684 12451 21696
rect 12523 22072 12569 22084
rect 12523 21696 12529 22072
rect 12563 21696 12569 22072
rect 12523 21684 12569 21696
rect 12641 22072 12687 22084
rect 12641 21696 12647 22072
rect 12681 21696 12687 22072
rect 12641 21684 12687 21696
rect 12759 22072 12805 22084
rect 12759 21696 12765 22072
rect 12799 21696 12805 22072
rect 12759 21684 12805 21696
rect 12877 22072 12923 22084
rect 12877 21696 12883 22072
rect 12917 21696 12923 22072
rect 12877 21684 12923 21696
rect 12995 22072 13041 22084
rect 12995 21696 13001 22072
rect 13035 21696 13041 22072
rect 12995 21684 13041 21696
rect 13113 22072 13159 22084
rect 13240 22080 13411 22096
rect 13552 22142 13823 22170
rect 13552 22080 13587 22142
rect 13789 22080 13823 22142
rect 13907 22142 14177 22170
rect 13907 22080 13941 22142
rect 14143 22080 14177 22142
rect 13113 21696 13119 22072
rect 13153 21696 13159 22072
rect 13113 21684 13159 21696
rect 8727 21563 9360 21575
rect 8727 21550 9320 21563
rect 6920 21447 7029 21501
rect 6920 21301 6954 21447
rect 7093 21433 7103 21530
rect 7202 21433 7212 21530
rect 7674 21444 7709 21536
rect 7104 21432 7201 21433
rect 7144 21365 7201 21432
rect 7482 21408 7709 21444
rect 7482 21374 7548 21408
rect 7038 21329 7307 21365
rect 7482 21340 7498 21374
rect 7532 21340 7548 21374
rect 7482 21334 7548 21340
rect 7038 21301 7071 21329
rect 7274 21301 7307 21329
rect 7674 21301 7709 21408
rect 9314 21387 9320 21550
rect 9354 21387 9360 21563
rect 9314 21375 9360 21387
rect 9432 21563 9478 21575
rect 9432 21387 9438 21563
rect 9472 21387 9478 21563
rect 9432 21375 9478 21387
rect 9549 21563 9595 21575
rect 6914 21289 6960 21301
rect 6914 21113 6920 21289
rect 6954 21113 6960 21289
rect 6914 21101 6960 21113
rect 7032 21289 7078 21301
rect 7032 21113 7038 21289
rect 7072 21113 7078 21289
rect 7032 21101 7078 21113
rect 7150 21289 7196 21301
rect 7150 21113 7156 21289
rect 7190 21113 7196 21289
rect 7150 21101 7196 21113
rect 7268 21289 7314 21301
rect 7268 21113 7274 21289
rect 7308 21234 7314 21289
rect 7433 21289 7479 21301
rect 7433 21234 7439 21289
rect 7308 21146 7439 21234
rect 7308 21113 7314 21146
rect 7268 21101 7314 21113
rect 7433 21113 7439 21146
rect 7473 21113 7479 21289
rect 7433 21101 7479 21113
rect 7551 21289 7597 21301
rect 7551 21113 7557 21289
rect 7591 21113 7597 21289
rect 7551 21101 7597 21113
rect 7669 21289 7715 21301
rect 7669 21113 7675 21289
rect 7709 21113 7715 21289
rect 7669 21101 7715 21113
rect 7787 21289 7833 21301
rect 7787 21113 7793 21289
rect 7827 21113 7833 21289
rect 9233 21259 9341 21269
rect 9437 21259 9472 21375
rect 9341 21211 9472 21259
rect 9549 21211 9555 21563
rect 9341 21187 9555 21211
rect 9589 21187 9595 21563
rect 9341 21175 9595 21187
rect 9667 21563 9713 21575
rect 9667 21187 9673 21563
rect 9707 21187 9713 21563
rect 9667 21175 9713 21187
rect 9785 21563 9831 21575
rect 9785 21187 9791 21563
rect 9825 21187 9831 21563
rect 11341 21515 11440 21517
rect 11341 21440 11441 21515
rect 11509 21440 11519 21515
rect 12411 21501 12445 21684
rect 12529 21643 12563 21684
rect 12765 21643 12799 21684
rect 12529 21614 12799 21643
rect 12883 21642 12917 21684
rect 13119 21642 13153 21684
rect 12883 21614 13153 21642
rect 13119 21566 13153 21614
rect 13090 21536 13153 21566
rect 12336 21447 12445 21501
rect 12518 21506 12618 21527
rect 12518 21452 12539 21506
rect 12604 21452 12618 21506
rect 12518 21447 12618 21452
rect 11341 21439 11492 21440
rect 9785 21175 9831 21187
rect 10714 21219 11003 21238
rect 9341 21171 9589 21175
rect 9341 21127 9415 21171
rect 10714 21170 10755 21219
rect 9953 21143 10755 21170
rect 9598 21137 9664 21143
rect 9233 21117 9341 21127
rect 7787 21101 7833 21113
rect 9598 21103 9614 21137
rect 9648 21103 9664 21137
rect 6921 21063 6954 21101
rect 7157 21063 7190 21101
rect 6921 21027 7190 21063
rect 7557 21062 7591 21101
rect 7793 21062 7827 21101
rect 7557 21027 7827 21062
rect 7557 21026 7793 21027
rect 7661 20952 7793 21026
rect 9598 21007 9664 21103
rect 9716 21137 10755 21143
rect 9716 21103 9732 21137
rect 9766 21103 10755 21137
rect 9716 21087 10755 21103
rect 9953 21083 10755 21087
rect 10979 21083 11003 21219
rect 9953 21071 11003 21083
rect 10016 21070 11003 21071
rect 10481 21066 11003 21070
rect 9952 21007 10418 21029
rect 9598 20959 10418 21007
rect 7651 20844 7661 20952
rect 7793 20844 7803 20952
rect 9952 20928 10418 20959
rect 10313 20672 10418 20928
rect 6790 20496 6853 20513
rect 9431 20648 9651 20668
rect 9431 20540 9475 20648
rect 9607 20540 9651 20648
rect 10233 20566 10243 20672
rect 10355 20566 10418 20672
rect 10269 20555 10418 20566
rect 9431 20498 9651 20540
rect 6790 20492 6928 20496
rect 6790 20458 8760 20492
rect 9070 20468 10047 20498
rect 6790 20429 8762 20458
rect 6790 20427 6928 20429
rect 8716 20413 8762 20429
rect 5754 20197 5764 20305
rect 5896 20197 5906 20305
rect 7652 20197 7662 20305
rect 7794 20197 7804 20305
rect 5764 20157 5896 20197
rect 7662 20157 7794 20197
rect 5764 20091 5897 20157
rect 7662 20091 7795 20157
rect 5095 20048 6568 20091
rect 5095 19745 5129 20048
rect 5460 19945 5494 20048
rect 5696 19945 5730 20048
rect 5932 19945 5966 20048
rect 6168 19945 6202 20048
rect 5454 19933 5500 19945
rect 4971 19733 5017 19745
rect 4971 19557 4977 19733
rect 5011 19557 5017 19733
rect 4971 19545 5017 19557
rect 5089 19733 5135 19745
rect 5089 19557 5095 19733
rect 5129 19557 5135 19733
rect 5089 19545 5135 19557
rect 5207 19733 5253 19745
rect 5207 19557 5213 19733
rect 5247 19557 5253 19733
rect 5207 19545 5253 19557
rect 5325 19733 5371 19745
rect 5454 19733 5460 19933
rect 5325 19557 5331 19733
rect 5365 19557 5460 19733
rect 5494 19557 5500 19933
rect 5325 19545 5371 19557
rect 5454 19545 5500 19557
rect 5572 19933 5618 19945
rect 5572 19557 5578 19933
rect 5612 19557 5618 19933
rect 5572 19545 5618 19557
rect 5690 19933 5736 19945
rect 5690 19557 5696 19933
rect 5730 19557 5736 19933
rect 5690 19545 5736 19557
rect 5808 19933 5854 19945
rect 5808 19557 5814 19933
rect 5848 19557 5854 19933
rect 5808 19545 5854 19557
rect 5926 19933 5972 19945
rect 5926 19557 5932 19933
rect 5966 19557 5972 19933
rect 5926 19545 5972 19557
rect 6044 19933 6090 19945
rect 6044 19557 6050 19933
rect 6084 19557 6090 19933
rect 6044 19545 6090 19557
rect 6162 19933 6208 19945
rect 6162 19557 6168 19933
rect 6202 19733 6208 19933
rect 6534 19745 6568 20048
rect 6993 20048 8466 20091
rect 6993 19745 7027 20048
rect 7358 19945 7392 20048
rect 7594 19945 7628 20048
rect 7830 19945 7864 20048
rect 8066 19945 8100 20048
rect 7352 19933 7398 19945
rect 6292 19733 6338 19745
rect 6202 19557 6298 19733
rect 6332 19557 6338 19733
rect 6162 19545 6208 19557
rect 6292 19545 6338 19557
rect 6410 19733 6456 19745
rect 6410 19557 6416 19733
rect 6450 19557 6456 19733
rect 6410 19545 6456 19557
rect 6528 19733 6574 19745
rect 6528 19557 6534 19733
rect 6568 19557 6574 19733
rect 6528 19545 6574 19557
rect 6646 19733 6692 19745
rect 6646 19557 6652 19733
rect 6686 19557 6692 19733
rect 6646 19545 6692 19557
rect 6869 19733 6915 19745
rect 6869 19557 6875 19733
rect 6909 19557 6915 19733
rect 6869 19545 6915 19557
rect 6987 19733 7033 19745
rect 6987 19557 6993 19733
rect 7027 19557 7033 19733
rect 6987 19545 7033 19557
rect 7105 19733 7151 19745
rect 7105 19557 7111 19733
rect 7145 19557 7151 19733
rect 7105 19545 7151 19557
rect 7223 19733 7269 19745
rect 7352 19733 7358 19933
rect 7223 19557 7229 19733
rect 7263 19557 7358 19733
rect 7392 19557 7398 19933
rect 7223 19545 7269 19557
rect 7352 19545 7398 19557
rect 7470 19933 7516 19945
rect 7470 19557 7476 19933
rect 7510 19557 7516 19933
rect 7470 19545 7516 19557
rect 7588 19933 7634 19945
rect 7588 19557 7594 19933
rect 7628 19557 7634 19933
rect 7588 19545 7634 19557
rect 7706 19933 7752 19945
rect 7706 19557 7712 19933
rect 7746 19557 7752 19933
rect 7706 19545 7752 19557
rect 7824 19933 7870 19945
rect 7824 19557 7830 19933
rect 7864 19557 7870 19933
rect 7824 19545 7870 19557
rect 7942 19933 7988 19945
rect 7942 19557 7948 19933
rect 7982 19557 7988 19933
rect 7942 19545 7988 19557
rect 8060 19933 8106 19945
rect 8060 19557 8066 19933
rect 8100 19733 8106 19933
rect 8432 19745 8466 20048
rect 8716 19961 8763 20413
rect 9070 20362 9104 20468
rect 9307 20362 9339 20468
rect 9543 20362 9575 20468
rect 9779 20362 9811 20468
rect 10015 20362 10047 20468
rect 8946 20350 8992 20362
rect 8946 20174 8952 20350
rect 8986 20174 8992 20350
rect 8946 20162 8992 20174
rect 9064 20350 9110 20362
rect 9064 20174 9070 20350
rect 9104 20174 9110 20350
rect 9064 20162 9110 20174
rect 9182 20350 9228 20362
rect 9182 20174 9188 20350
rect 9222 20174 9228 20350
rect 9182 20162 9228 20174
rect 9300 20350 9346 20362
rect 9300 20174 9306 20350
rect 9340 20174 9346 20350
rect 9300 20162 9346 20174
rect 9418 20350 9464 20362
rect 9418 20174 9424 20350
rect 9458 20174 9464 20350
rect 9418 20162 9464 20174
rect 9536 20350 9582 20362
rect 9536 20174 9542 20350
rect 9576 20174 9582 20350
rect 9536 20162 9582 20174
rect 9654 20350 9700 20362
rect 9654 20174 9660 20350
rect 9694 20174 9700 20350
rect 9654 20162 9700 20174
rect 9772 20350 9818 20362
rect 9772 20174 9778 20350
rect 9812 20174 9818 20350
rect 9772 20162 9818 20174
rect 9890 20350 9936 20362
rect 9890 20174 9896 20350
rect 9930 20174 9936 20350
rect 9890 20162 9936 20174
rect 10008 20350 10054 20362
rect 10008 20174 10014 20350
rect 10048 20174 10054 20350
rect 10008 20162 10054 20174
rect 8717 19945 8763 19961
rect 8717 19944 8798 19945
rect 8952 19944 8987 20162
rect 9231 20114 9297 20121
rect 9231 20080 9247 20114
rect 9281 20080 9297 20114
rect 9231 20069 9297 20080
rect 9423 20069 9459 20162
rect 9231 20068 9459 20069
rect 9659 20068 9695 20162
rect 9895 20068 9931 20162
rect 9231 20039 9931 20068
rect 9349 20038 9931 20039
rect 9349 19997 9415 20038
rect 9349 19963 9365 19997
rect 9399 19963 9415 19997
rect 9349 19956 9415 19963
rect 8717 19929 8987 19944
rect 8717 19925 9341 19929
rect 9777 19925 9811 20038
rect 8717 19913 9346 19925
rect 8717 19901 9306 19913
rect 8717 19899 8798 19901
rect 9064 19900 9306 19901
rect 8190 19733 8236 19745
rect 8100 19557 8196 19733
rect 8230 19557 8236 19733
rect 8060 19545 8106 19557
rect 8190 19545 8236 19557
rect 8308 19733 8354 19745
rect 8308 19557 8314 19733
rect 8348 19557 8354 19733
rect 8308 19545 8354 19557
rect 8426 19733 8472 19745
rect 8426 19557 8432 19733
rect 8466 19557 8472 19733
rect 8426 19545 8472 19557
rect 8544 19733 8590 19745
rect 8544 19557 8550 19733
rect 8584 19557 8590 19733
rect 9300 19737 9306 19900
rect 9340 19737 9346 19913
rect 9300 19725 9346 19737
rect 9418 19913 9464 19925
rect 9418 19737 9424 19913
rect 9458 19737 9464 19913
rect 9418 19725 9464 19737
rect 9535 19913 9581 19925
rect 8544 19545 8590 19557
rect 9219 19609 9327 19619
rect 9423 19609 9458 19725
rect 4977 19511 5011 19545
rect 5213 19511 5247 19545
rect 4977 19476 5247 19511
rect 5814 19511 5848 19545
rect 6050 19511 6084 19545
rect 6652 19511 6686 19545
rect 5814 19476 6084 19511
rect 6527 19476 6686 19511
rect 6875 19511 6909 19545
rect 7111 19511 7145 19545
rect 6875 19476 7145 19511
rect 7712 19511 7746 19545
rect 7948 19511 7982 19545
rect 8550 19511 8584 19545
rect 7712 19476 7982 19511
rect 8425 19476 8584 19511
rect 9327 19561 9458 19609
rect 9535 19561 9541 19913
rect 9327 19537 9541 19561
rect 9575 19537 9581 19913
rect 9327 19525 9581 19537
rect 9653 19913 9699 19925
rect 9653 19537 9659 19913
rect 9693 19537 9699 19913
rect 9653 19525 9699 19537
rect 9771 19913 9817 19925
rect 9771 19537 9777 19913
rect 9811 19537 9817 19913
rect 9771 19525 9817 19537
rect 9327 19521 9575 19525
rect 9944 19521 9954 19553
rect 9327 19477 9401 19521
rect 9939 19493 9954 19521
rect 9584 19487 9650 19493
rect 4963 19298 5030 19322
rect 4963 19264 4979 19298
rect 5013 19264 5030 19298
rect 4747 18841 4902 18849
rect 4746 18835 4902 18841
rect 4746 18737 4758 18835
rect 4890 18737 4902 18835
rect 4746 16739 4902 18737
rect 4963 17881 5030 19264
rect 5111 18693 5145 19476
rect 5814 19414 5848 19476
rect 5517 19376 6259 19414
rect 5517 19252 5551 19376
rect 5753 19252 5787 19376
rect 5989 19252 6023 19376
rect 6225 19252 6259 19376
rect 5511 19240 5557 19252
rect 5511 18864 5517 19240
rect 5551 18864 5557 19240
rect 5511 18852 5557 18864
rect 5629 19240 5675 19252
rect 5629 18864 5635 19240
rect 5669 18864 5675 19240
rect 5629 18852 5675 18864
rect 5747 19240 5793 19252
rect 5747 18864 5753 19240
rect 5787 18864 5793 19240
rect 5747 18852 5793 18864
rect 5865 19240 5911 19252
rect 5865 18864 5871 19240
rect 5905 18864 5911 19240
rect 5865 18852 5911 18864
rect 5983 19240 6029 19252
rect 5983 18864 5989 19240
rect 6023 18864 6029 19240
rect 5983 18852 6029 18864
rect 6101 19240 6147 19252
rect 6101 18864 6107 19240
rect 6141 18864 6147 19240
rect 6101 18852 6147 18864
rect 6219 19240 6265 19252
rect 6219 18864 6225 19240
rect 6259 18864 6265 19240
rect 6219 18852 6265 18864
rect 5111 18692 5418 18693
rect 5464 18692 5533 18693
rect 6527 18692 6561 19476
rect 5111 18688 5533 18692
rect 5111 18677 5600 18688
rect 6245 18687 6561 18692
rect 5111 18649 5549 18677
rect 5111 18648 5418 18649
rect 5111 18520 5145 18648
rect 5533 18643 5549 18649
rect 5583 18643 5600 18677
rect 5533 18637 5600 18643
rect 6178 18676 6561 18687
rect 6178 18642 6195 18676
rect 6229 18649 6561 18676
rect 6229 18642 6245 18649
rect 6178 18636 6245 18642
rect 5251 18608 5307 18620
rect 6364 18609 6420 18621
rect 6364 18608 6380 18609
rect 5251 18574 5257 18608
rect 5291 18593 5861 18608
rect 5291 18574 5811 18593
rect 5251 18559 5811 18574
rect 5845 18559 5861 18593
rect 5251 18558 5307 18559
rect 5794 18549 5861 18559
rect 5913 18592 6380 18608
rect 5913 18558 5929 18592
rect 5963 18575 6380 18592
rect 6414 18575 6420 18609
rect 5963 18559 6420 18575
rect 5963 18558 5979 18559
rect 5913 18551 5979 18558
rect 6527 18520 6561 18649
rect 7009 18693 7043 19476
rect 7712 19414 7746 19476
rect 7415 19376 8157 19414
rect 7076 19269 7086 19335
rect 7149 19269 7159 19335
rect 7415 19252 7449 19376
rect 7651 19252 7685 19376
rect 7887 19252 7921 19376
rect 8123 19252 8157 19376
rect 7409 19240 7455 19252
rect 7409 18864 7415 19240
rect 7449 18864 7455 19240
rect 7409 18852 7455 18864
rect 7527 19240 7573 19252
rect 7527 18864 7533 19240
rect 7567 18864 7573 19240
rect 7527 18852 7573 18864
rect 7645 19240 7691 19252
rect 7645 18864 7651 19240
rect 7685 18864 7691 19240
rect 7645 18852 7691 18864
rect 7763 19240 7809 19252
rect 7763 18864 7769 19240
rect 7803 18864 7809 19240
rect 7763 18852 7809 18864
rect 7881 19240 7927 19252
rect 7881 18864 7887 19240
rect 7921 18864 7927 19240
rect 7881 18852 7927 18864
rect 7999 19240 8045 19252
rect 7999 18864 8005 19240
rect 8039 18864 8045 19240
rect 7999 18852 8045 18864
rect 8117 19240 8163 19252
rect 8117 18864 8123 19240
rect 8157 18864 8163 19240
rect 8117 18852 8163 18864
rect 7009 18692 7316 18693
rect 8425 18692 8459 19476
rect 9219 19467 9327 19477
rect 9584 19453 9600 19487
rect 9634 19453 9650 19487
rect 9584 19357 9650 19453
rect 9702 19487 9954 19493
rect 9702 19453 9718 19487
rect 9752 19453 9954 19487
rect 9702 19437 9954 19453
rect 9939 19435 9954 19437
rect 10072 19435 10082 19553
rect 9939 19421 10039 19435
rect 9939 19378 10039 19379
rect 10313 19378 10418 20555
rect 9939 19357 10418 19378
rect 9584 19309 10418 19357
rect 9939 19280 10418 19309
rect 9939 19279 10039 19280
rect 10313 19278 10418 19280
rect 10481 19172 10574 21066
rect 10714 21065 11003 21066
rect 10697 20658 10864 20705
rect 10697 20655 10738 20658
rect 10697 20642 10737 20655
rect 10695 20549 10737 20642
rect 10849 20549 10864 20658
rect 10695 20538 10864 20549
rect 10697 20537 10864 20538
rect 11341 19705 11440 21439
rect 12336 21301 12370 21447
rect 12520 21432 12617 21447
rect 13090 21444 13125 21536
rect 12560 21365 12617 21432
rect 12898 21408 13125 21444
rect 12898 21374 12964 21408
rect 12454 21329 12723 21365
rect 12898 21340 12914 21374
rect 12948 21340 12964 21374
rect 12898 21334 12964 21340
rect 12454 21301 12487 21329
rect 12690 21301 12723 21329
rect 13090 21301 13125 21408
rect 12330 21289 12376 21301
rect 12330 21113 12336 21289
rect 12370 21113 12376 21289
rect 12330 21101 12376 21113
rect 12448 21289 12494 21301
rect 12448 21113 12454 21289
rect 12488 21113 12494 21289
rect 12448 21101 12494 21113
rect 12566 21289 12612 21301
rect 12566 21113 12572 21289
rect 12606 21113 12612 21289
rect 12566 21101 12612 21113
rect 12684 21289 12730 21301
rect 12684 21113 12690 21289
rect 12724 21234 12730 21289
rect 12849 21289 12895 21301
rect 12849 21234 12855 21289
rect 12724 21146 12855 21234
rect 12724 21113 12730 21146
rect 12684 21101 12730 21113
rect 12849 21113 12855 21146
rect 12889 21113 12895 21289
rect 12849 21101 12895 21113
rect 12967 21289 13013 21301
rect 12967 21113 12973 21289
rect 13007 21113 13013 21289
rect 12967 21101 13013 21113
rect 13085 21289 13131 21301
rect 13085 21113 13091 21289
rect 13125 21113 13131 21289
rect 13085 21101 13131 21113
rect 13203 21289 13249 21301
rect 13203 21113 13209 21289
rect 13243 21113 13249 21289
rect 13203 21101 13249 21113
rect 12337 21063 12370 21101
rect 12573 21063 12606 21101
rect 12337 21027 12606 21063
rect 12973 21062 13007 21101
rect 13209 21062 13243 21101
rect 12973 21026 13243 21062
rect 13077 21025 13243 21026
rect 13077 20946 13209 21025
rect 13067 20838 13077 20946
rect 13209 20838 13219 20946
rect 13349 20509 13411 22080
rect 13547 22068 13593 22080
rect 13547 21692 13553 22068
rect 13587 21692 13593 22068
rect 13547 21680 13593 21692
rect 13665 22068 13711 22080
rect 13665 21692 13671 22068
rect 13705 21692 13711 22068
rect 13665 21680 13711 21692
rect 13783 22068 13829 22080
rect 13783 21692 13789 22068
rect 13823 21692 13829 22068
rect 13783 21680 13829 21692
rect 13901 22068 13947 22080
rect 13901 21692 13907 22068
rect 13941 21692 13947 22068
rect 13901 21680 13947 21692
rect 14019 22068 14065 22080
rect 14019 21692 14025 22068
rect 14059 21692 14065 22068
rect 14019 21680 14065 21692
rect 14137 22068 14183 22080
rect 14137 21692 14143 22068
rect 14177 21692 14183 22068
rect 14137 21680 14183 21692
rect 14255 22068 14301 22080
rect 14350 22076 14360 22142
rect 14426 22076 14436 22142
rect 14255 21692 14261 22068
rect 14295 21692 14301 22068
rect 14255 21680 14301 21692
rect 13553 21497 13587 21680
rect 13671 21639 13705 21680
rect 13907 21639 13941 21680
rect 13671 21610 13941 21639
rect 14025 21638 14059 21680
rect 14261 21638 14295 21680
rect 14025 21610 14295 21638
rect 14261 21562 14295 21610
rect 14232 21532 14295 21562
rect 15285 21603 15352 22193
rect 16003 22186 16047 22294
rect 16179 22186 16223 22294
rect 18942 22290 18952 22353
rect 18940 22279 18952 22290
rect 16003 22144 16223 22186
rect 18939 22245 18952 22279
rect 19084 22245 19094 22353
rect 20089 22290 20099 22353
rect 20087 22279 20099 22290
rect 19774 22269 19830 22271
rect 18939 22207 19084 22245
rect 18939 22179 18980 22207
rect 19764 22203 19774 22269
rect 19830 22203 19840 22269
rect 20086 22245 20099 22279
rect 20231 22245 20241 22353
rect 22537 22299 22757 22319
rect 20904 22257 20960 22265
rect 20904 22249 21886 22257
rect 20086 22207 20231 22245
rect 20904 22215 20910 22249
rect 20944 22215 21886 22249
rect 18939 22151 19215 22179
rect 15642 22114 16619 22144
rect 15642 22008 15676 22114
rect 15879 22008 15911 22114
rect 16115 22008 16147 22114
rect 16351 22008 16383 22114
rect 16587 22008 16619 22114
rect 18939 22089 18979 22151
rect 19181 22089 19215 22151
rect 19299 22151 19569 22179
rect 20086 22175 20127 22207
rect 20904 22199 21886 22215
rect 20907 22198 21886 22199
rect 19299 22089 19333 22151
rect 19535 22089 19569 22151
rect 19774 22135 19945 22151
rect 19774 22101 19780 22135
rect 19814 22101 19945 22135
rect 18939 22077 18985 22089
rect 15518 21996 15564 22008
rect 15518 21820 15524 21996
rect 15558 21820 15564 21996
rect 15518 21808 15564 21820
rect 15636 21996 15682 22008
rect 15636 21820 15642 21996
rect 15676 21820 15682 21996
rect 15636 21808 15682 21820
rect 15754 21996 15800 22008
rect 15754 21820 15760 21996
rect 15794 21820 15800 21996
rect 15754 21808 15800 21820
rect 15872 21996 15918 22008
rect 15872 21820 15878 21996
rect 15912 21820 15918 21996
rect 15872 21808 15918 21820
rect 15990 21996 16036 22008
rect 15990 21820 15996 21996
rect 16030 21820 16036 21996
rect 15990 21808 16036 21820
rect 16108 21996 16154 22008
rect 16108 21820 16114 21996
rect 16148 21820 16154 21996
rect 16108 21808 16154 21820
rect 16226 21996 16272 22008
rect 16226 21820 16232 21996
rect 16266 21820 16272 21996
rect 16226 21808 16272 21820
rect 16344 21996 16390 22008
rect 16344 21820 16350 21996
rect 16384 21820 16390 21996
rect 16344 21808 16390 21820
rect 16462 21996 16508 22008
rect 16462 21820 16468 21996
rect 16502 21820 16508 21996
rect 16462 21808 16508 21820
rect 16580 21996 16626 22008
rect 16580 21820 16586 21996
rect 16620 21820 16626 21996
rect 16580 21808 16626 21820
rect 15524 21603 15559 21808
rect 15803 21760 15869 21767
rect 15803 21726 15819 21760
rect 15853 21726 15869 21760
rect 15803 21715 15869 21726
rect 15995 21715 16031 21808
rect 15803 21714 16031 21715
rect 16231 21714 16267 21808
rect 16467 21714 16503 21808
rect 15803 21685 16503 21714
rect 18939 21701 18945 22077
rect 18979 21701 18985 22077
rect 18939 21689 18985 21701
rect 19057 22077 19103 22089
rect 19057 21701 19063 22077
rect 19097 21701 19103 22077
rect 19057 21689 19103 21701
rect 19175 22077 19221 22089
rect 19175 21701 19181 22077
rect 19215 21701 19221 22077
rect 19175 21689 19221 21701
rect 19293 22077 19339 22089
rect 19293 21701 19299 22077
rect 19333 21701 19339 22077
rect 19293 21689 19339 21701
rect 19411 22077 19457 22089
rect 19411 21701 19417 22077
rect 19451 21701 19457 22077
rect 19411 21689 19457 21701
rect 19529 22077 19575 22089
rect 19529 21701 19535 22077
rect 19569 21701 19575 22077
rect 19529 21689 19575 21701
rect 19647 22077 19693 22089
rect 19774 22085 19945 22101
rect 20086 22147 20357 22175
rect 20086 22085 20121 22147
rect 20323 22085 20357 22147
rect 20441 22147 20711 22175
rect 20441 22085 20475 22147
rect 20677 22085 20711 22147
rect 19647 21701 19653 22077
rect 19687 21701 19693 22077
rect 19647 21689 19693 21701
rect 15285 21575 15559 21603
rect 15921 21684 16503 21685
rect 15921 21643 15987 21684
rect 15921 21609 15937 21643
rect 15971 21609 15987 21643
rect 15921 21602 15987 21609
rect 15285 21571 15913 21575
rect 16349 21571 16383 21684
rect 15285 21559 15918 21571
rect 15285 21546 15878 21559
rect 13478 21443 13587 21497
rect 13478 21297 13512 21443
rect 13651 21429 13661 21526
rect 13760 21429 13770 21526
rect 14232 21440 14267 21532
rect 13662 21428 13759 21429
rect 13702 21361 13759 21428
rect 14040 21404 14267 21440
rect 14040 21370 14106 21404
rect 13596 21325 13865 21361
rect 14040 21336 14056 21370
rect 14090 21336 14106 21370
rect 14040 21330 14106 21336
rect 13596 21297 13629 21325
rect 13832 21297 13865 21325
rect 14232 21297 14267 21404
rect 15872 21383 15878 21546
rect 15912 21383 15918 21559
rect 15872 21371 15918 21383
rect 15990 21559 16036 21571
rect 15990 21383 15996 21559
rect 16030 21383 16036 21559
rect 15990 21371 16036 21383
rect 16107 21559 16153 21571
rect 13472 21285 13518 21297
rect 13472 21109 13478 21285
rect 13512 21109 13518 21285
rect 13472 21097 13518 21109
rect 13590 21285 13636 21297
rect 13590 21109 13596 21285
rect 13630 21109 13636 21285
rect 13590 21097 13636 21109
rect 13708 21285 13754 21297
rect 13708 21109 13714 21285
rect 13748 21109 13754 21285
rect 13708 21097 13754 21109
rect 13826 21285 13872 21297
rect 13826 21109 13832 21285
rect 13866 21230 13872 21285
rect 13991 21285 14037 21297
rect 13991 21230 13997 21285
rect 13866 21142 13997 21230
rect 13866 21109 13872 21142
rect 13826 21097 13872 21109
rect 13991 21109 13997 21142
rect 14031 21109 14037 21285
rect 13991 21097 14037 21109
rect 14109 21285 14155 21297
rect 14109 21109 14115 21285
rect 14149 21109 14155 21285
rect 14109 21097 14155 21109
rect 14227 21285 14273 21297
rect 14227 21109 14233 21285
rect 14267 21109 14273 21285
rect 14227 21097 14273 21109
rect 14345 21285 14391 21297
rect 14345 21109 14351 21285
rect 14385 21109 14391 21285
rect 15791 21255 15899 21265
rect 15995 21255 16030 21371
rect 15899 21207 16030 21255
rect 16107 21207 16113 21559
rect 15899 21183 16113 21207
rect 16147 21183 16153 21559
rect 15899 21171 16153 21183
rect 16225 21559 16271 21571
rect 16225 21183 16231 21559
rect 16265 21183 16271 21559
rect 16225 21171 16271 21183
rect 16343 21559 16389 21571
rect 16343 21183 16349 21559
rect 16383 21183 16389 21559
rect 17875 21503 17975 21520
rect 17873 21445 17975 21503
rect 18043 21445 18053 21520
rect 18945 21506 18979 21689
rect 19063 21648 19097 21689
rect 19299 21648 19333 21689
rect 19063 21619 19333 21648
rect 19417 21647 19451 21689
rect 19653 21647 19687 21689
rect 19417 21619 19687 21647
rect 19653 21571 19687 21619
rect 19624 21541 19687 21571
rect 18870 21452 18979 21506
rect 19052 21511 19152 21532
rect 19052 21457 19073 21511
rect 19138 21457 19152 21511
rect 19052 21452 19152 21457
rect 17873 21444 18026 21445
rect 16343 21171 16389 21183
rect 17272 21233 17561 21245
rect 15899 21167 16147 21171
rect 15899 21123 15973 21167
rect 17272 21166 17298 21233
rect 16511 21139 17298 21166
rect 16156 21133 16222 21139
rect 15791 21113 15899 21123
rect 14345 21097 14391 21109
rect 16156 21099 16172 21133
rect 16206 21099 16222 21133
rect 13479 21059 13512 21097
rect 13715 21059 13748 21097
rect 13479 21023 13748 21059
rect 14115 21058 14149 21097
rect 14351 21058 14385 21097
rect 14115 21023 14385 21058
rect 14115 21022 14351 21023
rect 14219 20948 14351 21022
rect 16156 21003 16222 21099
rect 16274 21133 17298 21139
rect 16274 21099 16290 21133
rect 16324 21099 17298 21133
rect 16274 21083 17298 21099
rect 16511 21077 17298 21083
rect 17548 21077 17561 21233
rect 16511 21067 17561 21077
rect 16574 21066 17561 21067
rect 17039 21062 17561 21066
rect 16510 21003 16976 21025
rect 16156 20955 16976 21003
rect 14209 20840 14219 20948
rect 14351 20840 14361 20948
rect 16510 20924 16976 20955
rect 16871 20668 16976 20924
rect 13348 20492 13411 20509
rect 15989 20644 16209 20664
rect 15989 20536 16033 20644
rect 16165 20536 16209 20644
rect 16791 20562 16801 20668
rect 16913 20562 16976 20668
rect 16827 20551 16976 20562
rect 15989 20494 16209 20536
rect 13348 20488 13486 20492
rect 13348 20454 15318 20488
rect 15628 20464 16605 20494
rect 13348 20425 15320 20454
rect 13348 20423 13486 20425
rect 15274 20409 15320 20425
rect 12312 20193 12322 20301
rect 12454 20193 12464 20301
rect 14210 20193 14220 20301
rect 14352 20193 14362 20301
rect 12322 20153 12454 20193
rect 14220 20153 14352 20193
rect 12322 20087 12455 20153
rect 14220 20087 14353 20153
rect 11653 20044 13126 20087
rect 11653 19741 11687 20044
rect 12018 19941 12052 20044
rect 12254 19941 12288 20044
rect 12490 19941 12524 20044
rect 12726 19941 12760 20044
rect 12012 19929 12058 19941
rect 10698 19602 11440 19705
rect 11529 19729 11575 19741
rect 10698 19543 10986 19602
rect 10698 19541 10738 19543
rect 10698 19530 10732 19541
rect 10697 19435 10732 19530
rect 10850 19437 10986 19543
rect 11529 19553 11535 19729
rect 11569 19553 11575 19729
rect 11529 19541 11575 19553
rect 11647 19729 11693 19741
rect 11647 19553 11653 19729
rect 11687 19553 11693 19729
rect 11647 19541 11693 19553
rect 11765 19729 11811 19741
rect 11765 19553 11771 19729
rect 11805 19553 11811 19729
rect 11765 19541 11811 19553
rect 11883 19729 11929 19741
rect 12012 19729 12018 19929
rect 11883 19553 11889 19729
rect 11923 19553 12018 19729
rect 12052 19553 12058 19929
rect 11883 19541 11929 19553
rect 12012 19541 12058 19553
rect 12130 19929 12176 19941
rect 12130 19553 12136 19929
rect 12170 19553 12176 19929
rect 12130 19541 12176 19553
rect 12248 19929 12294 19941
rect 12248 19553 12254 19929
rect 12288 19553 12294 19929
rect 12248 19541 12294 19553
rect 12366 19929 12412 19941
rect 12366 19553 12372 19929
rect 12406 19553 12412 19929
rect 12366 19541 12412 19553
rect 12484 19929 12530 19941
rect 12484 19553 12490 19929
rect 12524 19553 12530 19929
rect 12484 19541 12530 19553
rect 12602 19929 12648 19941
rect 12602 19553 12608 19929
rect 12642 19553 12648 19929
rect 12602 19541 12648 19553
rect 12720 19929 12766 19941
rect 12720 19553 12726 19929
rect 12760 19729 12766 19929
rect 13092 19741 13126 20044
rect 13551 20044 15024 20087
rect 13551 19741 13585 20044
rect 13916 19941 13950 20044
rect 14152 19941 14186 20044
rect 14388 19941 14422 20044
rect 14624 19941 14658 20044
rect 13910 19929 13956 19941
rect 12850 19729 12896 19741
rect 12760 19553 12856 19729
rect 12890 19553 12896 19729
rect 12720 19541 12766 19553
rect 12850 19541 12896 19553
rect 12968 19729 13014 19741
rect 12968 19553 12974 19729
rect 13008 19553 13014 19729
rect 12968 19541 13014 19553
rect 13086 19729 13132 19741
rect 13086 19553 13092 19729
rect 13126 19553 13132 19729
rect 13086 19541 13132 19553
rect 13204 19729 13250 19741
rect 13204 19553 13210 19729
rect 13244 19553 13250 19729
rect 13204 19541 13250 19553
rect 13427 19729 13473 19741
rect 13427 19553 13433 19729
rect 13467 19553 13473 19729
rect 13427 19541 13473 19553
rect 13545 19729 13591 19741
rect 13545 19553 13551 19729
rect 13585 19553 13591 19729
rect 13545 19541 13591 19553
rect 13663 19729 13709 19741
rect 13663 19553 13669 19729
rect 13703 19553 13709 19729
rect 13663 19541 13709 19553
rect 13781 19729 13827 19741
rect 13910 19729 13916 19929
rect 13781 19553 13787 19729
rect 13821 19553 13916 19729
rect 13950 19553 13956 19929
rect 13781 19541 13827 19553
rect 13910 19541 13956 19553
rect 14028 19929 14074 19941
rect 14028 19553 14034 19929
rect 14068 19553 14074 19929
rect 14028 19541 14074 19553
rect 14146 19929 14192 19941
rect 14146 19553 14152 19929
rect 14186 19553 14192 19929
rect 14146 19541 14192 19553
rect 14264 19929 14310 19941
rect 14264 19553 14270 19929
rect 14304 19553 14310 19929
rect 14264 19541 14310 19553
rect 14382 19929 14428 19941
rect 14382 19553 14388 19929
rect 14422 19553 14428 19929
rect 14382 19541 14428 19553
rect 14500 19929 14546 19941
rect 14500 19553 14506 19929
rect 14540 19553 14546 19929
rect 14500 19541 14546 19553
rect 14618 19929 14664 19941
rect 14618 19553 14624 19929
rect 14658 19729 14664 19929
rect 14990 19741 15024 20044
rect 15274 19957 15321 20409
rect 15628 20358 15662 20464
rect 15865 20358 15897 20464
rect 16101 20358 16133 20464
rect 16337 20358 16369 20464
rect 16573 20358 16605 20464
rect 15504 20346 15550 20358
rect 15504 20170 15510 20346
rect 15544 20170 15550 20346
rect 15504 20158 15550 20170
rect 15622 20346 15668 20358
rect 15622 20170 15628 20346
rect 15662 20170 15668 20346
rect 15622 20158 15668 20170
rect 15740 20346 15786 20358
rect 15740 20170 15746 20346
rect 15780 20170 15786 20346
rect 15740 20158 15786 20170
rect 15858 20346 15904 20358
rect 15858 20170 15864 20346
rect 15898 20170 15904 20346
rect 15858 20158 15904 20170
rect 15976 20346 16022 20358
rect 15976 20170 15982 20346
rect 16016 20170 16022 20346
rect 15976 20158 16022 20170
rect 16094 20346 16140 20358
rect 16094 20170 16100 20346
rect 16134 20170 16140 20346
rect 16094 20158 16140 20170
rect 16212 20346 16258 20358
rect 16212 20170 16218 20346
rect 16252 20170 16258 20346
rect 16212 20158 16258 20170
rect 16330 20346 16376 20358
rect 16330 20170 16336 20346
rect 16370 20170 16376 20346
rect 16330 20158 16376 20170
rect 16448 20346 16494 20358
rect 16448 20170 16454 20346
rect 16488 20170 16494 20346
rect 16448 20158 16494 20170
rect 16566 20346 16612 20358
rect 16566 20170 16572 20346
rect 16606 20170 16612 20346
rect 16566 20158 16612 20170
rect 15275 19941 15321 19957
rect 15275 19940 15356 19941
rect 15510 19940 15545 20158
rect 15789 20110 15855 20117
rect 15789 20076 15805 20110
rect 15839 20076 15855 20110
rect 15789 20065 15855 20076
rect 15981 20065 16017 20158
rect 15789 20064 16017 20065
rect 16217 20064 16253 20158
rect 16453 20064 16489 20158
rect 15789 20035 16489 20064
rect 15907 20034 16489 20035
rect 15907 19993 15973 20034
rect 15907 19959 15923 19993
rect 15957 19959 15973 19993
rect 15907 19952 15973 19959
rect 15275 19925 15545 19940
rect 15275 19921 15899 19925
rect 16335 19921 16369 20034
rect 15275 19909 15904 19921
rect 15275 19897 15864 19909
rect 15275 19895 15356 19897
rect 15622 19896 15864 19897
rect 14748 19729 14794 19741
rect 14658 19553 14754 19729
rect 14788 19553 14794 19729
rect 14618 19541 14664 19553
rect 14748 19541 14794 19553
rect 14866 19729 14912 19741
rect 14866 19553 14872 19729
rect 14906 19553 14912 19729
rect 14866 19541 14912 19553
rect 14984 19729 15030 19741
rect 14984 19553 14990 19729
rect 15024 19553 15030 19729
rect 14984 19541 15030 19553
rect 15102 19729 15148 19741
rect 15102 19553 15108 19729
rect 15142 19553 15148 19729
rect 15858 19733 15864 19896
rect 15898 19733 15904 19909
rect 15858 19721 15904 19733
rect 15976 19909 16022 19921
rect 15976 19733 15982 19909
rect 16016 19733 16022 19909
rect 15976 19721 16022 19733
rect 16093 19909 16139 19921
rect 15102 19541 15148 19553
rect 15777 19605 15885 19615
rect 15981 19605 16016 19721
rect 11535 19507 11569 19541
rect 11771 19507 11805 19541
rect 11535 19472 11805 19507
rect 12372 19507 12406 19541
rect 12608 19507 12642 19541
rect 13210 19507 13244 19541
rect 12372 19472 12642 19507
rect 13085 19472 13244 19507
rect 13433 19507 13467 19541
rect 13669 19507 13703 19541
rect 13433 19472 13703 19507
rect 14270 19507 14304 19541
rect 14506 19507 14540 19541
rect 15108 19507 15142 19541
rect 14270 19472 14540 19507
rect 14983 19472 15142 19507
rect 15885 19557 16016 19605
rect 16093 19557 16099 19909
rect 15885 19533 16099 19557
rect 16133 19533 16139 19909
rect 15885 19521 16139 19533
rect 16211 19909 16257 19921
rect 16211 19533 16217 19909
rect 16251 19533 16257 19909
rect 16211 19521 16257 19533
rect 16329 19909 16375 19921
rect 16329 19533 16335 19909
rect 16369 19533 16375 19909
rect 16329 19521 16375 19533
rect 15885 19517 16133 19521
rect 16502 19517 16512 19549
rect 15885 19473 15959 19517
rect 16497 19489 16512 19517
rect 16142 19483 16208 19489
rect 10844 19435 10986 19437
rect 10697 19426 10986 19435
rect 10698 19425 10986 19426
rect 10730 19424 10986 19425
rect 11521 19294 11588 19318
rect 11521 19260 11537 19294
rect 11571 19260 11588 19294
rect 10472 19093 10482 19172
rect 10575 19093 10585 19172
rect 9436 19044 9656 19064
rect 9436 18936 9480 19044
rect 9612 18936 9656 19044
rect 9436 18894 9656 18936
rect 9075 18864 10052 18894
rect 9075 18758 9109 18864
rect 9312 18758 9344 18864
rect 9548 18758 9580 18864
rect 9784 18758 9816 18864
rect 10020 18758 10052 18864
rect 7009 18687 7429 18692
rect 8143 18687 8459 18692
rect 7009 18676 7496 18687
rect 7009 18649 7445 18676
rect 7009 18648 7316 18649
rect 7009 18520 7043 18648
rect 7429 18642 7445 18649
rect 7479 18642 7496 18676
rect 7429 18636 7496 18642
rect 8076 18676 8459 18687
rect 8076 18642 8093 18676
rect 8127 18649 8459 18676
rect 8127 18642 8143 18649
rect 8076 18636 8143 18642
rect 7149 18608 7205 18620
rect 8262 18609 8318 18621
rect 8262 18608 8278 18609
rect 7149 18574 7155 18608
rect 7189 18593 7759 18608
rect 7189 18574 7709 18593
rect 7149 18559 7709 18574
rect 7743 18559 7759 18593
rect 7149 18558 7205 18559
rect 7692 18549 7759 18559
rect 7811 18592 8278 18608
rect 7811 18558 7827 18592
rect 7861 18575 8278 18592
rect 8312 18575 8318 18609
rect 7861 18559 8318 18575
rect 7861 18558 7877 18559
rect 7811 18551 7877 18558
rect 8425 18520 8459 18649
rect 8951 18746 8997 18758
rect 8951 18570 8957 18746
rect 8991 18570 8997 18746
rect 8951 18558 8997 18570
rect 9069 18746 9115 18758
rect 9069 18570 9075 18746
rect 9109 18570 9115 18746
rect 9069 18558 9115 18570
rect 9187 18746 9233 18758
rect 9187 18570 9193 18746
rect 9227 18570 9233 18746
rect 9187 18558 9233 18570
rect 9305 18746 9351 18758
rect 9305 18570 9311 18746
rect 9345 18570 9351 18746
rect 9305 18558 9351 18570
rect 9423 18746 9469 18758
rect 9423 18570 9429 18746
rect 9463 18570 9469 18746
rect 9423 18558 9469 18570
rect 9541 18746 9587 18758
rect 9541 18570 9547 18746
rect 9581 18570 9587 18746
rect 9541 18558 9587 18570
rect 9659 18746 9705 18758
rect 9659 18570 9665 18746
rect 9699 18570 9705 18746
rect 9659 18558 9705 18570
rect 9777 18746 9823 18758
rect 9777 18570 9783 18746
rect 9817 18570 9823 18746
rect 9777 18558 9823 18570
rect 9895 18746 9941 18758
rect 9895 18570 9901 18746
rect 9935 18570 9941 18746
rect 9895 18558 9941 18570
rect 10013 18746 10059 18758
rect 10013 18570 10019 18746
rect 10053 18570 10059 18746
rect 10013 18558 10059 18570
rect 5105 18508 5151 18520
rect 5105 18332 5111 18508
rect 5145 18332 5151 18508
rect 5105 18320 5151 18332
rect 5223 18508 5269 18520
rect 5223 18332 5229 18508
rect 5263 18332 5269 18508
rect 5223 18320 5269 18332
rect 5629 18508 5675 18520
rect 5230 18026 5263 18320
rect 5629 18132 5635 18508
rect 5669 18132 5675 18508
rect 5629 18120 5675 18132
rect 5747 18508 5793 18520
rect 5747 18132 5753 18508
rect 5787 18132 5793 18508
rect 5747 18120 5793 18132
rect 5865 18508 5911 18520
rect 5865 18132 5871 18508
rect 5905 18132 5911 18508
rect 5865 18120 5911 18132
rect 5983 18508 6029 18520
rect 5983 18132 5989 18508
rect 6023 18132 6029 18508
rect 5983 18120 6029 18132
rect 6101 18508 6147 18520
rect 6101 18132 6107 18508
rect 6141 18132 6147 18508
rect 6403 18508 6449 18520
rect 6403 18332 6409 18508
rect 6443 18332 6449 18508
rect 6403 18320 6449 18332
rect 6521 18508 6567 18520
rect 6521 18332 6527 18508
rect 6561 18332 6567 18508
rect 6521 18320 6567 18332
rect 7003 18508 7049 18520
rect 7003 18332 7009 18508
rect 7043 18332 7049 18508
rect 7003 18320 7049 18332
rect 7121 18508 7167 18520
rect 7121 18332 7127 18508
rect 7161 18332 7167 18508
rect 7121 18320 7167 18332
rect 7527 18508 7573 18520
rect 6101 18120 6147 18132
rect 5753 18026 5787 18120
rect 6410 18026 6444 18320
rect 5230 17994 6444 18026
rect 7128 18026 7161 18320
rect 7527 18132 7533 18508
rect 7567 18132 7573 18508
rect 7527 18120 7573 18132
rect 7645 18508 7691 18520
rect 7645 18132 7651 18508
rect 7685 18132 7691 18508
rect 7645 18120 7691 18132
rect 7763 18508 7809 18520
rect 7763 18132 7769 18508
rect 7803 18132 7809 18508
rect 7763 18120 7809 18132
rect 7881 18508 7927 18520
rect 7881 18132 7887 18508
rect 7921 18132 7927 18508
rect 7881 18120 7927 18132
rect 7999 18508 8045 18520
rect 7999 18132 8005 18508
rect 8039 18132 8045 18508
rect 8301 18508 8347 18520
rect 8301 18332 8307 18508
rect 8341 18332 8347 18508
rect 8301 18320 8347 18332
rect 8419 18508 8465 18520
rect 8419 18332 8425 18508
rect 8459 18332 8465 18508
rect 8419 18320 8465 18332
rect 8957 18325 8992 18558
rect 9236 18510 9302 18517
rect 9236 18476 9252 18510
rect 9286 18476 9302 18510
rect 9236 18465 9302 18476
rect 9428 18465 9464 18558
rect 9236 18464 9464 18465
rect 9664 18464 9700 18558
rect 9900 18464 9936 18558
rect 9236 18435 9936 18464
rect 9354 18434 9936 18435
rect 9354 18393 9420 18434
rect 9354 18359 9370 18393
rect 9404 18359 9420 18393
rect 9354 18352 9420 18359
rect 8957 18321 9346 18325
rect 9782 18321 9816 18434
rect 7999 18120 8045 18132
rect 7651 18026 7685 18120
rect 8308 18026 8342 18320
rect 8957 18309 9351 18321
rect 8957 18296 9311 18309
rect 8957 18293 9035 18296
rect 8952 18241 8962 18293
rect 9025 18241 9035 18293
rect 8957 18235 9030 18241
rect 9305 18133 9311 18296
rect 9345 18133 9351 18309
rect 9305 18121 9351 18133
rect 9423 18309 9469 18321
rect 9423 18133 9429 18309
rect 9463 18133 9469 18309
rect 9423 18121 9469 18133
rect 9540 18309 9586 18321
rect 7128 17994 8342 18026
rect 9224 18005 9332 18015
rect 9428 18005 9463 18121
rect 5819 17909 5951 17994
rect 7717 17909 7849 17994
rect 4964 17602 5030 17881
rect 5809 17801 5819 17909
rect 5951 17801 5961 17909
rect 7707 17801 7717 17909
rect 7849 17801 7859 17909
rect 9332 17957 9463 18005
rect 9540 17957 9546 18309
rect 9332 17933 9546 17957
rect 9580 17933 9586 18309
rect 9332 17921 9586 17933
rect 9658 18309 9704 18321
rect 9658 17933 9664 18309
rect 9698 17933 9704 18309
rect 9658 17921 9704 17933
rect 9776 18309 9822 18321
rect 9776 17933 9782 18309
rect 9816 17933 9822 18309
rect 9776 17921 9822 17933
rect 9332 17917 9580 17921
rect 10481 17919 10574 19093
rect 9989 17917 10574 17919
rect 9332 17873 9406 17917
rect 9944 17889 10574 17917
rect 9589 17883 9655 17889
rect 9224 17863 9332 17873
rect 9589 17849 9605 17883
rect 9639 17849 9655 17883
rect 9589 17753 9655 17849
rect 9707 17883 10574 17889
rect 9707 17849 9723 17883
rect 9757 17849 10574 17883
rect 9707 17833 10574 17849
rect 9944 17817 10574 17833
rect 9989 17813 10574 17817
rect 10473 17812 10574 17813
rect 11304 18831 11460 18837
rect 11304 18733 11316 18831
rect 11448 18733 11460 18831
rect 9944 17764 10044 17775
rect 9944 17753 9958 17764
rect 9589 17705 9958 17753
rect 9590 17602 9656 17705
rect 9944 17675 9958 17705
rect 9948 17658 9958 17675
rect 10070 17658 10080 17764
rect 4964 17522 9658 17602
rect 11304 16842 11460 18733
rect 11521 17877 11588 19260
rect 11669 18689 11703 19472
rect 12372 19410 12406 19472
rect 12075 19372 12817 19410
rect 12075 19248 12109 19372
rect 12311 19248 12345 19372
rect 12547 19248 12581 19372
rect 12783 19248 12817 19372
rect 12069 19236 12115 19248
rect 12069 18860 12075 19236
rect 12109 18860 12115 19236
rect 12069 18848 12115 18860
rect 12187 19236 12233 19248
rect 12187 18860 12193 19236
rect 12227 18860 12233 19236
rect 12187 18848 12233 18860
rect 12305 19236 12351 19248
rect 12305 18860 12311 19236
rect 12345 18860 12351 19236
rect 12305 18848 12351 18860
rect 12423 19236 12469 19248
rect 12423 18860 12429 19236
rect 12463 18860 12469 19236
rect 12423 18848 12469 18860
rect 12541 19236 12587 19248
rect 12541 18860 12547 19236
rect 12581 18860 12587 19236
rect 12541 18848 12587 18860
rect 12659 19236 12705 19248
rect 12659 18860 12665 19236
rect 12699 18860 12705 19236
rect 12659 18848 12705 18860
rect 12777 19236 12823 19248
rect 12777 18860 12783 19236
rect 12817 18860 12823 19236
rect 12777 18848 12823 18860
rect 11669 18688 11976 18689
rect 12022 18688 12091 18689
rect 13085 18688 13119 19472
rect 11669 18684 12091 18688
rect 11669 18673 12158 18684
rect 12803 18683 13119 18688
rect 11669 18645 12107 18673
rect 11669 18644 11976 18645
rect 11669 18516 11703 18644
rect 12091 18639 12107 18645
rect 12141 18639 12158 18673
rect 12091 18633 12158 18639
rect 12736 18672 13119 18683
rect 12736 18638 12753 18672
rect 12787 18645 13119 18672
rect 12787 18638 12803 18645
rect 12736 18632 12803 18638
rect 11809 18604 11865 18616
rect 12922 18605 12978 18617
rect 12922 18604 12938 18605
rect 11809 18570 11815 18604
rect 11849 18589 12419 18604
rect 11849 18570 12369 18589
rect 11809 18555 12369 18570
rect 12403 18555 12419 18589
rect 11809 18554 11865 18555
rect 12352 18545 12419 18555
rect 12471 18588 12938 18604
rect 12471 18554 12487 18588
rect 12521 18571 12938 18588
rect 12972 18571 12978 18605
rect 12521 18555 12978 18571
rect 12521 18554 12537 18555
rect 12471 18547 12537 18554
rect 13085 18516 13119 18645
rect 13567 18689 13601 19472
rect 14270 19410 14304 19472
rect 13973 19372 14715 19410
rect 13634 19265 13644 19331
rect 13707 19265 13717 19331
rect 13973 19248 14007 19372
rect 14209 19248 14243 19372
rect 14445 19248 14479 19372
rect 14681 19248 14715 19372
rect 13967 19236 14013 19248
rect 13967 18860 13973 19236
rect 14007 18860 14013 19236
rect 13967 18848 14013 18860
rect 14085 19236 14131 19248
rect 14085 18860 14091 19236
rect 14125 18860 14131 19236
rect 14085 18848 14131 18860
rect 14203 19236 14249 19248
rect 14203 18860 14209 19236
rect 14243 18860 14249 19236
rect 14203 18848 14249 18860
rect 14321 19236 14367 19248
rect 14321 18860 14327 19236
rect 14361 18860 14367 19236
rect 14321 18848 14367 18860
rect 14439 19236 14485 19248
rect 14439 18860 14445 19236
rect 14479 18860 14485 19236
rect 14439 18848 14485 18860
rect 14557 19236 14603 19248
rect 14557 18860 14563 19236
rect 14597 18860 14603 19236
rect 14557 18848 14603 18860
rect 14675 19236 14721 19248
rect 14675 18860 14681 19236
rect 14715 18860 14721 19236
rect 14675 18848 14721 18860
rect 13567 18688 13874 18689
rect 14983 18688 15017 19472
rect 15777 19463 15885 19473
rect 16142 19449 16158 19483
rect 16192 19449 16208 19483
rect 16142 19353 16208 19449
rect 16260 19483 16512 19489
rect 16260 19449 16276 19483
rect 16310 19449 16512 19483
rect 16260 19433 16512 19449
rect 16497 19431 16512 19433
rect 16630 19431 16640 19549
rect 16497 19417 16597 19431
rect 16497 19374 16597 19375
rect 16871 19374 16976 20551
rect 16497 19353 16976 19374
rect 16142 19305 16976 19353
rect 16497 19276 16976 19305
rect 16497 19275 16597 19276
rect 16871 19274 16976 19276
rect 17039 19168 17132 21062
rect 17272 21061 17561 21062
rect 17255 20651 17425 20704
rect 17255 20638 17295 20651
rect 17253 20545 17295 20638
rect 17407 20545 17425 20651
rect 17253 20534 17425 20545
rect 17255 20533 17425 20534
rect 17873 19704 17973 21444
rect 18870 21306 18904 21452
rect 19054 21437 19151 21452
rect 19624 21449 19659 21541
rect 19094 21370 19151 21437
rect 19432 21413 19659 21449
rect 19432 21379 19498 21413
rect 18988 21334 19257 21370
rect 19432 21345 19448 21379
rect 19482 21345 19498 21379
rect 19432 21339 19498 21345
rect 18988 21306 19021 21334
rect 19224 21306 19257 21334
rect 19624 21306 19659 21413
rect 18864 21294 18910 21306
rect 18864 21118 18870 21294
rect 18904 21118 18910 21294
rect 18864 21106 18910 21118
rect 18982 21294 19028 21306
rect 18982 21118 18988 21294
rect 19022 21118 19028 21294
rect 18982 21106 19028 21118
rect 19100 21294 19146 21306
rect 19100 21118 19106 21294
rect 19140 21118 19146 21294
rect 19100 21106 19146 21118
rect 19218 21294 19264 21306
rect 19218 21118 19224 21294
rect 19258 21239 19264 21294
rect 19383 21294 19429 21306
rect 19383 21239 19389 21294
rect 19258 21151 19389 21239
rect 19258 21118 19264 21151
rect 19218 21106 19264 21118
rect 19383 21118 19389 21151
rect 19423 21118 19429 21294
rect 19383 21106 19429 21118
rect 19501 21294 19547 21306
rect 19501 21118 19507 21294
rect 19541 21118 19547 21294
rect 19501 21106 19547 21118
rect 19619 21294 19665 21306
rect 19619 21118 19625 21294
rect 19659 21118 19665 21294
rect 19619 21106 19665 21118
rect 19737 21294 19783 21306
rect 19737 21118 19743 21294
rect 19777 21118 19783 21294
rect 19737 21106 19783 21118
rect 18871 21068 18904 21106
rect 19107 21068 19140 21106
rect 18871 21032 19140 21068
rect 19507 21067 19541 21106
rect 19743 21067 19777 21106
rect 19507 21031 19777 21067
rect 19611 21030 19777 21031
rect 19611 20951 19743 21030
rect 19601 20843 19611 20951
rect 19743 20843 19753 20951
rect 19883 20514 19945 22085
rect 20081 22073 20127 22085
rect 20081 21697 20087 22073
rect 20121 21697 20127 22073
rect 20081 21685 20127 21697
rect 20199 22073 20245 22085
rect 20199 21697 20205 22073
rect 20239 21697 20245 22073
rect 20199 21685 20245 21697
rect 20317 22073 20363 22085
rect 20317 21697 20323 22073
rect 20357 21697 20363 22073
rect 20317 21685 20363 21697
rect 20435 22073 20481 22085
rect 20435 21697 20441 22073
rect 20475 21697 20481 22073
rect 20435 21685 20481 21697
rect 20553 22073 20599 22085
rect 20553 21697 20559 22073
rect 20593 21697 20599 22073
rect 20553 21685 20599 21697
rect 20671 22073 20717 22085
rect 20671 21697 20677 22073
rect 20711 21697 20717 22073
rect 20671 21685 20717 21697
rect 20789 22073 20835 22085
rect 20884 22081 20894 22147
rect 20960 22081 20970 22147
rect 20789 21697 20795 22073
rect 20829 21697 20835 22073
rect 20789 21685 20835 21697
rect 20087 21502 20121 21685
rect 20205 21644 20239 21685
rect 20441 21644 20475 21685
rect 20205 21615 20475 21644
rect 20559 21643 20593 21685
rect 20795 21643 20829 21685
rect 20559 21615 20829 21643
rect 20795 21567 20829 21615
rect 20766 21537 20829 21567
rect 21819 21608 21886 22198
rect 22537 22191 22581 22299
rect 22713 22191 22757 22299
rect 25455 22293 25465 22356
rect 25453 22282 25465 22293
rect 22537 22149 22757 22191
rect 25452 22248 25465 22282
rect 25597 22248 25607 22356
rect 26602 22293 26612 22356
rect 26600 22282 26612 22293
rect 26287 22272 26343 22274
rect 25452 22210 25597 22248
rect 25452 22182 25493 22210
rect 26277 22206 26287 22272
rect 26343 22206 26353 22272
rect 26599 22248 26612 22282
rect 26744 22248 26754 22356
rect 29050 22302 29270 22322
rect 27417 22260 27473 22268
rect 27417 22252 28399 22260
rect 26599 22210 26744 22248
rect 27417 22218 27423 22252
rect 27457 22218 28399 22252
rect 25452 22154 25728 22182
rect 22176 22119 23153 22149
rect 22176 22013 22210 22119
rect 22413 22013 22445 22119
rect 22649 22013 22681 22119
rect 22885 22013 22917 22119
rect 23121 22013 23153 22119
rect 25452 22092 25492 22154
rect 25694 22092 25728 22154
rect 25812 22154 26082 22182
rect 26599 22178 26640 22210
rect 27417 22202 28399 22218
rect 27420 22201 28399 22202
rect 25812 22092 25846 22154
rect 26048 22092 26082 22154
rect 26287 22138 26458 22154
rect 26287 22104 26293 22138
rect 26327 22104 26458 22138
rect 25452 22080 25498 22092
rect 22052 22001 22098 22013
rect 22052 21825 22058 22001
rect 22092 21825 22098 22001
rect 22052 21813 22098 21825
rect 22170 22001 22216 22013
rect 22170 21825 22176 22001
rect 22210 21825 22216 22001
rect 22170 21813 22216 21825
rect 22288 22001 22334 22013
rect 22288 21825 22294 22001
rect 22328 21825 22334 22001
rect 22288 21813 22334 21825
rect 22406 22001 22452 22013
rect 22406 21825 22412 22001
rect 22446 21825 22452 22001
rect 22406 21813 22452 21825
rect 22524 22001 22570 22013
rect 22524 21825 22530 22001
rect 22564 21825 22570 22001
rect 22524 21813 22570 21825
rect 22642 22001 22688 22013
rect 22642 21825 22648 22001
rect 22682 21825 22688 22001
rect 22642 21813 22688 21825
rect 22760 22001 22806 22013
rect 22760 21825 22766 22001
rect 22800 21825 22806 22001
rect 22760 21813 22806 21825
rect 22878 22001 22924 22013
rect 22878 21825 22884 22001
rect 22918 21825 22924 22001
rect 22878 21813 22924 21825
rect 22996 22001 23042 22013
rect 22996 21825 23002 22001
rect 23036 21825 23042 22001
rect 22996 21813 23042 21825
rect 23114 22001 23160 22013
rect 23114 21825 23120 22001
rect 23154 21825 23160 22001
rect 23114 21813 23160 21825
rect 22058 21608 22093 21813
rect 22337 21765 22403 21772
rect 22337 21731 22353 21765
rect 22387 21731 22403 21765
rect 22337 21720 22403 21731
rect 22529 21720 22565 21813
rect 22337 21719 22565 21720
rect 22765 21719 22801 21813
rect 23001 21719 23037 21813
rect 22337 21690 23037 21719
rect 25452 21704 25458 22080
rect 25492 21704 25498 22080
rect 25452 21692 25498 21704
rect 25570 22080 25616 22092
rect 25570 21704 25576 22080
rect 25610 21704 25616 22080
rect 25570 21692 25616 21704
rect 25688 22080 25734 22092
rect 25688 21704 25694 22080
rect 25728 21704 25734 22080
rect 25688 21692 25734 21704
rect 25806 22080 25852 22092
rect 25806 21704 25812 22080
rect 25846 21704 25852 22080
rect 25806 21692 25852 21704
rect 25924 22080 25970 22092
rect 25924 21704 25930 22080
rect 25964 21704 25970 22080
rect 25924 21692 25970 21704
rect 26042 22080 26088 22092
rect 26042 21704 26048 22080
rect 26082 21704 26088 22080
rect 26042 21692 26088 21704
rect 26160 22080 26206 22092
rect 26287 22088 26458 22104
rect 26599 22150 26870 22178
rect 26599 22088 26634 22150
rect 26836 22088 26870 22150
rect 26954 22150 27224 22178
rect 26954 22088 26988 22150
rect 27190 22088 27224 22150
rect 26160 21704 26166 22080
rect 26200 21704 26206 22080
rect 26160 21692 26206 21704
rect 21819 21580 22093 21608
rect 22455 21689 23037 21690
rect 22455 21648 22521 21689
rect 22455 21614 22471 21648
rect 22505 21614 22521 21648
rect 22455 21607 22521 21614
rect 21819 21576 22447 21580
rect 22883 21576 22917 21689
rect 21819 21564 22452 21576
rect 21819 21551 22412 21564
rect 20012 21448 20121 21502
rect 20012 21302 20046 21448
rect 20185 21434 20195 21531
rect 20294 21434 20304 21531
rect 20766 21445 20801 21537
rect 20196 21433 20293 21434
rect 20236 21366 20293 21433
rect 20574 21409 20801 21445
rect 20574 21375 20640 21409
rect 20130 21330 20399 21366
rect 20574 21341 20590 21375
rect 20624 21341 20640 21375
rect 20574 21335 20640 21341
rect 20130 21302 20163 21330
rect 20366 21302 20399 21330
rect 20766 21302 20801 21409
rect 22406 21388 22412 21551
rect 22446 21388 22452 21564
rect 22406 21376 22452 21388
rect 22524 21564 22570 21576
rect 22524 21388 22530 21564
rect 22564 21388 22570 21564
rect 22524 21376 22570 21388
rect 22641 21564 22687 21576
rect 20006 21290 20052 21302
rect 20006 21114 20012 21290
rect 20046 21114 20052 21290
rect 20006 21102 20052 21114
rect 20124 21290 20170 21302
rect 20124 21114 20130 21290
rect 20164 21114 20170 21290
rect 20124 21102 20170 21114
rect 20242 21290 20288 21302
rect 20242 21114 20248 21290
rect 20282 21114 20288 21290
rect 20242 21102 20288 21114
rect 20360 21290 20406 21302
rect 20360 21114 20366 21290
rect 20400 21235 20406 21290
rect 20525 21290 20571 21302
rect 20525 21235 20531 21290
rect 20400 21147 20531 21235
rect 20400 21114 20406 21147
rect 20360 21102 20406 21114
rect 20525 21114 20531 21147
rect 20565 21114 20571 21290
rect 20525 21102 20571 21114
rect 20643 21290 20689 21302
rect 20643 21114 20649 21290
rect 20683 21114 20689 21290
rect 20643 21102 20689 21114
rect 20761 21290 20807 21302
rect 20761 21114 20767 21290
rect 20801 21114 20807 21290
rect 20761 21102 20807 21114
rect 20879 21290 20925 21302
rect 20879 21114 20885 21290
rect 20919 21114 20925 21290
rect 22325 21260 22433 21270
rect 22529 21260 22564 21376
rect 22433 21212 22564 21260
rect 22641 21212 22647 21564
rect 22433 21188 22647 21212
rect 22681 21188 22687 21564
rect 22433 21176 22687 21188
rect 22759 21564 22805 21576
rect 22759 21188 22765 21564
rect 22799 21188 22805 21564
rect 22759 21176 22805 21188
rect 22877 21564 22923 21576
rect 22877 21188 22883 21564
rect 22917 21188 22923 21564
rect 24388 21448 24488 21523
rect 24556 21448 24566 21523
rect 25458 21509 25492 21692
rect 25576 21651 25610 21692
rect 25812 21651 25846 21692
rect 25576 21622 25846 21651
rect 25930 21650 25964 21692
rect 26166 21650 26200 21692
rect 25930 21622 26200 21650
rect 26166 21574 26200 21622
rect 26137 21544 26200 21574
rect 25383 21455 25492 21509
rect 25565 21514 25665 21535
rect 25565 21460 25586 21514
rect 25651 21460 25665 21514
rect 25565 21455 25665 21460
rect 24388 21447 24539 21448
rect 22877 21176 22923 21188
rect 23806 21222 24095 21240
rect 22433 21172 22681 21176
rect 22433 21128 22507 21172
rect 23806 21171 23847 21222
rect 23045 21144 23847 21171
rect 22690 21138 22756 21144
rect 22325 21118 22433 21128
rect 20879 21102 20925 21114
rect 22690 21104 22706 21138
rect 22740 21104 22756 21138
rect 20013 21064 20046 21102
rect 20249 21064 20282 21102
rect 20013 21028 20282 21064
rect 20649 21063 20683 21102
rect 20885 21063 20919 21102
rect 20649 21028 20919 21063
rect 20649 21027 20885 21028
rect 20753 20953 20885 21027
rect 22690 21008 22756 21104
rect 22808 21138 23847 21144
rect 22808 21104 22824 21138
rect 22858 21104 23847 21138
rect 22808 21088 23847 21104
rect 23045 21085 23847 21088
rect 24075 21085 24095 21222
rect 23045 21072 24095 21085
rect 23108 21071 24095 21072
rect 23573 21067 24095 21071
rect 23044 21008 23510 21030
rect 22690 20960 23510 21008
rect 20743 20845 20753 20953
rect 20885 20845 20895 20953
rect 23044 20929 23510 20960
rect 23405 20673 23510 20929
rect 19882 20497 19945 20514
rect 22523 20649 22743 20669
rect 22523 20541 22567 20649
rect 22699 20541 22743 20649
rect 23325 20567 23335 20673
rect 23447 20567 23510 20673
rect 23361 20556 23510 20567
rect 22523 20499 22743 20541
rect 19882 20493 20020 20497
rect 19882 20459 21852 20493
rect 22162 20469 23139 20499
rect 19882 20430 21854 20459
rect 19882 20428 20020 20430
rect 21808 20414 21854 20430
rect 18846 20198 18856 20306
rect 18988 20198 18998 20306
rect 20744 20198 20754 20306
rect 20886 20198 20896 20306
rect 18856 20158 18988 20198
rect 20754 20158 20886 20198
rect 18856 20092 18989 20158
rect 20754 20092 20887 20158
rect 18187 20049 19660 20092
rect 18187 19746 18221 20049
rect 18552 19946 18586 20049
rect 18788 19946 18822 20049
rect 19024 19946 19058 20049
rect 19260 19946 19294 20049
rect 18546 19934 18592 19946
rect 17288 19701 17973 19704
rect 17256 19603 17973 19701
rect 18063 19734 18109 19746
rect 17256 19602 17731 19603
rect 17256 19539 17544 19602
rect 18063 19558 18069 19734
rect 18103 19558 18109 19734
rect 18063 19546 18109 19558
rect 18181 19734 18227 19746
rect 18181 19558 18187 19734
rect 18221 19558 18227 19734
rect 18181 19546 18227 19558
rect 18299 19734 18345 19746
rect 18299 19558 18305 19734
rect 18339 19558 18345 19734
rect 18299 19546 18345 19558
rect 18417 19734 18463 19746
rect 18546 19734 18552 19934
rect 18417 19558 18423 19734
rect 18457 19558 18552 19734
rect 18586 19558 18592 19934
rect 18417 19546 18463 19558
rect 18546 19546 18592 19558
rect 18664 19934 18710 19946
rect 18664 19558 18670 19934
rect 18704 19558 18710 19934
rect 18664 19546 18710 19558
rect 18782 19934 18828 19946
rect 18782 19558 18788 19934
rect 18822 19558 18828 19934
rect 18782 19546 18828 19558
rect 18900 19934 18946 19946
rect 18900 19558 18906 19934
rect 18940 19558 18946 19934
rect 18900 19546 18946 19558
rect 19018 19934 19064 19946
rect 19018 19558 19024 19934
rect 19058 19558 19064 19934
rect 19018 19546 19064 19558
rect 19136 19934 19182 19946
rect 19136 19558 19142 19934
rect 19176 19558 19182 19934
rect 19136 19546 19182 19558
rect 19254 19934 19300 19946
rect 19254 19558 19260 19934
rect 19294 19734 19300 19934
rect 19626 19746 19660 20049
rect 20085 20049 21558 20092
rect 20085 19746 20119 20049
rect 20450 19946 20484 20049
rect 20686 19946 20720 20049
rect 20922 19946 20956 20049
rect 21158 19946 21192 20049
rect 20444 19934 20490 19946
rect 19384 19734 19430 19746
rect 19294 19558 19390 19734
rect 19424 19558 19430 19734
rect 19254 19546 19300 19558
rect 19384 19546 19430 19558
rect 19502 19734 19548 19746
rect 19502 19558 19508 19734
rect 19542 19558 19548 19734
rect 19502 19546 19548 19558
rect 19620 19734 19666 19746
rect 19620 19558 19626 19734
rect 19660 19558 19666 19734
rect 19620 19546 19666 19558
rect 19738 19734 19784 19746
rect 19738 19558 19744 19734
rect 19778 19558 19784 19734
rect 19738 19546 19784 19558
rect 19961 19734 20007 19746
rect 19961 19558 19967 19734
rect 20001 19558 20007 19734
rect 19961 19546 20007 19558
rect 20079 19734 20125 19746
rect 20079 19558 20085 19734
rect 20119 19558 20125 19734
rect 20079 19546 20125 19558
rect 20197 19734 20243 19746
rect 20197 19558 20203 19734
rect 20237 19558 20243 19734
rect 20197 19546 20243 19558
rect 20315 19734 20361 19746
rect 20444 19734 20450 19934
rect 20315 19558 20321 19734
rect 20355 19558 20450 19734
rect 20484 19558 20490 19934
rect 20315 19546 20361 19558
rect 20444 19546 20490 19558
rect 20562 19934 20608 19946
rect 20562 19558 20568 19934
rect 20602 19558 20608 19934
rect 20562 19546 20608 19558
rect 20680 19934 20726 19946
rect 20680 19558 20686 19934
rect 20720 19558 20726 19934
rect 20680 19546 20726 19558
rect 20798 19934 20844 19946
rect 20798 19558 20804 19934
rect 20838 19558 20844 19934
rect 20798 19546 20844 19558
rect 20916 19934 20962 19946
rect 20916 19558 20922 19934
rect 20956 19558 20962 19934
rect 20916 19546 20962 19558
rect 21034 19934 21080 19946
rect 21034 19558 21040 19934
rect 21074 19558 21080 19934
rect 21034 19546 21080 19558
rect 21152 19934 21198 19946
rect 21152 19558 21158 19934
rect 21192 19734 21198 19934
rect 21524 19746 21558 20049
rect 21808 19962 21855 20414
rect 22162 20363 22196 20469
rect 22399 20363 22431 20469
rect 22635 20363 22667 20469
rect 22871 20363 22903 20469
rect 23107 20363 23139 20469
rect 22038 20351 22084 20363
rect 22038 20175 22044 20351
rect 22078 20175 22084 20351
rect 22038 20163 22084 20175
rect 22156 20351 22202 20363
rect 22156 20175 22162 20351
rect 22196 20175 22202 20351
rect 22156 20163 22202 20175
rect 22274 20351 22320 20363
rect 22274 20175 22280 20351
rect 22314 20175 22320 20351
rect 22274 20163 22320 20175
rect 22392 20351 22438 20363
rect 22392 20175 22398 20351
rect 22432 20175 22438 20351
rect 22392 20163 22438 20175
rect 22510 20351 22556 20363
rect 22510 20175 22516 20351
rect 22550 20175 22556 20351
rect 22510 20163 22556 20175
rect 22628 20351 22674 20363
rect 22628 20175 22634 20351
rect 22668 20175 22674 20351
rect 22628 20163 22674 20175
rect 22746 20351 22792 20363
rect 22746 20175 22752 20351
rect 22786 20175 22792 20351
rect 22746 20163 22792 20175
rect 22864 20351 22910 20363
rect 22864 20175 22870 20351
rect 22904 20175 22910 20351
rect 22864 20163 22910 20175
rect 22982 20351 23028 20363
rect 22982 20175 22988 20351
rect 23022 20175 23028 20351
rect 22982 20163 23028 20175
rect 23100 20351 23146 20363
rect 23100 20175 23106 20351
rect 23140 20175 23146 20351
rect 23100 20163 23146 20175
rect 21809 19946 21855 19962
rect 21809 19945 21890 19946
rect 22044 19945 22079 20163
rect 22323 20115 22389 20122
rect 22323 20081 22339 20115
rect 22373 20081 22389 20115
rect 22323 20070 22389 20081
rect 22515 20070 22551 20163
rect 22323 20069 22551 20070
rect 22751 20069 22787 20163
rect 22987 20069 23023 20163
rect 22323 20040 23023 20069
rect 22441 20039 23023 20040
rect 22441 19998 22507 20039
rect 22441 19964 22457 19998
rect 22491 19964 22507 19998
rect 22441 19957 22507 19964
rect 21809 19930 22079 19945
rect 21809 19926 22433 19930
rect 22869 19926 22903 20039
rect 21809 19914 22438 19926
rect 21809 19902 22398 19914
rect 21809 19900 21890 19902
rect 22156 19901 22398 19902
rect 21282 19734 21328 19746
rect 21192 19558 21288 19734
rect 21322 19558 21328 19734
rect 21152 19546 21198 19558
rect 21282 19546 21328 19558
rect 21400 19734 21446 19746
rect 21400 19558 21406 19734
rect 21440 19558 21446 19734
rect 21400 19546 21446 19558
rect 21518 19734 21564 19746
rect 21518 19558 21524 19734
rect 21558 19558 21564 19734
rect 21518 19546 21564 19558
rect 21636 19734 21682 19746
rect 21636 19558 21642 19734
rect 21676 19558 21682 19734
rect 22392 19738 22398 19901
rect 22432 19738 22438 19914
rect 22392 19726 22438 19738
rect 22510 19914 22556 19926
rect 22510 19738 22516 19914
rect 22550 19738 22556 19914
rect 22510 19726 22556 19738
rect 22627 19914 22673 19926
rect 21636 19546 21682 19558
rect 22311 19610 22419 19620
rect 22515 19610 22550 19726
rect 17256 19537 17296 19539
rect 17256 19526 17290 19537
rect 17255 19431 17290 19526
rect 17408 19433 17544 19539
rect 18069 19512 18103 19546
rect 18305 19512 18339 19546
rect 18069 19477 18339 19512
rect 18906 19512 18940 19546
rect 19142 19512 19176 19546
rect 19744 19512 19778 19546
rect 18906 19477 19176 19512
rect 19619 19477 19778 19512
rect 19967 19512 20001 19546
rect 20203 19512 20237 19546
rect 19967 19477 20237 19512
rect 20804 19512 20838 19546
rect 21040 19512 21074 19546
rect 21642 19512 21676 19546
rect 20804 19477 21074 19512
rect 21517 19477 21676 19512
rect 22419 19562 22550 19610
rect 22627 19562 22633 19914
rect 22419 19538 22633 19562
rect 22667 19538 22673 19914
rect 22419 19526 22673 19538
rect 22745 19914 22791 19926
rect 22745 19538 22751 19914
rect 22785 19538 22791 19914
rect 22745 19526 22791 19538
rect 22863 19914 22909 19926
rect 22863 19538 22869 19914
rect 22903 19538 22909 19914
rect 22863 19526 22909 19538
rect 22419 19522 22667 19526
rect 23036 19522 23046 19554
rect 22419 19478 22493 19522
rect 23031 19494 23046 19522
rect 22676 19488 22742 19494
rect 17402 19431 17544 19433
rect 17255 19422 17544 19431
rect 17256 19421 17544 19422
rect 17288 19420 17544 19421
rect 18055 19299 18122 19323
rect 18055 19265 18071 19299
rect 18105 19265 18122 19299
rect 17030 19089 17040 19168
rect 17133 19089 17143 19168
rect 15994 19040 16214 19060
rect 15994 18932 16038 19040
rect 16170 18932 16214 19040
rect 15994 18890 16214 18932
rect 15633 18860 16610 18890
rect 15633 18754 15667 18860
rect 15870 18754 15902 18860
rect 16106 18754 16138 18860
rect 16342 18754 16374 18860
rect 16578 18754 16610 18860
rect 13567 18683 13987 18688
rect 14701 18683 15017 18688
rect 13567 18672 14054 18683
rect 13567 18645 14003 18672
rect 13567 18644 13874 18645
rect 13567 18516 13601 18644
rect 13987 18638 14003 18645
rect 14037 18638 14054 18672
rect 13987 18632 14054 18638
rect 14634 18672 15017 18683
rect 14634 18638 14651 18672
rect 14685 18645 15017 18672
rect 14685 18638 14701 18645
rect 14634 18632 14701 18638
rect 13707 18604 13763 18616
rect 14820 18605 14876 18617
rect 14820 18604 14836 18605
rect 13707 18570 13713 18604
rect 13747 18589 14317 18604
rect 13747 18570 14267 18589
rect 13707 18555 14267 18570
rect 14301 18555 14317 18589
rect 13707 18554 13763 18555
rect 14250 18545 14317 18555
rect 14369 18588 14836 18604
rect 14369 18554 14385 18588
rect 14419 18571 14836 18588
rect 14870 18571 14876 18605
rect 14419 18555 14876 18571
rect 14419 18554 14435 18555
rect 14369 18547 14435 18554
rect 14983 18516 15017 18645
rect 15509 18742 15555 18754
rect 15509 18566 15515 18742
rect 15549 18566 15555 18742
rect 15509 18554 15555 18566
rect 15627 18742 15673 18754
rect 15627 18566 15633 18742
rect 15667 18566 15673 18742
rect 15627 18554 15673 18566
rect 15745 18742 15791 18754
rect 15745 18566 15751 18742
rect 15785 18566 15791 18742
rect 15745 18554 15791 18566
rect 15863 18742 15909 18754
rect 15863 18566 15869 18742
rect 15903 18566 15909 18742
rect 15863 18554 15909 18566
rect 15981 18742 16027 18754
rect 15981 18566 15987 18742
rect 16021 18566 16027 18742
rect 15981 18554 16027 18566
rect 16099 18742 16145 18754
rect 16099 18566 16105 18742
rect 16139 18566 16145 18742
rect 16099 18554 16145 18566
rect 16217 18742 16263 18754
rect 16217 18566 16223 18742
rect 16257 18566 16263 18742
rect 16217 18554 16263 18566
rect 16335 18742 16381 18754
rect 16335 18566 16341 18742
rect 16375 18566 16381 18742
rect 16335 18554 16381 18566
rect 16453 18742 16499 18754
rect 16453 18566 16459 18742
rect 16493 18566 16499 18742
rect 16453 18554 16499 18566
rect 16571 18742 16617 18754
rect 16571 18566 16577 18742
rect 16611 18566 16617 18742
rect 16571 18554 16617 18566
rect 11663 18504 11709 18516
rect 11663 18328 11669 18504
rect 11703 18328 11709 18504
rect 11663 18316 11709 18328
rect 11781 18504 11827 18516
rect 11781 18328 11787 18504
rect 11821 18328 11827 18504
rect 11781 18316 11827 18328
rect 12187 18504 12233 18516
rect 11788 18022 11821 18316
rect 12187 18128 12193 18504
rect 12227 18128 12233 18504
rect 12187 18116 12233 18128
rect 12305 18504 12351 18516
rect 12305 18128 12311 18504
rect 12345 18128 12351 18504
rect 12305 18116 12351 18128
rect 12423 18504 12469 18516
rect 12423 18128 12429 18504
rect 12463 18128 12469 18504
rect 12423 18116 12469 18128
rect 12541 18504 12587 18516
rect 12541 18128 12547 18504
rect 12581 18128 12587 18504
rect 12541 18116 12587 18128
rect 12659 18504 12705 18516
rect 12659 18128 12665 18504
rect 12699 18128 12705 18504
rect 12961 18504 13007 18516
rect 12961 18328 12967 18504
rect 13001 18328 13007 18504
rect 12961 18316 13007 18328
rect 13079 18504 13125 18516
rect 13079 18328 13085 18504
rect 13119 18328 13125 18504
rect 13079 18316 13125 18328
rect 13561 18504 13607 18516
rect 13561 18328 13567 18504
rect 13601 18328 13607 18504
rect 13561 18316 13607 18328
rect 13679 18504 13725 18516
rect 13679 18328 13685 18504
rect 13719 18328 13725 18504
rect 13679 18316 13725 18328
rect 14085 18504 14131 18516
rect 12659 18116 12705 18128
rect 12311 18022 12345 18116
rect 12968 18022 13002 18316
rect 11788 17990 13002 18022
rect 13686 18022 13719 18316
rect 14085 18128 14091 18504
rect 14125 18128 14131 18504
rect 14085 18116 14131 18128
rect 14203 18504 14249 18516
rect 14203 18128 14209 18504
rect 14243 18128 14249 18504
rect 14203 18116 14249 18128
rect 14321 18504 14367 18516
rect 14321 18128 14327 18504
rect 14361 18128 14367 18504
rect 14321 18116 14367 18128
rect 14439 18504 14485 18516
rect 14439 18128 14445 18504
rect 14479 18128 14485 18504
rect 14439 18116 14485 18128
rect 14557 18504 14603 18516
rect 14557 18128 14563 18504
rect 14597 18128 14603 18504
rect 14859 18504 14905 18516
rect 14859 18328 14865 18504
rect 14899 18328 14905 18504
rect 14859 18316 14905 18328
rect 14977 18504 15023 18516
rect 14977 18328 14983 18504
rect 15017 18328 15023 18504
rect 14977 18316 15023 18328
rect 15515 18321 15550 18554
rect 15794 18506 15860 18513
rect 15794 18472 15810 18506
rect 15844 18472 15860 18506
rect 15794 18461 15860 18472
rect 15986 18461 16022 18554
rect 15794 18460 16022 18461
rect 16222 18460 16258 18554
rect 16458 18460 16494 18554
rect 15794 18431 16494 18460
rect 15912 18430 16494 18431
rect 15912 18389 15978 18430
rect 15912 18355 15928 18389
rect 15962 18355 15978 18389
rect 15912 18348 15978 18355
rect 15515 18317 15904 18321
rect 16340 18317 16374 18430
rect 14557 18116 14603 18128
rect 14209 18022 14243 18116
rect 14866 18022 14900 18316
rect 15515 18305 15909 18317
rect 15515 18292 15869 18305
rect 15515 18289 15593 18292
rect 15510 18237 15520 18289
rect 15583 18237 15593 18289
rect 15515 18231 15588 18237
rect 15863 18129 15869 18292
rect 15903 18129 15909 18305
rect 15863 18117 15909 18129
rect 15981 18305 16027 18317
rect 15981 18129 15987 18305
rect 16021 18129 16027 18305
rect 15981 18117 16027 18129
rect 16098 18305 16144 18317
rect 13686 17990 14900 18022
rect 15782 18001 15890 18011
rect 15986 18001 16021 18117
rect 12377 17905 12509 17990
rect 14275 17905 14407 17990
rect 11522 17598 11588 17877
rect 12367 17797 12377 17905
rect 12509 17797 12519 17905
rect 14265 17797 14275 17905
rect 14407 17797 14417 17905
rect 15890 17953 16021 18001
rect 16098 17953 16104 18305
rect 15890 17929 16104 17953
rect 16138 17929 16144 18305
rect 15890 17917 16144 17929
rect 16216 18305 16262 18317
rect 16216 17929 16222 18305
rect 16256 17929 16262 18305
rect 16216 17917 16262 17929
rect 16334 18305 16380 18317
rect 16334 17929 16340 18305
rect 16374 17929 16380 18305
rect 16334 17917 16380 17929
rect 15890 17913 16138 17917
rect 17039 17915 17132 19089
rect 16547 17913 17132 17915
rect 15890 17869 15964 17913
rect 16502 17885 17132 17913
rect 16147 17879 16213 17885
rect 15782 17859 15890 17869
rect 16147 17845 16163 17879
rect 16197 17845 16213 17879
rect 16147 17749 16213 17845
rect 16265 17879 17132 17885
rect 16265 17845 16281 17879
rect 16315 17845 17132 17879
rect 16265 17829 17132 17845
rect 16502 17813 17132 17829
rect 16547 17809 17132 17813
rect 17031 17808 17132 17809
rect 17838 18836 17994 18842
rect 17838 18738 17850 18836
rect 17982 18793 17994 18836
rect 17982 18738 17995 18793
rect 16502 17760 16602 17771
rect 16502 17749 16516 17760
rect 16147 17701 16516 17749
rect 16148 17598 16214 17701
rect 16502 17671 16516 17701
rect 16506 17654 16516 17671
rect 16628 17654 16638 17760
rect 11522 17518 16216 17598
rect 17838 16953 17995 18738
rect 18055 17882 18122 19265
rect 18203 18694 18237 19477
rect 18906 19415 18940 19477
rect 18609 19377 19351 19415
rect 18609 19253 18643 19377
rect 18845 19253 18879 19377
rect 19081 19253 19115 19377
rect 19317 19253 19351 19377
rect 18603 19241 18649 19253
rect 18603 18865 18609 19241
rect 18643 18865 18649 19241
rect 18603 18853 18649 18865
rect 18721 19241 18767 19253
rect 18721 18865 18727 19241
rect 18761 18865 18767 19241
rect 18721 18853 18767 18865
rect 18839 19241 18885 19253
rect 18839 18865 18845 19241
rect 18879 18865 18885 19241
rect 18839 18853 18885 18865
rect 18957 19241 19003 19253
rect 18957 18865 18963 19241
rect 18997 18865 19003 19241
rect 18957 18853 19003 18865
rect 19075 19241 19121 19253
rect 19075 18865 19081 19241
rect 19115 18865 19121 19241
rect 19075 18853 19121 18865
rect 19193 19241 19239 19253
rect 19193 18865 19199 19241
rect 19233 18865 19239 19241
rect 19193 18853 19239 18865
rect 19311 19241 19357 19253
rect 19311 18865 19317 19241
rect 19351 18865 19357 19241
rect 19311 18853 19357 18865
rect 18203 18693 18510 18694
rect 18556 18693 18625 18694
rect 19619 18693 19653 19477
rect 18203 18689 18625 18693
rect 18203 18678 18692 18689
rect 19337 18688 19653 18693
rect 18203 18650 18641 18678
rect 18203 18649 18510 18650
rect 18203 18521 18237 18649
rect 18625 18644 18641 18650
rect 18675 18644 18692 18678
rect 18625 18638 18692 18644
rect 19270 18677 19653 18688
rect 19270 18643 19287 18677
rect 19321 18650 19653 18677
rect 19321 18643 19337 18650
rect 19270 18637 19337 18643
rect 18343 18609 18399 18621
rect 19456 18610 19512 18622
rect 19456 18609 19472 18610
rect 18343 18575 18349 18609
rect 18383 18594 18953 18609
rect 18383 18575 18903 18594
rect 18343 18560 18903 18575
rect 18937 18560 18953 18594
rect 18343 18559 18399 18560
rect 18886 18550 18953 18560
rect 19005 18593 19472 18609
rect 19005 18559 19021 18593
rect 19055 18576 19472 18593
rect 19506 18576 19512 18610
rect 19055 18560 19512 18576
rect 19055 18559 19071 18560
rect 19005 18552 19071 18559
rect 19619 18521 19653 18650
rect 20101 18694 20135 19477
rect 20804 19415 20838 19477
rect 20507 19377 21249 19415
rect 20168 19270 20178 19336
rect 20241 19270 20251 19336
rect 20507 19253 20541 19377
rect 20743 19253 20777 19377
rect 20979 19253 21013 19377
rect 21215 19253 21249 19377
rect 20501 19241 20547 19253
rect 20501 18865 20507 19241
rect 20541 18865 20547 19241
rect 20501 18853 20547 18865
rect 20619 19241 20665 19253
rect 20619 18865 20625 19241
rect 20659 18865 20665 19241
rect 20619 18853 20665 18865
rect 20737 19241 20783 19253
rect 20737 18865 20743 19241
rect 20777 18865 20783 19241
rect 20737 18853 20783 18865
rect 20855 19241 20901 19253
rect 20855 18865 20861 19241
rect 20895 18865 20901 19241
rect 20855 18853 20901 18865
rect 20973 19241 21019 19253
rect 20973 18865 20979 19241
rect 21013 18865 21019 19241
rect 20973 18853 21019 18865
rect 21091 19241 21137 19253
rect 21091 18865 21097 19241
rect 21131 18865 21137 19241
rect 21091 18853 21137 18865
rect 21209 19241 21255 19253
rect 21209 18865 21215 19241
rect 21249 18865 21255 19241
rect 21209 18853 21255 18865
rect 20101 18693 20408 18694
rect 21517 18693 21551 19477
rect 22311 19468 22419 19478
rect 22676 19454 22692 19488
rect 22726 19454 22742 19488
rect 22676 19358 22742 19454
rect 22794 19488 23046 19494
rect 22794 19454 22810 19488
rect 22844 19454 23046 19488
rect 22794 19438 23046 19454
rect 23031 19436 23046 19438
rect 23164 19436 23174 19554
rect 23031 19422 23131 19436
rect 23031 19379 23131 19380
rect 23405 19379 23510 20556
rect 23031 19358 23510 19379
rect 22676 19310 23510 19358
rect 23031 19281 23510 19310
rect 23031 19280 23131 19281
rect 23405 19279 23510 19281
rect 23573 19173 23666 21067
rect 23806 21066 24095 21067
rect 23789 20656 23966 20703
rect 23789 20643 23829 20656
rect 23787 20550 23829 20643
rect 23941 20550 23966 20656
rect 23787 20539 23966 20550
rect 23789 20538 23966 20539
rect 24388 19706 24489 21447
rect 25383 21309 25417 21455
rect 25567 21440 25664 21455
rect 26137 21452 26172 21544
rect 25607 21373 25664 21440
rect 25945 21416 26172 21452
rect 25945 21382 26011 21416
rect 25501 21337 25770 21373
rect 25945 21348 25961 21382
rect 25995 21348 26011 21382
rect 25945 21342 26011 21348
rect 25501 21309 25534 21337
rect 25737 21309 25770 21337
rect 26137 21309 26172 21416
rect 25377 21297 25423 21309
rect 25377 21121 25383 21297
rect 25417 21121 25423 21297
rect 25377 21109 25423 21121
rect 25495 21297 25541 21309
rect 25495 21121 25501 21297
rect 25535 21121 25541 21297
rect 25495 21109 25541 21121
rect 25613 21297 25659 21309
rect 25613 21121 25619 21297
rect 25653 21121 25659 21297
rect 25613 21109 25659 21121
rect 25731 21297 25777 21309
rect 25731 21121 25737 21297
rect 25771 21242 25777 21297
rect 25896 21297 25942 21309
rect 25896 21242 25902 21297
rect 25771 21154 25902 21242
rect 25771 21121 25777 21154
rect 25731 21109 25777 21121
rect 25896 21121 25902 21154
rect 25936 21121 25942 21297
rect 25896 21109 25942 21121
rect 26014 21297 26060 21309
rect 26014 21121 26020 21297
rect 26054 21121 26060 21297
rect 26014 21109 26060 21121
rect 26132 21297 26178 21309
rect 26132 21121 26138 21297
rect 26172 21121 26178 21297
rect 26132 21109 26178 21121
rect 26250 21297 26296 21309
rect 26250 21121 26256 21297
rect 26290 21121 26296 21297
rect 26250 21109 26296 21121
rect 25384 21071 25417 21109
rect 25620 21071 25653 21109
rect 25384 21035 25653 21071
rect 26020 21070 26054 21109
rect 26256 21070 26290 21109
rect 26020 21034 26290 21070
rect 26124 21033 26290 21034
rect 26124 20954 26256 21033
rect 26114 20846 26124 20954
rect 26256 20846 26266 20954
rect 26396 20517 26458 22088
rect 26594 22076 26640 22088
rect 26594 21700 26600 22076
rect 26634 21700 26640 22076
rect 26594 21688 26640 21700
rect 26712 22076 26758 22088
rect 26712 21700 26718 22076
rect 26752 21700 26758 22076
rect 26712 21688 26758 21700
rect 26830 22076 26876 22088
rect 26830 21700 26836 22076
rect 26870 21700 26876 22076
rect 26830 21688 26876 21700
rect 26948 22076 26994 22088
rect 26948 21700 26954 22076
rect 26988 21700 26994 22076
rect 26948 21688 26994 21700
rect 27066 22076 27112 22088
rect 27066 21700 27072 22076
rect 27106 21700 27112 22076
rect 27066 21688 27112 21700
rect 27184 22076 27230 22088
rect 27184 21700 27190 22076
rect 27224 21700 27230 22076
rect 27184 21688 27230 21700
rect 27302 22076 27348 22088
rect 27397 22084 27407 22150
rect 27473 22084 27483 22150
rect 27302 21700 27308 22076
rect 27342 21700 27348 22076
rect 27302 21688 27348 21700
rect 26600 21505 26634 21688
rect 26718 21647 26752 21688
rect 26954 21647 26988 21688
rect 26718 21618 26988 21647
rect 27072 21646 27106 21688
rect 27308 21646 27342 21688
rect 27072 21618 27342 21646
rect 27308 21570 27342 21618
rect 27279 21540 27342 21570
rect 28332 21611 28399 22201
rect 29050 22194 29094 22302
rect 29226 22194 29270 22302
rect 29050 22152 29270 22194
rect 28689 22122 29666 22152
rect 28689 22016 28723 22122
rect 28926 22016 28958 22122
rect 29162 22016 29194 22122
rect 29398 22016 29430 22122
rect 29634 22016 29666 22122
rect 28565 22004 28611 22016
rect 28565 21828 28571 22004
rect 28605 21828 28611 22004
rect 28565 21816 28611 21828
rect 28683 22004 28729 22016
rect 28683 21828 28689 22004
rect 28723 21828 28729 22004
rect 28683 21816 28729 21828
rect 28801 22004 28847 22016
rect 28801 21828 28807 22004
rect 28841 21828 28847 22004
rect 28801 21816 28847 21828
rect 28919 22004 28965 22016
rect 28919 21828 28925 22004
rect 28959 21828 28965 22004
rect 28919 21816 28965 21828
rect 29037 22004 29083 22016
rect 29037 21828 29043 22004
rect 29077 21828 29083 22004
rect 29037 21816 29083 21828
rect 29155 22004 29201 22016
rect 29155 21828 29161 22004
rect 29195 21828 29201 22004
rect 29155 21816 29201 21828
rect 29273 22004 29319 22016
rect 29273 21828 29279 22004
rect 29313 21828 29319 22004
rect 29273 21816 29319 21828
rect 29391 22004 29437 22016
rect 29391 21828 29397 22004
rect 29431 21828 29437 22004
rect 29391 21816 29437 21828
rect 29509 22004 29555 22016
rect 29509 21828 29515 22004
rect 29549 21828 29555 22004
rect 29509 21816 29555 21828
rect 29627 22004 29673 22016
rect 29627 21828 29633 22004
rect 29667 21828 29673 22004
rect 29627 21816 29673 21828
rect 28571 21611 28606 21816
rect 28850 21768 28916 21775
rect 28850 21734 28866 21768
rect 28900 21734 28916 21768
rect 28850 21723 28916 21734
rect 29042 21723 29078 21816
rect 28850 21722 29078 21723
rect 29278 21722 29314 21816
rect 29514 21722 29550 21816
rect 28850 21693 29550 21722
rect 28332 21583 28606 21611
rect 28968 21692 29550 21693
rect 28968 21651 29034 21692
rect 28968 21617 28984 21651
rect 29018 21617 29034 21651
rect 28968 21610 29034 21617
rect 28332 21579 28960 21583
rect 29396 21579 29430 21692
rect 28332 21567 28965 21579
rect 28332 21554 28925 21567
rect 26525 21451 26634 21505
rect 26525 21305 26559 21451
rect 26698 21437 26708 21534
rect 26807 21437 26817 21534
rect 27279 21448 27314 21540
rect 26709 21436 26806 21437
rect 26749 21369 26806 21436
rect 27087 21412 27314 21448
rect 27087 21378 27153 21412
rect 26643 21333 26912 21369
rect 27087 21344 27103 21378
rect 27137 21344 27153 21378
rect 27087 21338 27153 21344
rect 26643 21305 26676 21333
rect 26879 21305 26912 21333
rect 27279 21305 27314 21412
rect 28919 21391 28925 21554
rect 28959 21391 28965 21567
rect 28919 21379 28965 21391
rect 29037 21567 29083 21579
rect 29037 21391 29043 21567
rect 29077 21391 29083 21567
rect 29037 21379 29083 21391
rect 29154 21567 29200 21579
rect 26519 21293 26565 21305
rect 26519 21117 26525 21293
rect 26559 21117 26565 21293
rect 26519 21105 26565 21117
rect 26637 21293 26683 21305
rect 26637 21117 26643 21293
rect 26677 21117 26683 21293
rect 26637 21105 26683 21117
rect 26755 21293 26801 21305
rect 26755 21117 26761 21293
rect 26795 21117 26801 21293
rect 26755 21105 26801 21117
rect 26873 21293 26919 21305
rect 26873 21117 26879 21293
rect 26913 21238 26919 21293
rect 27038 21293 27084 21305
rect 27038 21238 27044 21293
rect 26913 21150 27044 21238
rect 26913 21117 26919 21150
rect 26873 21105 26919 21117
rect 27038 21117 27044 21150
rect 27078 21117 27084 21293
rect 27038 21105 27084 21117
rect 27156 21293 27202 21305
rect 27156 21117 27162 21293
rect 27196 21117 27202 21293
rect 27156 21105 27202 21117
rect 27274 21293 27320 21305
rect 27274 21117 27280 21293
rect 27314 21117 27320 21293
rect 27274 21105 27320 21117
rect 27392 21293 27438 21305
rect 27392 21117 27398 21293
rect 27432 21117 27438 21293
rect 28838 21263 28946 21273
rect 29042 21263 29077 21379
rect 28946 21215 29077 21263
rect 29154 21215 29160 21567
rect 28946 21191 29160 21215
rect 29194 21191 29200 21567
rect 28946 21179 29200 21191
rect 29272 21567 29318 21579
rect 29272 21191 29278 21567
rect 29312 21191 29318 21567
rect 29272 21179 29318 21191
rect 29390 21567 29436 21579
rect 29390 21191 29396 21567
rect 29430 21191 29436 21567
rect 29390 21179 29436 21191
rect 30319 21216 30608 21237
rect 28946 21175 29194 21179
rect 28946 21131 29020 21175
rect 30319 21174 30360 21216
rect 29558 21147 30360 21174
rect 29203 21141 29269 21147
rect 28838 21121 28946 21131
rect 27392 21105 27438 21117
rect 29203 21107 29219 21141
rect 29253 21107 29269 21141
rect 26526 21067 26559 21105
rect 26762 21067 26795 21105
rect 26526 21031 26795 21067
rect 27162 21066 27196 21105
rect 27398 21066 27432 21105
rect 27162 21031 27432 21066
rect 27162 21030 27398 21031
rect 27266 20956 27398 21030
rect 29203 21011 29269 21107
rect 29321 21141 30360 21147
rect 29321 21107 29337 21141
rect 29371 21107 30360 21141
rect 29321 21091 30360 21107
rect 29558 21085 30360 21091
rect 30592 21085 30608 21216
rect 29558 21075 30608 21085
rect 29621 21074 30608 21075
rect 30086 21070 30608 21074
rect 29557 21011 30023 21033
rect 29203 20963 30023 21011
rect 27256 20848 27266 20956
rect 27398 20848 27408 20956
rect 29557 20932 30023 20963
rect 29918 20676 30023 20932
rect 26395 20500 26458 20517
rect 29036 20652 29256 20672
rect 29036 20544 29080 20652
rect 29212 20544 29256 20652
rect 29838 20570 29848 20676
rect 29960 20570 30023 20676
rect 29874 20559 30023 20570
rect 29036 20502 29256 20544
rect 26395 20496 26533 20500
rect 26395 20462 28365 20496
rect 28675 20472 29652 20502
rect 26395 20433 28367 20462
rect 26395 20431 26533 20433
rect 28321 20417 28367 20433
rect 25359 20201 25369 20309
rect 25501 20201 25511 20309
rect 27257 20201 27267 20309
rect 27399 20201 27409 20309
rect 25369 20161 25501 20201
rect 27267 20161 27399 20201
rect 25369 20095 25502 20161
rect 27267 20095 27400 20161
rect 24700 20052 26173 20095
rect 24700 19749 24734 20052
rect 25065 19949 25099 20052
rect 25301 19949 25335 20052
rect 25537 19949 25571 20052
rect 25773 19949 25807 20052
rect 25059 19937 25105 19949
rect 23790 19604 24489 19706
rect 24576 19737 24622 19749
rect 23790 19544 24078 19604
rect 24576 19561 24582 19737
rect 24616 19561 24622 19737
rect 24576 19549 24622 19561
rect 24694 19737 24740 19749
rect 24694 19561 24700 19737
rect 24734 19561 24740 19737
rect 24694 19549 24740 19561
rect 24812 19737 24858 19749
rect 24812 19561 24818 19737
rect 24852 19561 24858 19737
rect 24812 19549 24858 19561
rect 24930 19737 24976 19749
rect 25059 19737 25065 19937
rect 24930 19561 24936 19737
rect 24970 19561 25065 19737
rect 25099 19561 25105 19937
rect 24930 19549 24976 19561
rect 25059 19549 25105 19561
rect 25177 19937 25223 19949
rect 25177 19561 25183 19937
rect 25217 19561 25223 19937
rect 25177 19549 25223 19561
rect 25295 19937 25341 19949
rect 25295 19561 25301 19937
rect 25335 19561 25341 19937
rect 25295 19549 25341 19561
rect 25413 19937 25459 19949
rect 25413 19561 25419 19937
rect 25453 19561 25459 19937
rect 25413 19549 25459 19561
rect 25531 19937 25577 19949
rect 25531 19561 25537 19937
rect 25571 19561 25577 19937
rect 25531 19549 25577 19561
rect 25649 19937 25695 19949
rect 25649 19561 25655 19937
rect 25689 19561 25695 19937
rect 25649 19549 25695 19561
rect 25767 19937 25813 19949
rect 25767 19561 25773 19937
rect 25807 19737 25813 19937
rect 26139 19749 26173 20052
rect 26598 20052 28071 20095
rect 26598 19749 26632 20052
rect 26963 19949 26997 20052
rect 27199 19949 27233 20052
rect 27435 19949 27469 20052
rect 27671 19949 27705 20052
rect 26957 19937 27003 19949
rect 25897 19737 25943 19749
rect 25807 19561 25903 19737
rect 25937 19561 25943 19737
rect 25767 19549 25813 19561
rect 25897 19549 25943 19561
rect 26015 19737 26061 19749
rect 26015 19561 26021 19737
rect 26055 19561 26061 19737
rect 26015 19549 26061 19561
rect 26133 19737 26179 19749
rect 26133 19561 26139 19737
rect 26173 19561 26179 19737
rect 26133 19549 26179 19561
rect 26251 19737 26297 19749
rect 26251 19561 26257 19737
rect 26291 19561 26297 19737
rect 26251 19549 26297 19561
rect 26474 19737 26520 19749
rect 26474 19561 26480 19737
rect 26514 19561 26520 19737
rect 26474 19549 26520 19561
rect 26592 19737 26638 19749
rect 26592 19561 26598 19737
rect 26632 19561 26638 19737
rect 26592 19549 26638 19561
rect 26710 19737 26756 19749
rect 26710 19561 26716 19737
rect 26750 19561 26756 19737
rect 26710 19549 26756 19561
rect 26828 19737 26874 19749
rect 26957 19737 26963 19937
rect 26828 19561 26834 19737
rect 26868 19561 26963 19737
rect 26997 19561 27003 19937
rect 26828 19549 26874 19561
rect 26957 19549 27003 19561
rect 27075 19937 27121 19949
rect 27075 19561 27081 19937
rect 27115 19561 27121 19937
rect 27075 19549 27121 19561
rect 27193 19937 27239 19949
rect 27193 19561 27199 19937
rect 27233 19561 27239 19937
rect 27193 19549 27239 19561
rect 27311 19937 27357 19949
rect 27311 19561 27317 19937
rect 27351 19561 27357 19937
rect 27311 19549 27357 19561
rect 27429 19937 27475 19949
rect 27429 19561 27435 19937
rect 27469 19561 27475 19937
rect 27429 19549 27475 19561
rect 27547 19937 27593 19949
rect 27547 19561 27553 19937
rect 27587 19561 27593 19937
rect 27547 19549 27593 19561
rect 27665 19937 27711 19949
rect 27665 19561 27671 19937
rect 27705 19737 27711 19937
rect 28037 19749 28071 20052
rect 28321 19965 28368 20417
rect 28675 20366 28709 20472
rect 28912 20366 28944 20472
rect 29148 20366 29180 20472
rect 29384 20366 29416 20472
rect 29620 20366 29652 20472
rect 28551 20354 28597 20366
rect 28551 20178 28557 20354
rect 28591 20178 28597 20354
rect 28551 20166 28597 20178
rect 28669 20354 28715 20366
rect 28669 20178 28675 20354
rect 28709 20178 28715 20354
rect 28669 20166 28715 20178
rect 28787 20354 28833 20366
rect 28787 20178 28793 20354
rect 28827 20178 28833 20354
rect 28787 20166 28833 20178
rect 28905 20354 28951 20366
rect 28905 20178 28911 20354
rect 28945 20178 28951 20354
rect 28905 20166 28951 20178
rect 29023 20354 29069 20366
rect 29023 20178 29029 20354
rect 29063 20178 29069 20354
rect 29023 20166 29069 20178
rect 29141 20354 29187 20366
rect 29141 20178 29147 20354
rect 29181 20178 29187 20354
rect 29141 20166 29187 20178
rect 29259 20354 29305 20366
rect 29259 20178 29265 20354
rect 29299 20178 29305 20354
rect 29259 20166 29305 20178
rect 29377 20354 29423 20366
rect 29377 20178 29383 20354
rect 29417 20178 29423 20354
rect 29377 20166 29423 20178
rect 29495 20354 29541 20366
rect 29495 20178 29501 20354
rect 29535 20178 29541 20354
rect 29495 20166 29541 20178
rect 29613 20354 29659 20366
rect 29613 20178 29619 20354
rect 29653 20178 29659 20354
rect 29613 20166 29659 20178
rect 28322 19949 28368 19965
rect 28322 19948 28403 19949
rect 28557 19948 28592 20166
rect 28836 20118 28902 20125
rect 28836 20084 28852 20118
rect 28886 20084 28902 20118
rect 28836 20073 28902 20084
rect 29028 20073 29064 20166
rect 28836 20072 29064 20073
rect 29264 20072 29300 20166
rect 29500 20072 29536 20166
rect 28836 20043 29536 20072
rect 28954 20042 29536 20043
rect 28954 20001 29020 20042
rect 28954 19967 28970 20001
rect 29004 19967 29020 20001
rect 28954 19960 29020 19967
rect 28322 19933 28592 19948
rect 28322 19929 28946 19933
rect 29382 19929 29416 20042
rect 28322 19917 28951 19929
rect 28322 19905 28911 19917
rect 28322 19903 28403 19905
rect 28669 19904 28911 19905
rect 27795 19737 27841 19749
rect 27705 19561 27801 19737
rect 27835 19561 27841 19737
rect 27665 19549 27711 19561
rect 27795 19549 27841 19561
rect 27913 19737 27959 19749
rect 27913 19561 27919 19737
rect 27953 19561 27959 19737
rect 27913 19549 27959 19561
rect 28031 19737 28077 19749
rect 28031 19561 28037 19737
rect 28071 19561 28077 19737
rect 28031 19549 28077 19561
rect 28149 19737 28195 19749
rect 28149 19561 28155 19737
rect 28189 19561 28195 19737
rect 28905 19741 28911 19904
rect 28945 19741 28951 19917
rect 28905 19729 28951 19741
rect 29023 19917 29069 19929
rect 29023 19741 29029 19917
rect 29063 19741 29069 19917
rect 29023 19729 29069 19741
rect 29140 19917 29186 19929
rect 28149 19549 28195 19561
rect 28824 19613 28932 19623
rect 29028 19613 29063 19729
rect 23790 19542 23830 19544
rect 23790 19531 23824 19542
rect 23789 19436 23824 19531
rect 23942 19438 24078 19544
rect 24582 19515 24616 19549
rect 24818 19515 24852 19549
rect 24582 19480 24852 19515
rect 25419 19515 25453 19549
rect 25655 19515 25689 19549
rect 26257 19515 26291 19549
rect 25419 19480 25689 19515
rect 26132 19480 26291 19515
rect 26480 19515 26514 19549
rect 26716 19515 26750 19549
rect 26480 19480 26750 19515
rect 27317 19515 27351 19549
rect 27553 19515 27587 19549
rect 28155 19515 28189 19549
rect 27317 19480 27587 19515
rect 28030 19480 28189 19515
rect 28932 19565 29063 19613
rect 29140 19565 29146 19917
rect 28932 19541 29146 19565
rect 29180 19541 29186 19917
rect 28932 19529 29186 19541
rect 29258 19917 29304 19929
rect 29258 19541 29264 19917
rect 29298 19541 29304 19917
rect 29258 19529 29304 19541
rect 29376 19917 29422 19929
rect 29376 19541 29382 19917
rect 29416 19541 29422 19917
rect 29376 19529 29422 19541
rect 28932 19525 29180 19529
rect 29549 19525 29559 19557
rect 28932 19481 29006 19525
rect 29544 19497 29559 19525
rect 29189 19491 29255 19497
rect 23936 19436 24078 19438
rect 23789 19427 24078 19436
rect 23790 19426 24078 19427
rect 23822 19425 24078 19426
rect 24568 19302 24635 19326
rect 24568 19268 24584 19302
rect 24618 19268 24635 19302
rect 23564 19094 23574 19173
rect 23667 19094 23677 19173
rect 22528 19045 22748 19065
rect 22528 18937 22572 19045
rect 22704 18937 22748 19045
rect 22528 18895 22748 18937
rect 22167 18865 23144 18895
rect 22167 18759 22201 18865
rect 22404 18759 22436 18865
rect 22640 18759 22672 18865
rect 22876 18759 22908 18865
rect 23112 18759 23144 18865
rect 20101 18688 20521 18693
rect 21235 18688 21551 18693
rect 20101 18677 20588 18688
rect 20101 18650 20537 18677
rect 20101 18649 20408 18650
rect 20101 18521 20135 18649
rect 20521 18643 20537 18650
rect 20571 18643 20588 18677
rect 20521 18637 20588 18643
rect 21168 18677 21551 18688
rect 21168 18643 21185 18677
rect 21219 18650 21551 18677
rect 21219 18643 21235 18650
rect 21168 18637 21235 18643
rect 20241 18609 20297 18621
rect 21354 18610 21410 18622
rect 21354 18609 21370 18610
rect 20241 18575 20247 18609
rect 20281 18594 20851 18609
rect 20281 18575 20801 18594
rect 20241 18560 20801 18575
rect 20835 18560 20851 18594
rect 20241 18559 20297 18560
rect 20784 18550 20851 18560
rect 20903 18593 21370 18609
rect 20903 18559 20919 18593
rect 20953 18576 21370 18593
rect 21404 18576 21410 18610
rect 20953 18560 21410 18576
rect 20953 18559 20969 18560
rect 20903 18552 20969 18559
rect 21517 18521 21551 18650
rect 22043 18747 22089 18759
rect 22043 18571 22049 18747
rect 22083 18571 22089 18747
rect 22043 18559 22089 18571
rect 22161 18747 22207 18759
rect 22161 18571 22167 18747
rect 22201 18571 22207 18747
rect 22161 18559 22207 18571
rect 22279 18747 22325 18759
rect 22279 18571 22285 18747
rect 22319 18571 22325 18747
rect 22279 18559 22325 18571
rect 22397 18747 22443 18759
rect 22397 18571 22403 18747
rect 22437 18571 22443 18747
rect 22397 18559 22443 18571
rect 22515 18747 22561 18759
rect 22515 18571 22521 18747
rect 22555 18571 22561 18747
rect 22515 18559 22561 18571
rect 22633 18747 22679 18759
rect 22633 18571 22639 18747
rect 22673 18571 22679 18747
rect 22633 18559 22679 18571
rect 22751 18747 22797 18759
rect 22751 18571 22757 18747
rect 22791 18571 22797 18747
rect 22751 18559 22797 18571
rect 22869 18747 22915 18759
rect 22869 18571 22875 18747
rect 22909 18571 22915 18747
rect 22869 18559 22915 18571
rect 22987 18747 23033 18759
rect 22987 18571 22993 18747
rect 23027 18571 23033 18747
rect 22987 18559 23033 18571
rect 23105 18747 23151 18759
rect 23105 18571 23111 18747
rect 23145 18571 23151 18747
rect 23105 18559 23151 18571
rect 18197 18509 18243 18521
rect 18197 18333 18203 18509
rect 18237 18333 18243 18509
rect 18197 18321 18243 18333
rect 18315 18509 18361 18521
rect 18315 18333 18321 18509
rect 18355 18333 18361 18509
rect 18315 18321 18361 18333
rect 18721 18509 18767 18521
rect 18322 18027 18355 18321
rect 18721 18133 18727 18509
rect 18761 18133 18767 18509
rect 18721 18121 18767 18133
rect 18839 18509 18885 18521
rect 18839 18133 18845 18509
rect 18879 18133 18885 18509
rect 18839 18121 18885 18133
rect 18957 18509 19003 18521
rect 18957 18133 18963 18509
rect 18997 18133 19003 18509
rect 18957 18121 19003 18133
rect 19075 18509 19121 18521
rect 19075 18133 19081 18509
rect 19115 18133 19121 18509
rect 19075 18121 19121 18133
rect 19193 18509 19239 18521
rect 19193 18133 19199 18509
rect 19233 18133 19239 18509
rect 19495 18509 19541 18521
rect 19495 18333 19501 18509
rect 19535 18333 19541 18509
rect 19495 18321 19541 18333
rect 19613 18509 19659 18521
rect 19613 18333 19619 18509
rect 19653 18333 19659 18509
rect 19613 18321 19659 18333
rect 20095 18509 20141 18521
rect 20095 18333 20101 18509
rect 20135 18333 20141 18509
rect 20095 18321 20141 18333
rect 20213 18509 20259 18521
rect 20213 18333 20219 18509
rect 20253 18333 20259 18509
rect 20213 18321 20259 18333
rect 20619 18509 20665 18521
rect 19193 18121 19239 18133
rect 18845 18027 18879 18121
rect 19502 18027 19536 18321
rect 18322 17995 19536 18027
rect 20220 18027 20253 18321
rect 20619 18133 20625 18509
rect 20659 18133 20665 18509
rect 20619 18121 20665 18133
rect 20737 18509 20783 18521
rect 20737 18133 20743 18509
rect 20777 18133 20783 18509
rect 20737 18121 20783 18133
rect 20855 18509 20901 18521
rect 20855 18133 20861 18509
rect 20895 18133 20901 18509
rect 20855 18121 20901 18133
rect 20973 18509 21019 18521
rect 20973 18133 20979 18509
rect 21013 18133 21019 18509
rect 20973 18121 21019 18133
rect 21091 18509 21137 18521
rect 21091 18133 21097 18509
rect 21131 18133 21137 18509
rect 21393 18509 21439 18521
rect 21393 18333 21399 18509
rect 21433 18333 21439 18509
rect 21393 18321 21439 18333
rect 21511 18509 21557 18521
rect 21511 18333 21517 18509
rect 21551 18333 21557 18509
rect 21511 18321 21557 18333
rect 22049 18326 22084 18559
rect 22328 18511 22394 18518
rect 22328 18477 22344 18511
rect 22378 18477 22394 18511
rect 22328 18466 22394 18477
rect 22520 18466 22556 18559
rect 22328 18465 22556 18466
rect 22756 18465 22792 18559
rect 22992 18465 23028 18559
rect 22328 18436 23028 18465
rect 22446 18435 23028 18436
rect 22446 18394 22512 18435
rect 22446 18360 22462 18394
rect 22496 18360 22512 18394
rect 22446 18353 22512 18360
rect 22049 18322 22438 18326
rect 22874 18322 22908 18435
rect 21091 18121 21137 18133
rect 20743 18027 20777 18121
rect 21400 18027 21434 18321
rect 22049 18310 22443 18322
rect 22049 18297 22403 18310
rect 22049 18294 22127 18297
rect 22044 18242 22054 18294
rect 22117 18242 22127 18294
rect 22049 18236 22122 18242
rect 22397 18134 22403 18297
rect 22437 18134 22443 18310
rect 22397 18122 22443 18134
rect 22515 18310 22561 18322
rect 22515 18134 22521 18310
rect 22555 18134 22561 18310
rect 22515 18122 22561 18134
rect 22632 18310 22678 18322
rect 20220 17995 21434 18027
rect 22316 18006 22424 18016
rect 22520 18006 22555 18122
rect 18911 17910 19043 17995
rect 20809 17910 20941 17995
rect 18056 17603 18122 17882
rect 18901 17802 18911 17910
rect 19043 17802 19053 17910
rect 20799 17802 20809 17910
rect 20941 17802 20951 17910
rect 22424 17958 22555 18006
rect 22632 17958 22638 18310
rect 22424 17934 22638 17958
rect 22672 17934 22678 18310
rect 22424 17922 22678 17934
rect 22750 18310 22796 18322
rect 22750 17934 22756 18310
rect 22790 17934 22796 18310
rect 22750 17922 22796 17934
rect 22868 18310 22914 18322
rect 22868 17934 22874 18310
rect 22908 17934 22914 18310
rect 22868 17922 22914 17934
rect 22424 17918 22672 17922
rect 23573 17920 23666 19094
rect 23081 17918 23666 17920
rect 22424 17874 22498 17918
rect 23036 17890 23666 17918
rect 22681 17884 22747 17890
rect 22316 17864 22424 17874
rect 22681 17850 22697 17884
rect 22731 17850 22747 17884
rect 22681 17754 22747 17850
rect 22799 17884 23666 17890
rect 22799 17850 22815 17884
rect 22849 17850 23666 17884
rect 22799 17834 23666 17850
rect 23036 17818 23666 17834
rect 23081 17814 23666 17818
rect 23565 17813 23666 17814
rect 24351 18839 24507 18845
rect 24351 18741 24363 18839
rect 24495 18741 24507 18839
rect 23036 17765 23136 17776
rect 23036 17754 23050 17765
rect 22681 17706 23050 17754
rect 22682 17603 22748 17706
rect 23036 17676 23050 17706
rect 23040 17659 23050 17676
rect 23162 17659 23172 17765
rect 18056 17523 22750 17603
rect 24351 17068 24507 18741
rect 24568 17885 24635 19268
rect 24716 18697 24750 19480
rect 25419 19418 25453 19480
rect 25122 19380 25864 19418
rect 25122 19256 25156 19380
rect 25358 19256 25392 19380
rect 25594 19256 25628 19380
rect 25830 19256 25864 19380
rect 25116 19244 25162 19256
rect 25116 18868 25122 19244
rect 25156 18868 25162 19244
rect 25116 18856 25162 18868
rect 25234 19244 25280 19256
rect 25234 18868 25240 19244
rect 25274 18868 25280 19244
rect 25234 18856 25280 18868
rect 25352 19244 25398 19256
rect 25352 18868 25358 19244
rect 25392 18868 25398 19244
rect 25352 18856 25398 18868
rect 25470 19244 25516 19256
rect 25470 18868 25476 19244
rect 25510 18868 25516 19244
rect 25470 18856 25516 18868
rect 25588 19244 25634 19256
rect 25588 18868 25594 19244
rect 25628 18868 25634 19244
rect 25588 18856 25634 18868
rect 25706 19244 25752 19256
rect 25706 18868 25712 19244
rect 25746 18868 25752 19244
rect 25706 18856 25752 18868
rect 25824 19244 25870 19256
rect 25824 18868 25830 19244
rect 25864 18868 25870 19244
rect 25824 18856 25870 18868
rect 24716 18696 25023 18697
rect 25069 18696 25138 18697
rect 26132 18696 26166 19480
rect 24716 18692 25138 18696
rect 24716 18681 25205 18692
rect 25850 18691 26166 18696
rect 24716 18653 25154 18681
rect 24716 18652 25023 18653
rect 24716 18524 24750 18652
rect 25138 18647 25154 18653
rect 25188 18647 25205 18681
rect 25138 18641 25205 18647
rect 25783 18680 26166 18691
rect 25783 18646 25800 18680
rect 25834 18653 26166 18680
rect 25834 18646 25850 18653
rect 25783 18640 25850 18646
rect 24856 18612 24912 18624
rect 25969 18613 26025 18625
rect 25969 18612 25985 18613
rect 24856 18578 24862 18612
rect 24896 18597 25466 18612
rect 24896 18578 25416 18597
rect 24856 18563 25416 18578
rect 25450 18563 25466 18597
rect 24856 18562 24912 18563
rect 25399 18553 25466 18563
rect 25518 18596 25985 18612
rect 25518 18562 25534 18596
rect 25568 18579 25985 18596
rect 26019 18579 26025 18613
rect 25568 18563 26025 18579
rect 25568 18562 25584 18563
rect 25518 18555 25584 18562
rect 26132 18524 26166 18653
rect 26614 18697 26648 19480
rect 27317 19418 27351 19480
rect 27020 19380 27762 19418
rect 26681 19273 26691 19339
rect 26754 19273 26764 19339
rect 27020 19256 27054 19380
rect 27256 19256 27290 19380
rect 27492 19256 27526 19380
rect 27728 19256 27762 19380
rect 27014 19244 27060 19256
rect 27014 18868 27020 19244
rect 27054 18868 27060 19244
rect 27014 18856 27060 18868
rect 27132 19244 27178 19256
rect 27132 18868 27138 19244
rect 27172 18868 27178 19244
rect 27132 18856 27178 18868
rect 27250 19244 27296 19256
rect 27250 18868 27256 19244
rect 27290 18868 27296 19244
rect 27250 18856 27296 18868
rect 27368 19244 27414 19256
rect 27368 18868 27374 19244
rect 27408 18868 27414 19244
rect 27368 18856 27414 18868
rect 27486 19244 27532 19256
rect 27486 18868 27492 19244
rect 27526 18868 27532 19244
rect 27486 18856 27532 18868
rect 27604 19244 27650 19256
rect 27604 18868 27610 19244
rect 27644 18868 27650 19244
rect 27604 18856 27650 18868
rect 27722 19244 27768 19256
rect 27722 18868 27728 19244
rect 27762 18868 27768 19244
rect 27722 18856 27768 18868
rect 26614 18696 26921 18697
rect 28030 18696 28064 19480
rect 28824 19471 28932 19481
rect 29189 19457 29205 19491
rect 29239 19457 29255 19491
rect 29189 19361 29255 19457
rect 29307 19491 29559 19497
rect 29307 19457 29323 19491
rect 29357 19457 29559 19491
rect 29307 19441 29559 19457
rect 29544 19439 29559 19441
rect 29677 19439 29687 19557
rect 29544 19425 29644 19439
rect 29544 19382 29644 19383
rect 29918 19382 30023 20559
rect 29544 19361 30023 19382
rect 29189 19313 30023 19361
rect 29544 19284 30023 19313
rect 29544 19283 29644 19284
rect 29918 19282 30023 19284
rect 30086 19176 30179 21070
rect 30895 19711 31022 26018
rect 34841 25402 37548 25403
rect 34841 25387 37645 25402
rect 34841 25322 34860 25387
rect 34943 25322 37645 25387
rect 34841 25309 37645 25322
rect 37561 25291 37645 25309
rect 37561 25234 37569 25291
rect 37637 25234 37645 25291
rect 37561 25232 37645 25234
rect 37729 25291 37813 25312
rect 37729 25234 37737 25291
rect 37805 25234 37813 25291
rect 37729 25232 37813 25234
rect 37569 25224 37637 25232
rect 37737 25224 37805 25232
rect 36955 25149 37155 25154
rect 36955 25148 37965 25149
rect 36955 25114 36967 25148
rect 37143 25114 37965 25148
rect 36955 25108 37155 25114
rect 36955 25030 37155 25036
rect 36955 24996 36967 25030
rect 37143 24996 37155 25030
rect 36955 24990 37155 24996
rect 36955 24912 37155 24918
rect 36955 24878 36967 24912
rect 37143 24878 37155 24912
rect 36955 24872 37155 24878
rect 36955 24794 37155 24800
rect 36955 24760 36967 24794
rect 37143 24760 37155 24794
rect 36955 24713 37155 24760
rect 36755 24707 37155 24713
rect 36611 24673 36767 24707
rect 37143 24673 37155 24707
rect 30514 19709 31022 19711
rect 30303 19555 31022 19709
rect 32144 24429 32318 24440
rect 32144 24351 32159 24429
rect 32304 24351 32318 24429
rect 30303 19547 30591 19555
rect 30303 19545 30343 19547
rect 30303 19534 30337 19545
rect 30302 19439 30337 19534
rect 30455 19441 30591 19547
rect 30449 19439 30591 19441
rect 30302 19430 30591 19439
rect 30303 19429 30591 19430
rect 30335 19428 30591 19429
rect 30077 19097 30087 19176
rect 30180 19097 30190 19176
rect 29041 19048 29261 19068
rect 29041 18940 29085 19048
rect 29217 18940 29261 19048
rect 29041 18898 29261 18940
rect 28680 18868 29657 18898
rect 28680 18762 28714 18868
rect 28917 18762 28949 18868
rect 29153 18762 29185 18868
rect 29389 18762 29421 18868
rect 29625 18762 29657 18868
rect 26614 18691 27034 18696
rect 27748 18691 28064 18696
rect 26614 18680 27101 18691
rect 26614 18653 27050 18680
rect 26614 18652 26921 18653
rect 26614 18524 26648 18652
rect 27034 18646 27050 18653
rect 27084 18646 27101 18680
rect 27034 18640 27101 18646
rect 27681 18680 28064 18691
rect 27681 18646 27698 18680
rect 27732 18653 28064 18680
rect 27732 18646 27748 18653
rect 27681 18640 27748 18646
rect 26754 18612 26810 18624
rect 27867 18613 27923 18625
rect 27867 18612 27883 18613
rect 26754 18578 26760 18612
rect 26794 18597 27364 18612
rect 26794 18578 27314 18597
rect 26754 18563 27314 18578
rect 27348 18563 27364 18597
rect 26754 18562 26810 18563
rect 27297 18553 27364 18563
rect 27416 18596 27883 18612
rect 27416 18562 27432 18596
rect 27466 18579 27883 18596
rect 27917 18579 27923 18613
rect 27466 18563 27923 18579
rect 27466 18562 27482 18563
rect 27416 18555 27482 18562
rect 28030 18524 28064 18653
rect 28556 18750 28602 18762
rect 28556 18574 28562 18750
rect 28596 18574 28602 18750
rect 28556 18562 28602 18574
rect 28674 18750 28720 18762
rect 28674 18574 28680 18750
rect 28714 18574 28720 18750
rect 28674 18562 28720 18574
rect 28792 18750 28838 18762
rect 28792 18574 28798 18750
rect 28832 18574 28838 18750
rect 28792 18562 28838 18574
rect 28910 18750 28956 18762
rect 28910 18574 28916 18750
rect 28950 18574 28956 18750
rect 28910 18562 28956 18574
rect 29028 18750 29074 18762
rect 29028 18574 29034 18750
rect 29068 18574 29074 18750
rect 29028 18562 29074 18574
rect 29146 18750 29192 18762
rect 29146 18574 29152 18750
rect 29186 18574 29192 18750
rect 29146 18562 29192 18574
rect 29264 18750 29310 18762
rect 29264 18574 29270 18750
rect 29304 18574 29310 18750
rect 29264 18562 29310 18574
rect 29382 18750 29428 18762
rect 29382 18574 29388 18750
rect 29422 18574 29428 18750
rect 29382 18562 29428 18574
rect 29500 18750 29546 18762
rect 29500 18574 29506 18750
rect 29540 18574 29546 18750
rect 29500 18562 29546 18574
rect 29618 18750 29664 18762
rect 29618 18574 29624 18750
rect 29658 18574 29664 18750
rect 29618 18562 29664 18574
rect 24710 18512 24756 18524
rect 24710 18336 24716 18512
rect 24750 18336 24756 18512
rect 24710 18324 24756 18336
rect 24828 18512 24874 18524
rect 24828 18336 24834 18512
rect 24868 18336 24874 18512
rect 24828 18324 24874 18336
rect 25234 18512 25280 18524
rect 24835 18030 24868 18324
rect 25234 18136 25240 18512
rect 25274 18136 25280 18512
rect 25234 18124 25280 18136
rect 25352 18512 25398 18524
rect 25352 18136 25358 18512
rect 25392 18136 25398 18512
rect 25352 18124 25398 18136
rect 25470 18512 25516 18524
rect 25470 18136 25476 18512
rect 25510 18136 25516 18512
rect 25470 18124 25516 18136
rect 25588 18512 25634 18524
rect 25588 18136 25594 18512
rect 25628 18136 25634 18512
rect 25588 18124 25634 18136
rect 25706 18512 25752 18524
rect 25706 18136 25712 18512
rect 25746 18136 25752 18512
rect 26008 18512 26054 18524
rect 26008 18336 26014 18512
rect 26048 18336 26054 18512
rect 26008 18324 26054 18336
rect 26126 18512 26172 18524
rect 26126 18336 26132 18512
rect 26166 18336 26172 18512
rect 26126 18324 26172 18336
rect 26608 18512 26654 18524
rect 26608 18336 26614 18512
rect 26648 18336 26654 18512
rect 26608 18324 26654 18336
rect 26726 18512 26772 18524
rect 26726 18336 26732 18512
rect 26766 18336 26772 18512
rect 26726 18324 26772 18336
rect 27132 18512 27178 18524
rect 25706 18124 25752 18136
rect 25358 18030 25392 18124
rect 26015 18030 26049 18324
rect 24835 17998 26049 18030
rect 26733 18030 26766 18324
rect 27132 18136 27138 18512
rect 27172 18136 27178 18512
rect 27132 18124 27178 18136
rect 27250 18512 27296 18524
rect 27250 18136 27256 18512
rect 27290 18136 27296 18512
rect 27250 18124 27296 18136
rect 27368 18512 27414 18524
rect 27368 18136 27374 18512
rect 27408 18136 27414 18512
rect 27368 18124 27414 18136
rect 27486 18512 27532 18524
rect 27486 18136 27492 18512
rect 27526 18136 27532 18512
rect 27486 18124 27532 18136
rect 27604 18512 27650 18524
rect 27604 18136 27610 18512
rect 27644 18136 27650 18512
rect 27906 18512 27952 18524
rect 27906 18336 27912 18512
rect 27946 18336 27952 18512
rect 27906 18324 27952 18336
rect 28024 18512 28070 18524
rect 28024 18336 28030 18512
rect 28064 18336 28070 18512
rect 28024 18324 28070 18336
rect 28562 18329 28597 18562
rect 28841 18514 28907 18521
rect 28841 18480 28857 18514
rect 28891 18480 28907 18514
rect 28841 18469 28907 18480
rect 29033 18469 29069 18562
rect 28841 18468 29069 18469
rect 29269 18468 29305 18562
rect 29505 18468 29541 18562
rect 28841 18439 29541 18468
rect 28959 18438 29541 18439
rect 28959 18397 29025 18438
rect 28959 18363 28975 18397
rect 29009 18363 29025 18397
rect 28959 18356 29025 18363
rect 28562 18325 28951 18329
rect 29387 18325 29421 18438
rect 27604 18124 27650 18136
rect 27256 18030 27290 18124
rect 27913 18030 27947 18324
rect 28562 18313 28956 18325
rect 28562 18300 28916 18313
rect 28562 18297 28640 18300
rect 28557 18245 28567 18297
rect 28630 18245 28640 18297
rect 28562 18239 28635 18245
rect 28910 18137 28916 18300
rect 28950 18137 28956 18313
rect 28910 18125 28956 18137
rect 29028 18313 29074 18325
rect 29028 18137 29034 18313
rect 29068 18137 29074 18313
rect 29028 18125 29074 18137
rect 29145 18313 29191 18325
rect 26733 17998 27947 18030
rect 28829 18009 28937 18019
rect 29033 18009 29068 18125
rect 25424 17913 25556 17998
rect 27322 17913 27454 17998
rect 24569 17606 24635 17885
rect 25414 17805 25424 17913
rect 25556 17805 25566 17913
rect 27312 17805 27322 17913
rect 27454 17805 27464 17913
rect 28937 17961 29068 18009
rect 29145 17961 29151 18313
rect 28937 17937 29151 17961
rect 29185 17937 29191 18313
rect 28937 17925 29191 17937
rect 29263 18313 29309 18325
rect 29263 17937 29269 18313
rect 29303 17937 29309 18313
rect 29263 17925 29309 17937
rect 29381 18313 29427 18325
rect 29381 17937 29387 18313
rect 29421 17937 29427 18313
rect 29381 17925 29427 17937
rect 28937 17921 29185 17925
rect 30086 17923 30179 19097
rect 32144 18662 32318 24351
rect 36611 23910 36668 24673
rect 36755 24667 37155 24673
rect 36755 24589 37155 24595
rect 36755 24555 36767 24589
rect 37143 24555 37155 24589
rect 36755 24549 37155 24555
rect 36755 24471 37155 24477
rect 36755 24437 36767 24471
rect 37143 24437 37155 24471
rect 36755 24431 37155 24437
rect 36755 24353 37155 24359
rect 36755 24319 36767 24353
rect 37143 24319 37155 24353
rect 36755 24313 37155 24319
rect 36755 24240 37155 24246
rect 36755 24206 36767 24240
rect 37143 24206 37281 24240
rect 36755 24200 37155 24206
rect 36755 24122 37155 24128
rect 36755 24088 36767 24122
rect 37143 24088 37155 24122
rect 36755 24082 37155 24088
rect 36755 24004 37155 24010
rect 36755 23970 36767 24004
rect 37143 23970 37155 24004
rect 36755 23964 37155 23970
rect 36511 23900 36668 23910
rect 36571 23820 36668 23900
rect 36755 23886 37155 23892
rect 36755 23852 36767 23886
rect 37143 23852 37155 23886
rect 36755 23846 37155 23852
rect 36511 23810 36668 23820
rect 36611 23532 36668 23810
rect 36755 23768 37155 23774
rect 36755 23734 36767 23768
rect 37143 23734 37155 23768
rect 36755 23728 37155 23734
rect 36755 23650 37155 23656
rect 36755 23616 36767 23650
rect 37143 23616 37155 23650
rect 36755 23610 37155 23616
rect 36755 23532 37155 23538
rect 36611 23498 36767 23532
rect 37143 23498 37155 23532
rect 32661 23049 32831 23063
rect 32661 22977 32676 23049
rect 32811 22977 32831 23049
rect 32661 22969 32831 22977
rect 32661 19132 32829 22969
rect 36611 22941 36668 23498
rect 36755 23492 37155 23498
rect 36755 23413 37155 23419
rect 36755 23379 36767 23413
rect 37143 23379 37155 23413
rect 36755 23373 37155 23379
rect 36755 23295 37155 23301
rect 36755 23261 36767 23295
rect 37143 23261 37155 23295
rect 36755 23255 37155 23261
rect 36755 23177 37155 23183
rect 36755 23143 36767 23177
rect 37143 23143 37155 23177
rect 36755 23137 37155 23143
rect 36755 23059 37155 23065
rect 37239 23059 37281 24206
rect 37341 24062 37408 25114
rect 37441 25047 37526 25059
rect 37441 24976 37454 25047
rect 37517 24976 37526 25047
rect 37441 24967 37526 24976
rect 37918 24315 37965 25114
rect 38088 24315 38288 24320
rect 37918 24314 38288 24315
rect 37918 24281 38100 24314
rect 37341 24028 37358 24062
rect 37392 24028 37408 24062
rect 37341 24012 37408 24028
rect 37729 24080 37814 24092
rect 37729 24012 37737 24080
rect 37802 24012 37814 24080
rect 37729 24000 37814 24012
rect 37444 23962 37529 23974
rect 37444 23892 37454 23962
rect 37516 23892 37529 23962
rect 37444 23882 37529 23892
rect 37918 23843 37965 24281
rect 38088 24280 38100 24281
rect 38276 24280 38288 24314
rect 38088 24274 38288 24280
rect 38088 24196 38288 24202
rect 38088 24162 38100 24196
rect 38276 24162 38707 24196
rect 38088 24128 38288 24162
rect 38088 24122 38488 24128
rect 38088 24088 38100 24122
rect 38476 24088 38488 24122
rect 38088 24082 38488 24088
rect 38088 24004 38488 24010
rect 38088 23970 38100 24004
rect 38476 23970 38488 24004
rect 38088 23964 38488 23970
rect 38088 23886 38488 23892
rect 38561 23886 38627 23901
rect 38088 23852 38100 23886
rect 38476 23885 38627 23886
rect 38476 23852 38577 23885
rect 38088 23846 38488 23852
rect 38561 23851 38577 23852
rect 38611 23851 38627 23885
rect 37918 23827 38028 23843
rect 38561 23835 38627 23851
rect 38655 23898 38707 24162
rect 38655 23886 38785 23898
rect 37918 23793 37978 23827
rect 38012 23793 38028 23827
rect 37918 23777 38028 23793
rect 38655 23820 38729 23886
rect 38781 23820 38785 23886
rect 38655 23806 38785 23820
rect 38088 23768 38488 23774
rect 38088 23734 38100 23768
rect 38476 23734 38488 23768
rect 38088 23728 38488 23734
rect 37568 23721 37640 23727
rect 37568 23662 37574 23721
rect 37634 23662 37640 23721
rect 37571 23658 37638 23662
rect 37574 23652 37634 23658
rect 38088 23650 38488 23656
rect 38088 23616 38100 23650
rect 38476 23616 38488 23650
rect 38088 23610 38488 23616
rect 38088 23572 38288 23610
rect 38655 23572 38707 23806
rect 38088 23538 38100 23572
rect 38276 23538 38707 23572
rect 38088 23532 38288 23538
rect 37917 23454 37964 23455
rect 38088 23454 38288 23460
rect 37917 23420 38100 23454
rect 38276 23420 38288 23454
rect 36755 23025 36767 23059
rect 37143 23025 37367 23059
rect 36755 23019 37155 23025
rect 36955 22941 37155 22946
rect 36611 22940 37155 22941
rect 35893 22917 36018 22918
rect 33301 22916 36018 22917
rect 33230 22899 36018 22916
rect 36611 22906 36967 22940
rect 37143 22906 37155 22940
rect 36611 22904 37155 22906
rect 36955 22900 37155 22904
rect 33230 22809 33244 22899
rect 33374 22809 36018 22899
rect 33230 22790 36018 22809
rect 33301 22788 36018 22790
rect 35893 22257 36018 22788
rect 36955 22822 37155 22828
rect 36955 22788 36967 22822
rect 37143 22788 37155 22822
rect 36955 22782 37155 22788
rect 37301 22752 37367 23025
rect 37301 22718 37317 22752
rect 37351 22718 37367 22752
rect 36955 22704 37155 22710
rect 36955 22670 36967 22704
rect 37143 22670 37155 22704
rect 37301 22702 37367 22718
rect 36955 22664 37155 22670
rect 36955 22586 37155 22592
rect 37917 22586 37964 23420
rect 38088 23414 38288 23420
rect 36955 22552 36967 22586
rect 37143 22554 37964 22586
rect 37143 22553 38044 22554
rect 39204 22553 39596 22677
rect 37143 22552 39596 22553
rect 36955 22551 39596 22552
rect 36955 22546 37155 22551
rect 37509 22405 39596 22551
rect 37605 22403 39596 22405
rect 39204 22308 39596 22403
rect 34496 22246 34557 22248
rect 34480 22163 34490 22246
rect 34558 22163 34568 22246
rect 35893 22170 37645 22257
rect 34496 22161 34557 22163
rect 37561 22147 37645 22170
rect 37561 22090 37569 22147
rect 37637 22090 37645 22147
rect 37561 22088 37645 22090
rect 37729 22147 37813 22169
rect 37729 22090 37737 22147
rect 37805 22090 37813 22147
rect 37729 22088 37813 22090
rect 37569 22080 37637 22088
rect 37737 22080 37805 22088
rect 36955 22005 37155 22010
rect 36955 22004 37965 22005
rect 36955 21970 36967 22004
rect 37143 21970 37965 22004
rect 36955 21964 37155 21970
rect 36955 21886 37155 21892
rect 36955 21852 36967 21886
rect 37143 21852 37155 21886
rect 36955 21846 37155 21852
rect 36955 21768 37155 21774
rect 36955 21734 36967 21768
rect 37143 21734 37155 21768
rect 36955 21728 37155 21734
rect 36955 21650 37155 21656
rect 36955 21616 36967 21650
rect 37143 21616 37155 21650
rect 36955 21569 37155 21616
rect 36755 21563 37155 21569
rect 36611 21529 36767 21563
rect 37143 21529 37155 21563
rect 36611 20766 36668 21529
rect 36755 21523 37155 21529
rect 36755 21445 37155 21451
rect 36755 21411 36767 21445
rect 37143 21411 37155 21445
rect 36755 21405 37155 21411
rect 36755 21327 37155 21333
rect 36755 21293 36767 21327
rect 37143 21293 37155 21327
rect 36755 21287 37155 21293
rect 36755 21209 37155 21215
rect 36755 21175 36767 21209
rect 37143 21175 37155 21209
rect 36755 21169 37155 21175
rect 36755 21096 37155 21102
rect 36755 21062 36767 21096
rect 37143 21062 37281 21096
rect 36755 21056 37155 21062
rect 36755 20978 37155 20984
rect 36755 20944 36767 20978
rect 37143 20944 37155 20978
rect 36755 20938 37155 20944
rect 36755 20860 37155 20866
rect 36755 20826 36767 20860
rect 37143 20826 37155 20860
rect 36755 20820 37155 20826
rect 36511 20756 36668 20766
rect 36571 20676 36668 20756
rect 36755 20742 37155 20748
rect 36755 20708 36767 20742
rect 37143 20708 37155 20742
rect 36755 20702 37155 20708
rect 36511 20666 36668 20676
rect 36611 20388 36668 20666
rect 36755 20624 37155 20630
rect 36755 20590 36767 20624
rect 37143 20590 37155 20624
rect 36755 20584 37155 20590
rect 36755 20506 37155 20512
rect 36755 20472 36767 20506
rect 37143 20472 37155 20506
rect 36755 20466 37155 20472
rect 36755 20388 37155 20394
rect 36611 20354 36767 20388
rect 37143 20354 37155 20388
rect 36611 19797 36668 20354
rect 36755 20348 37155 20354
rect 36755 20269 37155 20275
rect 36755 20235 36767 20269
rect 37143 20235 37155 20269
rect 36755 20229 37155 20235
rect 36755 20151 37155 20157
rect 36755 20117 36767 20151
rect 37143 20117 37155 20151
rect 36755 20111 37155 20117
rect 36755 20033 37155 20039
rect 36755 19999 36767 20033
rect 37143 19999 37155 20033
rect 36755 19993 37155 19999
rect 36755 19915 37155 19921
rect 37239 19915 37281 21062
rect 37341 20918 37408 21970
rect 37441 21903 37526 21915
rect 37441 21832 37454 21903
rect 37517 21832 37526 21903
rect 37441 21823 37526 21832
rect 37918 21171 37965 21970
rect 38088 21171 38288 21176
rect 37918 21170 38288 21171
rect 37918 21137 38100 21170
rect 37341 20884 37358 20918
rect 37392 20884 37408 20918
rect 37341 20868 37408 20884
rect 37729 20936 37814 20948
rect 37729 20868 37737 20936
rect 37802 20868 37814 20936
rect 37729 20856 37814 20868
rect 37444 20818 37529 20830
rect 37444 20748 37454 20818
rect 37516 20748 37529 20818
rect 37444 20738 37529 20748
rect 37918 20699 37965 21137
rect 38088 21136 38100 21137
rect 38276 21136 38288 21170
rect 38088 21130 38288 21136
rect 38088 21052 38288 21058
rect 38088 21018 38100 21052
rect 38276 21018 38707 21052
rect 38088 20984 38288 21018
rect 38088 20978 38488 20984
rect 38088 20944 38100 20978
rect 38476 20944 38488 20978
rect 38088 20938 38488 20944
rect 38088 20860 38488 20866
rect 38088 20826 38100 20860
rect 38476 20826 38488 20860
rect 38088 20820 38488 20826
rect 38088 20742 38488 20748
rect 38561 20742 38627 20757
rect 38088 20708 38100 20742
rect 38476 20741 38627 20742
rect 38476 20708 38577 20741
rect 38088 20702 38488 20708
rect 38561 20707 38577 20708
rect 38611 20707 38627 20741
rect 37918 20683 38028 20699
rect 38561 20691 38627 20707
rect 38655 20754 38707 21018
rect 38655 20742 38785 20754
rect 37918 20649 37978 20683
rect 38012 20649 38028 20683
rect 37918 20633 38028 20649
rect 38655 20676 38729 20742
rect 38781 20676 38785 20742
rect 38655 20662 38785 20676
rect 38088 20624 38488 20630
rect 38088 20590 38100 20624
rect 38476 20590 38488 20624
rect 38088 20584 38488 20590
rect 37568 20577 37640 20583
rect 37568 20518 37574 20577
rect 37634 20518 37640 20577
rect 37571 20514 37638 20518
rect 37574 20508 37634 20514
rect 38088 20506 38488 20512
rect 38088 20472 38100 20506
rect 38476 20472 38488 20506
rect 38088 20466 38488 20472
rect 38088 20428 38288 20466
rect 38655 20428 38707 20662
rect 38088 20394 38100 20428
rect 38276 20394 38707 20428
rect 38088 20388 38288 20394
rect 37917 20310 37964 20311
rect 38088 20310 38288 20316
rect 37917 20276 38100 20310
rect 38276 20276 38288 20310
rect 36755 19881 36767 19915
rect 37143 19881 37367 19915
rect 36755 19875 37155 19881
rect 36955 19797 37155 19802
rect 36611 19796 37155 19797
rect 36611 19762 36967 19796
rect 37143 19762 37155 19796
rect 36611 19760 37155 19762
rect 36955 19756 37155 19760
rect 36955 19678 37155 19684
rect 36955 19644 36967 19678
rect 37143 19644 37155 19678
rect 36955 19638 37155 19644
rect 37301 19608 37367 19881
rect 37301 19574 37317 19608
rect 37351 19574 37367 19608
rect 36955 19560 37155 19566
rect 36955 19526 36967 19560
rect 37143 19526 37155 19560
rect 37301 19558 37367 19574
rect 36955 19520 37155 19526
rect 36955 19442 37155 19448
rect 37917 19442 37964 20276
rect 38088 20270 38288 20276
rect 36955 19408 36967 19442
rect 37143 19412 37964 19442
rect 37143 19411 38054 19412
rect 39205 19411 39597 19535
rect 37143 19408 39597 19411
rect 36955 19407 39597 19408
rect 36955 19402 37155 19407
rect 37509 19262 39597 19407
rect 37509 19261 37655 19262
rect 37965 19261 39597 19262
rect 39205 19166 39597 19261
rect 32661 19054 37642 19132
rect 32662 19032 37642 19054
rect 32662 19030 33541 19032
rect 37557 19015 37641 19032
rect 37557 18958 37565 19015
rect 37633 18958 37641 19015
rect 37557 18956 37641 18958
rect 37725 19015 37809 19033
rect 37725 18958 37733 19015
rect 37801 18958 37809 19015
rect 37725 18956 37809 18958
rect 37565 18948 37633 18956
rect 37733 18948 37801 18956
rect 36951 18873 37151 18878
rect 36951 18872 37961 18873
rect 36951 18838 36963 18872
rect 37139 18838 37961 18872
rect 36951 18832 37151 18838
rect 36951 18754 37151 18760
rect 36951 18720 36963 18754
rect 37139 18720 37151 18754
rect 36951 18714 37151 18720
rect 32144 18509 35897 18662
rect 36951 18636 37151 18642
rect 36951 18602 36963 18636
rect 37139 18602 37151 18636
rect 36951 18596 37151 18602
rect 32250 18508 35897 18509
rect 29594 17921 30179 17923
rect 28937 17877 29011 17921
rect 29549 17893 30179 17921
rect 29194 17887 29260 17893
rect 28829 17867 28937 17877
rect 29194 17853 29210 17887
rect 29244 17853 29260 17887
rect 29194 17757 29260 17853
rect 29312 17887 30179 17893
rect 29312 17853 29328 17887
rect 29362 17853 30179 17887
rect 29312 17837 30179 17853
rect 29549 17821 30179 17837
rect 29594 17817 30179 17821
rect 30078 17816 30179 17817
rect 29549 17768 29649 17779
rect 29549 17757 29563 17768
rect 29194 17709 29563 17757
rect 29195 17606 29261 17709
rect 29549 17679 29563 17709
rect 29553 17662 29563 17679
rect 29675 17662 29685 17768
rect 24569 17526 29263 17606
rect 24351 16988 35434 17068
rect 35218 16953 35298 16954
rect 17838 16870 35298 16953
rect 11304 16769 35176 16842
rect 4746 16633 35045 16739
rect 4794 16632 35045 16633
rect 32275 16629 35045 16632
rect 30657 16600 30780 16601
rect 30476 16599 30780 16600
rect 52 16592 30780 16599
rect 52 16591 30617 16592
rect 52 16502 30607 16591
rect 52 16501 30617 16502
rect 30768 16501 30780 16592
rect 52 16488 30780 16501
rect 30657 16486 30780 16488
rect 34956 16594 35045 16629
rect -86 16446 22331 16447
rect -86 16433 24261 16446
rect -86 16345 24097 16433
rect 24246 16345 24261 16433
rect -86 16336 24261 16345
rect 20247 16335 24261 16336
rect 23841 16333 24261 16335
rect -216 16286 17738 16296
rect -216 16198 17570 16286
rect 17726 16198 17738 16286
rect -216 16185 17738 16198
rect 23963 16176 23973 16251
rect 24059 16176 24069 16251
rect -349 16126 11143 16140
rect -349 16029 11000 16126
rect 11129 16029 11143 16126
rect 17440 16060 17450 16130
rect 17537 16060 17547 16130
rect -349 16019 11143 16029
rect 2300 15963 34901 15964
rect -514 15952 34901 15963
rect -514 15871 34744 15952
rect 34888 15871 34901 15952
rect -514 15861 34901 15871
rect -514 15860 32183 15861
rect 10865 15736 10875 15797
rect 10968 15736 10978 15797
rect 28928 15686 34897 15794
rect 28928 15532 29041 15686
rect 34778 15675 34897 15686
rect 29111 15590 34737 15658
rect 21320 15482 21456 15502
rect 8117 15462 8253 15482
rect 8117 15400 8153 15462
rect 8213 15400 8253 15462
rect 8117 15372 8253 15400
rect 14666 15461 14802 15481
rect 14666 15399 14702 15461
rect 14762 15399 14802 15461
rect 7813 15342 8790 15372
rect 14666 15371 14802 15399
rect 21320 15420 21356 15482
rect 21416 15420 21456 15482
rect 21320 15392 21456 15420
rect 7813 15236 7845 15342
rect 8049 15236 8081 15342
rect 8285 15236 8317 15342
rect 8521 15236 8553 15342
rect 8756 15236 8790 15342
rect 14362 15341 15339 15371
rect 7806 15224 7852 15236
rect 7806 15048 7812 15224
rect 7846 15048 7852 15224
rect 7806 15036 7852 15048
rect 7924 15224 7970 15236
rect 7924 15048 7930 15224
rect 7964 15048 7970 15224
rect 7924 15036 7970 15048
rect 8042 15224 8088 15236
rect 8042 15048 8048 15224
rect 8082 15048 8088 15224
rect 8042 15036 8088 15048
rect 8160 15224 8206 15236
rect 8160 15048 8166 15224
rect 8200 15048 8206 15224
rect 8160 15036 8206 15048
rect 8278 15224 8324 15236
rect 8278 15048 8284 15224
rect 8318 15048 8324 15224
rect 8278 15036 8324 15048
rect 8396 15224 8442 15236
rect 8396 15048 8402 15224
rect 8436 15048 8442 15224
rect 8396 15036 8442 15048
rect 8514 15224 8560 15236
rect 8514 15048 8520 15224
rect 8554 15048 8560 15224
rect 8514 15036 8560 15048
rect 8632 15224 8678 15236
rect 8632 15048 8638 15224
rect 8672 15048 8678 15224
rect 8632 15036 8678 15048
rect 8750 15224 8796 15236
rect 8750 15048 8756 15224
rect 8790 15048 8796 15224
rect 8750 15036 8796 15048
rect 8868 15224 8914 15236
rect 14362 15235 14394 15341
rect 14598 15235 14630 15341
rect 14834 15235 14866 15341
rect 15070 15235 15102 15341
rect 15305 15235 15339 15341
rect 21016 15362 21993 15392
rect 21016 15256 21048 15362
rect 21252 15256 21284 15362
rect 21488 15256 21520 15362
rect 21724 15256 21756 15362
rect 21959 15256 21993 15362
rect 21009 15244 21055 15256
rect 8868 15048 8874 15224
rect 8908 15048 8914 15224
rect 8868 15036 8914 15048
rect 14355 15223 14401 15235
rect 14355 15047 14361 15223
rect 14395 15047 14401 15223
rect 7929 14942 7965 15036
rect 8165 14942 8201 15036
rect 8401 14943 8437 15036
rect 8563 14988 8629 14995
rect 8563 14954 8579 14988
rect 8613 14954 8629 14988
rect 8563 14943 8629 14954
rect 8401 14942 8629 14943
rect 7929 14913 8629 14942
rect 7929 14912 8511 14913
rect 8049 14799 8083 14912
rect 8445 14871 8511 14912
rect 8445 14837 8461 14871
rect 8495 14837 8511 14871
rect 8445 14830 8511 14837
rect 8873 14805 8908 15036
rect 14355 15035 14401 15047
rect 14473 15223 14519 15235
rect 14473 15047 14479 15223
rect 14513 15047 14519 15223
rect 14473 15035 14519 15047
rect 14591 15223 14637 15235
rect 14591 15047 14597 15223
rect 14631 15047 14637 15223
rect 14591 15035 14637 15047
rect 14709 15223 14755 15235
rect 14709 15047 14715 15223
rect 14749 15047 14755 15223
rect 14709 15035 14755 15047
rect 14827 15223 14873 15235
rect 14827 15047 14833 15223
rect 14867 15047 14873 15223
rect 14827 15035 14873 15047
rect 14945 15223 14991 15235
rect 14945 15047 14951 15223
rect 14985 15047 14991 15223
rect 14945 15035 14991 15047
rect 15063 15223 15109 15235
rect 15063 15047 15069 15223
rect 15103 15047 15109 15223
rect 15063 15035 15109 15047
rect 15181 15223 15227 15235
rect 15181 15047 15187 15223
rect 15221 15047 15227 15223
rect 15181 15035 15227 15047
rect 15299 15223 15345 15235
rect 15299 15047 15305 15223
rect 15339 15047 15345 15223
rect 15299 15035 15345 15047
rect 15417 15223 15463 15235
rect 15417 15047 15423 15223
rect 15457 15047 15463 15223
rect 21009 15068 21015 15244
rect 21049 15068 21055 15244
rect 21009 15056 21055 15068
rect 21127 15244 21173 15256
rect 21127 15068 21133 15244
rect 21167 15068 21173 15244
rect 21127 15056 21173 15068
rect 21245 15244 21291 15256
rect 21245 15068 21251 15244
rect 21285 15068 21291 15244
rect 21245 15056 21291 15068
rect 21363 15244 21409 15256
rect 21363 15068 21369 15244
rect 21403 15068 21409 15244
rect 21363 15056 21409 15068
rect 21481 15244 21527 15256
rect 21481 15068 21487 15244
rect 21521 15068 21527 15244
rect 21481 15056 21527 15068
rect 21599 15244 21645 15256
rect 21599 15068 21605 15244
rect 21639 15068 21645 15244
rect 21599 15056 21645 15068
rect 21717 15244 21763 15256
rect 21717 15068 21723 15244
rect 21757 15068 21763 15244
rect 21717 15056 21763 15068
rect 21835 15244 21881 15256
rect 21835 15068 21841 15244
rect 21875 15068 21881 15244
rect 21835 15056 21881 15068
rect 21953 15244 21999 15256
rect 21953 15068 21959 15244
rect 21993 15068 21999 15244
rect 21953 15056 21999 15068
rect 22071 15244 22117 15256
rect 22071 15068 22077 15244
rect 22111 15068 22117 15244
rect 22071 15056 22117 15068
rect 15417 15035 15463 15047
rect 14478 14941 14514 15035
rect 14714 14941 14750 15035
rect 14950 14942 14986 15035
rect 15112 14987 15178 14994
rect 15112 14953 15128 14987
rect 15162 14953 15178 14987
rect 15112 14942 15178 14953
rect 14950 14941 15178 14942
rect 14478 14912 15178 14941
rect 14478 14911 15060 14912
rect 8803 14803 10120 14805
rect 8519 14799 10120 14803
rect 8043 14787 8089 14799
rect 8043 14411 8049 14787
rect 8083 14411 8089 14787
rect 8043 14399 8089 14411
rect 8161 14787 8207 14799
rect 8161 14411 8167 14787
rect 8201 14411 8207 14787
rect 8161 14399 8207 14411
rect 8279 14787 8325 14799
rect 8279 14411 8285 14787
rect 8319 14438 8325 14787
rect 8396 14787 8442 14799
rect 8396 14611 8402 14787
rect 8436 14611 8442 14787
rect 8396 14604 8442 14611
rect 8514 14787 10120 14799
rect 14598 14798 14632 14911
rect 14994 14870 15060 14911
rect 14994 14836 15010 14870
rect 15044 14836 15060 14870
rect 14994 14829 15060 14836
rect 15422 14837 15457 15035
rect 21132 14962 21168 15056
rect 21368 14962 21404 15056
rect 21604 14963 21640 15056
rect 21766 15008 21832 15015
rect 21766 14974 21782 15008
rect 21816 14974 21832 15008
rect 21766 14963 21832 14974
rect 21604 14962 21832 14963
rect 21132 14933 21832 14962
rect 21132 14932 21714 14933
rect 15422 14802 15458 14837
rect 21252 14819 21286 14932
rect 21648 14891 21714 14932
rect 21648 14857 21664 14891
rect 21698 14857 21714 14891
rect 21648 14850 21714 14857
rect 22076 14823 22111 15056
rect 21722 14819 23396 14823
rect 21246 14807 21292 14819
rect 15068 14798 16770 14802
rect 8514 14611 8520 14787
rect 8554 14774 10120 14787
rect 8554 14611 8560 14774
rect 8803 14693 10120 14774
rect 8396 14599 8445 14604
rect 8514 14599 8560 14611
rect 8402 14438 8445 14599
rect 8319 14411 8445 14438
rect 8279 14399 8445 14411
rect 8285 14395 8445 14399
rect 7790 14361 8158 14367
rect 7790 14327 8108 14361
rect 8142 14327 8158 14361
rect 7790 14311 8158 14327
rect 8210 14361 8276 14367
rect 8210 14327 8226 14361
rect 8260 14327 8276 14361
rect -661 14192 -651 14246
rect -594 14192 -584 14246
rect -661 12190 -586 14192
rect 7790 14119 7869 14311
rect 8210 14282 8276 14327
rect 203 14109 7869 14119
rect 203 14059 227 14109
rect 288 14059 7869 14109
rect 203 14049 7869 14059
rect 7927 14274 8276 14282
rect 7927 14242 8277 14274
rect 8369 14258 8445 14395
rect 7927 13948 7981 14242
rect 8365 14198 8375 14258
rect 8437 14198 8447 14258
rect 7924 13936 7985 13948
rect 54 13927 229 13933
rect 54 13871 66 13927
rect 125 13924 229 13927
rect 125 13871 135 13924
rect 54 13866 135 13871
rect 219 13866 229 13924
rect 7924 13882 7930 13936
rect 7979 13882 7985 13936
rect 7924 13870 7985 13882
rect 54 13865 229 13866
rect 1453 13562 1589 13582
rect 368 13539 449 13542
rect 363 13487 373 13539
rect 441 13487 451 13539
rect 1453 13500 1489 13562
rect 1549 13500 1589 13562
rect 368 13485 449 13487
rect 1453 13472 1589 13500
rect 6989 13522 7068 13534
rect 4507 13472 4586 13484
rect 1149 13442 2126 13472
rect 1149 13336 1181 13442
rect 1385 13336 1417 13442
rect 1621 13336 1653 13442
rect 1857 13336 1889 13442
rect 2092 13336 2126 13442
rect 4507 13375 4513 13472
rect 4435 13355 4513 13375
rect 4580 13375 4586 13472
rect 6989 13409 6995 13522
rect 7062 13409 7068 13522
rect 8131 13524 8210 13536
rect 8131 13409 8137 13524
rect 8204 13409 8210 13524
rect 4580 13355 4655 13375
rect 1142 13324 1188 13336
rect 1142 13148 1148 13324
rect 1182 13148 1188 13324
rect 1142 13136 1188 13148
rect 1260 13324 1306 13336
rect 1260 13148 1266 13324
rect 1300 13148 1306 13324
rect 1260 13136 1306 13148
rect 1378 13324 1424 13336
rect 1378 13148 1384 13324
rect 1418 13148 1424 13324
rect 1378 13136 1424 13148
rect 1496 13324 1542 13336
rect 1496 13148 1502 13324
rect 1536 13148 1542 13324
rect 1496 13136 1542 13148
rect 1614 13324 1660 13336
rect 1614 13148 1620 13324
rect 1654 13148 1660 13324
rect 1614 13136 1660 13148
rect 1732 13324 1778 13336
rect 1732 13148 1738 13324
rect 1772 13148 1778 13324
rect 1732 13136 1778 13148
rect 1850 13324 1896 13336
rect 1850 13148 1856 13324
rect 1890 13148 1896 13324
rect 1850 13136 1896 13148
rect 1968 13324 2014 13336
rect 1968 13148 1974 13324
rect 2008 13148 2014 13324
rect 1968 13136 2014 13148
rect 2086 13324 2132 13336
rect 2086 13148 2092 13324
rect 2126 13148 2132 13324
rect 2086 13136 2132 13148
rect 2204 13324 2250 13336
rect 2204 13148 2210 13324
rect 2244 13148 2250 13324
rect 4435 13247 4479 13355
rect 4611 13247 4655 13355
rect 6232 13313 6288 13321
rect 4435 13205 4655 13247
rect 5306 13305 6288 13313
rect 5306 13271 6248 13305
rect 6282 13271 6288 13305
rect 6951 13301 6961 13409
rect 7093 13346 7103 13409
rect 7093 13335 7105 13346
rect 7093 13301 7106 13335
rect 7362 13325 7418 13327
rect 5306 13255 6288 13271
rect 6961 13263 7106 13301
rect 5306 13254 6285 13255
rect 2204 13136 2250 13148
rect 4039 13175 5016 13205
rect 1265 13042 1301 13136
rect 1501 13042 1537 13136
rect 1737 13043 1773 13136
rect 1899 13088 1965 13095
rect 1899 13054 1915 13088
rect 1949 13054 1965 13088
rect 1899 13043 1965 13054
rect 1737 13042 1965 13043
rect 1265 13013 1965 13042
rect 1265 13012 1847 13013
rect 1385 12899 1419 13012
rect 1781 12971 1847 13012
rect 1781 12937 1797 12971
rect 1831 12937 1847 12971
rect 1781 12930 1847 12937
rect 2209 12903 2244 13136
rect 4039 13069 4071 13175
rect 4275 13069 4307 13175
rect 4511 13069 4543 13175
rect 4747 13069 4779 13175
rect 4982 13069 5016 13175
rect 1855 12899 2244 12903
rect 1379 12887 1425 12899
rect 5 12582 1339 12597
rect 5 12512 23 12582
rect 97 12580 1339 12582
rect 97 12512 645 12580
rect 5 12504 645 12512
rect 734 12504 1339 12580
rect 5 12497 1339 12504
rect 1379 12511 1385 12887
rect 1419 12511 1425 12887
rect 1379 12499 1425 12511
rect 1497 12887 1543 12899
rect 1497 12511 1503 12887
rect 1537 12511 1543 12887
rect 1497 12499 1543 12511
rect 1615 12887 1661 12899
rect 1615 12511 1621 12887
rect 1655 12538 1661 12887
rect 1732 12887 1778 12899
rect 1732 12711 1738 12887
rect 1772 12711 1778 12887
rect 1732 12704 1778 12711
rect 1850 12887 2244 12899
rect 1850 12711 1856 12887
rect 1890 12874 2244 12887
rect 1890 12711 1896 12874
rect 1732 12699 1781 12704
rect 1850 12699 1896 12711
rect 1738 12538 1781 12699
rect 1655 12511 1781 12538
rect 1615 12499 1781 12511
rect 1263 12467 1317 12497
rect 1621 12495 1781 12499
rect 1263 12461 1494 12467
rect 1263 12427 1444 12461
rect 1478 12427 1494 12461
rect 4 12405 1207 12417
rect 1263 12411 1494 12427
rect 1546 12461 1612 12467
rect 1546 12427 1562 12461
rect 1596 12427 1612 12461
rect 4 12326 17 12405
rect 5 12313 17 12326
rect 107 12402 1207 12405
rect 107 12318 207 12402
rect 320 12386 1207 12402
rect 320 12342 1139 12386
rect 1195 12382 1207 12386
rect 1546 12382 1612 12427
rect 1195 12374 1612 12382
rect 1195 12342 1613 12374
rect 1705 12358 1781 12495
rect 320 12318 1208 12342
rect 107 12313 1208 12318
rect 5 12306 1208 12313
rect 1701 12298 1711 12358
rect 1773 12298 1783 12358
rect 2140 12230 2244 12874
rect 4032 13057 4078 13069
rect 4032 12881 4038 13057
rect 4072 12881 4078 13057
rect 4032 12869 4078 12881
rect 4150 13057 4196 13069
rect 4150 12881 4156 13057
rect 4190 12881 4196 13057
rect 4150 12869 4196 12881
rect 4268 13057 4314 13069
rect 4268 12881 4274 13057
rect 4308 12881 4314 13057
rect 4268 12869 4314 12881
rect 4386 13057 4432 13069
rect 4386 12881 4392 13057
rect 4426 12881 4432 13057
rect 4386 12869 4432 12881
rect 4504 13057 4550 13069
rect 4504 12881 4510 13057
rect 4544 12881 4550 13057
rect 4504 12869 4550 12881
rect 4622 13057 4668 13069
rect 4622 12881 4628 13057
rect 4662 12881 4668 13057
rect 4622 12869 4668 12881
rect 4740 13057 4786 13069
rect 4740 12881 4746 13057
rect 4780 12881 4786 13057
rect 4740 12869 4786 12881
rect 4858 13057 4904 13069
rect 4858 12881 4864 13057
rect 4898 12881 4904 13057
rect 4858 12869 4904 12881
rect 4976 13057 5022 13069
rect 4976 12881 4982 13057
rect 5016 12881 5022 13057
rect 4976 12869 5022 12881
rect 5094 13057 5140 13069
rect 5094 12881 5100 13057
rect 5134 12881 5140 13057
rect 5094 12869 5140 12881
rect 4155 12775 4191 12869
rect 4391 12775 4427 12869
rect 4627 12776 4663 12869
rect 4789 12821 4855 12828
rect 4789 12787 4805 12821
rect 4839 12787 4855 12821
rect 4789 12776 4855 12787
rect 4627 12775 4855 12776
rect 4155 12746 4855 12775
rect 4155 12745 4737 12746
rect 4275 12632 4309 12745
rect 4671 12704 4737 12745
rect 4671 12670 4687 12704
rect 4721 12670 4737 12704
rect 4671 12663 4737 12670
rect 5099 12664 5134 12869
rect 5306 12664 5373 13254
rect 7065 13231 7106 13263
rect 7352 13259 7362 13325
rect 7418 13259 7428 13325
rect 8098 13301 8108 13409
rect 8240 13346 8250 13409
rect 8240 13335 8252 13346
rect 8240 13301 8253 13335
rect 8108 13263 8253 13301
rect 8212 13235 8253 13263
rect 6481 13203 6751 13231
rect 6222 13137 6232 13203
rect 6298 13137 6308 13203
rect 6481 13141 6515 13203
rect 6717 13141 6751 13203
rect 6835 13203 7106 13231
rect 7623 13207 7893 13235
rect 6835 13141 6869 13203
rect 7071 13141 7106 13203
rect 7247 13191 7418 13207
rect 7247 13157 7378 13191
rect 7412 13157 7418 13191
rect 7247 13141 7418 13157
rect 7623 13145 7657 13207
rect 7859 13145 7893 13207
rect 7977 13207 8253 13235
rect 7977 13145 8011 13207
rect 8213 13145 8253 13207
rect 6357 13129 6403 13141
rect 6357 12753 6363 13129
rect 6397 12753 6403 13129
rect 6357 12741 6403 12753
rect 6475 13129 6521 13141
rect 6475 12753 6481 13129
rect 6515 12753 6521 13129
rect 6475 12741 6521 12753
rect 6593 13129 6639 13141
rect 6593 12753 6599 13129
rect 6633 12753 6639 13129
rect 6593 12741 6639 12753
rect 6711 13129 6757 13141
rect 6711 12753 6717 13129
rect 6751 12753 6757 13129
rect 6711 12741 6757 12753
rect 6829 13129 6875 13141
rect 6829 12753 6835 13129
rect 6869 12753 6875 13129
rect 6829 12741 6875 12753
rect 6947 13129 6993 13141
rect 6947 12753 6953 13129
rect 6987 12753 6993 13129
rect 6947 12741 6993 12753
rect 7065 13129 7111 13141
rect 7065 12753 7071 13129
rect 7105 12753 7111 13129
rect 7065 12741 7111 12753
rect 5099 12636 5373 12664
rect 4745 12632 5373 12636
rect 4269 12620 4315 12632
rect 4269 12244 4275 12620
rect 4309 12244 4315 12620
rect 4269 12232 4315 12244
rect 4387 12620 4433 12632
rect 4387 12244 4393 12620
rect 4427 12244 4433 12620
rect 4387 12232 4433 12244
rect 4505 12620 4551 12632
rect 4505 12244 4511 12620
rect 4545 12268 4551 12620
rect 4622 12620 4668 12632
rect 4622 12444 4628 12620
rect 4662 12444 4668 12620
rect 4622 12432 4668 12444
rect 4740 12620 5373 12632
rect 4740 12444 4746 12620
rect 4780 12607 5373 12620
rect 6363 12699 6397 12741
rect 6599 12699 6633 12741
rect 6363 12671 6633 12699
rect 6717 12700 6751 12741
rect 6953 12700 6987 12741
rect 6717 12671 6987 12700
rect 6363 12623 6397 12671
rect 4780 12444 4786 12607
rect 6363 12593 6426 12623
rect 4740 12432 4786 12444
rect 6391 12501 6426 12593
rect 6391 12465 6618 12501
rect 6888 12490 6898 12587
rect 6997 12490 7007 12587
rect 7071 12558 7105 12741
rect 7071 12504 7180 12558
rect 4628 12316 4663 12432
rect 6391 12358 6426 12465
rect 6552 12431 6618 12465
rect 6552 12397 6568 12431
rect 6602 12397 6618 12431
rect 6899 12489 6996 12490
rect 6899 12422 6956 12489
rect 6552 12391 6618 12397
rect 6793 12386 7062 12422
rect 6793 12358 6826 12386
rect 7029 12358 7062 12386
rect 7146 12358 7180 12504
rect 6267 12346 6313 12358
rect 4759 12316 4867 12326
rect 4628 12268 4759 12316
rect 4867 12283 5015 12289
rect 4545 12244 4759 12268
rect 4505 12232 4759 12244
rect 2140 12229 2247 12230
rect 2140 12228 2836 12229
rect 4511 12228 4759 12232
rect 2140 12227 3386 12228
rect 2140 12200 4147 12227
rect 2140 12194 4384 12200
rect -665 12129 -655 12190
rect -592 12129 -582 12190
rect 2140 12160 4334 12194
rect 4368 12160 4384 12194
rect 2140 12144 4384 12160
rect 4436 12194 4502 12200
rect 4436 12160 4452 12194
rect 4486 12160 4502 12194
rect 4685 12184 4759 12228
rect 5003 12216 5015 12283
rect 4867 12210 5015 12216
rect 4759 12174 4867 12184
rect -661 10126 -586 12129
rect 2140 12128 4147 12144
rect 2140 12127 4084 12128
rect 2140 12123 3619 12127
rect 2140 12122 3386 12123
rect 2140 12120 3227 12122
rect 2429 11712 3403 11741
rect 2429 11606 3251 11712
rect 3363 11699 3403 11712
rect 3363 11606 3405 11699
rect 2429 11595 3405 11606
rect 2429 11594 3403 11595
rect 1445 10977 1581 10997
rect 1445 10915 1481 10977
rect 1541 10915 1581 10977
rect 1445 10887 1581 10915
rect 1141 10857 2118 10887
rect 1141 10751 1173 10857
rect 1377 10751 1409 10857
rect 1613 10751 1645 10857
rect 1849 10751 1881 10857
rect 2084 10751 2118 10857
rect 1134 10739 1180 10751
rect 1134 10563 1140 10739
rect 1174 10563 1180 10739
rect 1134 10551 1180 10563
rect 1252 10739 1298 10751
rect 1252 10563 1258 10739
rect 1292 10563 1298 10739
rect 1252 10551 1298 10563
rect 1370 10739 1416 10751
rect 1370 10563 1376 10739
rect 1410 10563 1416 10739
rect 1370 10551 1416 10563
rect 1488 10739 1534 10751
rect 1488 10563 1494 10739
rect 1528 10563 1534 10739
rect 1488 10551 1534 10563
rect 1606 10739 1652 10751
rect 1606 10563 1612 10739
rect 1646 10563 1652 10739
rect 1606 10551 1652 10563
rect 1724 10739 1770 10751
rect 1724 10563 1730 10739
rect 1764 10563 1770 10739
rect 1724 10551 1770 10563
rect 1842 10739 1888 10751
rect 1842 10563 1848 10739
rect 1882 10563 1888 10739
rect 1842 10551 1888 10563
rect 1960 10739 2006 10751
rect 1960 10563 1966 10739
rect 2000 10563 2006 10739
rect 1960 10551 2006 10563
rect 2078 10739 2124 10751
rect 2078 10563 2084 10739
rect 2118 10563 2124 10739
rect 2078 10551 2124 10563
rect 2196 10739 2242 10751
rect 2196 10563 2202 10739
rect 2236 10563 2242 10739
rect 2196 10551 2242 10563
rect 1257 10457 1293 10551
rect 1493 10457 1529 10551
rect 1729 10458 1765 10551
rect 1891 10503 1957 10510
rect 1891 10469 1907 10503
rect 1941 10469 1957 10503
rect 1891 10458 1957 10469
rect 1729 10457 1957 10458
rect 1257 10428 1957 10457
rect 1257 10427 1839 10428
rect 1377 10314 1411 10427
rect 1773 10386 1839 10427
rect 1773 10352 1789 10386
rect 1823 10352 1839 10386
rect 1773 10345 1839 10352
rect 2201 10318 2236 10551
rect 2429 10318 2549 11594
rect 3221 10601 3402 10631
rect 3221 10491 3250 10601
rect 3368 10587 3402 10601
rect 3368 10491 3403 10587
rect 3221 10483 3403 10491
rect 3221 10481 3402 10483
rect 1847 10314 2549 10318
rect 1371 10302 1417 10314
rect -665 10065 -655 10126
rect -592 10065 -582 10126
rect -661 8061 -586 10065
rect 1371 9926 1377 10302
rect 1411 9926 1417 10302
rect 1371 9914 1417 9926
rect 1489 10302 1535 10314
rect 1489 9926 1495 10302
rect 1529 9926 1535 10302
rect 1489 9914 1535 9926
rect 1607 10302 1653 10314
rect 1607 9926 1613 10302
rect 1647 9953 1653 10302
rect 1724 10302 1770 10314
rect 1724 10126 1730 10302
rect 1764 10126 1770 10302
rect 1724 10119 1770 10126
rect 1842 10302 2549 10314
rect 1842 10126 1848 10302
rect 1882 10289 2549 10302
rect 1882 10126 1888 10289
rect 2132 10210 2549 10289
rect 3526 10229 3619 12123
rect 3682 12064 4148 12086
rect 4436 12064 4502 12160
rect 6267 12170 6273 12346
rect 6307 12170 6313 12346
rect 6267 12158 6313 12170
rect 6385 12346 6431 12358
rect 6385 12170 6391 12346
rect 6425 12170 6431 12346
rect 6385 12158 6431 12170
rect 6503 12346 6549 12358
rect 6503 12170 6509 12346
rect 6543 12170 6549 12346
rect 6503 12158 6549 12170
rect 6621 12346 6667 12358
rect 6621 12170 6627 12346
rect 6661 12291 6667 12346
rect 6786 12346 6832 12358
rect 6786 12291 6792 12346
rect 6661 12203 6792 12291
rect 6661 12170 6667 12203
rect 6621 12158 6667 12170
rect 6786 12170 6792 12203
rect 6826 12170 6832 12346
rect 6786 12158 6832 12170
rect 6904 12346 6950 12358
rect 6904 12170 6910 12346
rect 6944 12170 6950 12346
rect 6904 12158 6950 12170
rect 7022 12346 7068 12358
rect 7022 12170 7028 12346
rect 7062 12170 7068 12346
rect 7022 12158 7068 12170
rect 7140 12346 7186 12358
rect 7140 12170 7146 12346
rect 7180 12170 7186 12346
rect 7140 12158 7186 12170
rect 6273 12119 6307 12158
rect 6509 12119 6543 12158
rect 6273 12084 6543 12119
rect 6910 12120 6943 12158
rect 7146 12120 7179 12158
rect 6910 12084 7179 12120
rect 3682 12016 4502 12064
rect 6307 12083 6543 12084
rect 3682 11985 4148 12016
rect 6307 12009 6439 12083
rect 3682 11729 3787 11985
rect 6297 11901 6307 12009
rect 6439 11901 6449 12009
rect 4519 11821 4598 11833
rect 3682 11623 3745 11729
rect 3857 11623 3867 11729
rect 4519 11725 4525 11821
rect 4449 11705 4525 11725
rect 4592 11725 4598 11821
rect 6334 11763 6340 11901
rect 6407 11763 6413 11901
rect 6334 11751 6413 11763
rect 4592 11705 4669 11725
rect 3682 11612 3831 11623
rect 3682 10435 3787 11612
rect 4449 11597 4493 11705
rect 4625 11597 4669 11705
rect 4449 11555 4669 11597
rect 7247 11570 7309 13141
rect 7499 13133 7545 13145
rect 7499 12757 7505 13133
rect 7539 12757 7545 13133
rect 7499 12745 7545 12757
rect 7617 13133 7663 13145
rect 7617 12757 7623 13133
rect 7657 12757 7663 13133
rect 7617 12745 7663 12757
rect 7735 13133 7781 13145
rect 7735 12757 7741 13133
rect 7775 12757 7781 13133
rect 7735 12745 7781 12757
rect 7853 13133 7899 13145
rect 7853 12757 7859 13133
rect 7893 12757 7899 13133
rect 7853 12745 7899 12757
rect 7971 13133 8017 13145
rect 7971 12757 7977 13133
rect 8011 12757 8017 13133
rect 7971 12745 8017 12757
rect 8089 13133 8135 13145
rect 8089 12757 8095 13133
rect 8129 12757 8135 13133
rect 8089 12745 8135 12757
rect 8207 13133 8253 13145
rect 8207 12757 8213 13133
rect 8247 12757 8253 13133
rect 8207 12745 8253 12757
rect 7505 12703 7539 12745
rect 7741 12703 7775 12745
rect 7505 12675 7775 12703
rect 7859 12704 7893 12745
rect 8095 12704 8129 12745
rect 7859 12675 8129 12704
rect 7505 12627 7539 12675
rect 7505 12597 7568 12627
rect 7533 12505 7568 12597
rect 8040 12567 8140 12588
rect 8040 12513 8054 12567
rect 8119 12513 8140 12567
rect 8040 12508 8140 12513
rect 8213 12562 8247 12745
rect 8213 12508 8322 12562
rect 9939 12523 10120 14693
rect 14592 14786 14638 14798
rect 14592 14410 14598 14786
rect 14632 14410 14638 14786
rect 14592 14398 14638 14410
rect 14710 14786 14756 14798
rect 14710 14410 14716 14786
rect 14750 14410 14756 14786
rect 14710 14398 14756 14410
rect 14828 14786 14874 14798
rect 14828 14410 14834 14786
rect 14868 14437 14874 14786
rect 14945 14786 14991 14798
rect 14945 14610 14951 14786
rect 14985 14610 14991 14786
rect 14945 14603 14991 14610
rect 15063 14786 16770 14798
rect 15063 14610 15069 14786
rect 15103 14773 16770 14786
rect 15103 14610 15109 14773
rect 15353 14693 16770 14773
rect 15357 14692 16770 14693
rect 14945 14598 14994 14603
rect 15063 14598 15109 14610
rect 14951 14437 14994 14598
rect 14868 14410 14994 14437
rect 14828 14398 14994 14410
rect 14834 14394 14994 14398
rect 14499 14366 14572 14367
rect 14499 14361 14707 14366
rect 14499 14315 14511 14361
rect 14560 14360 14707 14361
rect 14560 14326 14657 14360
rect 14691 14326 14707 14360
rect 14560 14315 14707 14326
rect 14499 14310 14707 14315
rect 14759 14360 14825 14366
rect 14759 14326 14775 14360
rect 14809 14326 14825 14360
rect 14499 14309 14572 14310
rect 14759 14281 14825 14326
rect 14362 14273 14825 14281
rect 14362 14241 14826 14273
rect 14918 14257 14994 14394
rect 14362 13822 14408 14241
rect 14914 14197 14924 14257
rect 14986 14197 14996 14257
rect 14348 13768 14358 13822
rect 14415 13768 14425 13822
rect 16589 13784 16770 14692
rect 21246 14431 21252 14807
rect 21286 14431 21292 14807
rect 21246 14419 21292 14431
rect 21364 14807 21410 14819
rect 21364 14431 21370 14807
rect 21404 14431 21410 14807
rect 21364 14419 21410 14431
rect 21482 14807 21528 14819
rect 21482 14431 21488 14807
rect 21522 14458 21528 14807
rect 21599 14807 21645 14819
rect 21599 14631 21605 14807
rect 21639 14631 21645 14807
rect 21599 14624 21645 14631
rect 21717 14807 23396 14819
rect 21717 14631 21723 14807
rect 21757 14794 23396 14807
rect 21757 14631 21763 14794
rect 22007 14713 23396 14794
rect 21599 14619 21648 14624
rect 21717 14619 21763 14631
rect 21605 14458 21648 14619
rect 21522 14431 21648 14458
rect 21482 14419 21648 14431
rect 21488 14415 21648 14419
rect 21106 14387 21191 14389
rect 21106 14383 21361 14387
rect 21106 14335 21118 14383
rect 21179 14381 21361 14383
rect 21179 14347 21311 14381
rect 21345 14347 21361 14381
rect 21179 14335 21361 14347
rect 21106 14331 21361 14335
rect 21413 14381 21479 14387
rect 21413 14347 21429 14381
rect 21463 14347 21479 14381
rect 21106 14329 21191 14331
rect 21413 14301 21479 14347
rect 21207 14294 21479 14301
rect 21207 14293 21480 14294
rect 21207 14255 21220 14293
rect 21265 14262 21480 14293
rect 21572 14278 21648 14415
rect 21265 14255 21279 14262
rect 21207 14246 21279 14255
rect 21568 14218 21578 14278
rect 21640 14218 21650 14278
rect 23215 13852 23396 14713
rect 13539 13611 13618 13623
rect 11056 13560 11135 13572
rect 11056 13463 11062 13560
rect 10984 13443 11062 13463
rect 11129 13463 11135 13560
rect 13539 13497 13545 13611
rect 13612 13497 13618 13611
rect 14683 13613 14762 13625
rect 14683 13497 14689 13613
rect 14756 13497 14762 13613
rect 11129 13443 11204 13463
rect 10984 13335 11028 13443
rect 11160 13335 11204 13443
rect 12781 13401 12837 13409
rect 10984 13293 11204 13335
rect 11855 13393 12837 13401
rect 11855 13359 12797 13393
rect 12831 13359 12837 13393
rect 13500 13389 13510 13497
rect 13642 13434 13652 13497
rect 13642 13423 13654 13434
rect 13642 13389 13655 13423
rect 13911 13413 13967 13415
rect 11855 13343 12837 13359
rect 13510 13351 13655 13389
rect 11855 13342 12834 13343
rect 10588 13263 11565 13293
rect 10588 13157 10620 13263
rect 10824 13157 10856 13263
rect 11060 13157 11092 13263
rect 11296 13157 11328 13263
rect 11531 13157 11565 13263
rect 10581 13145 10627 13157
rect 10581 12969 10587 13145
rect 10621 12969 10627 13145
rect 10581 12957 10627 12969
rect 10699 13145 10745 13157
rect 10699 12969 10705 13145
rect 10739 12969 10745 13145
rect 10699 12957 10745 12969
rect 10817 13145 10863 13157
rect 10817 12969 10823 13145
rect 10857 12969 10863 13145
rect 10817 12957 10863 12969
rect 10935 13145 10981 13157
rect 10935 12969 10941 13145
rect 10975 12969 10981 13145
rect 10935 12957 10981 12969
rect 11053 13145 11099 13157
rect 11053 12969 11059 13145
rect 11093 12969 11099 13145
rect 11053 12957 11099 12969
rect 11171 13145 11217 13157
rect 11171 12969 11177 13145
rect 11211 12969 11217 13145
rect 11171 12957 11217 12969
rect 11289 13145 11335 13157
rect 11289 12969 11295 13145
rect 11329 12969 11335 13145
rect 11289 12957 11335 12969
rect 11407 13145 11453 13157
rect 11407 12969 11413 13145
rect 11447 12969 11453 13145
rect 11407 12957 11453 12969
rect 11525 13145 11571 13157
rect 11525 12969 11531 13145
rect 11565 12969 11571 13145
rect 11525 12957 11571 12969
rect 11643 13145 11689 13157
rect 11643 12969 11649 13145
rect 11683 12969 11689 13145
rect 11643 12957 11689 12969
rect 10704 12863 10740 12957
rect 10940 12863 10976 12957
rect 11176 12864 11212 12957
rect 11338 12909 11404 12916
rect 11338 12875 11354 12909
rect 11388 12875 11404 12909
rect 11338 12864 11404 12875
rect 11176 12863 11404 12864
rect 10704 12834 11404 12863
rect 10704 12833 11286 12834
rect 10824 12720 10858 12833
rect 11220 12792 11286 12833
rect 11220 12758 11236 12792
rect 11270 12758 11286 12792
rect 11220 12751 11286 12758
rect 11648 12752 11683 12957
rect 11855 12752 11922 13342
rect 13614 13319 13655 13351
rect 13901 13347 13911 13413
rect 13967 13347 13977 13413
rect 14647 13389 14657 13497
rect 14789 13434 14799 13497
rect 14789 13423 14801 13434
rect 14789 13389 14802 13423
rect 14657 13351 14802 13389
rect 14761 13323 14802 13351
rect 13030 13291 13300 13319
rect 12771 13225 12781 13291
rect 12847 13225 12857 13291
rect 13030 13229 13064 13291
rect 13266 13229 13300 13291
rect 13384 13291 13655 13319
rect 14172 13295 14442 13323
rect 13384 13229 13418 13291
rect 13620 13229 13655 13291
rect 13796 13279 13967 13295
rect 13796 13245 13927 13279
rect 13961 13245 13967 13279
rect 13796 13229 13967 13245
rect 14172 13233 14206 13295
rect 14408 13233 14442 13295
rect 14526 13295 14802 13323
rect 14526 13233 14560 13295
rect 14762 13233 14802 13295
rect 12906 13217 12952 13229
rect 12906 12841 12912 13217
rect 12946 12841 12952 13217
rect 12906 12829 12952 12841
rect 13024 13217 13070 13229
rect 13024 12841 13030 13217
rect 13064 12841 13070 13217
rect 13024 12829 13070 12841
rect 13142 13217 13188 13229
rect 13142 12841 13148 13217
rect 13182 12841 13188 13217
rect 13142 12829 13188 12841
rect 13260 13217 13306 13229
rect 13260 12841 13266 13217
rect 13300 12841 13306 13217
rect 13260 12829 13306 12841
rect 13378 13217 13424 13229
rect 13378 12841 13384 13217
rect 13418 12841 13424 13217
rect 13378 12829 13424 12841
rect 13496 13217 13542 13229
rect 13496 12841 13502 13217
rect 13536 12841 13542 13217
rect 13496 12829 13542 12841
rect 13614 13217 13660 13229
rect 13614 12841 13620 13217
rect 13654 12841 13660 13217
rect 13614 12829 13660 12841
rect 11648 12724 11922 12752
rect 11294 12720 11922 12724
rect 7533 12469 7760 12505
rect 7533 12362 7568 12469
rect 7694 12435 7760 12469
rect 7694 12401 7710 12435
rect 7744 12401 7760 12435
rect 8041 12493 8138 12508
rect 8041 12426 8098 12493
rect 7694 12395 7760 12401
rect 7935 12390 8204 12426
rect 7935 12362 7968 12390
rect 8171 12362 8204 12390
rect 8288 12362 8322 12508
rect 7409 12350 7455 12362
rect 7409 12174 7415 12350
rect 7449 12174 7455 12350
rect 7409 12162 7455 12174
rect 7527 12350 7573 12362
rect 7527 12174 7533 12350
rect 7567 12174 7573 12350
rect 7527 12162 7573 12174
rect 7645 12350 7691 12362
rect 7645 12174 7651 12350
rect 7685 12174 7691 12350
rect 7645 12162 7691 12174
rect 7763 12350 7809 12362
rect 7763 12174 7769 12350
rect 7803 12295 7809 12350
rect 7928 12350 7974 12362
rect 7928 12295 7934 12350
rect 7803 12207 7934 12295
rect 7803 12174 7809 12207
rect 7763 12162 7809 12174
rect 7928 12174 7934 12207
rect 7968 12174 7974 12350
rect 7928 12162 7974 12174
rect 8046 12350 8092 12362
rect 8046 12174 8052 12350
rect 8086 12174 8092 12350
rect 8046 12162 8092 12174
rect 8164 12350 8210 12362
rect 8164 12174 8170 12350
rect 8204 12174 8210 12350
rect 8164 12162 8210 12174
rect 8282 12350 8328 12362
rect 8282 12174 8288 12350
rect 8322 12174 8328 12350
rect 9940 12315 10120 12523
rect 10818 12708 10864 12720
rect 10818 12332 10824 12708
rect 10858 12332 10864 12708
rect 10818 12320 10864 12332
rect 10936 12708 10982 12720
rect 10936 12332 10942 12708
rect 10976 12332 10982 12708
rect 10936 12320 10982 12332
rect 11054 12708 11100 12720
rect 11054 12332 11060 12708
rect 11094 12356 11100 12708
rect 11171 12708 11217 12720
rect 11171 12532 11177 12708
rect 11211 12532 11217 12708
rect 11171 12520 11217 12532
rect 11289 12708 11922 12720
rect 11289 12532 11295 12708
rect 11329 12695 11922 12708
rect 12912 12787 12946 12829
rect 13148 12787 13182 12829
rect 12912 12759 13182 12787
rect 13266 12788 13300 12829
rect 13502 12788 13536 12829
rect 13266 12759 13536 12788
rect 12912 12711 12946 12759
rect 11329 12532 11335 12695
rect 12912 12681 12975 12711
rect 11289 12520 11335 12532
rect 12940 12589 12975 12681
rect 12940 12553 13167 12589
rect 13437 12578 13447 12675
rect 13546 12578 13556 12675
rect 13620 12646 13654 12829
rect 13620 12592 13729 12646
rect 11177 12404 11212 12520
rect 12940 12446 12975 12553
rect 13101 12519 13167 12553
rect 13101 12485 13117 12519
rect 13151 12485 13167 12519
rect 13448 12577 13545 12578
rect 13448 12510 13505 12577
rect 13101 12479 13167 12485
rect 13342 12474 13611 12510
rect 13342 12446 13375 12474
rect 13578 12446 13611 12474
rect 13695 12446 13729 12592
rect 12816 12434 12862 12446
rect 11308 12404 11416 12414
rect 11177 12356 11308 12404
rect 11416 12365 11561 12371
rect 11094 12332 11308 12356
rect 11054 12320 11308 12332
rect 11060 12316 11308 12320
rect 9940 12288 10696 12315
rect 9940 12282 10933 12288
rect 9940 12248 10883 12282
rect 10917 12248 10933 12282
rect 9940 12232 10933 12248
rect 10985 12282 11051 12288
rect 10985 12248 11001 12282
rect 11035 12248 11051 12282
rect 11234 12272 11308 12316
rect 11549 12298 11561 12365
rect 11416 12292 11561 12298
rect 11308 12262 11416 12272
rect 9940 12216 10696 12232
rect 9940 12215 10633 12216
rect 9940 12211 10168 12215
rect 8282 12162 8328 12174
rect 7415 12123 7449 12162
rect 7651 12123 7685 12162
rect 7415 12087 7685 12123
rect 8052 12124 8085 12162
rect 8288 12124 8321 12162
rect 8052 12088 8321 12124
rect 7415 12086 7581 12087
rect 7449 12007 7581 12086
rect 7439 11899 7449 12007
rect 7581 11899 7591 12007
rect 7472 11765 7478 11899
rect 7545 11765 7551 11899
rect 7472 11753 7551 11765
rect 9439 11800 9952 11832
rect 9439 11694 9800 11800
rect 9912 11787 9952 11800
rect 9912 11694 9954 11787
rect 9439 11683 9954 11694
rect 9439 11682 9952 11683
rect 4053 11525 5030 11555
rect 7247 11553 7310 11570
rect 7172 11549 7310 11553
rect 4053 11419 4085 11525
rect 4289 11419 4321 11525
rect 4525 11419 4557 11525
rect 4761 11419 4793 11525
rect 4996 11419 5030 11525
rect 5340 11515 7310 11549
rect 5338 11486 7310 11515
rect 5338 11470 5384 11486
rect 7172 11484 7310 11486
rect 4046 11407 4092 11419
rect 4046 11231 4052 11407
rect 4086 11231 4092 11407
rect 4046 11219 4092 11231
rect 4164 11407 4210 11419
rect 4164 11231 4170 11407
rect 4204 11231 4210 11407
rect 4164 11219 4210 11231
rect 4282 11407 4328 11419
rect 4282 11231 4288 11407
rect 4322 11231 4328 11407
rect 4282 11219 4328 11231
rect 4400 11407 4446 11419
rect 4400 11231 4406 11407
rect 4440 11231 4446 11407
rect 4400 11219 4446 11231
rect 4518 11407 4564 11419
rect 4518 11231 4524 11407
rect 4558 11231 4564 11407
rect 4518 11219 4564 11231
rect 4636 11407 4682 11419
rect 4636 11231 4642 11407
rect 4676 11231 4682 11407
rect 4636 11219 4682 11231
rect 4754 11407 4800 11419
rect 4754 11231 4760 11407
rect 4794 11231 4800 11407
rect 4754 11219 4800 11231
rect 4872 11407 4918 11419
rect 4872 11231 4878 11407
rect 4912 11231 4918 11407
rect 4872 11219 4918 11231
rect 4990 11407 5036 11419
rect 4990 11231 4996 11407
rect 5030 11231 5036 11407
rect 4990 11219 5036 11231
rect 5108 11407 5154 11419
rect 5108 11231 5114 11407
rect 5148 11231 5154 11407
rect 5108 11219 5154 11231
rect 4169 11125 4205 11219
rect 4405 11125 4441 11219
rect 4641 11126 4677 11219
rect 4803 11171 4869 11178
rect 4803 11137 4819 11171
rect 4853 11137 4869 11171
rect 4803 11126 4869 11137
rect 4641 11125 4869 11126
rect 4169 11096 4869 11125
rect 4169 11095 4751 11096
rect 4289 10982 4323 11095
rect 4685 11054 4751 11095
rect 4685 11020 4701 11054
rect 4735 11020 4751 11054
rect 4685 11013 4751 11020
rect 5113 11001 5148 11219
rect 5337 11018 5384 11470
rect 8231 11479 8310 11491
rect 8231 11362 8237 11479
rect 8304 11362 8310 11479
rect 6296 11254 6306 11362
rect 6438 11254 6448 11362
rect 8194 11254 8204 11362
rect 8336 11254 8346 11362
rect 6306 11214 6438 11254
rect 8204 11214 8336 11254
rect 6305 11148 6438 11214
rect 8203 11148 8336 11214
rect 5634 11105 7107 11148
rect 5337 11002 5383 11018
rect 5302 11001 5383 11002
rect 5113 10986 5383 11001
rect 4759 10982 5383 10986
rect 4283 10970 4329 10982
rect 4018 10492 4028 10610
rect 4146 10578 4156 10610
rect 4283 10594 4289 10970
rect 4323 10594 4329 10970
rect 4283 10582 4329 10594
rect 4401 10970 4447 10982
rect 4401 10594 4407 10970
rect 4441 10594 4447 10970
rect 4401 10582 4447 10594
rect 4519 10970 4565 10982
rect 4519 10594 4525 10970
rect 4559 10618 4565 10970
rect 4636 10970 4682 10982
rect 4636 10794 4642 10970
rect 4676 10794 4682 10970
rect 4636 10782 4682 10794
rect 4754 10970 5383 10982
rect 4754 10794 4760 10970
rect 4794 10958 5383 10970
rect 4794 10957 5036 10958
rect 4794 10794 4800 10957
rect 5302 10956 5383 10958
rect 5634 10802 5668 11105
rect 6000 11002 6034 11105
rect 6236 11002 6270 11105
rect 6472 11002 6506 11105
rect 6708 11002 6742 11105
rect 5994 10990 6040 11002
rect 4754 10782 4800 10794
rect 5510 10790 5556 10802
rect 4642 10666 4677 10782
rect 4773 10666 4881 10676
rect 4642 10618 4773 10666
rect 4881 10633 5030 10639
rect 4559 10594 4773 10618
rect 4519 10582 4773 10594
rect 4525 10578 4773 10582
rect 4146 10550 4161 10578
rect 4146 10544 4398 10550
rect 4146 10510 4348 10544
rect 4382 10510 4398 10544
rect 4146 10494 4398 10510
rect 4450 10544 4516 10550
rect 4450 10510 4466 10544
rect 4500 10510 4516 10544
rect 4699 10534 4773 10578
rect 5018 10566 5030 10633
rect 5510 10614 5516 10790
rect 5550 10614 5556 10790
rect 5510 10602 5556 10614
rect 5628 10790 5674 10802
rect 5628 10614 5634 10790
rect 5668 10614 5674 10790
rect 5628 10602 5674 10614
rect 5746 10790 5792 10802
rect 5746 10614 5752 10790
rect 5786 10614 5792 10790
rect 5746 10602 5792 10614
rect 5864 10790 5910 10802
rect 5994 10790 6000 10990
rect 5864 10614 5870 10790
rect 5904 10614 6000 10790
rect 6034 10614 6040 10990
rect 5864 10602 5910 10614
rect 5994 10602 6040 10614
rect 6112 10990 6158 11002
rect 6112 10614 6118 10990
rect 6152 10614 6158 10990
rect 6112 10602 6158 10614
rect 6230 10990 6276 11002
rect 6230 10614 6236 10990
rect 6270 10614 6276 10990
rect 6230 10602 6276 10614
rect 6348 10990 6394 11002
rect 6348 10614 6354 10990
rect 6388 10614 6394 10990
rect 6348 10602 6394 10614
rect 6466 10990 6512 11002
rect 6466 10614 6472 10990
rect 6506 10614 6512 10990
rect 6466 10602 6512 10614
rect 6584 10990 6630 11002
rect 6584 10614 6590 10990
rect 6624 10614 6630 10990
rect 6584 10602 6630 10614
rect 6702 10990 6748 11002
rect 6702 10614 6708 10990
rect 6742 10790 6748 10990
rect 7073 10802 7107 11105
rect 7532 11105 9005 11148
rect 7532 10802 7566 11105
rect 7898 11002 7932 11105
rect 8134 11002 8168 11105
rect 8370 11002 8404 11105
rect 8606 11002 8640 11105
rect 7892 10990 7938 11002
rect 6831 10790 6877 10802
rect 6742 10614 6837 10790
rect 6871 10614 6877 10790
rect 6702 10602 6748 10614
rect 6831 10602 6877 10614
rect 6949 10790 6995 10802
rect 6949 10614 6955 10790
rect 6989 10614 6995 10790
rect 6949 10602 6995 10614
rect 7067 10790 7113 10802
rect 7067 10614 7073 10790
rect 7107 10614 7113 10790
rect 7067 10602 7113 10614
rect 7185 10790 7231 10802
rect 7185 10614 7191 10790
rect 7225 10614 7231 10790
rect 7185 10602 7231 10614
rect 7408 10790 7454 10802
rect 7408 10614 7414 10790
rect 7448 10614 7454 10790
rect 7408 10602 7454 10614
rect 7526 10790 7572 10802
rect 7526 10614 7532 10790
rect 7566 10614 7572 10790
rect 7526 10602 7572 10614
rect 7644 10790 7690 10802
rect 7644 10614 7650 10790
rect 7684 10614 7690 10790
rect 7644 10602 7690 10614
rect 7762 10790 7808 10802
rect 7892 10790 7898 10990
rect 7762 10614 7768 10790
rect 7802 10614 7898 10790
rect 7932 10614 7938 10990
rect 7762 10602 7808 10614
rect 7892 10602 7938 10614
rect 8010 10990 8056 11002
rect 8010 10614 8016 10990
rect 8050 10614 8056 10990
rect 8010 10602 8056 10614
rect 8128 10990 8174 11002
rect 8128 10614 8134 10990
rect 8168 10614 8174 10990
rect 8128 10602 8174 10614
rect 8246 10990 8292 11002
rect 8246 10614 8252 10990
rect 8286 10614 8292 10990
rect 8246 10602 8292 10614
rect 8364 10990 8410 11002
rect 8364 10614 8370 10990
rect 8404 10614 8410 10990
rect 8364 10602 8410 10614
rect 8482 10990 8528 11002
rect 8482 10614 8488 10990
rect 8522 10614 8528 10990
rect 8482 10602 8528 10614
rect 8600 10990 8646 11002
rect 8600 10614 8606 10990
rect 8640 10790 8646 10990
rect 8971 10802 9005 11105
rect 8729 10790 8775 10802
rect 8640 10614 8735 10790
rect 8769 10614 8775 10790
rect 8600 10602 8646 10614
rect 8729 10602 8775 10614
rect 8847 10790 8893 10802
rect 8847 10614 8853 10790
rect 8887 10614 8893 10790
rect 8847 10602 8893 10614
rect 8965 10790 9011 10802
rect 8965 10614 8971 10790
rect 9005 10614 9011 10790
rect 8965 10602 9011 10614
rect 9083 10790 9129 10802
rect 9083 10614 9089 10790
rect 9123 10614 9129 10790
rect 9083 10602 9129 10614
rect 4881 10560 5030 10566
rect 5516 10568 5550 10602
rect 6118 10568 6152 10602
rect 6354 10568 6388 10602
rect 4773 10524 4881 10534
rect 5516 10533 5675 10568
rect 6118 10533 6388 10568
rect 6955 10568 6989 10602
rect 7191 10568 7225 10602
rect 6955 10533 7225 10568
rect 7414 10568 7448 10602
rect 8016 10568 8050 10602
rect 8252 10568 8286 10602
rect 7414 10533 7573 10568
rect 8016 10533 8286 10568
rect 8853 10568 8887 10602
rect 9089 10568 9123 10602
rect 8853 10533 9123 10568
rect 4146 10492 4161 10494
rect 4061 10478 4161 10492
rect 4061 10435 4161 10436
rect 3682 10414 4161 10435
rect 4450 10414 4516 10510
rect 3682 10366 4516 10414
rect 3682 10337 4161 10366
rect 3682 10335 3787 10337
rect 4061 10336 4161 10337
rect 3515 10150 3525 10229
rect 3618 10150 3628 10229
rect 4517 10215 4596 10227
rect 1724 10114 1773 10119
rect 1842 10114 1888 10126
rect 1730 9953 1773 10114
rect 1647 9926 1773 9953
rect 1607 9914 1773 9926
rect 1613 9910 1773 9914
rect 777 9876 1486 9882
rect 777 9842 1436 9876
rect 1470 9842 1486 9876
rect 777 9826 1486 9842
rect 1538 9876 1604 9882
rect 1538 9842 1554 9876
rect 1588 9842 1604 9876
rect 5 9788 272 9793
rect 5 9775 174 9788
rect 5 9694 20 9775
rect 114 9694 174 9775
rect 5 9684 174 9694
rect 261 9684 272 9788
rect 5 9678 272 9684
rect -666 7994 -656 8061
rect -589 7994 -579 8061
rect -3257 1874 -723 1940
rect -661 5987 -586 7994
rect -661 5933 -650 5987
rect -594 5933 -584 5987
rect -661 3919 -586 5933
rect 777 4136 882 9826
rect 1538 9797 1604 9842
rect 940 9789 1604 9797
rect 940 9783 1605 9789
rect 940 9687 971 9783
rect 1048 9757 1605 9783
rect 1697 9773 1773 9910
rect 1048 9687 1058 9757
rect 1693 9713 1703 9773
rect 1765 9713 1775 9773
rect 940 6896 1058 9687
rect 3526 8976 3619 10150
rect 4517 10121 4523 10215
rect 4444 10101 4523 10121
rect 4590 10121 4596 10215
rect 4590 10101 4664 10121
rect 4444 9993 4488 10101
rect 4620 9993 4664 10101
rect 4444 9951 4664 9993
rect 4048 9921 5025 9951
rect 4048 9815 4080 9921
rect 4284 9815 4316 9921
rect 4520 9815 4552 9921
rect 4756 9815 4788 9921
rect 4991 9815 5025 9921
rect 4041 9803 4087 9815
rect 4041 9627 4047 9803
rect 4081 9627 4087 9803
rect 4041 9615 4087 9627
rect 4159 9803 4205 9815
rect 4159 9627 4165 9803
rect 4199 9627 4205 9803
rect 4159 9615 4205 9627
rect 4277 9803 4323 9815
rect 4277 9627 4283 9803
rect 4317 9627 4323 9803
rect 4277 9615 4323 9627
rect 4395 9803 4441 9815
rect 4395 9627 4401 9803
rect 4435 9627 4441 9803
rect 4395 9615 4441 9627
rect 4513 9803 4559 9815
rect 4513 9627 4519 9803
rect 4553 9627 4559 9803
rect 4513 9615 4559 9627
rect 4631 9803 4677 9815
rect 4631 9627 4637 9803
rect 4671 9627 4677 9803
rect 4631 9615 4677 9627
rect 4749 9803 4795 9815
rect 4749 9627 4755 9803
rect 4789 9627 4795 9803
rect 4749 9615 4795 9627
rect 4867 9803 4913 9815
rect 4867 9627 4873 9803
rect 4907 9627 4913 9803
rect 4867 9615 4913 9627
rect 4985 9803 5031 9815
rect 4985 9627 4991 9803
rect 5025 9627 5031 9803
rect 4985 9615 5031 9627
rect 5103 9803 5149 9815
rect 5103 9627 5109 9803
rect 5143 9627 5149 9803
rect 5103 9615 5149 9627
rect 5641 9749 5675 10533
rect 6354 10471 6388 10533
rect 5943 10433 6685 10471
rect 5943 10309 5977 10433
rect 6179 10309 6213 10433
rect 6415 10309 6449 10433
rect 6651 10309 6685 10433
rect 6941 10326 6951 10392
rect 7014 10326 7024 10392
rect 5937 10297 5983 10309
rect 5937 9921 5943 10297
rect 5977 9921 5983 10297
rect 5937 9909 5983 9921
rect 6055 10297 6101 10309
rect 6055 9921 6061 10297
rect 6095 9921 6101 10297
rect 6055 9909 6101 9921
rect 6173 10297 6219 10309
rect 6173 9921 6179 10297
rect 6213 9921 6219 10297
rect 6173 9909 6219 9921
rect 6291 10297 6337 10309
rect 6291 9921 6297 10297
rect 6331 9921 6337 10297
rect 6291 9909 6337 9921
rect 6409 10297 6455 10309
rect 6409 9921 6415 10297
rect 6449 9921 6455 10297
rect 6409 9909 6455 9921
rect 6527 10297 6573 10309
rect 6527 9921 6533 10297
rect 6567 9921 6573 10297
rect 6527 9909 6573 9921
rect 6645 10297 6691 10309
rect 6645 9921 6651 10297
rect 6685 9921 6691 10297
rect 6645 9909 6691 9921
rect 7057 9750 7091 10533
rect 6784 9749 7091 9750
rect 5641 9744 5957 9749
rect 6671 9744 7091 9749
rect 5641 9733 6024 9744
rect 5641 9706 5973 9733
rect 4164 9521 4200 9615
rect 4400 9521 4436 9615
rect 4636 9522 4672 9615
rect 4798 9567 4864 9574
rect 4798 9533 4814 9567
rect 4848 9533 4864 9567
rect 4798 9522 4864 9533
rect 4636 9521 4864 9522
rect 4164 9492 4864 9521
rect 4164 9491 4746 9492
rect 4284 9378 4318 9491
rect 4680 9450 4746 9491
rect 4680 9416 4696 9450
rect 4730 9416 4746 9450
rect 4680 9409 4746 9416
rect 5108 9382 5143 9615
rect 5641 9577 5675 9706
rect 5957 9699 5973 9706
rect 6007 9699 6024 9733
rect 5957 9693 6024 9699
rect 6604 9733 7091 9744
rect 6604 9699 6621 9733
rect 6655 9706 7091 9733
rect 6655 9699 6671 9706
rect 6784 9705 7091 9706
rect 6604 9693 6671 9699
rect 5782 9666 5838 9678
rect 5782 9632 5788 9666
rect 5822 9665 5838 9666
rect 6895 9665 6951 9677
rect 5822 9649 6289 9665
rect 5822 9632 6239 9649
rect 5782 9616 6239 9632
rect 6223 9615 6239 9616
rect 6273 9615 6289 9649
rect 6223 9608 6289 9615
rect 6341 9650 6911 9665
rect 6341 9616 6357 9650
rect 6391 9631 6911 9650
rect 6945 9631 6951 9665
rect 6391 9616 6951 9631
rect 6341 9606 6408 9616
rect 6895 9615 6951 9616
rect 7057 9577 7091 9705
rect 7539 9749 7573 10533
rect 8252 10471 8286 10533
rect 7841 10433 8583 10471
rect 7841 10309 7875 10433
rect 8077 10309 8111 10433
rect 8313 10309 8347 10433
rect 8549 10309 8583 10433
rect 7835 10297 7881 10309
rect 7835 9921 7841 10297
rect 7875 9921 7881 10297
rect 7835 9909 7881 9921
rect 7953 10297 7999 10309
rect 7953 9921 7959 10297
rect 7993 9921 7999 10297
rect 7953 9909 7999 9921
rect 8071 10297 8117 10309
rect 8071 9921 8077 10297
rect 8111 9921 8117 10297
rect 8071 9909 8117 9921
rect 8189 10297 8235 10309
rect 8189 9921 8195 10297
rect 8229 9921 8235 10297
rect 8189 9909 8235 9921
rect 8307 10297 8353 10309
rect 8307 9921 8313 10297
rect 8347 9921 8353 10297
rect 8307 9909 8353 9921
rect 8425 10297 8471 10309
rect 8425 9921 8431 10297
rect 8465 9921 8471 10297
rect 8425 9909 8471 9921
rect 8543 10297 8589 10309
rect 8543 9921 8549 10297
rect 8583 9921 8589 10297
rect 8543 9909 8589 9921
rect 8955 9750 8989 10533
rect 8567 9749 8636 9750
rect 8682 9749 8989 9750
rect 7539 9744 7855 9749
rect 8567 9745 8989 9749
rect 7539 9733 7922 9744
rect 7539 9706 7871 9733
rect 7539 9577 7573 9706
rect 7855 9699 7871 9706
rect 7905 9699 7922 9733
rect 7855 9693 7922 9699
rect 8500 9734 8989 9745
rect 8500 9700 8517 9734
rect 8551 9706 8989 9734
rect 8551 9700 8567 9706
rect 8682 9705 8989 9706
rect 8500 9694 8567 9700
rect 7680 9666 7736 9678
rect 7680 9632 7686 9666
rect 7720 9665 7736 9666
rect 8793 9665 8849 9677
rect 7720 9649 8187 9665
rect 7720 9632 8137 9649
rect 7680 9616 8137 9632
rect 8121 9615 8137 9616
rect 8171 9615 8187 9649
rect 8121 9608 8187 9615
rect 8239 9650 8809 9665
rect 8239 9616 8255 9650
rect 8289 9631 8809 9650
rect 8843 9631 8849 9665
rect 8289 9616 8849 9631
rect 8239 9606 8306 9616
rect 8793 9615 8849 9616
rect 8955 9577 8989 9705
rect 9070 10355 9137 10379
rect 9070 10321 9087 10355
rect 9121 10321 9137 10355
rect 4754 9378 5143 9382
rect 4278 9366 4324 9378
rect 4278 8990 4284 9366
rect 4318 8990 4324 9366
rect 4278 8978 4324 8990
rect 4396 9366 4442 9378
rect 4396 8990 4402 9366
rect 4436 8990 4442 9366
rect 4396 8978 4442 8990
rect 4514 9366 4560 9378
rect 4514 8990 4520 9366
rect 4554 9014 4560 9366
rect 4631 9366 4677 9378
rect 4631 9190 4637 9366
rect 4671 9190 4677 9366
rect 4631 9178 4677 9190
rect 4749 9366 5143 9378
rect 5635 9565 5681 9577
rect 5635 9389 5641 9565
rect 5675 9389 5681 9565
rect 5635 9377 5681 9389
rect 5753 9565 5799 9577
rect 5753 9389 5759 9565
rect 5793 9389 5799 9565
rect 5753 9377 5799 9389
rect 6055 9565 6101 9577
rect 4749 9190 4755 9366
rect 4789 9353 5143 9366
rect 4789 9190 4795 9353
rect 5065 9350 5143 9353
rect 5065 9298 5075 9350
rect 5138 9298 5148 9350
rect 5070 9292 5143 9298
rect 4749 9178 4795 9190
rect 4637 9062 4672 9178
rect 5758 9083 5792 9377
rect 6055 9189 6061 9565
rect 6095 9189 6101 9565
rect 6055 9177 6101 9189
rect 6173 9565 6219 9577
rect 6173 9189 6179 9565
rect 6213 9189 6219 9565
rect 6173 9177 6219 9189
rect 6291 9565 6337 9577
rect 6291 9189 6297 9565
rect 6331 9189 6337 9565
rect 6291 9177 6337 9189
rect 6409 9565 6455 9577
rect 6409 9189 6415 9565
rect 6449 9189 6455 9565
rect 6409 9177 6455 9189
rect 6527 9565 6573 9577
rect 6527 9189 6533 9565
rect 6567 9189 6573 9565
rect 6933 9565 6979 9577
rect 6933 9389 6939 9565
rect 6973 9389 6979 9565
rect 6933 9377 6979 9389
rect 7051 9565 7097 9577
rect 7051 9389 7057 9565
rect 7091 9389 7097 9565
rect 7051 9377 7097 9389
rect 7533 9565 7579 9577
rect 7533 9389 7539 9565
rect 7573 9389 7579 9565
rect 7533 9377 7579 9389
rect 7651 9565 7697 9577
rect 7651 9389 7657 9565
rect 7691 9389 7697 9565
rect 7651 9377 7697 9389
rect 7953 9565 7999 9577
rect 6527 9177 6573 9189
rect 6415 9083 6449 9177
rect 6939 9083 6972 9377
rect 4768 9062 4876 9072
rect 4637 9014 4768 9062
rect 5758 9051 6972 9083
rect 7656 9083 7690 9377
rect 7953 9189 7959 9565
rect 7993 9189 7999 9565
rect 7953 9177 7999 9189
rect 8071 9565 8117 9577
rect 8071 9189 8077 9565
rect 8111 9189 8117 9565
rect 8071 9177 8117 9189
rect 8189 9565 8235 9577
rect 8189 9189 8195 9565
rect 8229 9189 8235 9565
rect 8189 9177 8235 9189
rect 8307 9565 8353 9577
rect 8307 9189 8313 9565
rect 8347 9189 8353 9565
rect 8307 9177 8353 9189
rect 8425 9565 8471 9577
rect 8425 9189 8431 9565
rect 8465 9189 8471 9565
rect 8831 9565 8877 9577
rect 8831 9389 8837 9565
rect 8871 9389 8877 9565
rect 8831 9377 8877 9389
rect 8949 9565 8995 9577
rect 8949 9389 8955 9565
rect 8989 9389 8995 9565
rect 8949 9377 8995 9389
rect 8425 9177 8471 9189
rect 8313 9083 8347 9177
rect 8837 9083 8870 9377
rect 7656 9051 8870 9083
rect 4876 9025 5028 9031
rect 4554 8990 4768 9014
rect 4514 8978 4768 8990
rect 3526 8974 4111 8976
rect 4520 8974 4768 8978
rect 3526 8946 4156 8974
rect 3526 8940 4393 8946
rect 3526 8906 4343 8940
rect 4377 8906 4393 8940
rect 3526 8890 4393 8906
rect 4445 8940 4511 8946
rect 4445 8906 4461 8940
rect 4495 8906 4511 8940
rect 4694 8930 4768 8974
rect 5016 8958 5028 9025
rect 6251 8966 6383 9051
rect 8149 8966 8281 9051
rect 4876 8952 5028 8958
rect 4768 8920 4876 8930
rect 3526 8874 4156 8890
rect 3526 8870 4111 8874
rect 3526 8869 3627 8870
rect 4056 8821 4156 8832
rect 4020 8715 4030 8821
rect 4142 8810 4156 8821
rect 4445 8810 4511 8906
rect 6241 8858 6251 8966
rect 6383 8858 6393 8966
rect 8139 8858 8149 8966
rect 8281 8858 8291 8966
rect 9070 8938 9137 10321
rect 4142 8762 4511 8810
rect 4142 8732 4156 8762
rect 4142 8715 4152 8732
rect 4444 8659 4510 8762
rect 6274 8723 6280 8858
rect 6347 8723 6353 8858
rect 6274 8711 6353 8723
rect 9070 8659 9136 8938
rect 4442 8579 9136 8659
rect 6975 7747 7054 7759
rect 1426 7699 1562 7719
rect 1426 7637 1462 7699
rect 1522 7637 1562 7699
rect 1426 7609 1562 7637
rect 4495 7692 4574 7704
rect 1122 7579 2099 7609
rect 4495 7595 4501 7692
rect 1122 7473 1154 7579
rect 1358 7473 1390 7579
rect 1594 7473 1626 7579
rect 1830 7473 1862 7579
rect 2065 7473 2099 7579
rect 4427 7575 4501 7595
rect 4568 7595 4574 7692
rect 6975 7629 6981 7747
rect 7048 7629 7054 7747
rect 8131 7744 8210 7756
rect 8131 7629 8137 7744
rect 8204 7629 8210 7744
rect 4568 7575 4647 7595
rect 1115 7461 1161 7473
rect 1115 7285 1121 7461
rect 1155 7285 1161 7461
rect 1115 7273 1161 7285
rect 1233 7461 1279 7473
rect 1233 7285 1239 7461
rect 1273 7285 1279 7461
rect 1233 7273 1279 7285
rect 1351 7461 1397 7473
rect 1351 7285 1357 7461
rect 1391 7285 1397 7461
rect 1351 7273 1397 7285
rect 1469 7461 1515 7473
rect 1469 7285 1475 7461
rect 1509 7285 1515 7461
rect 1469 7273 1515 7285
rect 1587 7461 1633 7473
rect 1587 7285 1593 7461
rect 1627 7285 1633 7461
rect 1587 7273 1633 7285
rect 1705 7461 1751 7473
rect 1705 7285 1711 7461
rect 1745 7285 1751 7461
rect 1705 7273 1751 7285
rect 1823 7461 1869 7473
rect 1823 7285 1829 7461
rect 1863 7285 1869 7461
rect 1823 7273 1869 7285
rect 1941 7461 1987 7473
rect 1941 7285 1947 7461
rect 1981 7285 1987 7461
rect 1941 7273 1987 7285
rect 2059 7461 2105 7473
rect 2059 7285 2065 7461
rect 2099 7285 2105 7461
rect 2059 7273 2105 7285
rect 2177 7461 2223 7473
rect 2177 7285 2183 7461
rect 2217 7285 2223 7461
rect 4427 7467 4471 7575
rect 4603 7467 4647 7575
rect 6224 7533 6280 7541
rect 4427 7425 4647 7467
rect 5298 7525 6280 7533
rect 5298 7491 6240 7525
rect 6274 7491 6280 7525
rect 6943 7521 6953 7629
rect 7085 7566 7095 7629
rect 7085 7555 7097 7566
rect 7085 7521 7098 7555
rect 7354 7545 7410 7547
rect 5298 7475 6280 7491
rect 6953 7483 7098 7521
rect 5298 7474 6277 7475
rect 4031 7395 5008 7425
rect 4031 7289 4063 7395
rect 4267 7289 4299 7395
rect 4503 7289 4535 7395
rect 4739 7289 4771 7395
rect 4974 7289 5008 7395
rect 2177 7273 2223 7285
rect 4024 7277 4070 7289
rect 1238 7179 1274 7273
rect 1474 7179 1510 7273
rect 1710 7180 1746 7273
rect 1872 7225 1938 7232
rect 1872 7191 1888 7225
rect 1922 7191 1938 7225
rect 1872 7180 1938 7191
rect 1710 7179 1938 7180
rect 1238 7150 1938 7179
rect 1238 7149 1820 7150
rect 1358 7036 1392 7149
rect 1754 7108 1820 7149
rect 1754 7074 1770 7108
rect 1804 7074 1820 7108
rect 1754 7067 1820 7074
rect 2182 7040 2217 7273
rect 4024 7101 4030 7277
rect 4064 7101 4070 7277
rect 4024 7089 4070 7101
rect 4142 7277 4188 7289
rect 4142 7101 4148 7277
rect 4182 7101 4188 7277
rect 4142 7089 4188 7101
rect 4260 7277 4306 7289
rect 4260 7101 4266 7277
rect 4300 7101 4306 7277
rect 4260 7089 4306 7101
rect 4378 7277 4424 7289
rect 4378 7101 4384 7277
rect 4418 7101 4424 7277
rect 4378 7089 4424 7101
rect 4496 7277 4542 7289
rect 4496 7101 4502 7277
rect 4536 7101 4542 7277
rect 4496 7089 4542 7101
rect 4614 7277 4660 7289
rect 4614 7101 4620 7277
rect 4654 7101 4660 7277
rect 4614 7089 4660 7101
rect 4732 7277 4778 7289
rect 4732 7101 4738 7277
rect 4772 7101 4778 7277
rect 4732 7089 4778 7101
rect 4850 7277 4896 7289
rect 4850 7101 4856 7277
rect 4890 7101 4896 7277
rect 4850 7089 4896 7101
rect 4968 7277 5014 7289
rect 4968 7101 4974 7277
rect 5008 7101 5014 7277
rect 4968 7089 5014 7101
rect 5086 7277 5132 7289
rect 5086 7101 5092 7277
rect 5126 7101 5132 7277
rect 5086 7089 5132 7101
rect 1828 7036 2217 7040
rect 1352 7024 1398 7036
rect 940 6796 1312 6896
rect 1236 6604 1290 6796
rect 1352 6648 1358 7024
rect 1392 6648 1398 7024
rect 1352 6636 1398 6648
rect 1470 7024 1516 7036
rect 1470 6648 1476 7024
rect 1510 6648 1516 7024
rect 1470 6636 1516 6648
rect 1588 7024 1634 7036
rect 1588 6648 1594 7024
rect 1628 6675 1634 7024
rect 1705 7024 1751 7036
rect 1705 6848 1711 7024
rect 1745 6848 1751 7024
rect 1705 6841 1751 6848
rect 1823 7024 2217 7036
rect 1823 6848 1829 7024
rect 1863 7015 2217 7024
rect 1863 7011 2219 7015
rect 1863 6848 1869 7011
rect 1705 6836 1754 6841
rect 1823 6836 1869 6848
rect 1711 6675 1754 6836
rect 1628 6648 1754 6675
rect 1588 6636 1754 6648
rect 1594 6632 1754 6636
rect 1236 6598 1467 6604
rect 1236 6564 1417 6598
rect 1451 6564 1467 6598
rect 1236 6548 1467 6564
rect 1519 6598 1585 6604
rect 1519 6564 1535 6598
rect 1569 6564 1585 6598
rect 1071 6527 1155 6533
rect 1071 6474 1083 6527
rect 1143 6519 1155 6527
rect 1519 6519 1585 6564
rect 1143 6511 1585 6519
rect 1143 6479 1586 6511
rect 1678 6495 1754 6632
rect 2112 6535 2219 7011
rect 4147 6995 4183 7089
rect 4383 6995 4419 7089
rect 4619 6996 4655 7089
rect 4781 7041 4847 7048
rect 4781 7007 4797 7041
rect 4831 7007 4847 7041
rect 4781 6996 4847 7007
rect 4619 6995 4847 6996
rect 4147 6966 4847 6995
rect 4147 6965 4729 6966
rect 4267 6852 4301 6965
rect 4663 6924 4729 6965
rect 4663 6890 4679 6924
rect 4713 6890 4729 6924
rect 4663 6883 4729 6890
rect 5091 6884 5126 7089
rect 5298 6884 5365 7474
rect 7057 7451 7098 7483
rect 7344 7479 7354 7545
rect 7410 7479 7420 7545
rect 8090 7521 8100 7629
rect 8232 7566 8242 7629
rect 8232 7555 8244 7566
rect 8232 7521 8245 7555
rect 8100 7483 8245 7521
rect 8204 7455 8245 7483
rect 6473 7423 6743 7451
rect 6214 7357 6224 7423
rect 6290 7357 6300 7423
rect 6473 7361 6507 7423
rect 6709 7361 6743 7423
rect 6827 7423 7098 7451
rect 7615 7427 7885 7455
rect 6827 7361 6861 7423
rect 7063 7361 7098 7423
rect 7239 7411 7410 7427
rect 7239 7377 7370 7411
rect 7404 7377 7410 7411
rect 7239 7361 7410 7377
rect 7615 7365 7649 7427
rect 7851 7365 7885 7427
rect 7969 7427 8245 7455
rect 7969 7365 8003 7427
rect 8205 7365 8245 7427
rect 6349 7349 6395 7361
rect 6349 6973 6355 7349
rect 6389 6973 6395 7349
rect 6349 6961 6395 6973
rect 6467 7349 6513 7361
rect 6467 6973 6473 7349
rect 6507 6973 6513 7349
rect 6467 6961 6513 6973
rect 6585 7349 6631 7361
rect 6585 6973 6591 7349
rect 6625 6973 6631 7349
rect 6585 6961 6631 6973
rect 6703 7349 6749 7361
rect 6703 6973 6709 7349
rect 6743 6973 6749 7349
rect 6703 6961 6749 6973
rect 6821 7349 6867 7361
rect 6821 6973 6827 7349
rect 6861 6973 6867 7349
rect 6821 6961 6867 6973
rect 6939 7349 6985 7361
rect 6939 6973 6945 7349
rect 6979 6973 6985 7349
rect 6939 6961 6985 6973
rect 7057 7349 7103 7361
rect 7057 6973 7063 7349
rect 7097 6973 7103 7349
rect 7057 6961 7103 6973
rect 5091 6856 5365 6884
rect 4737 6852 5365 6856
rect 1143 6474 1155 6479
rect 1071 6468 1155 6474
rect 1674 6435 1684 6495
rect 1746 6435 1756 6495
rect 2111 6447 2219 6535
rect 4261 6840 4307 6852
rect 4261 6464 4267 6840
rect 4301 6464 4307 6840
rect 4261 6452 4307 6464
rect 4379 6840 4425 6852
rect 4379 6464 4385 6840
rect 4419 6464 4425 6840
rect 4379 6452 4425 6464
rect 4497 6840 4543 6852
rect 4497 6464 4503 6840
rect 4537 6488 4543 6840
rect 4614 6840 4660 6852
rect 4614 6664 4620 6840
rect 4654 6664 4660 6840
rect 4614 6652 4660 6664
rect 4732 6840 5365 6852
rect 4732 6664 4738 6840
rect 4772 6827 5365 6840
rect 6355 6919 6389 6961
rect 6591 6919 6625 6961
rect 6355 6891 6625 6919
rect 6709 6920 6743 6961
rect 6945 6920 6979 6961
rect 6709 6891 6979 6920
rect 6355 6843 6389 6891
rect 4772 6664 4778 6827
rect 6355 6813 6418 6843
rect 4732 6652 4778 6664
rect 6383 6721 6418 6813
rect 6383 6685 6610 6721
rect 6880 6710 6890 6807
rect 6989 6710 6999 6807
rect 7063 6778 7097 6961
rect 7063 6724 7172 6778
rect 4620 6536 4655 6652
rect 6383 6578 6418 6685
rect 6544 6651 6610 6685
rect 6544 6617 6560 6651
rect 6594 6617 6610 6651
rect 6891 6709 6988 6710
rect 6891 6642 6948 6709
rect 6544 6611 6610 6617
rect 6785 6606 7054 6642
rect 6785 6578 6818 6606
rect 7021 6578 7054 6606
rect 7138 6578 7172 6724
rect 6259 6566 6305 6578
rect 4751 6536 4859 6546
rect 4620 6488 4751 6536
rect 4859 6496 5005 6502
rect 4537 6464 4751 6488
rect 4497 6452 4751 6464
rect 4503 6448 4751 6452
rect 2111 6420 4139 6447
rect 2111 6414 4376 6420
rect 2111 6380 4326 6414
rect 4360 6380 4376 6414
rect 2111 6364 4376 6380
rect 4428 6414 4494 6420
rect 4428 6380 4444 6414
rect 4478 6380 4494 6414
rect 4677 6404 4751 6448
rect 4993 6429 5005 6496
rect 4859 6423 5005 6429
rect 4751 6394 4859 6404
rect 2111 6348 4139 6364
rect 2111 6347 4076 6348
rect 2111 6346 3611 6347
rect 3106 5959 3395 5960
rect 2610 5958 3395 5959
rect 2427 5932 3395 5958
rect 2427 5826 3243 5932
rect 3355 5919 3395 5932
rect 3355 5826 3397 5919
rect 2427 5815 3397 5826
rect 2427 5814 3395 5815
rect 1442 4939 1578 4959
rect 1442 4877 1478 4939
rect 1538 4877 1578 4939
rect 1442 4849 1578 4877
rect 1138 4819 2115 4849
rect 1138 4713 1170 4819
rect 1374 4713 1406 4819
rect 1610 4713 1642 4819
rect 1846 4713 1878 4819
rect 2081 4713 2115 4819
rect 1131 4701 1177 4713
rect 1131 4525 1137 4701
rect 1171 4525 1177 4701
rect 1131 4513 1177 4525
rect 1249 4701 1295 4713
rect 1249 4525 1255 4701
rect 1289 4525 1295 4701
rect 1249 4513 1295 4525
rect 1367 4701 1413 4713
rect 1367 4525 1373 4701
rect 1407 4525 1413 4701
rect 1367 4513 1413 4525
rect 1485 4701 1531 4713
rect 1485 4525 1491 4701
rect 1525 4525 1531 4701
rect 1485 4513 1531 4525
rect 1603 4701 1649 4713
rect 1603 4525 1609 4701
rect 1643 4525 1649 4701
rect 1603 4513 1649 4525
rect 1721 4701 1767 4713
rect 1721 4525 1727 4701
rect 1761 4525 1767 4701
rect 1721 4513 1767 4525
rect 1839 4701 1885 4713
rect 1839 4525 1845 4701
rect 1879 4525 1885 4701
rect 1839 4513 1885 4525
rect 1957 4701 2003 4713
rect 1957 4525 1963 4701
rect 1997 4525 2003 4701
rect 1957 4513 2003 4525
rect 2075 4701 2121 4713
rect 2075 4525 2081 4701
rect 2115 4525 2121 4701
rect 2075 4513 2121 4525
rect 2193 4701 2239 4713
rect 2193 4525 2199 4701
rect 2233 4525 2239 4701
rect 2193 4513 2239 4525
rect 1254 4419 1290 4513
rect 1490 4419 1526 4513
rect 1726 4420 1762 4513
rect 1888 4465 1954 4472
rect 1888 4431 1904 4465
rect 1938 4431 1954 4465
rect 1888 4420 1954 4431
rect 1726 4419 1954 4420
rect 1254 4390 1954 4419
rect 1254 4389 1836 4390
rect 1374 4276 1408 4389
rect 1770 4348 1836 4389
rect 1770 4314 1786 4348
rect 1820 4314 1836 4348
rect 1770 4307 1836 4314
rect 2198 4280 2233 4513
rect 2427 4280 2550 5814
rect 3518 4449 3611 6346
rect 3674 6284 4140 6306
rect 4428 6284 4494 6380
rect 6259 6390 6265 6566
rect 6299 6390 6305 6566
rect 6259 6378 6305 6390
rect 6377 6566 6423 6578
rect 6377 6390 6383 6566
rect 6417 6390 6423 6566
rect 6377 6378 6423 6390
rect 6495 6566 6541 6578
rect 6495 6390 6501 6566
rect 6535 6390 6541 6566
rect 6495 6378 6541 6390
rect 6613 6566 6659 6578
rect 6613 6390 6619 6566
rect 6653 6511 6659 6566
rect 6778 6566 6824 6578
rect 6778 6511 6784 6566
rect 6653 6423 6784 6511
rect 6653 6390 6659 6423
rect 6613 6378 6659 6390
rect 6778 6390 6784 6423
rect 6818 6390 6824 6566
rect 6778 6378 6824 6390
rect 6896 6566 6942 6578
rect 6896 6390 6902 6566
rect 6936 6390 6942 6566
rect 6896 6378 6942 6390
rect 7014 6566 7060 6578
rect 7014 6390 7020 6566
rect 7054 6390 7060 6566
rect 7014 6378 7060 6390
rect 7132 6566 7178 6578
rect 7132 6390 7138 6566
rect 7172 6390 7178 6566
rect 7132 6378 7178 6390
rect 6265 6339 6299 6378
rect 6501 6339 6535 6378
rect 6265 6304 6535 6339
rect 6902 6340 6935 6378
rect 7138 6340 7171 6378
rect 6902 6304 7171 6340
rect 3674 6236 4494 6284
rect 6299 6303 6535 6304
rect 3674 6205 4140 6236
rect 6299 6229 6431 6303
rect 3674 5949 3779 6205
rect 6289 6121 6299 6229
rect 6431 6121 6441 6229
rect 4516 6039 4595 6051
rect 3674 5843 3737 5949
rect 3849 5843 3859 5949
rect 4516 5945 4522 6039
rect 4441 5925 4522 5945
rect 4589 5945 4595 6039
rect 6315 5986 6321 6121
rect 6388 5986 6394 6121
rect 6315 5974 6394 5986
rect 4589 5925 4661 5945
rect 3674 5832 3823 5843
rect 3674 4655 3779 5832
rect 4441 5817 4485 5925
rect 4617 5817 4661 5925
rect 4441 5775 4661 5817
rect 7239 5790 7301 7361
rect 7491 7353 7537 7365
rect 7491 6977 7497 7353
rect 7531 6977 7537 7353
rect 7491 6965 7537 6977
rect 7609 7353 7655 7365
rect 7609 6977 7615 7353
rect 7649 6977 7655 7353
rect 7609 6965 7655 6977
rect 7727 7353 7773 7365
rect 7727 6977 7733 7353
rect 7767 6977 7773 7353
rect 7727 6965 7773 6977
rect 7845 7353 7891 7365
rect 7845 6977 7851 7353
rect 7885 6977 7891 7353
rect 7845 6965 7891 6977
rect 7963 7353 8009 7365
rect 7963 6977 7969 7353
rect 8003 6977 8009 7353
rect 7963 6965 8009 6977
rect 8081 7353 8127 7365
rect 8081 6977 8087 7353
rect 8121 6977 8127 7353
rect 8081 6965 8127 6977
rect 8199 7353 8245 7365
rect 8199 6977 8205 7353
rect 8239 6977 8245 7353
rect 8199 6965 8245 6977
rect 7497 6923 7531 6965
rect 7733 6923 7767 6965
rect 7497 6895 7767 6923
rect 7851 6924 7885 6965
rect 8087 6924 8121 6965
rect 7851 6895 8121 6924
rect 7497 6847 7531 6895
rect 7497 6817 7560 6847
rect 7525 6725 7560 6817
rect 8032 6787 8132 6808
rect 8032 6733 8046 6787
rect 8111 6733 8132 6787
rect 8032 6728 8132 6733
rect 8205 6782 8239 6965
rect 9439 6797 9551 11682
rect 10075 10317 10168 12211
rect 10231 12152 10697 12174
rect 10985 12152 11051 12248
rect 12816 12258 12822 12434
rect 12856 12258 12862 12434
rect 12816 12246 12862 12258
rect 12934 12434 12980 12446
rect 12934 12258 12940 12434
rect 12974 12258 12980 12434
rect 12934 12246 12980 12258
rect 13052 12434 13098 12446
rect 13052 12258 13058 12434
rect 13092 12258 13098 12434
rect 13052 12246 13098 12258
rect 13170 12434 13216 12446
rect 13170 12258 13176 12434
rect 13210 12379 13216 12434
rect 13335 12434 13381 12446
rect 13335 12379 13341 12434
rect 13210 12291 13341 12379
rect 13210 12258 13216 12291
rect 13170 12246 13216 12258
rect 13335 12258 13341 12291
rect 13375 12258 13381 12434
rect 13335 12246 13381 12258
rect 13453 12434 13499 12446
rect 13453 12258 13459 12434
rect 13493 12258 13499 12434
rect 13453 12246 13499 12258
rect 13571 12434 13617 12446
rect 13571 12258 13577 12434
rect 13611 12258 13617 12434
rect 13571 12246 13617 12258
rect 13689 12434 13735 12446
rect 13689 12258 13695 12434
rect 13729 12258 13735 12434
rect 13689 12246 13735 12258
rect 12822 12207 12856 12246
rect 13058 12207 13092 12246
rect 12822 12172 13092 12207
rect 13459 12208 13492 12246
rect 13695 12208 13728 12246
rect 13459 12172 13728 12208
rect 10231 12104 11051 12152
rect 12856 12171 13092 12172
rect 10231 12073 10697 12104
rect 12856 12097 12988 12171
rect 10231 11817 10336 12073
rect 12846 11989 12856 12097
rect 12988 11989 12998 12097
rect 11070 11908 11149 11920
rect 10231 11711 10294 11817
rect 10406 11711 10416 11817
rect 11070 11813 11076 11908
rect 10998 11793 11076 11813
rect 11143 11813 11149 11908
rect 12879 11859 12885 11989
rect 12952 11859 12958 11989
rect 12879 11847 12958 11859
rect 11143 11793 11218 11813
rect 10231 11700 10380 11711
rect 10231 10523 10336 11700
rect 10998 11685 11042 11793
rect 11174 11685 11218 11793
rect 10998 11643 11218 11685
rect 13796 11658 13858 13229
rect 14048 13221 14094 13233
rect 14048 12845 14054 13221
rect 14088 12845 14094 13221
rect 14048 12833 14094 12845
rect 14166 13221 14212 13233
rect 14166 12845 14172 13221
rect 14206 12845 14212 13221
rect 14166 12833 14212 12845
rect 14284 13221 14330 13233
rect 14284 12845 14290 13221
rect 14324 12845 14330 13221
rect 14284 12833 14330 12845
rect 14402 13221 14448 13233
rect 14402 12845 14408 13221
rect 14442 12845 14448 13221
rect 14402 12833 14448 12845
rect 14520 13221 14566 13233
rect 14520 12845 14526 13221
rect 14560 12845 14566 13221
rect 14520 12833 14566 12845
rect 14638 13221 14684 13233
rect 14638 12845 14644 13221
rect 14678 12845 14684 13221
rect 14638 12833 14684 12845
rect 14756 13221 14802 13233
rect 14756 12845 14762 13221
rect 14796 12845 14802 13221
rect 14756 12833 14802 12845
rect 14054 12791 14088 12833
rect 14290 12791 14324 12833
rect 14054 12763 14324 12791
rect 14408 12792 14442 12833
rect 14644 12792 14678 12833
rect 14408 12763 14678 12792
rect 14054 12715 14088 12763
rect 14054 12685 14117 12715
rect 14082 12593 14117 12685
rect 14589 12655 14689 12676
rect 14589 12601 14603 12655
rect 14668 12601 14689 12655
rect 14589 12596 14689 12601
rect 14762 12650 14796 12833
rect 14762 12596 14871 12650
rect 14082 12557 14309 12593
rect 14082 12450 14117 12557
rect 14243 12523 14309 12557
rect 14243 12489 14259 12523
rect 14293 12489 14309 12523
rect 14590 12581 14687 12596
rect 14590 12514 14647 12581
rect 14243 12483 14309 12489
rect 14484 12478 14753 12514
rect 14484 12450 14517 12478
rect 14720 12450 14753 12478
rect 14837 12450 14871 12596
rect 15688 12589 15698 12664
rect 15766 12589 16160 12664
rect 15715 12588 16160 12589
rect 13958 12438 14004 12450
rect 13958 12262 13964 12438
rect 13998 12262 14004 12438
rect 13958 12250 14004 12262
rect 14076 12438 14122 12450
rect 14076 12262 14082 12438
rect 14116 12262 14122 12438
rect 14076 12250 14122 12262
rect 14194 12438 14240 12450
rect 14194 12262 14200 12438
rect 14234 12262 14240 12438
rect 14194 12250 14240 12262
rect 14312 12438 14358 12450
rect 14312 12262 14318 12438
rect 14352 12383 14358 12438
rect 14477 12438 14523 12450
rect 14477 12383 14483 12438
rect 14352 12295 14483 12383
rect 14352 12262 14358 12295
rect 14312 12250 14358 12262
rect 14477 12262 14483 12295
rect 14517 12262 14523 12438
rect 14477 12250 14523 12262
rect 14595 12438 14641 12450
rect 14595 12262 14601 12438
rect 14635 12262 14641 12438
rect 14595 12250 14641 12262
rect 14713 12438 14759 12450
rect 14713 12262 14719 12438
rect 14753 12262 14759 12438
rect 14713 12250 14759 12262
rect 14831 12438 14877 12450
rect 14831 12262 14837 12438
rect 14871 12262 14877 12438
rect 14831 12250 14877 12262
rect 13964 12211 13998 12250
rect 14200 12211 14234 12250
rect 13964 12175 14234 12211
rect 14601 12212 14634 12250
rect 14837 12212 14870 12250
rect 14601 12176 14870 12212
rect 13964 12174 14130 12175
rect 13998 12095 14130 12174
rect 13988 11987 13998 12095
rect 14130 11987 14140 12095
rect 14018 11851 14024 11987
rect 14091 11851 14097 11987
rect 14018 11839 14097 11851
rect 10602 11613 11579 11643
rect 13796 11641 13859 11658
rect 13721 11637 13859 11641
rect 10602 11507 10634 11613
rect 10838 11507 10870 11613
rect 11074 11507 11106 11613
rect 11310 11507 11342 11613
rect 11545 11507 11579 11613
rect 11889 11603 13859 11637
rect 11887 11574 13859 11603
rect 11887 11558 11933 11574
rect 13721 11572 13859 11574
rect 10595 11495 10641 11507
rect 10595 11319 10601 11495
rect 10635 11319 10641 11495
rect 10595 11307 10641 11319
rect 10713 11495 10759 11507
rect 10713 11319 10719 11495
rect 10753 11319 10759 11495
rect 10713 11307 10759 11319
rect 10831 11495 10877 11507
rect 10831 11319 10837 11495
rect 10871 11319 10877 11495
rect 10831 11307 10877 11319
rect 10949 11495 10995 11507
rect 10949 11319 10955 11495
rect 10989 11319 10995 11495
rect 10949 11307 10995 11319
rect 11067 11495 11113 11507
rect 11067 11319 11073 11495
rect 11107 11319 11113 11495
rect 11067 11307 11113 11319
rect 11185 11495 11231 11507
rect 11185 11319 11191 11495
rect 11225 11319 11231 11495
rect 11185 11307 11231 11319
rect 11303 11495 11349 11507
rect 11303 11319 11309 11495
rect 11343 11319 11349 11495
rect 11303 11307 11349 11319
rect 11421 11495 11467 11507
rect 11421 11319 11427 11495
rect 11461 11319 11467 11495
rect 11421 11307 11467 11319
rect 11539 11495 11585 11507
rect 11539 11319 11545 11495
rect 11579 11319 11585 11495
rect 11539 11307 11585 11319
rect 11657 11495 11703 11507
rect 11657 11319 11663 11495
rect 11697 11319 11703 11495
rect 11657 11307 11703 11319
rect 10718 11213 10754 11307
rect 10954 11213 10990 11307
rect 11190 11214 11226 11307
rect 11352 11259 11418 11266
rect 11352 11225 11368 11259
rect 11402 11225 11418 11259
rect 11352 11214 11418 11225
rect 11190 11213 11418 11214
rect 10718 11184 11418 11213
rect 10718 11183 11300 11184
rect 10838 11070 10872 11183
rect 11234 11142 11300 11183
rect 11234 11108 11250 11142
rect 11284 11108 11300 11142
rect 11234 11101 11300 11108
rect 11662 11089 11697 11307
rect 11886 11106 11933 11558
rect 14785 11566 14864 11578
rect 14785 11450 14791 11566
rect 14858 11450 14864 11566
rect 12845 11342 12855 11450
rect 12987 11342 12997 11450
rect 14743 11342 14753 11450
rect 14885 11342 14895 11450
rect 12855 11302 12987 11342
rect 14753 11302 14885 11342
rect 12854 11236 12987 11302
rect 14752 11236 14885 11302
rect 12183 11193 13656 11236
rect 11886 11090 11932 11106
rect 11851 11089 11932 11090
rect 11662 11074 11932 11089
rect 11308 11070 11932 11074
rect 10832 11058 10878 11070
rect 10567 10580 10577 10698
rect 10695 10666 10705 10698
rect 10832 10682 10838 11058
rect 10872 10682 10878 11058
rect 10832 10670 10878 10682
rect 10950 11058 10996 11070
rect 10950 10682 10956 11058
rect 10990 10682 10996 11058
rect 10950 10670 10996 10682
rect 11068 11058 11114 11070
rect 11068 10682 11074 11058
rect 11108 10706 11114 11058
rect 11185 11058 11231 11070
rect 11185 10882 11191 11058
rect 11225 10882 11231 11058
rect 11185 10870 11231 10882
rect 11303 11058 11932 11070
rect 11303 10882 11309 11058
rect 11343 11046 11932 11058
rect 11343 11045 11585 11046
rect 11343 10882 11349 11045
rect 11851 11044 11932 11046
rect 12183 10890 12217 11193
rect 12549 11090 12583 11193
rect 12785 11090 12819 11193
rect 13021 11090 13055 11193
rect 13257 11090 13291 11193
rect 12543 11078 12589 11090
rect 11303 10870 11349 10882
rect 12059 10878 12105 10890
rect 11191 10754 11226 10870
rect 11322 10754 11430 10764
rect 11191 10706 11322 10754
rect 11430 10715 11579 10721
rect 11108 10682 11322 10706
rect 11068 10670 11322 10682
rect 11074 10666 11322 10670
rect 10695 10638 10710 10666
rect 10695 10632 10947 10638
rect 10695 10598 10897 10632
rect 10931 10598 10947 10632
rect 10695 10582 10947 10598
rect 10999 10632 11065 10638
rect 10999 10598 11015 10632
rect 11049 10598 11065 10632
rect 11248 10622 11322 10666
rect 11567 10648 11579 10715
rect 12059 10702 12065 10878
rect 12099 10702 12105 10878
rect 12059 10690 12105 10702
rect 12177 10878 12223 10890
rect 12177 10702 12183 10878
rect 12217 10702 12223 10878
rect 12177 10690 12223 10702
rect 12295 10878 12341 10890
rect 12295 10702 12301 10878
rect 12335 10702 12341 10878
rect 12295 10690 12341 10702
rect 12413 10878 12459 10890
rect 12543 10878 12549 11078
rect 12413 10702 12419 10878
rect 12453 10702 12549 10878
rect 12583 10702 12589 11078
rect 12413 10690 12459 10702
rect 12543 10690 12589 10702
rect 12661 11078 12707 11090
rect 12661 10702 12667 11078
rect 12701 10702 12707 11078
rect 12661 10690 12707 10702
rect 12779 11078 12825 11090
rect 12779 10702 12785 11078
rect 12819 10702 12825 11078
rect 12779 10690 12825 10702
rect 12897 11078 12943 11090
rect 12897 10702 12903 11078
rect 12937 10702 12943 11078
rect 12897 10690 12943 10702
rect 13015 11078 13061 11090
rect 13015 10702 13021 11078
rect 13055 10702 13061 11078
rect 13015 10690 13061 10702
rect 13133 11078 13179 11090
rect 13133 10702 13139 11078
rect 13173 10702 13179 11078
rect 13133 10690 13179 10702
rect 13251 11078 13297 11090
rect 13251 10702 13257 11078
rect 13291 10878 13297 11078
rect 13622 10890 13656 11193
rect 14081 11193 15554 11236
rect 14081 10890 14115 11193
rect 14447 11090 14481 11193
rect 14683 11090 14717 11193
rect 14919 11090 14953 11193
rect 15155 11090 15189 11193
rect 14441 11078 14487 11090
rect 13380 10878 13426 10890
rect 13291 10702 13386 10878
rect 13420 10702 13426 10878
rect 13251 10690 13297 10702
rect 13380 10690 13426 10702
rect 13498 10878 13544 10890
rect 13498 10702 13504 10878
rect 13538 10702 13544 10878
rect 13498 10690 13544 10702
rect 13616 10878 13662 10890
rect 13616 10702 13622 10878
rect 13656 10702 13662 10878
rect 13616 10690 13662 10702
rect 13734 10878 13780 10890
rect 13734 10702 13740 10878
rect 13774 10702 13780 10878
rect 13734 10690 13780 10702
rect 13957 10878 14003 10890
rect 13957 10702 13963 10878
rect 13997 10702 14003 10878
rect 13957 10690 14003 10702
rect 14075 10878 14121 10890
rect 14075 10702 14081 10878
rect 14115 10702 14121 10878
rect 14075 10690 14121 10702
rect 14193 10878 14239 10890
rect 14193 10702 14199 10878
rect 14233 10702 14239 10878
rect 14193 10690 14239 10702
rect 14311 10878 14357 10890
rect 14441 10878 14447 11078
rect 14311 10702 14317 10878
rect 14351 10702 14447 10878
rect 14481 10702 14487 11078
rect 14311 10690 14357 10702
rect 14441 10690 14487 10702
rect 14559 11078 14605 11090
rect 14559 10702 14565 11078
rect 14599 10702 14605 11078
rect 14559 10690 14605 10702
rect 14677 11078 14723 11090
rect 14677 10702 14683 11078
rect 14717 10702 14723 11078
rect 14677 10690 14723 10702
rect 14795 11078 14841 11090
rect 14795 10702 14801 11078
rect 14835 10702 14841 11078
rect 14795 10690 14841 10702
rect 14913 11078 14959 11090
rect 14913 10702 14919 11078
rect 14953 10702 14959 11078
rect 14913 10690 14959 10702
rect 15031 11078 15077 11090
rect 15031 10702 15037 11078
rect 15071 10702 15077 11078
rect 15031 10690 15077 10702
rect 15149 11078 15195 11090
rect 15149 10702 15155 11078
rect 15189 10878 15195 11078
rect 15520 10890 15554 11193
rect 15278 10878 15324 10890
rect 15189 10702 15284 10878
rect 15318 10702 15324 10878
rect 15149 10690 15195 10702
rect 15278 10690 15324 10702
rect 15396 10878 15442 10890
rect 15396 10702 15402 10878
rect 15436 10702 15442 10878
rect 15396 10690 15442 10702
rect 15514 10878 15560 10890
rect 15514 10702 15520 10878
rect 15554 10702 15560 10878
rect 15514 10690 15560 10702
rect 15632 10878 15678 10890
rect 15632 10702 15638 10878
rect 15672 10702 15678 10878
rect 15632 10690 15678 10702
rect 11430 10642 11579 10648
rect 12065 10656 12099 10690
rect 12667 10656 12701 10690
rect 12903 10656 12937 10690
rect 11322 10612 11430 10622
rect 12065 10621 12224 10656
rect 12667 10621 12937 10656
rect 13504 10656 13538 10690
rect 13740 10656 13774 10690
rect 13504 10621 13774 10656
rect 13963 10656 13997 10690
rect 14565 10656 14599 10690
rect 14801 10656 14835 10690
rect 13963 10621 14122 10656
rect 14565 10621 14835 10656
rect 15402 10656 15436 10690
rect 15638 10656 15672 10690
rect 15402 10621 15672 10656
rect 10695 10580 10710 10582
rect 10610 10566 10710 10580
rect 10610 10523 10710 10524
rect 10231 10502 10710 10523
rect 10999 10502 11065 10598
rect 10231 10454 11065 10502
rect 10231 10425 10710 10454
rect 10231 10423 10336 10425
rect 10610 10424 10710 10425
rect 10064 10238 10074 10317
rect 10167 10238 10177 10317
rect 11062 10308 11141 10320
rect 10075 9064 10168 10238
rect 11062 10209 11068 10308
rect 10993 10189 11068 10209
rect 11135 10209 11141 10308
rect 11135 10189 11213 10209
rect 10993 10081 11037 10189
rect 11169 10081 11213 10189
rect 10993 10039 11213 10081
rect 10597 10009 11574 10039
rect 10597 9903 10629 10009
rect 10833 9903 10865 10009
rect 11069 9903 11101 10009
rect 11305 9903 11337 10009
rect 11540 9903 11574 10009
rect 10590 9891 10636 9903
rect 10590 9715 10596 9891
rect 10630 9715 10636 9891
rect 10590 9703 10636 9715
rect 10708 9891 10754 9903
rect 10708 9715 10714 9891
rect 10748 9715 10754 9891
rect 10708 9703 10754 9715
rect 10826 9891 10872 9903
rect 10826 9715 10832 9891
rect 10866 9715 10872 9891
rect 10826 9703 10872 9715
rect 10944 9891 10990 9903
rect 10944 9715 10950 9891
rect 10984 9715 10990 9891
rect 10944 9703 10990 9715
rect 11062 9891 11108 9903
rect 11062 9715 11068 9891
rect 11102 9715 11108 9891
rect 11062 9703 11108 9715
rect 11180 9891 11226 9903
rect 11180 9715 11186 9891
rect 11220 9715 11226 9891
rect 11180 9703 11226 9715
rect 11298 9891 11344 9903
rect 11298 9715 11304 9891
rect 11338 9715 11344 9891
rect 11298 9703 11344 9715
rect 11416 9891 11462 9903
rect 11416 9715 11422 9891
rect 11456 9715 11462 9891
rect 11416 9703 11462 9715
rect 11534 9891 11580 9903
rect 11534 9715 11540 9891
rect 11574 9715 11580 9891
rect 11534 9703 11580 9715
rect 11652 9891 11698 9903
rect 11652 9715 11658 9891
rect 11692 9715 11698 9891
rect 11652 9703 11698 9715
rect 12190 9837 12224 10621
rect 12903 10559 12937 10621
rect 12492 10521 13234 10559
rect 12492 10397 12526 10521
rect 12728 10397 12762 10521
rect 12964 10397 12998 10521
rect 13200 10397 13234 10521
rect 13490 10414 13500 10480
rect 13563 10414 13573 10480
rect 12486 10385 12532 10397
rect 12486 10009 12492 10385
rect 12526 10009 12532 10385
rect 12486 9997 12532 10009
rect 12604 10385 12650 10397
rect 12604 10009 12610 10385
rect 12644 10009 12650 10385
rect 12604 9997 12650 10009
rect 12722 10385 12768 10397
rect 12722 10009 12728 10385
rect 12762 10009 12768 10385
rect 12722 9997 12768 10009
rect 12840 10385 12886 10397
rect 12840 10009 12846 10385
rect 12880 10009 12886 10385
rect 12840 9997 12886 10009
rect 12958 10385 13004 10397
rect 12958 10009 12964 10385
rect 12998 10009 13004 10385
rect 12958 9997 13004 10009
rect 13076 10385 13122 10397
rect 13076 10009 13082 10385
rect 13116 10009 13122 10385
rect 13076 9997 13122 10009
rect 13194 10385 13240 10397
rect 13194 10009 13200 10385
rect 13234 10009 13240 10385
rect 13194 9997 13240 10009
rect 13606 9838 13640 10621
rect 13333 9837 13640 9838
rect 12190 9832 12506 9837
rect 13220 9832 13640 9837
rect 12190 9821 12573 9832
rect 12190 9794 12522 9821
rect 10713 9609 10749 9703
rect 10949 9609 10985 9703
rect 11185 9610 11221 9703
rect 11347 9655 11413 9662
rect 11347 9621 11363 9655
rect 11397 9621 11413 9655
rect 11347 9610 11413 9621
rect 11185 9609 11413 9610
rect 10713 9580 11413 9609
rect 10713 9579 11295 9580
rect 10833 9466 10867 9579
rect 11229 9538 11295 9579
rect 11229 9504 11245 9538
rect 11279 9504 11295 9538
rect 11229 9497 11295 9504
rect 11657 9470 11692 9703
rect 12190 9665 12224 9794
rect 12506 9787 12522 9794
rect 12556 9787 12573 9821
rect 12506 9781 12573 9787
rect 13153 9821 13640 9832
rect 13153 9787 13170 9821
rect 13204 9794 13640 9821
rect 13204 9787 13220 9794
rect 13333 9793 13640 9794
rect 13153 9781 13220 9787
rect 12331 9754 12387 9766
rect 12331 9720 12337 9754
rect 12371 9753 12387 9754
rect 13444 9753 13500 9765
rect 12371 9737 12838 9753
rect 12371 9720 12788 9737
rect 12331 9704 12788 9720
rect 12772 9703 12788 9704
rect 12822 9703 12838 9737
rect 12772 9696 12838 9703
rect 12890 9738 13460 9753
rect 12890 9704 12906 9738
rect 12940 9719 13460 9738
rect 13494 9719 13500 9753
rect 12940 9704 13500 9719
rect 12890 9694 12957 9704
rect 13444 9703 13500 9704
rect 13606 9665 13640 9793
rect 14088 9837 14122 10621
rect 14801 10559 14835 10621
rect 14390 10521 15132 10559
rect 14390 10397 14424 10521
rect 14626 10397 14660 10521
rect 14862 10397 14896 10521
rect 15098 10397 15132 10521
rect 14384 10385 14430 10397
rect 14384 10009 14390 10385
rect 14424 10009 14430 10385
rect 14384 9997 14430 10009
rect 14502 10385 14548 10397
rect 14502 10009 14508 10385
rect 14542 10009 14548 10385
rect 14502 9997 14548 10009
rect 14620 10385 14666 10397
rect 14620 10009 14626 10385
rect 14660 10009 14666 10385
rect 14620 9997 14666 10009
rect 14738 10385 14784 10397
rect 14738 10009 14744 10385
rect 14778 10009 14784 10385
rect 14738 9997 14784 10009
rect 14856 10385 14902 10397
rect 14856 10009 14862 10385
rect 14896 10009 14902 10385
rect 14856 9997 14902 10009
rect 14974 10385 15020 10397
rect 14974 10009 14980 10385
rect 15014 10009 15020 10385
rect 14974 9997 15020 10009
rect 15092 10385 15138 10397
rect 15092 10009 15098 10385
rect 15132 10009 15138 10385
rect 15092 9997 15138 10009
rect 15504 9838 15538 10621
rect 15116 9837 15185 9838
rect 15231 9837 15538 9838
rect 14088 9832 14404 9837
rect 15116 9833 15538 9837
rect 14088 9821 14471 9832
rect 14088 9794 14420 9821
rect 14088 9665 14122 9794
rect 14404 9787 14420 9794
rect 14454 9787 14471 9821
rect 14404 9781 14471 9787
rect 15049 9822 15538 9833
rect 15049 9788 15066 9822
rect 15100 9794 15538 9822
rect 15100 9788 15116 9794
rect 15231 9793 15538 9794
rect 15049 9782 15116 9788
rect 14229 9754 14285 9766
rect 14229 9720 14235 9754
rect 14269 9753 14285 9754
rect 15342 9753 15398 9765
rect 14269 9737 14736 9753
rect 14269 9720 14686 9737
rect 14229 9704 14686 9720
rect 14670 9703 14686 9704
rect 14720 9703 14736 9737
rect 14670 9696 14736 9703
rect 14788 9738 15358 9753
rect 14788 9704 14804 9738
rect 14838 9719 15358 9738
rect 15392 9719 15398 9753
rect 14838 9704 15398 9719
rect 14788 9694 14855 9704
rect 15342 9703 15398 9704
rect 15504 9665 15538 9793
rect 15619 10443 15686 10467
rect 15619 10409 15636 10443
rect 15670 10409 15686 10443
rect 11303 9466 11692 9470
rect 10827 9454 10873 9466
rect 10827 9078 10833 9454
rect 10867 9078 10873 9454
rect 10827 9066 10873 9078
rect 10945 9454 10991 9466
rect 10945 9078 10951 9454
rect 10985 9078 10991 9454
rect 10945 9066 10991 9078
rect 11063 9454 11109 9466
rect 11063 9078 11069 9454
rect 11103 9102 11109 9454
rect 11180 9454 11226 9466
rect 11180 9278 11186 9454
rect 11220 9278 11226 9454
rect 11180 9266 11226 9278
rect 11298 9454 11692 9466
rect 12184 9653 12230 9665
rect 12184 9477 12190 9653
rect 12224 9477 12230 9653
rect 12184 9465 12230 9477
rect 12302 9653 12348 9665
rect 12302 9477 12308 9653
rect 12342 9477 12348 9653
rect 12302 9465 12348 9477
rect 12604 9653 12650 9665
rect 11298 9278 11304 9454
rect 11338 9441 11692 9454
rect 11338 9278 11344 9441
rect 11614 9438 11692 9441
rect 11614 9386 11624 9438
rect 11687 9386 11697 9438
rect 11619 9380 11692 9386
rect 11298 9266 11344 9278
rect 11186 9150 11221 9266
rect 12307 9171 12341 9465
rect 12604 9277 12610 9653
rect 12644 9277 12650 9653
rect 12604 9265 12650 9277
rect 12722 9653 12768 9665
rect 12722 9277 12728 9653
rect 12762 9277 12768 9653
rect 12722 9265 12768 9277
rect 12840 9653 12886 9665
rect 12840 9277 12846 9653
rect 12880 9277 12886 9653
rect 12840 9265 12886 9277
rect 12958 9653 13004 9665
rect 12958 9277 12964 9653
rect 12998 9277 13004 9653
rect 12958 9265 13004 9277
rect 13076 9653 13122 9665
rect 13076 9277 13082 9653
rect 13116 9277 13122 9653
rect 13482 9653 13528 9665
rect 13482 9477 13488 9653
rect 13522 9477 13528 9653
rect 13482 9465 13528 9477
rect 13600 9653 13646 9665
rect 13600 9477 13606 9653
rect 13640 9477 13646 9653
rect 13600 9465 13646 9477
rect 14082 9653 14128 9665
rect 14082 9477 14088 9653
rect 14122 9477 14128 9653
rect 14082 9465 14128 9477
rect 14200 9653 14246 9665
rect 14200 9477 14206 9653
rect 14240 9477 14246 9653
rect 14200 9465 14246 9477
rect 14502 9653 14548 9665
rect 13076 9265 13122 9277
rect 12964 9171 12998 9265
rect 13488 9171 13521 9465
rect 11317 9150 11425 9160
rect 11186 9102 11317 9150
rect 12307 9139 13521 9171
rect 14205 9171 14239 9465
rect 14502 9277 14508 9653
rect 14542 9277 14548 9653
rect 14502 9265 14548 9277
rect 14620 9653 14666 9665
rect 14620 9277 14626 9653
rect 14660 9277 14666 9653
rect 14620 9265 14666 9277
rect 14738 9653 14784 9665
rect 14738 9277 14744 9653
rect 14778 9277 14784 9653
rect 14738 9265 14784 9277
rect 14856 9653 14902 9665
rect 14856 9277 14862 9653
rect 14896 9277 14902 9653
rect 14856 9265 14902 9277
rect 14974 9653 15020 9665
rect 14974 9277 14980 9653
rect 15014 9277 15020 9653
rect 15380 9653 15426 9665
rect 15380 9477 15386 9653
rect 15420 9477 15426 9653
rect 15380 9465 15426 9477
rect 15498 9653 15544 9665
rect 15498 9477 15504 9653
rect 15538 9477 15544 9653
rect 15498 9465 15544 9477
rect 14974 9265 15020 9277
rect 14862 9171 14896 9265
rect 15386 9171 15419 9465
rect 14205 9139 15419 9171
rect 11425 9114 11576 9120
rect 11103 9078 11317 9102
rect 11063 9066 11317 9078
rect 10075 9062 10660 9064
rect 11069 9062 11317 9066
rect 10075 9034 10705 9062
rect 10075 9028 10942 9034
rect 10075 8994 10892 9028
rect 10926 8994 10942 9028
rect 10075 8978 10942 8994
rect 10994 9028 11060 9034
rect 10994 8994 11010 9028
rect 11044 8994 11060 9028
rect 11243 9018 11317 9062
rect 11564 9047 11576 9114
rect 12800 9054 12932 9139
rect 14698 9054 14830 9139
rect 11425 9041 11576 9047
rect 11317 9008 11425 9018
rect 10075 8962 10705 8978
rect 10075 8958 10660 8962
rect 10075 8957 10176 8958
rect 10605 8909 10705 8920
rect 10569 8803 10579 8909
rect 10691 8898 10705 8909
rect 10994 8898 11060 8994
rect 12790 8946 12800 9054
rect 12932 8946 12942 9054
rect 14688 8946 14698 9054
rect 14830 8946 14840 9054
rect 15619 9026 15686 10409
rect 15747 9980 15903 9986
rect 15747 9882 15759 9980
rect 15891 9882 15903 9980
rect 15747 9876 15903 9882
rect 10691 8850 11060 8898
rect 10691 8820 10705 8850
rect 10691 8803 10701 8820
rect 10993 8747 11059 8850
rect 12823 8808 12829 8946
rect 12896 8808 12902 8946
rect 12823 8796 12902 8808
rect 15619 8747 15685 9026
rect 10991 8667 15685 8747
rect 13531 7743 13610 7755
rect 11050 7690 11129 7702
rect 11050 7593 11056 7690
rect 10978 7573 11056 7593
rect 11123 7593 11129 7690
rect 13531 7627 13537 7743
rect 13604 7627 13610 7743
rect 14679 7743 14758 7755
rect 14679 7627 14685 7743
rect 14752 7627 14758 7743
rect 11123 7573 11198 7593
rect 10978 7465 11022 7573
rect 11154 7465 11198 7573
rect 12775 7531 12831 7539
rect 10978 7423 11198 7465
rect 11849 7523 12831 7531
rect 11849 7489 12791 7523
rect 12825 7489 12831 7523
rect 13494 7519 13504 7627
rect 13636 7564 13646 7627
rect 13636 7553 13648 7564
rect 13636 7519 13649 7553
rect 13905 7543 13961 7545
rect 11849 7473 12831 7489
rect 13504 7481 13649 7519
rect 11849 7472 12828 7473
rect 10582 7393 11559 7423
rect 10582 7287 10614 7393
rect 10818 7287 10850 7393
rect 11054 7287 11086 7393
rect 11290 7287 11322 7393
rect 11525 7287 11559 7393
rect 10575 7275 10621 7287
rect 10575 7099 10581 7275
rect 10615 7099 10621 7275
rect 10575 7087 10621 7099
rect 10693 7275 10739 7287
rect 10693 7099 10699 7275
rect 10733 7099 10739 7275
rect 10693 7087 10739 7099
rect 10811 7275 10857 7287
rect 10811 7099 10817 7275
rect 10851 7099 10857 7275
rect 10811 7087 10857 7099
rect 10929 7275 10975 7287
rect 10929 7099 10935 7275
rect 10969 7099 10975 7275
rect 10929 7087 10975 7099
rect 11047 7275 11093 7287
rect 11047 7099 11053 7275
rect 11087 7099 11093 7275
rect 11047 7087 11093 7099
rect 11165 7275 11211 7287
rect 11165 7099 11171 7275
rect 11205 7099 11211 7275
rect 11165 7087 11211 7099
rect 11283 7275 11329 7287
rect 11283 7099 11289 7275
rect 11323 7099 11329 7275
rect 11283 7087 11329 7099
rect 11401 7275 11447 7287
rect 11401 7099 11407 7275
rect 11441 7099 11447 7275
rect 11401 7087 11447 7099
rect 11519 7275 11565 7287
rect 11519 7099 11525 7275
rect 11559 7099 11565 7275
rect 11519 7087 11565 7099
rect 11637 7275 11683 7287
rect 11637 7099 11643 7275
rect 11677 7099 11683 7275
rect 11637 7087 11683 7099
rect 10698 6993 10734 7087
rect 10934 6993 10970 7087
rect 11170 6994 11206 7087
rect 11332 7039 11398 7046
rect 11332 7005 11348 7039
rect 11382 7005 11398 7039
rect 11332 6994 11398 7005
rect 11170 6993 11398 6994
rect 10698 6964 11398 6993
rect 10698 6963 11280 6964
rect 10818 6850 10852 6963
rect 11214 6922 11280 6963
rect 11214 6888 11230 6922
rect 11264 6888 11280 6922
rect 11214 6881 11280 6888
rect 11642 6882 11677 7087
rect 11849 6882 11916 7472
rect 13608 7449 13649 7481
rect 13895 7477 13905 7543
rect 13961 7477 13971 7543
rect 14641 7519 14651 7627
rect 14783 7564 14793 7627
rect 14783 7553 14795 7564
rect 14783 7519 14796 7553
rect 14651 7481 14796 7519
rect 14755 7453 14796 7481
rect 13024 7421 13294 7449
rect 12765 7355 12775 7421
rect 12841 7355 12851 7421
rect 13024 7359 13058 7421
rect 13260 7359 13294 7421
rect 13378 7421 13649 7449
rect 14166 7425 14436 7453
rect 13378 7359 13412 7421
rect 13614 7359 13649 7421
rect 13790 7409 13961 7425
rect 13790 7375 13921 7409
rect 13955 7375 13961 7409
rect 13790 7359 13961 7375
rect 14166 7363 14200 7425
rect 14402 7363 14436 7425
rect 14520 7425 14796 7453
rect 14520 7363 14554 7425
rect 14756 7363 14796 7425
rect 12900 7347 12946 7359
rect 12900 6971 12906 7347
rect 12940 6971 12946 7347
rect 12900 6959 12946 6971
rect 13018 7347 13064 7359
rect 13018 6971 13024 7347
rect 13058 6971 13064 7347
rect 13018 6959 13064 6971
rect 13136 7347 13182 7359
rect 13136 6971 13142 7347
rect 13176 6971 13182 7347
rect 13136 6959 13182 6971
rect 13254 7347 13300 7359
rect 13254 6971 13260 7347
rect 13294 6971 13300 7347
rect 13254 6959 13300 6971
rect 13372 7347 13418 7359
rect 13372 6971 13378 7347
rect 13412 6971 13418 7347
rect 13372 6959 13418 6971
rect 13490 7347 13536 7359
rect 13490 6971 13496 7347
rect 13530 6971 13536 7347
rect 13490 6959 13536 6971
rect 13608 7347 13654 7359
rect 13608 6971 13614 7347
rect 13648 6971 13654 7347
rect 13608 6959 13654 6971
rect 11642 6854 11916 6882
rect 11288 6850 11916 6854
rect 9196 6796 9551 6797
rect 8205 6728 8314 6782
rect 7525 6689 7752 6725
rect 7525 6582 7560 6689
rect 7686 6655 7752 6689
rect 7686 6621 7702 6655
rect 7736 6621 7752 6655
rect 8033 6713 8130 6728
rect 8033 6646 8090 6713
rect 7686 6615 7752 6621
rect 7927 6610 8196 6646
rect 7927 6582 7960 6610
rect 8163 6582 8196 6610
rect 8280 6582 8314 6728
rect 9131 6721 9141 6796
rect 9209 6721 9551 6796
rect 9158 6720 9551 6721
rect 9196 6719 9551 6720
rect 10812 6838 10858 6850
rect 7401 6570 7447 6582
rect 7401 6394 7407 6570
rect 7441 6394 7447 6570
rect 7401 6382 7447 6394
rect 7519 6570 7565 6582
rect 7519 6394 7525 6570
rect 7559 6394 7565 6570
rect 7519 6382 7565 6394
rect 7637 6570 7683 6582
rect 7637 6394 7643 6570
rect 7677 6394 7683 6570
rect 7637 6382 7683 6394
rect 7755 6570 7801 6582
rect 7755 6394 7761 6570
rect 7795 6515 7801 6570
rect 7920 6570 7966 6582
rect 7920 6515 7926 6570
rect 7795 6427 7926 6515
rect 7795 6394 7801 6427
rect 7755 6382 7801 6394
rect 7920 6394 7926 6427
rect 7960 6394 7966 6570
rect 7920 6382 7966 6394
rect 8038 6570 8084 6582
rect 8038 6394 8044 6570
rect 8078 6394 8084 6570
rect 8038 6382 8084 6394
rect 8156 6570 8202 6582
rect 8156 6394 8162 6570
rect 8196 6394 8202 6570
rect 8156 6382 8202 6394
rect 8274 6570 8320 6582
rect 8274 6394 8280 6570
rect 8314 6394 8320 6570
rect 10812 6462 10818 6838
rect 10852 6462 10858 6838
rect 10812 6450 10858 6462
rect 10930 6838 10976 6850
rect 10930 6462 10936 6838
rect 10970 6462 10976 6838
rect 10930 6450 10976 6462
rect 11048 6838 11094 6850
rect 11048 6462 11054 6838
rect 11088 6486 11094 6838
rect 11165 6838 11211 6850
rect 11165 6662 11171 6838
rect 11205 6662 11211 6838
rect 11165 6650 11211 6662
rect 11283 6838 11916 6850
rect 11283 6662 11289 6838
rect 11323 6825 11916 6838
rect 12906 6917 12940 6959
rect 13142 6917 13176 6959
rect 12906 6889 13176 6917
rect 13260 6918 13294 6959
rect 13496 6918 13530 6959
rect 13260 6889 13530 6918
rect 12906 6841 12940 6889
rect 11323 6662 11329 6825
rect 12906 6811 12969 6841
rect 11283 6650 11329 6662
rect 12934 6719 12969 6811
rect 12934 6683 13161 6719
rect 13431 6708 13441 6805
rect 13540 6708 13550 6805
rect 13614 6776 13648 6959
rect 13614 6722 13723 6776
rect 11171 6534 11206 6650
rect 12934 6576 12969 6683
rect 13095 6649 13161 6683
rect 13095 6615 13111 6649
rect 13145 6615 13161 6649
rect 13442 6707 13539 6708
rect 13442 6640 13499 6707
rect 13095 6609 13161 6615
rect 13336 6604 13605 6640
rect 13336 6576 13369 6604
rect 13572 6576 13605 6604
rect 13689 6576 13723 6722
rect 12810 6564 12856 6576
rect 11302 6534 11410 6544
rect 11171 6486 11302 6534
rect 11410 6490 11555 6496
rect 11088 6462 11302 6486
rect 11048 6450 11302 6462
rect 11054 6446 11302 6450
rect 8274 6382 8320 6394
rect 9190 6418 10690 6445
rect 9190 6412 10927 6418
rect 7407 6343 7441 6382
rect 7643 6343 7677 6382
rect 7407 6307 7677 6343
rect 8044 6344 8077 6382
rect 8280 6344 8313 6382
rect 8044 6308 8313 6344
rect 9190 6378 10877 6412
rect 10911 6378 10927 6412
rect 9190 6362 10927 6378
rect 10979 6412 11045 6418
rect 10979 6378 10995 6412
rect 11029 6378 11045 6412
rect 11228 6402 11302 6446
rect 11543 6423 11555 6490
rect 11410 6417 11555 6423
rect 11302 6392 11410 6402
rect 9190 6346 10690 6362
rect 9190 6345 10627 6346
rect 9190 6339 10162 6345
rect 7407 6306 7573 6307
rect 7441 6227 7573 6306
rect 7431 6119 7441 6227
rect 7573 6119 7583 6227
rect 7468 5981 7474 6119
rect 7541 5981 7547 6119
rect 7468 5969 7547 5981
rect 4045 5745 5022 5775
rect 7239 5773 7302 5790
rect 7164 5769 7302 5773
rect 4045 5639 4077 5745
rect 4281 5639 4313 5745
rect 4517 5639 4549 5745
rect 4753 5639 4785 5745
rect 4988 5639 5022 5745
rect 5332 5735 7302 5769
rect 5330 5706 7302 5735
rect 5330 5690 5376 5706
rect 7164 5704 7302 5706
rect 4038 5627 4084 5639
rect 4038 5451 4044 5627
rect 4078 5451 4084 5627
rect 4038 5439 4084 5451
rect 4156 5627 4202 5639
rect 4156 5451 4162 5627
rect 4196 5451 4202 5627
rect 4156 5439 4202 5451
rect 4274 5627 4320 5639
rect 4274 5451 4280 5627
rect 4314 5451 4320 5627
rect 4274 5439 4320 5451
rect 4392 5627 4438 5639
rect 4392 5451 4398 5627
rect 4432 5451 4438 5627
rect 4392 5439 4438 5451
rect 4510 5627 4556 5639
rect 4510 5451 4516 5627
rect 4550 5451 4556 5627
rect 4510 5439 4556 5451
rect 4628 5627 4674 5639
rect 4628 5451 4634 5627
rect 4668 5451 4674 5627
rect 4628 5439 4674 5451
rect 4746 5627 4792 5639
rect 4746 5451 4752 5627
rect 4786 5451 4792 5627
rect 4746 5439 4792 5451
rect 4864 5627 4910 5639
rect 4864 5451 4870 5627
rect 4904 5451 4910 5627
rect 4864 5439 4910 5451
rect 4982 5627 5028 5639
rect 4982 5451 4988 5627
rect 5022 5451 5028 5627
rect 4982 5439 5028 5451
rect 5100 5627 5146 5639
rect 5100 5451 5106 5627
rect 5140 5451 5146 5627
rect 5100 5439 5146 5451
rect 4161 5345 4197 5439
rect 4397 5345 4433 5439
rect 4633 5346 4669 5439
rect 4795 5391 4861 5398
rect 4795 5357 4811 5391
rect 4845 5357 4861 5391
rect 4795 5346 4861 5357
rect 4633 5345 4861 5346
rect 4161 5316 4861 5345
rect 4161 5315 4743 5316
rect 4281 5202 4315 5315
rect 4677 5274 4743 5315
rect 4677 5240 4693 5274
rect 4727 5240 4743 5274
rect 4677 5233 4743 5240
rect 5105 5221 5140 5439
rect 5329 5238 5376 5690
rect 8222 5698 8301 5710
rect 8222 5582 8228 5698
rect 8295 5582 8301 5698
rect 6288 5474 6298 5582
rect 6430 5474 6440 5582
rect 8186 5474 8196 5582
rect 8328 5474 8338 5582
rect 6298 5434 6430 5474
rect 8196 5434 8328 5474
rect 6297 5368 6430 5434
rect 8195 5368 8328 5434
rect 5626 5325 7099 5368
rect 5329 5222 5375 5238
rect 5294 5221 5375 5222
rect 5105 5206 5375 5221
rect 4751 5202 5375 5206
rect 4275 5190 4321 5202
rect 4010 4712 4020 4830
rect 4138 4798 4148 4830
rect 4275 4814 4281 5190
rect 4315 4814 4321 5190
rect 4275 4802 4321 4814
rect 4393 5190 4439 5202
rect 4393 4814 4399 5190
rect 4433 4814 4439 5190
rect 4393 4802 4439 4814
rect 4511 5190 4557 5202
rect 4511 4814 4517 5190
rect 4551 4838 4557 5190
rect 4628 5190 4674 5202
rect 4628 5014 4634 5190
rect 4668 5014 4674 5190
rect 4628 5002 4674 5014
rect 4746 5190 5375 5202
rect 4746 5014 4752 5190
rect 4786 5178 5375 5190
rect 4786 5177 5028 5178
rect 4786 5014 4792 5177
rect 5294 5176 5375 5178
rect 5626 5022 5660 5325
rect 5992 5222 6026 5325
rect 6228 5222 6262 5325
rect 6464 5222 6498 5325
rect 6700 5222 6734 5325
rect 5986 5210 6032 5222
rect 4746 5002 4792 5014
rect 5502 5010 5548 5022
rect 4634 4886 4669 5002
rect 4765 4886 4873 4896
rect 4634 4838 4765 4886
rect 4873 4846 5013 4852
rect 4551 4814 4765 4838
rect 4511 4802 4765 4814
rect 4517 4798 4765 4802
rect 4138 4770 4153 4798
rect 4138 4764 4390 4770
rect 4138 4730 4340 4764
rect 4374 4730 4390 4764
rect 4138 4714 4390 4730
rect 4442 4764 4508 4770
rect 4442 4730 4458 4764
rect 4492 4730 4508 4764
rect 4691 4754 4765 4798
rect 5001 4779 5013 4846
rect 5502 4834 5508 5010
rect 5542 4834 5548 5010
rect 5502 4822 5548 4834
rect 5620 5010 5666 5022
rect 5620 4834 5626 5010
rect 5660 4834 5666 5010
rect 5620 4822 5666 4834
rect 5738 5010 5784 5022
rect 5738 4834 5744 5010
rect 5778 4834 5784 5010
rect 5738 4822 5784 4834
rect 5856 5010 5902 5022
rect 5986 5010 5992 5210
rect 5856 4834 5862 5010
rect 5896 4834 5992 5010
rect 6026 4834 6032 5210
rect 5856 4822 5902 4834
rect 5986 4822 6032 4834
rect 6104 5210 6150 5222
rect 6104 4834 6110 5210
rect 6144 4834 6150 5210
rect 6104 4822 6150 4834
rect 6222 5210 6268 5222
rect 6222 4834 6228 5210
rect 6262 4834 6268 5210
rect 6222 4822 6268 4834
rect 6340 5210 6386 5222
rect 6340 4834 6346 5210
rect 6380 4834 6386 5210
rect 6340 4822 6386 4834
rect 6458 5210 6504 5222
rect 6458 4834 6464 5210
rect 6498 4834 6504 5210
rect 6458 4822 6504 4834
rect 6576 5210 6622 5222
rect 6576 4834 6582 5210
rect 6616 4834 6622 5210
rect 6576 4822 6622 4834
rect 6694 5210 6740 5222
rect 6694 4834 6700 5210
rect 6734 5010 6740 5210
rect 7065 5022 7099 5325
rect 7524 5325 8997 5368
rect 7524 5022 7558 5325
rect 7890 5222 7924 5325
rect 8126 5222 8160 5325
rect 8362 5222 8396 5325
rect 8598 5222 8632 5325
rect 7884 5210 7930 5222
rect 6823 5010 6869 5022
rect 6734 4834 6829 5010
rect 6863 4834 6869 5010
rect 6694 4822 6740 4834
rect 6823 4822 6869 4834
rect 6941 5010 6987 5022
rect 6941 4834 6947 5010
rect 6981 4834 6987 5010
rect 6941 4822 6987 4834
rect 7059 5010 7105 5022
rect 7059 4834 7065 5010
rect 7099 4834 7105 5010
rect 7059 4822 7105 4834
rect 7177 5010 7223 5022
rect 7177 4834 7183 5010
rect 7217 4834 7223 5010
rect 7177 4822 7223 4834
rect 7400 5010 7446 5022
rect 7400 4834 7406 5010
rect 7440 4834 7446 5010
rect 7400 4822 7446 4834
rect 7518 5010 7564 5022
rect 7518 4834 7524 5010
rect 7558 4834 7564 5010
rect 7518 4822 7564 4834
rect 7636 5010 7682 5022
rect 7636 4834 7642 5010
rect 7676 4834 7682 5010
rect 7636 4822 7682 4834
rect 7754 5010 7800 5022
rect 7884 5010 7890 5210
rect 7754 4834 7760 5010
rect 7794 4834 7890 5010
rect 7924 4834 7930 5210
rect 7754 4822 7800 4834
rect 7884 4822 7930 4834
rect 8002 5210 8048 5222
rect 8002 4834 8008 5210
rect 8042 4834 8048 5210
rect 8002 4822 8048 4834
rect 8120 5210 8166 5222
rect 8120 4834 8126 5210
rect 8160 4834 8166 5210
rect 8120 4822 8166 4834
rect 8238 5210 8284 5222
rect 8238 4834 8244 5210
rect 8278 4834 8284 5210
rect 8238 4822 8284 4834
rect 8356 5210 8402 5222
rect 8356 4834 8362 5210
rect 8396 4834 8402 5210
rect 8356 4822 8402 4834
rect 8474 5210 8520 5222
rect 8474 4834 8480 5210
rect 8514 4834 8520 5210
rect 8474 4822 8520 4834
rect 8592 5210 8638 5222
rect 8592 4834 8598 5210
rect 8632 5010 8638 5210
rect 8963 5022 8997 5325
rect 8721 5010 8767 5022
rect 8632 4834 8727 5010
rect 8761 4834 8767 5010
rect 8592 4822 8638 4834
rect 8721 4822 8767 4834
rect 8839 5010 8885 5022
rect 8839 4834 8845 5010
rect 8879 4834 8885 5010
rect 8839 4822 8885 4834
rect 8957 5010 9003 5022
rect 8957 4834 8963 5010
rect 8997 4834 9003 5010
rect 8957 4822 9003 4834
rect 9075 5010 9121 5022
rect 9075 4834 9081 5010
rect 9115 4834 9121 5010
rect 9075 4822 9121 4834
rect 4873 4773 5013 4779
rect 5508 4788 5542 4822
rect 6110 4788 6144 4822
rect 6346 4788 6380 4822
rect 4765 4744 4873 4754
rect 5508 4753 5667 4788
rect 6110 4753 6380 4788
rect 6947 4788 6981 4822
rect 7183 4788 7217 4822
rect 6947 4753 7217 4788
rect 7406 4788 7440 4822
rect 8008 4788 8042 4822
rect 8244 4788 8278 4822
rect 7406 4753 7565 4788
rect 8008 4753 8278 4788
rect 8845 4788 8879 4822
rect 9081 4788 9115 4822
rect 8845 4753 9115 4788
rect 4138 4712 4153 4714
rect 4053 4698 4153 4712
rect 4053 4655 4153 4656
rect 3674 4634 4153 4655
rect 4442 4634 4508 4730
rect 3674 4586 4508 4634
rect 3674 4557 4153 4586
rect 3674 4555 3779 4557
rect 4053 4556 4153 4557
rect 3507 4370 3517 4449
rect 3610 4370 3620 4449
rect 4505 4440 4584 4452
rect 1844 4276 2550 4280
rect 1368 4264 1414 4276
rect 5 4125 1328 4136
rect 5 4044 16 4125
rect 103 4119 1328 4125
rect 103 4056 369 4119
rect 450 4056 1328 4119
rect 103 4044 1328 4056
rect 5 4038 1328 4044
rect 1252 4036 1328 4038
rect 8 4008 1152 4009
rect 8 4001 1216 4008
rect 8 3919 21 4001
rect 103 4000 1216 4001
rect 103 3919 499 4000
rect 601 3919 1216 4000
rect -661 3865 -650 3919
rect -594 3865 -584 3919
rect 8 3908 1216 3919
rect -3608 1776 -3408 1782
rect -3608 1742 -3596 1776
rect -3420 1742 -3339 1776
rect -3608 1736 -3408 1742
rect -3608 1658 -3408 1664
rect -3954 1624 -3596 1658
rect -3420 1624 -3408 1658
rect -3954 1292 -3911 1624
rect -3608 1618 -3408 1624
rect -3374 1651 -3339 1742
rect -3257 1772 -3190 1874
rect -661 1857 -586 3865
rect -661 1803 -650 1857
rect -594 1803 -584 1857
rect -661 1791 -586 1803
rect -3257 1757 -3191 1772
rect -3067 1769 -2995 1787
rect -3070 1704 -3061 1769
rect -3001 1704 -2991 1769
rect -3067 1703 -3061 1704
rect -3001 1703 -2995 1704
rect -3067 1691 -2995 1703
rect -3257 1681 -3191 1691
rect -2383 1651 -2183 1657
rect -3374 1617 -2371 1651
rect -2195 1617 -2183 1651
rect -3608 1540 -3408 1546
rect -3608 1506 -3596 1540
rect -3420 1506 -3408 1540
rect -3608 1500 -3408 1506
rect -3608 1422 -3408 1428
rect -3608 1388 -3596 1422
rect -3420 1388 -3408 1422
rect -3608 1382 -3408 1388
rect -3596 1298 -3420 1382
rect -3115 1349 -2715 1355
rect -3277 1315 -3103 1349
rect -2727 1315 -2715 1349
rect -2555 1335 -2512 1617
rect -2383 1611 -2183 1617
rect -2383 1534 -2183 1539
rect -2383 1533 -1857 1534
rect -2484 1504 -2422 1510
rect -2484 1470 -2472 1504
rect -2438 1470 -2422 1504
rect -2383 1499 -2371 1533
rect -2195 1500 -1857 1533
rect -2195 1499 -2183 1500
rect -2383 1493 -2183 1499
rect -2484 1454 -2422 1470
rect -3808 1292 -3408 1298
rect -3954 1258 -3796 1292
rect -3420 1258 -3408 1292
rect -3954 1056 -3911 1258
rect -3808 1252 -3408 1258
rect -3808 1174 -3408 1180
rect -3808 1140 -3796 1174
rect -3420 1140 -3339 1174
rect -3808 1134 -3408 1140
rect -3808 1056 -3408 1062
rect -3954 1022 -3796 1056
rect -3420 1022 -3408 1056
rect -3954 987 -3911 1022
rect -3808 1016 -3408 1022
rect -4037 959 -3911 987
rect -4059 949 -3911 959
rect -4005 895 -3911 949
rect -3808 938 -3408 944
rect -3374 938 -3339 1140
rect -3277 1113 -3239 1315
rect -3115 1309 -2715 1315
rect -2550 1319 -2499 1335
rect -2550 1285 -2539 1319
rect -2505 1285 -2499 1319
rect -2550 1268 -2499 1285
rect -3115 1231 -2715 1237
rect -3115 1197 -3103 1231
rect -2727 1197 -2715 1231
rect -3115 1191 -2715 1197
rect -3115 1113 -2715 1119
rect -3277 1079 -3103 1113
rect -2727 1079 -2715 1113
rect -3277 938 -3239 1079
rect -3115 1073 -2715 1079
rect -2471 1069 -2422 1454
rect -2383 1231 -1983 1237
rect -2383 1197 -2371 1231
rect -1995 1197 -1983 1231
rect -2383 1191 -1983 1197
rect -2383 1113 -1983 1119
rect -2383 1079 -2371 1113
rect -1995 1079 -1983 1113
rect -2383 1073 -1983 1079
rect -2471 1053 -2414 1069
rect -2471 1019 -2455 1053
rect -2421 1019 -2414 1053
rect -2471 1003 -2414 1019
rect -1889 1041 -1857 1500
rect -1889 1007 -1772 1041
rect -3115 995 -2715 1001
rect -3115 961 -3103 995
rect -2727 961 -2715 995
rect -3115 955 -2715 961
rect -2383 995 -1983 1001
rect -2383 961 -2371 995
rect -1995 961 -1983 995
rect -2383 955 -1983 961
rect -3808 904 -3796 938
rect -3420 904 -3239 938
rect -3808 898 -3408 904
rect -4059 885 -3911 895
rect -4037 853 -3911 885
rect -3954 820 -3911 853
rect -3277 877 -3239 904
rect -2471 935 -2412 951
rect -2471 901 -2456 935
rect -2422 901 -2412 935
rect -2471 884 -2412 901
rect -1889 945 -1835 1007
rect -1777 945 -1772 1007
rect -1889 909 -1772 945
rect 772 1028 890 3908
rect 1138 3759 1192 3908
rect 1252 3844 1306 4036
rect 1368 3888 1374 4264
rect 1408 3888 1414 4264
rect 1368 3876 1414 3888
rect 1486 4264 1532 4276
rect 1486 3888 1492 4264
rect 1526 3888 1532 4264
rect 1486 3876 1532 3888
rect 1604 4264 1650 4276
rect 1604 3888 1610 4264
rect 1644 3915 1650 4264
rect 1721 4264 1767 4276
rect 1721 4088 1727 4264
rect 1761 4088 1767 4264
rect 1721 4081 1767 4088
rect 1839 4264 2550 4276
rect 1839 4088 1845 4264
rect 1879 4251 2550 4264
rect 1879 4088 1885 4251
rect 2129 4172 2550 4251
rect 2129 4171 2233 4172
rect 1721 4076 1770 4081
rect 1839 4076 1885 4088
rect 1727 3915 1770 4076
rect 1644 3888 1770 3915
rect 1604 3876 1770 3888
rect 1610 3872 1770 3876
rect 1252 3838 1483 3844
rect 1252 3804 1433 3838
rect 1467 3804 1483 3838
rect 1252 3788 1483 3804
rect 1535 3838 1601 3844
rect 1535 3804 1551 3838
rect 1585 3804 1601 3838
rect 1535 3759 1601 3804
rect 1138 3751 1601 3759
rect 1138 3719 1602 3751
rect 1694 3735 1770 3872
rect 1690 3675 1700 3735
rect 1762 3675 1772 3735
rect 3518 3196 3611 4370
rect 4505 4341 4511 4440
rect 4436 4321 4511 4341
rect 4578 4341 4584 4440
rect 4578 4321 4656 4341
rect 4436 4213 4480 4321
rect 4612 4213 4656 4321
rect 4436 4171 4656 4213
rect 4040 4141 5017 4171
rect 4040 4035 4072 4141
rect 4276 4035 4308 4141
rect 4512 4035 4544 4141
rect 4748 4035 4780 4141
rect 4983 4035 5017 4141
rect 4033 4023 4079 4035
rect 4033 3847 4039 4023
rect 4073 3847 4079 4023
rect 4033 3835 4079 3847
rect 4151 4023 4197 4035
rect 4151 3847 4157 4023
rect 4191 3847 4197 4023
rect 4151 3835 4197 3847
rect 4269 4023 4315 4035
rect 4269 3847 4275 4023
rect 4309 3847 4315 4023
rect 4269 3835 4315 3847
rect 4387 4023 4433 4035
rect 4387 3847 4393 4023
rect 4427 3847 4433 4023
rect 4387 3835 4433 3847
rect 4505 4023 4551 4035
rect 4505 3847 4511 4023
rect 4545 3847 4551 4023
rect 4505 3835 4551 3847
rect 4623 4023 4669 4035
rect 4623 3847 4629 4023
rect 4663 3847 4669 4023
rect 4623 3835 4669 3847
rect 4741 4023 4787 4035
rect 4741 3847 4747 4023
rect 4781 3847 4787 4023
rect 4741 3835 4787 3847
rect 4859 4023 4905 4035
rect 4859 3847 4865 4023
rect 4899 3847 4905 4023
rect 4859 3835 4905 3847
rect 4977 4023 5023 4035
rect 4977 3847 4983 4023
rect 5017 3847 5023 4023
rect 4977 3835 5023 3847
rect 5095 4023 5141 4035
rect 5095 3847 5101 4023
rect 5135 3847 5141 4023
rect 5095 3835 5141 3847
rect 5633 3969 5667 4753
rect 6346 4691 6380 4753
rect 5935 4653 6677 4691
rect 5935 4529 5969 4653
rect 6171 4529 6205 4653
rect 6407 4529 6441 4653
rect 6643 4529 6677 4653
rect 6933 4546 6943 4612
rect 7006 4546 7016 4612
rect 5929 4517 5975 4529
rect 5929 4141 5935 4517
rect 5969 4141 5975 4517
rect 5929 4129 5975 4141
rect 6047 4517 6093 4529
rect 6047 4141 6053 4517
rect 6087 4141 6093 4517
rect 6047 4129 6093 4141
rect 6165 4517 6211 4529
rect 6165 4141 6171 4517
rect 6205 4141 6211 4517
rect 6165 4129 6211 4141
rect 6283 4517 6329 4529
rect 6283 4141 6289 4517
rect 6323 4141 6329 4517
rect 6283 4129 6329 4141
rect 6401 4517 6447 4529
rect 6401 4141 6407 4517
rect 6441 4141 6447 4517
rect 6401 4129 6447 4141
rect 6519 4517 6565 4529
rect 6519 4141 6525 4517
rect 6559 4141 6565 4517
rect 6519 4129 6565 4141
rect 6637 4517 6683 4529
rect 6637 4141 6643 4517
rect 6677 4141 6683 4517
rect 6637 4129 6683 4141
rect 7049 3970 7083 4753
rect 6776 3969 7083 3970
rect 5633 3964 5949 3969
rect 6663 3964 7083 3969
rect 5633 3953 6016 3964
rect 5633 3926 5965 3953
rect 4156 3741 4192 3835
rect 4392 3741 4428 3835
rect 4628 3742 4664 3835
rect 4790 3787 4856 3794
rect 4790 3753 4806 3787
rect 4840 3753 4856 3787
rect 4790 3742 4856 3753
rect 4628 3741 4856 3742
rect 4156 3712 4856 3741
rect 4156 3711 4738 3712
rect 4276 3598 4310 3711
rect 4672 3670 4738 3711
rect 4672 3636 4688 3670
rect 4722 3636 4738 3670
rect 4672 3629 4738 3636
rect 5100 3602 5135 3835
rect 5633 3797 5667 3926
rect 5949 3919 5965 3926
rect 5999 3919 6016 3953
rect 5949 3913 6016 3919
rect 6596 3953 7083 3964
rect 6596 3919 6613 3953
rect 6647 3926 7083 3953
rect 6647 3919 6663 3926
rect 6776 3925 7083 3926
rect 6596 3913 6663 3919
rect 5774 3886 5830 3898
rect 5774 3852 5780 3886
rect 5814 3885 5830 3886
rect 6887 3885 6943 3897
rect 5814 3869 6281 3885
rect 5814 3852 6231 3869
rect 5774 3836 6231 3852
rect 6215 3835 6231 3836
rect 6265 3835 6281 3869
rect 6215 3828 6281 3835
rect 6333 3870 6903 3885
rect 6333 3836 6349 3870
rect 6383 3851 6903 3870
rect 6937 3851 6943 3885
rect 6383 3836 6943 3851
rect 6333 3826 6400 3836
rect 6887 3835 6943 3836
rect 7049 3797 7083 3925
rect 7531 3969 7565 4753
rect 8244 4691 8278 4753
rect 7833 4653 8575 4691
rect 7833 4529 7867 4653
rect 8069 4529 8103 4653
rect 8305 4529 8339 4653
rect 8541 4529 8575 4653
rect 7827 4517 7873 4529
rect 7827 4141 7833 4517
rect 7867 4141 7873 4517
rect 7827 4129 7873 4141
rect 7945 4517 7991 4529
rect 7945 4141 7951 4517
rect 7985 4141 7991 4517
rect 7945 4129 7991 4141
rect 8063 4517 8109 4529
rect 8063 4141 8069 4517
rect 8103 4141 8109 4517
rect 8063 4129 8109 4141
rect 8181 4517 8227 4529
rect 8181 4141 8187 4517
rect 8221 4141 8227 4517
rect 8181 4129 8227 4141
rect 8299 4517 8345 4529
rect 8299 4141 8305 4517
rect 8339 4141 8345 4517
rect 8299 4129 8345 4141
rect 8417 4517 8463 4529
rect 8417 4141 8423 4517
rect 8457 4141 8463 4517
rect 8417 4129 8463 4141
rect 8535 4517 8581 4529
rect 8535 4141 8541 4517
rect 8575 4141 8581 4517
rect 8535 4129 8581 4141
rect 8947 3970 8981 4753
rect 8559 3969 8628 3970
rect 8674 3969 8981 3970
rect 7531 3964 7847 3969
rect 8559 3965 8981 3969
rect 7531 3953 7914 3964
rect 7531 3926 7863 3953
rect 7531 3797 7565 3926
rect 7847 3919 7863 3926
rect 7897 3919 7914 3953
rect 7847 3913 7914 3919
rect 8492 3954 8981 3965
rect 8492 3920 8509 3954
rect 8543 3926 8981 3954
rect 8543 3920 8559 3926
rect 8674 3925 8981 3926
rect 8492 3914 8559 3920
rect 7672 3886 7728 3898
rect 7672 3852 7678 3886
rect 7712 3885 7728 3886
rect 8785 3885 8841 3897
rect 7712 3869 8179 3885
rect 7712 3852 8129 3869
rect 7672 3836 8129 3852
rect 8113 3835 8129 3836
rect 8163 3835 8179 3869
rect 8113 3828 8179 3835
rect 8231 3870 8801 3885
rect 8231 3836 8247 3870
rect 8281 3851 8801 3870
rect 8835 3851 8841 3885
rect 8281 3836 8841 3851
rect 8231 3826 8298 3836
rect 8785 3835 8841 3836
rect 8947 3797 8981 3925
rect 9062 4575 9129 4599
rect 9062 4541 9079 4575
rect 9113 4541 9129 4575
rect 4746 3598 5135 3602
rect 4270 3586 4316 3598
rect 4270 3210 4276 3586
rect 4310 3210 4316 3586
rect 4270 3198 4316 3210
rect 4388 3586 4434 3598
rect 4388 3210 4394 3586
rect 4428 3210 4434 3586
rect 4388 3198 4434 3210
rect 4506 3586 4552 3598
rect 4506 3210 4512 3586
rect 4546 3234 4552 3586
rect 4623 3586 4669 3598
rect 4623 3410 4629 3586
rect 4663 3410 4669 3586
rect 4623 3398 4669 3410
rect 4741 3586 5135 3598
rect 5627 3785 5673 3797
rect 5627 3609 5633 3785
rect 5667 3609 5673 3785
rect 5627 3597 5673 3609
rect 5745 3785 5791 3797
rect 5745 3609 5751 3785
rect 5785 3609 5791 3785
rect 5745 3597 5791 3609
rect 6047 3785 6093 3797
rect 4741 3410 4747 3586
rect 4781 3573 5135 3586
rect 4781 3410 4787 3573
rect 5057 3570 5135 3573
rect 5057 3518 5067 3570
rect 5130 3518 5140 3570
rect 5062 3512 5135 3518
rect 4741 3398 4787 3410
rect 4629 3282 4664 3398
rect 5750 3303 5784 3597
rect 6047 3409 6053 3785
rect 6087 3409 6093 3785
rect 6047 3397 6093 3409
rect 6165 3785 6211 3797
rect 6165 3409 6171 3785
rect 6205 3409 6211 3785
rect 6165 3397 6211 3409
rect 6283 3785 6329 3797
rect 6283 3409 6289 3785
rect 6323 3409 6329 3785
rect 6283 3397 6329 3409
rect 6401 3785 6447 3797
rect 6401 3409 6407 3785
rect 6441 3409 6447 3785
rect 6401 3397 6447 3409
rect 6519 3785 6565 3797
rect 6519 3409 6525 3785
rect 6559 3409 6565 3785
rect 6925 3785 6971 3797
rect 6925 3609 6931 3785
rect 6965 3609 6971 3785
rect 6925 3597 6971 3609
rect 7043 3785 7089 3797
rect 7043 3609 7049 3785
rect 7083 3609 7089 3785
rect 7043 3597 7089 3609
rect 7525 3785 7571 3797
rect 7525 3609 7531 3785
rect 7565 3609 7571 3785
rect 7525 3597 7571 3609
rect 7643 3785 7689 3797
rect 7643 3609 7649 3785
rect 7683 3609 7689 3785
rect 7643 3597 7689 3609
rect 7945 3785 7991 3797
rect 6519 3397 6565 3409
rect 6407 3303 6441 3397
rect 6931 3303 6964 3597
rect 4760 3282 4868 3292
rect 4629 3234 4760 3282
rect 5750 3271 6964 3303
rect 7648 3303 7682 3597
rect 7945 3409 7951 3785
rect 7985 3409 7991 3785
rect 7945 3397 7991 3409
rect 8063 3785 8109 3797
rect 8063 3409 8069 3785
rect 8103 3409 8109 3785
rect 8063 3397 8109 3409
rect 8181 3785 8227 3797
rect 8181 3409 8187 3785
rect 8221 3409 8227 3785
rect 8181 3397 8227 3409
rect 8299 3785 8345 3797
rect 8299 3409 8305 3785
rect 8339 3409 8345 3785
rect 8299 3397 8345 3409
rect 8417 3785 8463 3797
rect 8417 3409 8423 3785
rect 8457 3409 8463 3785
rect 8823 3785 8869 3797
rect 8823 3609 8829 3785
rect 8863 3609 8869 3785
rect 8823 3597 8869 3609
rect 8941 3785 8987 3797
rect 8941 3609 8947 3785
rect 8981 3609 8987 3785
rect 8941 3597 8987 3609
rect 8417 3397 8463 3409
rect 8305 3303 8339 3397
rect 8829 3303 8862 3597
rect 7648 3271 8862 3303
rect 4868 3254 5013 3260
rect 4546 3210 4760 3234
rect 4506 3198 4760 3210
rect 3518 3194 4103 3196
rect 4512 3194 4760 3198
rect 3518 3166 4148 3194
rect 3518 3160 4385 3166
rect 3518 3126 4335 3160
rect 4369 3126 4385 3160
rect 3518 3110 4385 3126
rect 4437 3160 4503 3166
rect 4437 3126 4453 3160
rect 4487 3126 4503 3160
rect 4686 3150 4760 3194
rect 5001 3187 5013 3254
rect 4868 3181 5013 3187
rect 6243 3186 6375 3271
rect 8141 3186 8273 3271
rect 4760 3140 4868 3150
rect 3518 3094 4148 3110
rect 3518 3090 4103 3094
rect 3518 3089 3619 3090
rect 4048 3041 4148 3052
rect 4012 2935 4022 3041
rect 4134 3030 4148 3041
rect 4437 3030 4503 3126
rect 6233 3078 6243 3186
rect 6375 3078 6385 3186
rect 8131 3078 8141 3186
rect 8273 3078 8283 3186
rect 9062 3158 9129 4541
rect 9190 4112 9348 6339
rect 9190 4014 9202 4112
rect 9334 4037 9348 4112
rect 9432 5930 9946 5954
rect 9432 5824 9794 5930
rect 9906 5917 9946 5930
rect 9906 5824 9948 5917
rect 9432 5813 9948 5824
rect 9432 5812 9946 5813
rect 9334 4014 9346 4037
rect 9190 4008 9346 4014
rect 4134 2982 4503 3030
rect 4134 2952 4148 2982
rect 4134 2935 4144 2952
rect 4436 2879 4502 2982
rect 6267 2937 6273 3078
rect 6340 2937 6346 3078
rect 6267 2925 6346 2937
rect 9062 2879 9128 3158
rect 4434 2799 9128 2879
rect 7848 2294 8312 2326
rect 8400 2310 8410 2370
rect 8472 2310 8482 2370
rect 7848 2286 8311 2294
rect 7848 2137 7902 2286
rect 7463 2131 7902 2137
rect 7461 2045 7471 2131
rect 7547 2045 7902 2131
rect 7463 2037 7902 2045
rect 7962 2241 8193 2257
rect 7962 2207 8143 2241
rect 8177 2207 8193 2241
rect 7962 2201 8193 2207
rect 8245 2241 8311 2286
rect 8245 2207 8261 2241
rect 8295 2207 8311 2241
rect 8245 2201 8311 2207
rect 7962 2009 8016 2201
rect 8404 2173 8480 2310
rect 8320 2169 8480 2173
rect 7698 2004 8016 2009
rect 7692 1913 7702 2004
rect 7831 1913 8016 2004
rect 7698 1909 8016 1913
rect 8078 2157 8124 2169
rect 8078 1781 8084 2157
rect 8118 1781 8124 2157
rect 8078 1769 8124 1781
rect 8196 2157 8242 2169
rect 8196 1781 8202 2157
rect 8236 1781 8242 2157
rect 8196 1769 8242 1781
rect 8314 2157 8480 2169
rect 8314 1781 8320 2157
rect 8354 2130 8480 2157
rect 8354 1781 8360 2130
rect 8437 1969 8480 2130
rect 8314 1769 8360 1781
rect 8431 1964 8480 1969
rect 8431 1957 8477 1964
rect 8431 1781 8437 1957
rect 8471 1781 8477 1957
rect 8431 1769 8477 1781
rect 8549 1957 8595 1969
rect 8549 1781 8555 1957
rect 8589 1794 8595 1957
rect 9432 1874 9568 5812
rect 10069 4447 10162 6339
rect 10225 6282 10691 6304
rect 10979 6282 11045 6378
rect 12810 6388 12816 6564
rect 12850 6388 12856 6564
rect 12810 6376 12856 6388
rect 12928 6564 12974 6576
rect 12928 6388 12934 6564
rect 12968 6388 12974 6564
rect 12928 6376 12974 6388
rect 13046 6564 13092 6576
rect 13046 6388 13052 6564
rect 13086 6388 13092 6564
rect 13046 6376 13092 6388
rect 13164 6564 13210 6576
rect 13164 6388 13170 6564
rect 13204 6509 13210 6564
rect 13329 6564 13375 6576
rect 13329 6509 13335 6564
rect 13204 6421 13335 6509
rect 13204 6388 13210 6421
rect 13164 6376 13210 6388
rect 13329 6388 13335 6421
rect 13369 6388 13375 6564
rect 13329 6376 13375 6388
rect 13447 6564 13493 6576
rect 13447 6388 13453 6564
rect 13487 6388 13493 6564
rect 13447 6376 13493 6388
rect 13565 6564 13611 6576
rect 13565 6388 13571 6564
rect 13605 6388 13611 6564
rect 13565 6376 13611 6388
rect 13683 6564 13729 6576
rect 13683 6388 13689 6564
rect 13723 6388 13729 6564
rect 13683 6376 13729 6388
rect 12816 6337 12850 6376
rect 13052 6337 13086 6376
rect 12816 6302 13086 6337
rect 13453 6338 13486 6376
rect 13689 6338 13722 6376
rect 13453 6302 13722 6338
rect 10225 6234 11045 6282
rect 12850 6301 13086 6302
rect 10225 6203 10691 6234
rect 12850 6227 12982 6301
rect 10225 5947 10330 6203
rect 12840 6119 12850 6227
rect 12982 6119 12992 6227
rect 11061 6046 11140 6058
rect 10225 5841 10288 5947
rect 10400 5841 10410 5947
rect 11061 5943 11067 6046
rect 10992 5923 11067 5943
rect 11134 5943 11140 6046
rect 12873 5983 12879 6119
rect 12946 5983 12952 6119
rect 12873 5971 12952 5983
rect 11134 5923 11212 5943
rect 10225 5830 10374 5841
rect 10225 4653 10330 5830
rect 10992 5815 11036 5923
rect 11168 5815 11212 5923
rect 10992 5773 11212 5815
rect 13790 5788 13852 7359
rect 14042 7351 14088 7363
rect 14042 6975 14048 7351
rect 14082 6975 14088 7351
rect 14042 6963 14088 6975
rect 14160 7351 14206 7363
rect 14160 6975 14166 7351
rect 14200 6975 14206 7351
rect 14160 6963 14206 6975
rect 14278 7351 14324 7363
rect 14278 6975 14284 7351
rect 14318 6975 14324 7351
rect 14278 6963 14324 6975
rect 14396 7351 14442 7363
rect 14396 6975 14402 7351
rect 14436 6975 14442 7351
rect 14396 6963 14442 6975
rect 14514 7351 14560 7363
rect 14514 6975 14520 7351
rect 14554 6975 14560 7351
rect 14514 6963 14560 6975
rect 14632 7351 14678 7363
rect 14632 6975 14638 7351
rect 14672 6975 14678 7351
rect 14632 6963 14678 6975
rect 14750 7351 14796 7363
rect 14750 6975 14756 7351
rect 14790 6975 14796 7351
rect 14750 6963 14796 6975
rect 14048 6921 14082 6963
rect 14284 6921 14318 6963
rect 14048 6893 14318 6921
rect 14402 6922 14436 6963
rect 14638 6922 14672 6963
rect 14402 6893 14672 6922
rect 14048 6845 14082 6893
rect 14048 6815 14111 6845
rect 14076 6723 14111 6815
rect 14583 6785 14683 6806
rect 14583 6731 14597 6785
rect 14662 6731 14683 6785
rect 14583 6726 14683 6731
rect 14756 6780 14790 6963
rect 14756 6726 14865 6780
rect 14076 6687 14303 6723
rect 14076 6580 14111 6687
rect 14237 6653 14303 6687
rect 14237 6619 14253 6653
rect 14287 6619 14303 6653
rect 14584 6711 14681 6726
rect 14584 6644 14641 6711
rect 14237 6613 14303 6619
rect 14478 6608 14747 6644
rect 14478 6580 14511 6608
rect 14714 6580 14747 6608
rect 14831 6580 14865 6726
rect 13952 6568 13998 6580
rect 13952 6392 13958 6568
rect 13992 6392 13998 6568
rect 13952 6380 13998 6392
rect 14070 6568 14116 6580
rect 14070 6392 14076 6568
rect 14110 6392 14116 6568
rect 14070 6380 14116 6392
rect 14188 6568 14234 6580
rect 14188 6392 14194 6568
rect 14228 6392 14234 6568
rect 14188 6380 14234 6392
rect 14306 6568 14352 6580
rect 14306 6392 14312 6568
rect 14346 6513 14352 6568
rect 14471 6568 14517 6580
rect 14471 6513 14477 6568
rect 14346 6425 14477 6513
rect 14346 6392 14352 6425
rect 14306 6380 14352 6392
rect 14471 6392 14477 6425
rect 14511 6392 14517 6568
rect 14471 6380 14517 6392
rect 14589 6568 14635 6580
rect 14589 6392 14595 6568
rect 14629 6392 14635 6568
rect 14589 6380 14635 6392
rect 14707 6568 14753 6580
rect 14707 6392 14713 6568
rect 14747 6392 14753 6568
rect 14707 6380 14753 6392
rect 14825 6568 14871 6580
rect 14825 6392 14831 6568
rect 14865 6392 14871 6568
rect 14825 6380 14871 6392
rect 16020 6447 16160 12588
rect 16589 12296 16771 13784
rect 20190 13546 20269 13558
rect 17709 13490 17788 13502
rect 17709 13395 17715 13490
rect 17638 13375 17715 13395
rect 17782 13395 17788 13490
rect 20190 13429 20196 13546
rect 20263 13429 20269 13546
rect 21337 13545 21416 13557
rect 21337 13429 21343 13545
rect 21410 13429 21416 13545
rect 17782 13375 17858 13395
rect 17638 13267 17682 13375
rect 17814 13267 17858 13375
rect 19435 13333 19491 13341
rect 17638 13225 17858 13267
rect 18509 13325 19491 13333
rect 18509 13291 19451 13325
rect 19485 13291 19491 13325
rect 20154 13321 20164 13429
rect 20296 13366 20306 13429
rect 20296 13355 20308 13366
rect 20296 13321 20309 13355
rect 20565 13345 20621 13347
rect 18509 13275 19491 13291
rect 20164 13283 20309 13321
rect 18509 13274 19488 13275
rect 17242 13195 18219 13225
rect 17242 13089 17274 13195
rect 17478 13089 17510 13195
rect 17714 13089 17746 13195
rect 17950 13089 17982 13195
rect 18185 13089 18219 13195
rect 17235 13077 17281 13089
rect 17235 12901 17241 13077
rect 17275 12901 17281 13077
rect 17235 12889 17281 12901
rect 17353 13077 17399 13089
rect 17353 12901 17359 13077
rect 17393 12901 17399 13077
rect 17353 12889 17399 12901
rect 17471 13077 17517 13089
rect 17471 12901 17477 13077
rect 17511 12901 17517 13077
rect 17471 12889 17517 12901
rect 17589 13077 17635 13089
rect 17589 12901 17595 13077
rect 17629 12901 17635 13077
rect 17589 12889 17635 12901
rect 17707 13077 17753 13089
rect 17707 12901 17713 13077
rect 17747 12901 17753 13077
rect 17707 12889 17753 12901
rect 17825 13077 17871 13089
rect 17825 12901 17831 13077
rect 17865 12901 17871 13077
rect 17825 12889 17871 12901
rect 17943 13077 17989 13089
rect 17943 12901 17949 13077
rect 17983 12901 17989 13077
rect 17943 12889 17989 12901
rect 18061 13077 18107 13089
rect 18061 12901 18067 13077
rect 18101 12901 18107 13077
rect 18061 12889 18107 12901
rect 18179 13077 18225 13089
rect 18179 12901 18185 13077
rect 18219 12901 18225 13077
rect 18179 12889 18225 12901
rect 18297 13077 18343 13089
rect 18297 12901 18303 13077
rect 18337 12901 18343 13077
rect 18297 12889 18343 12901
rect 17358 12795 17394 12889
rect 17594 12795 17630 12889
rect 17830 12796 17866 12889
rect 17992 12841 18058 12848
rect 17992 12807 18008 12841
rect 18042 12807 18058 12841
rect 17992 12796 18058 12807
rect 17830 12795 18058 12796
rect 17358 12766 18058 12795
rect 17358 12765 17940 12766
rect 17478 12652 17512 12765
rect 17874 12724 17940 12765
rect 17874 12690 17890 12724
rect 17924 12690 17940 12724
rect 17874 12683 17940 12690
rect 18302 12684 18337 12889
rect 18509 12684 18576 13274
rect 20268 13251 20309 13283
rect 20555 13279 20565 13345
rect 20621 13279 20631 13345
rect 21301 13321 21311 13429
rect 21443 13366 21453 13429
rect 21443 13355 21455 13366
rect 21443 13321 21456 13355
rect 21311 13283 21456 13321
rect 21415 13255 21456 13283
rect 19684 13223 19954 13251
rect 19425 13157 19435 13223
rect 19501 13157 19511 13223
rect 19684 13161 19718 13223
rect 19920 13161 19954 13223
rect 20038 13223 20309 13251
rect 20826 13227 21096 13255
rect 20038 13161 20072 13223
rect 20274 13161 20309 13223
rect 20450 13211 20621 13227
rect 20450 13177 20581 13211
rect 20615 13177 20621 13211
rect 20450 13161 20621 13177
rect 20826 13165 20860 13227
rect 21062 13165 21096 13227
rect 21180 13227 21456 13255
rect 21180 13165 21214 13227
rect 21416 13165 21456 13227
rect 19560 13149 19606 13161
rect 19560 12773 19566 13149
rect 19600 12773 19606 13149
rect 19560 12761 19606 12773
rect 19678 13149 19724 13161
rect 19678 12773 19684 13149
rect 19718 12773 19724 13149
rect 19678 12761 19724 12773
rect 19796 13149 19842 13161
rect 19796 12773 19802 13149
rect 19836 12773 19842 13149
rect 19796 12761 19842 12773
rect 19914 13149 19960 13161
rect 19914 12773 19920 13149
rect 19954 12773 19960 13149
rect 19914 12761 19960 12773
rect 20032 13149 20078 13161
rect 20032 12773 20038 13149
rect 20072 12773 20078 13149
rect 20032 12761 20078 12773
rect 20150 13149 20196 13161
rect 20150 12773 20156 13149
rect 20190 12773 20196 13149
rect 20150 12761 20196 12773
rect 20268 13149 20314 13161
rect 20268 12773 20274 13149
rect 20308 12773 20314 13149
rect 20268 12761 20314 12773
rect 18302 12656 18576 12684
rect 17948 12652 18576 12656
rect 16588 12247 16771 12296
rect 17472 12640 17518 12652
rect 17472 12264 17478 12640
rect 17512 12264 17518 12640
rect 17472 12252 17518 12264
rect 17590 12640 17636 12652
rect 17590 12264 17596 12640
rect 17630 12264 17636 12640
rect 17590 12252 17636 12264
rect 17708 12640 17754 12652
rect 17708 12264 17714 12640
rect 17748 12288 17754 12640
rect 17825 12640 17871 12652
rect 17825 12464 17831 12640
rect 17865 12464 17871 12640
rect 17825 12452 17871 12464
rect 17943 12640 18576 12652
rect 17943 12464 17949 12640
rect 17983 12627 18576 12640
rect 19566 12719 19600 12761
rect 19802 12719 19836 12761
rect 19566 12691 19836 12719
rect 19920 12720 19954 12761
rect 20156 12720 20190 12761
rect 19920 12691 20190 12720
rect 19566 12643 19600 12691
rect 17983 12464 17989 12627
rect 19566 12613 19629 12643
rect 17943 12452 17989 12464
rect 19594 12521 19629 12613
rect 19594 12485 19821 12521
rect 20091 12510 20101 12607
rect 20200 12510 20210 12607
rect 20274 12578 20308 12761
rect 20274 12524 20383 12578
rect 17831 12336 17866 12452
rect 19594 12378 19629 12485
rect 19755 12451 19821 12485
rect 19755 12417 19771 12451
rect 19805 12417 19821 12451
rect 20102 12509 20199 12510
rect 20102 12442 20159 12509
rect 19755 12411 19821 12417
rect 19996 12406 20265 12442
rect 19996 12378 20029 12406
rect 20232 12378 20265 12406
rect 20349 12378 20383 12524
rect 19470 12366 19516 12378
rect 17962 12336 18070 12346
rect 17831 12288 17962 12336
rect 18070 12299 18211 12305
rect 17748 12264 17962 12288
rect 17708 12252 17962 12264
rect 17714 12248 17962 12252
rect 16588 12220 17350 12247
rect 16588 12214 17587 12220
rect 16588 12180 17537 12214
rect 17571 12180 17587 12214
rect 16588 12164 17587 12180
rect 17639 12214 17705 12220
rect 17639 12180 17655 12214
rect 17689 12180 17705 12214
rect 17888 12204 17962 12248
rect 18199 12232 18211 12299
rect 18070 12226 18211 12232
rect 17962 12194 18070 12204
rect 16588 12148 17350 12164
rect 16588 12147 17287 12148
rect 16588 12143 16822 12147
rect 16440 10630 16605 10650
rect 16440 10513 16452 10630
rect 16591 10607 16605 10630
rect 16591 10513 16606 10607
rect 16440 10512 16459 10513
rect 16571 10512 16606 10513
rect 16440 10503 16606 10512
rect 16440 10502 16605 10503
rect 16440 10501 16573 10502
rect 16729 10249 16822 12143
rect 16885 12084 17351 12106
rect 17639 12084 17705 12180
rect 19470 12190 19476 12366
rect 19510 12190 19516 12366
rect 19470 12178 19516 12190
rect 19588 12366 19634 12378
rect 19588 12190 19594 12366
rect 19628 12190 19634 12366
rect 19588 12178 19634 12190
rect 19706 12366 19752 12378
rect 19706 12190 19712 12366
rect 19746 12190 19752 12366
rect 19706 12178 19752 12190
rect 19824 12366 19870 12378
rect 19824 12190 19830 12366
rect 19864 12311 19870 12366
rect 19989 12366 20035 12378
rect 19989 12311 19995 12366
rect 19864 12223 19995 12311
rect 19864 12190 19870 12223
rect 19824 12178 19870 12190
rect 19989 12190 19995 12223
rect 20029 12190 20035 12366
rect 19989 12178 20035 12190
rect 20107 12366 20153 12378
rect 20107 12190 20113 12366
rect 20147 12190 20153 12366
rect 20107 12178 20153 12190
rect 20225 12366 20271 12378
rect 20225 12190 20231 12366
rect 20265 12190 20271 12366
rect 20225 12178 20271 12190
rect 20343 12366 20389 12378
rect 20343 12190 20349 12366
rect 20383 12190 20389 12366
rect 20343 12178 20389 12190
rect 19476 12139 19510 12178
rect 19712 12139 19746 12178
rect 19476 12104 19746 12139
rect 20113 12140 20146 12178
rect 20349 12140 20382 12178
rect 20113 12104 20382 12140
rect 16885 12036 17705 12084
rect 19510 12103 19746 12104
rect 16885 12005 17351 12036
rect 19510 12029 19642 12103
rect 16885 11749 16990 12005
rect 19500 11921 19510 12029
rect 19642 11921 19652 12029
rect 17724 11842 17803 11854
rect 16885 11643 16948 11749
rect 17060 11643 17070 11749
rect 17724 11745 17730 11842
rect 17652 11725 17730 11745
rect 17797 11745 17803 11842
rect 19532 11787 19538 11921
rect 19605 11787 19611 11921
rect 19532 11775 19611 11787
rect 17797 11725 17872 11745
rect 16885 11632 17034 11643
rect 16885 10455 16990 11632
rect 17652 11617 17696 11725
rect 17828 11617 17872 11725
rect 17652 11575 17872 11617
rect 20450 11590 20512 13161
rect 20702 13153 20748 13165
rect 20702 12777 20708 13153
rect 20742 12777 20748 13153
rect 20702 12765 20748 12777
rect 20820 13153 20866 13165
rect 20820 12777 20826 13153
rect 20860 12777 20866 13153
rect 20820 12765 20866 12777
rect 20938 13153 20984 13165
rect 20938 12777 20944 13153
rect 20978 12777 20984 13153
rect 20938 12765 20984 12777
rect 21056 13153 21102 13165
rect 21056 12777 21062 13153
rect 21096 12777 21102 13153
rect 21056 12765 21102 12777
rect 21174 13153 21220 13165
rect 21174 12777 21180 13153
rect 21214 12777 21220 13153
rect 21174 12765 21220 12777
rect 21292 13153 21338 13165
rect 21292 12777 21298 13153
rect 21332 12777 21338 13153
rect 21292 12765 21338 12777
rect 21410 13153 21456 13165
rect 21410 12777 21416 13153
rect 21450 12777 21456 13153
rect 21410 12765 21456 12777
rect 20708 12723 20742 12765
rect 20944 12723 20978 12765
rect 20708 12695 20978 12723
rect 21062 12724 21096 12765
rect 21298 12724 21332 12765
rect 21062 12695 21332 12724
rect 20708 12647 20742 12695
rect 20708 12617 20771 12647
rect 20736 12525 20771 12617
rect 21243 12587 21343 12608
rect 21243 12533 21257 12587
rect 21322 12533 21343 12587
rect 21243 12528 21343 12533
rect 21416 12582 21450 12765
rect 21416 12528 21525 12582
rect 20736 12489 20963 12525
rect 20736 12382 20771 12489
rect 20897 12455 20963 12489
rect 20897 12421 20913 12455
rect 20947 12421 20963 12455
rect 21244 12513 21341 12528
rect 21244 12446 21301 12513
rect 20897 12415 20963 12421
rect 21138 12410 21407 12446
rect 21138 12382 21171 12410
rect 21374 12382 21407 12410
rect 21491 12382 21525 12528
rect 20612 12370 20658 12382
rect 20612 12194 20618 12370
rect 20652 12194 20658 12370
rect 20612 12182 20658 12194
rect 20730 12370 20776 12382
rect 20730 12194 20736 12370
rect 20770 12194 20776 12370
rect 20730 12182 20776 12194
rect 20848 12370 20894 12382
rect 20848 12194 20854 12370
rect 20888 12194 20894 12370
rect 20848 12182 20894 12194
rect 20966 12370 21012 12382
rect 20966 12194 20972 12370
rect 21006 12315 21012 12370
rect 21131 12370 21177 12382
rect 21131 12315 21137 12370
rect 21006 12227 21137 12315
rect 21006 12194 21012 12227
rect 20966 12182 21012 12194
rect 21131 12194 21137 12227
rect 21171 12194 21177 12370
rect 21131 12182 21177 12194
rect 21249 12370 21295 12382
rect 21249 12194 21255 12370
rect 21289 12194 21295 12370
rect 21249 12182 21295 12194
rect 21367 12370 21413 12382
rect 21367 12194 21373 12370
rect 21407 12194 21413 12370
rect 21367 12182 21413 12194
rect 21485 12370 21531 12382
rect 21485 12194 21491 12370
rect 21525 12194 21531 12370
rect 23215 12315 23397 13852
rect 26813 13611 26892 13623
rect 24329 13559 24408 13571
rect 24329 13463 24335 13559
rect 24263 13443 24335 13463
rect 24402 13463 24408 13559
rect 26813 13497 26819 13611
rect 26886 13497 26892 13611
rect 27962 13617 28041 13629
rect 27962 13497 27968 13617
rect 28035 13497 28041 13617
rect 24402 13443 24483 13463
rect 24263 13335 24307 13443
rect 24439 13335 24483 13443
rect 26060 13401 26116 13409
rect 24263 13293 24483 13335
rect 25134 13393 26116 13401
rect 25134 13359 26076 13393
rect 26110 13359 26116 13393
rect 26779 13389 26789 13497
rect 26921 13434 26931 13497
rect 26921 13423 26933 13434
rect 26921 13389 26934 13423
rect 27190 13413 27246 13415
rect 25134 13343 26116 13359
rect 26789 13351 26934 13389
rect 25134 13342 26113 13343
rect 23867 13263 24844 13293
rect 23867 13157 23899 13263
rect 24103 13157 24135 13263
rect 24339 13157 24371 13263
rect 24575 13157 24607 13263
rect 24810 13157 24844 13263
rect 23860 13145 23906 13157
rect 23860 12969 23866 13145
rect 23900 12969 23906 13145
rect 23860 12957 23906 12969
rect 23978 13145 24024 13157
rect 23978 12969 23984 13145
rect 24018 12969 24024 13145
rect 23978 12957 24024 12969
rect 24096 13145 24142 13157
rect 24096 12969 24102 13145
rect 24136 12969 24142 13145
rect 24096 12957 24142 12969
rect 24214 13145 24260 13157
rect 24214 12969 24220 13145
rect 24254 12969 24260 13145
rect 24214 12957 24260 12969
rect 24332 13145 24378 13157
rect 24332 12969 24338 13145
rect 24372 12969 24378 13145
rect 24332 12957 24378 12969
rect 24450 13145 24496 13157
rect 24450 12969 24456 13145
rect 24490 12969 24496 13145
rect 24450 12957 24496 12969
rect 24568 13145 24614 13157
rect 24568 12969 24574 13145
rect 24608 12969 24614 13145
rect 24568 12957 24614 12969
rect 24686 13145 24732 13157
rect 24686 12969 24692 13145
rect 24726 12969 24732 13145
rect 24686 12957 24732 12969
rect 24804 13145 24850 13157
rect 24804 12969 24810 13145
rect 24844 12969 24850 13145
rect 24804 12957 24850 12969
rect 24922 13145 24968 13157
rect 24922 12969 24928 13145
rect 24962 12969 24968 13145
rect 24922 12957 24968 12969
rect 23983 12863 24019 12957
rect 24219 12863 24255 12957
rect 24455 12864 24491 12957
rect 24617 12909 24683 12916
rect 24617 12875 24633 12909
rect 24667 12875 24683 12909
rect 24617 12864 24683 12875
rect 24455 12863 24683 12864
rect 23983 12834 24683 12863
rect 23983 12833 24565 12834
rect 24103 12720 24137 12833
rect 24499 12792 24565 12833
rect 24499 12758 24515 12792
rect 24549 12758 24565 12792
rect 24499 12751 24565 12758
rect 24927 12752 24962 12957
rect 25134 12752 25201 13342
rect 26893 13319 26934 13351
rect 27180 13347 27190 13413
rect 27246 13347 27256 13413
rect 27926 13389 27936 13497
rect 28068 13434 28078 13497
rect 28068 13423 28080 13434
rect 28068 13389 28081 13423
rect 27936 13351 28081 13389
rect 28040 13323 28081 13351
rect 26309 13291 26579 13319
rect 26050 13225 26060 13291
rect 26126 13225 26136 13291
rect 26309 13229 26343 13291
rect 26545 13229 26579 13291
rect 26663 13291 26934 13319
rect 27451 13295 27721 13323
rect 26663 13229 26697 13291
rect 26899 13229 26934 13291
rect 27075 13279 27246 13295
rect 27075 13245 27206 13279
rect 27240 13245 27246 13279
rect 27075 13229 27246 13245
rect 27451 13233 27485 13295
rect 27687 13233 27721 13295
rect 27805 13295 28081 13323
rect 27805 13233 27839 13295
rect 28041 13233 28081 13295
rect 26185 13217 26231 13229
rect 26185 12841 26191 13217
rect 26225 12841 26231 13217
rect 26185 12829 26231 12841
rect 26303 13217 26349 13229
rect 26303 12841 26309 13217
rect 26343 12841 26349 13217
rect 26303 12829 26349 12841
rect 26421 13217 26467 13229
rect 26421 12841 26427 13217
rect 26461 12841 26467 13217
rect 26421 12829 26467 12841
rect 26539 13217 26585 13229
rect 26539 12841 26545 13217
rect 26579 12841 26585 13217
rect 26539 12829 26585 12841
rect 26657 13217 26703 13229
rect 26657 12841 26663 13217
rect 26697 12841 26703 13217
rect 26657 12829 26703 12841
rect 26775 13217 26821 13229
rect 26775 12841 26781 13217
rect 26815 12841 26821 13217
rect 26775 12829 26821 12841
rect 26893 13217 26939 13229
rect 26893 12841 26899 13217
rect 26933 12841 26939 13217
rect 26893 12829 26939 12841
rect 24927 12724 25201 12752
rect 24573 12720 25201 12724
rect 24097 12708 24143 12720
rect 24097 12332 24103 12708
rect 24137 12332 24143 12708
rect 24097 12320 24143 12332
rect 24215 12708 24261 12720
rect 24215 12332 24221 12708
rect 24255 12332 24261 12708
rect 24215 12320 24261 12332
rect 24333 12708 24379 12720
rect 24333 12332 24339 12708
rect 24373 12356 24379 12708
rect 24450 12708 24496 12720
rect 24450 12532 24456 12708
rect 24490 12532 24496 12708
rect 24450 12520 24496 12532
rect 24568 12708 25201 12720
rect 24568 12532 24574 12708
rect 24608 12695 25201 12708
rect 26191 12787 26225 12829
rect 26427 12787 26461 12829
rect 26191 12759 26461 12787
rect 26545 12788 26579 12829
rect 26781 12788 26815 12829
rect 26545 12759 26815 12788
rect 26191 12711 26225 12759
rect 24608 12532 24614 12695
rect 26191 12681 26254 12711
rect 24568 12520 24614 12532
rect 26219 12589 26254 12681
rect 26219 12553 26446 12589
rect 26716 12578 26726 12675
rect 26825 12578 26835 12675
rect 26899 12646 26933 12829
rect 26899 12592 27008 12646
rect 24456 12404 24491 12520
rect 26219 12446 26254 12553
rect 26380 12519 26446 12553
rect 26380 12485 26396 12519
rect 26430 12485 26446 12519
rect 26727 12577 26824 12578
rect 26727 12510 26784 12577
rect 26380 12479 26446 12485
rect 26621 12474 26890 12510
rect 26621 12446 26654 12474
rect 26857 12446 26890 12474
rect 26974 12446 27008 12592
rect 26095 12434 26141 12446
rect 24587 12404 24695 12414
rect 24456 12356 24587 12404
rect 24695 12375 24843 12381
rect 24373 12332 24587 12356
rect 24333 12320 24587 12332
rect 24339 12316 24587 12320
rect 23215 12288 23975 12315
rect 23215 12282 24212 12288
rect 23215 12248 24162 12282
rect 24196 12248 24212 12282
rect 23215 12232 24212 12248
rect 24264 12282 24330 12288
rect 24264 12248 24280 12282
rect 24314 12248 24330 12282
rect 24513 12272 24587 12316
rect 24831 12308 24843 12375
rect 24695 12302 24843 12308
rect 24587 12262 24695 12272
rect 23215 12216 23975 12232
rect 23215 12215 23912 12216
rect 23215 12211 23447 12215
rect 21485 12182 21531 12194
rect 20618 12143 20652 12182
rect 20854 12143 20888 12182
rect 20618 12107 20888 12143
rect 21255 12144 21288 12182
rect 21491 12144 21524 12182
rect 21255 12108 21524 12144
rect 20618 12106 20784 12107
rect 20652 12027 20784 12106
rect 20642 11919 20652 12027
rect 20784 11919 20794 12027
rect 20678 11790 20684 11919
rect 20751 11790 20757 11919
rect 20678 11778 20757 11790
rect 22627 11800 23231 11828
rect 22627 11694 23079 11800
rect 23191 11787 23231 11800
rect 23191 11694 23233 11787
rect 22627 11683 23233 11694
rect 17256 11545 18233 11575
rect 20450 11573 20513 11590
rect 20375 11569 20513 11573
rect 17256 11439 17288 11545
rect 17492 11439 17524 11545
rect 17728 11439 17760 11545
rect 17964 11439 17996 11545
rect 18199 11439 18233 11545
rect 18543 11535 20513 11569
rect 18541 11506 20513 11535
rect 18541 11490 18587 11506
rect 20375 11504 20513 11506
rect 17249 11427 17295 11439
rect 17249 11251 17255 11427
rect 17289 11251 17295 11427
rect 17249 11239 17295 11251
rect 17367 11427 17413 11439
rect 17367 11251 17373 11427
rect 17407 11251 17413 11427
rect 17367 11239 17413 11251
rect 17485 11427 17531 11439
rect 17485 11251 17491 11427
rect 17525 11251 17531 11427
rect 17485 11239 17531 11251
rect 17603 11427 17649 11439
rect 17603 11251 17609 11427
rect 17643 11251 17649 11427
rect 17603 11239 17649 11251
rect 17721 11427 17767 11439
rect 17721 11251 17727 11427
rect 17761 11251 17767 11427
rect 17721 11239 17767 11251
rect 17839 11427 17885 11439
rect 17839 11251 17845 11427
rect 17879 11251 17885 11427
rect 17839 11239 17885 11251
rect 17957 11427 18003 11439
rect 17957 11251 17963 11427
rect 17997 11251 18003 11427
rect 17957 11239 18003 11251
rect 18075 11427 18121 11439
rect 18075 11251 18081 11427
rect 18115 11251 18121 11427
rect 18075 11239 18121 11251
rect 18193 11427 18239 11439
rect 18193 11251 18199 11427
rect 18233 11251 18239 11427
rect 18193 11239 18239 11251
rect 18311 11427 18357 11439
rect 18311 11251 18317 11427
rect 18351 11251 18357 11427
rect 18311 11239 18357 11251
rect 17372 11145 17408 11239
rect 17608 11145 17644 11239
rect 17844 11146 17880 11239
rect 18006 11191 18072 11198
rect 18006 11157 18022 11191
rect 18056 11157 18072 11191
rect 18006 11146 18072 11157
rect 17844 11145 18072 11146
rect 17372 11116 18072 11145
rect 17372 11115 17954 11116
rect 17492 11002 17526 11115
rect 17888 11074 17954 11115
rect 17888 11040 17904 11074
rect 17938 11040 17954 11074
rect 17888 11033 17954 11040
rect 18316 11021 18351 11239
rect 18540 11038 18587 11490
rect 21431 11494 21510 11506
rect 21431 11382 21437 11494
rect 21504 11382 21510 11494
rect 19499 11274 19509 11382
rect 19641 11274 19651 11382
rect 21397 11274 21407 11382
rect 21539 11274 21549 11382
rect 19509 11234 19641 11274
rect 21407 11234 21539 11274
rect 19508 11168 19641 11234
rect 21406 11168 21539 11234
rect 22627 11183 22777 11683
rect 22838 11682 23231 11683
rect 18837 11125 20310 11168
rect 18540 11022 18586 11038
rect 18505 11021 18586 11022
rect 18316 11006 18586 11021
rect 17962 11002 18586 11006
rect 17486 10990 17532 11002
rect 17221 10512 17231 10630
rect 17349 10598 17359 10630
rect 17486 10614 17492 10990
rect 17526 10614 17532 10990
rect 17486 10602 17532 10614
rect 17604 10990 17650 11002
rect 17604 10614 17610 10990
rect 17644 10614 17650 10990
rect 17604 10602 17650 10614
rect 17722 10990 17768 11002
rect 17722 10614 17728 10990
rect 17762 10638 17768 10990
rect 17839 10990 17885 11002
rect 17839 10814 17845 10990
rect 17879 10814 17885 10990
rect 17839 10802 17885 10814
rect 17957 10990 18586 11002
rect 17957 10814 17963 10990
rect 17997 10978 18586 10990
rect 17997 10977 18239 10978
rect 17997 10814 18003 10977
rect 18505 10976 18586 10978
rect 18837 10822 18871 11125
rect 19203 11022 19237 11125
rect 19439 11022 19473 11125
rect 19675 11022 19709 11125
rect 19911 11022 19945 11125
rect 19197 11010 19243 11022
rect 17957 10802 18003 10814
rect 18713 10810 18759 10822
rect 17845 10686 17880 10802
rect 17976 10686 18084 10696
rect 17845 10638 17976 10686
rect 18084 10648 18228 10654
rect 17762 10614 17976 10638
rect 17722 10602 17976 10614
rect 17728 10598 17976 10602
rect 17349 10570 17364 10598
rect 17349 10564 17601 10570
rect 17349 10530 17551 10564
rect 17585 10530 17601 10564
rect 17349 10514 17601 10530
rect 17653 10564 17719 10570
rect 17653 10530 17669 10564
rect 17703 10530 17719 10564
rect 17902 10554 17976 10598
rect 18216 10581 18228 10648
rect 18713 10634 18719 10810
rect 18753 10634 18759 10810
rect 18713 10622 18759 10634
rect 18831 10810 18877 10822
rect 18831 10634 18837 10810
rect 18871 10634 18877 10810
rect 18831 10622 18877 10634
rect 18949 10810 18995 10822
rect 18949 10634 18955 10810
rect 18989 10634 18995 10810
rect 18949 10622 18995 10634
rect 19067 10810 19113 10822
rect 19197 10810 19203 11010
rect 19067 10634 19073 10810
rect 19107 10634 19203 10810
rect 19237 10634 19243 11010
rect 19067 10622 19113 10634
rect 19197 10622 19243 10634
rect 19315 11010 19361 11022
rect 19315 10634 19321 11010
rect 19355 10634 19361 11010
rect 19315 10622 19361 10634
rect 19433 11010 19479 11022
rect 19433 10634 19439 11010
rect 19473 10634 19479 11010
rect 19433 10622 19479 10634
rect 19551 11010 19597 11022
rect 19551 10634 19557 11010
rect 19591 10634 19597 11010
rect 19551 10622 19597 10634
rect 19669 11010 19715 11022
rect 19669 10634 19675 11010
rect 19709 10634 19715 11010
rect 19669 10622 19715 10634
rect 19787 11010 19833 11022
rect 19787 10634 19793 11010
rect 19827 10634 19833 11010
rect 19787 10622 19833 10634
rect 19905 11010 19951 11022
rect 19905 10634 19911 11010
rect 19945 10810 19951 11010
rect 20276 10822 20310 11125
rect 20735 11125 22208 11168
rect 20735 10822 20769 11125
rect 21101 11022 21135 11125
rect 21337 11022 21371 11125
rect 21573 11022 21607 11125
rect 21809 11022 21843 11125
rect 21095 11010 21141 11022
rect 20034 10810 20080 10822
rect 19945 10634 20040 10810
rect 20074 10634 20080 10810
rect 19905 10622 19951 10634
rect 20034 10622 20080 10634
rect 20152 10810 20198 10822
rect 20152 10634 20158 10810
rect 20192 10634 20198 10810
rect 20152 10622 20198 10634
rect 20270 10810 20316 10822
rect 20270 10634 20276 10810
rect 20310 10634 20316 10810
rect 20270 10622 20316 10634
rect 20388 10810 20434 10822
rect 20388 10634 20394 10810
rect 20428 10634 20434 10810
rect 20388 10622 20434 10634
rect 20611 10810 20657 10822
rect 20611 10634 20617 10810
rect 20651 10634 20657 10810
rect 20611 10622 20657 10634
rect 20729 10810 20775 10822
rect 20729 10634 20735 10810
rect 20769 10634 20775 10810
rect 20729 10622 20775 10634
rect 20847 10810 20893 10822
rect 20847 10634 20853 10810
rect 20887 10634 20893 10810
rect 20847 10622 20893 10634
rect 20965 10810 21011 10822
rect 21095 10810 21101 11010
rect 20965 10634 20971 10810
rect 21005 10634 21101 10810
rect 21135 10634 21141 11010
rect 20965 10622 21011 10634
rect 21095 10622 21141 10634
rect 21213 11010 21259 11022
rect 21213 10634 21219 11010
rect 21253 10634 21259 11010
rect 21213 10622 21259 10634
rect 21331 11010 21377 11022
rect 21331 10634 21337 11010
rect 21371 10634 21377 11010
rect 21331 10622 21377 10634
rect 21449 11010 21495 11022
rect 21449 10634 21455 11010
rect 21489 10634 21495 11010
rect 21449 10622 21495 10634
rect 21567 11010 21613 11022
rect 21567 10634 21573 11010
rect 21607 10634 21613 11010
rect 21567 10622 21613 10634
rect 21685 11010 21731 11022
rect 21685 10634 21691 11010
rect 21725 10634 21731 11010
rect 21685 10622 21731 10634
rect 21803 11010 21849 11022
rect 21803 10634 21809 11010
rect 21843 10810 21849 11010
rect 22174 10822 22208 11125
rect 22626 11117 22777 11183
rect 21932 10810 21978 10822
rect 21843 10634 21938 10810
rect 21972 10634 21978 10810
rect 21803 10622 21849 10634
rect 21932 10622 21978 10634
rect 22050 10810 22096 10822
rect 22050 10634 22056 10810
rect 22090 10634 22096 10810
rect 22050 10622 22096 10634
rect 22168 10810 22214 10822
rect 22168 10634 22174 10810
rect 22208 10634 22214 10810
rect 22168 10622 22214 10634
rect 22286 10810 22332 10822
rect 22286 10634 22292 10810
rect 22326 10634 22332 10810
rect 22286 10622 22332 10634
rect 18084 10575 18228 10581
rect 18719 10588 18753 10622
rect 19321 10588 19355 10622
rect 19557 10588 19591 10622
rect 17976 10544 18084 10554
rect 18719 10553 18878 10588
rect 19321 10553 19591 10588
rect 20158 10588 20192 10622
rect 20394 10588 20428 10622
rect 20158 10553 20428 10588
rect 20617 10588 20651 10622
rect 21219 10588 21253 10622
rect 21455 10588 21489 10622
rect 20617 10553 20776 10588
rect 21219 10553 21489 10588
rect 22056 10588 22090 10622
rect 22292 10588 22326 10622
rect 22056 10553 22326 10588
rect 17349 10512 17364 10514
rect 17264 10498 17364 10512
rect 17264 10455 17364 10456
rect 16885 10434 17364 10455
rect 17653 10434 17719 10530
rect 16885 10386 17719 10434
rect 16885 10357 17364 10386
rect 16885 10355 16990 10357
rect 17264 10356 17364 10357
rect 16718 10170 16728 10249
rect 16821 10170 16831 10249
rect 17719 10239 17798 10251
rect 16729 8996 16822 10170
rect 17719 10141 17725 10239
rect 17647 10121 17725 10141
rect 17792 10141 17798 10239
rect 17792 10121 17867 10141
rect 17647 10013 17691 10121
rect 17823 10013 17867 10121
rect 17647 9971 17867 10013
rect 17251 9941 18228 9971
rect 17251 9835 17283 9941
rect 17487 9835 17519 9941
rect 17723 9835 17755 9941
rect 17959 9835 17991 9941
rect 18194 9835 18228 9941
rect 17244 9823 17290 9835
rect 17244 9647 17250 9823
rect 17284 9647 17290 9823
rect 17244 9635 17290 9647
rect 17362 9823 17408 9835
rect 17362 9647 17368 9823
rect 17402 9647 17408 9823
rect 17362 9635 17408 9647
rect 17480 9823 17526 9835
rect 17480 9647 17486 9823
rect 17520 9647 17526 9823
rect 17480 9635 17526 9647
rect 17598 9823 17644 9835
rect 17598 9647 17604 9823
rect 17638 9647 17644 9823
rect 17598 9635 17644 9647
rect 17716 9823 17762 9835
rect 17716 9647 17722 9823
rect 17756 9647 17762 9823
rect 17716 9635 17762 9647
rect 17834 9823 17880 9835
rect 17834 9647 17840 9823
rect 17874 9647 17880 9823
rect 17834 9635 17880 9647
rect 17952 9823 17998 9835
rect 17952 9647 17958 9823
rect 17992 9647 17998 9823
rect 17952 9635 17998 9647
rect 18070 9823 18116 9835
rect 18070 9647 18076 9823
rect 18110 9647 18116 9823
rect 18070 9635 18116 9647
rect 18188 9823 18234 9835
rect 18188 9647 18194 9823
rect 18228 9647 18234 9823
rect 18188 9635 18234 9647
rect 18306 9823 18352 9835
rect 18306 9647 18312 9823
rect 18346 9647 18352 9823
rect 18306 9635 18352 9647
rect 18844 9769 18878 10553
rect 19557 10491 19591 10553
rect 19146 10453 19888 10491
rect 19146 10329 19180 10453
rect 19382 10329 19416 10453
rect 19618 10329 19652 10453
rect 19854 10329 19888 10453
rect 20144 10346 20154 10412
rect 20217 10346 20227 10412
rect 19140 10317 19186 10329
rect 19140 9941 19146 10317
rect 19180 9941 19186 10317
rect 19140 9929 19186 9941
rect 19258 10317 19304 10329
rect 19258 9941 19264 10317
rect 19298 9941 19304 10317
rect 19258 9929 19304 9941
rect 19376 10317 19422 10329
rect 19376 9941 19382 10317
rect 19416 9941 19422 10317
rect 19376 9929 19422 9941
rect 19494 10317 19540 10329
rect 19494 9941 19500 10317
rect 19534 9941 19540 10317
rect 19494 9929 19540 9941
rect 19612 10317 19658 10329
rect 19612 9941 19618 10317
rect 19652 9941 19658 10317
rect 19612 9929 19658 9941
rect 19730 10317 19776 10329
rect 19730 9941 19736 10317
rect 19770 9941 19776 10317
rect 19730 9929 19776 9941
rect 19848 10317 19894 10329
rect 19848 9941 19854 10317
rect 19888 9941 19894 10317
rect 19848 9929 19894 9941
rect 20260 9770 20294 10553
rect 19987 9769 20294 9770
rect 18844 9764 19160 9769
rect 19874 9764 20294 9769
rect 18844 9753 19227 9764
rect 18844 9726 19176 9753
rect 17367 9541 17403 9635
rect 17603 9541 17639 9635
rect 17839 9542 17875 9635
rect 18001 9587 18067 9594
rect 18001 9553 18017 9587
rect 18051 9553 18067 9587
rect 18001 9542 18067 9553
rect 17839 9541 18067 9542
rect 17367 9512 18067 9541
rect 17367 9511 17949 9512
rect 17487 9398 17521 9511
rect 17883 9470 17949 9511
rect 17883 9436 17899 9470
rect 17933 9436 17949 9470
rect 17883 9429 17949 9436
rect 18311 9402 18346 9635
rect 18844 9597 18878 9726
rect 19160 9719 19176 9726
rect 19210 9719 19227 9753
rect 19160 9713 19227 9719
rect 19807 9753 20294 9764
rect 19807 9719 19824 9753
rect 19858 9726 20294 9753
rect 19858 9719 19874 9726
rect 19987 9725 20294 9726
rect 19807 9713 19874 9719
rect 18985 9686 19041 9698
rect 18985 9652 18991 9686
rect 19025 9685 19041 9686
rect 20098 9685 20154 9697
rect 19025 9669 19492 9685
rect 19025 9652 19442 9669
rect 18985 9636 19442 9652
rect 19426 9635 19442 9636
rect 19476 9635 19492 9669
rect 19426 9628 19492 9635
rect 19544 9670 20114 9685
rect 19544 9636 19560 9670
rect 19594 9651 20114 9670
rect 20148 9651 20154 9685
rect 19594 9636 20154 9651
rect 19544 9626 19611 9636
rect 20098 9635 20154 9636
rect 20260 9597 20294 9725
rect 20742 9769 20776 10553
rect 21455 10491 21489 10553
rect 21044 10453 21786 10491
rect 21044 10329 21078 10453
rect 21280 10329 21314 10453
rect 21516 10329 21550 10453
rect 21752 10329 21786 10453
rect 21038 10317 21084 10329
rect 21038 9941 21044 10317
rect 21078 9941 21084 10317
rect 21038 9929 21084 9941
rect 21156 10317 21202 10329
rect 21156 9941 21162 10317
rect 21196 9941 21202 10317
rect 21156 9929 21202 9941
rect 21274 10317 21320 10329
rect 21274 9941 21280 10317
rect 21314 9941 21320 10317
rect 21274 9929 21320 9941
rect 21392 10317 21438 10329
rect 21392 9941 21398 10317
rect 21432 9941 21438 10317
rect 21392 9929 21438 9941
rect 21510 10317 21556 10329
rect 21510 9941 21516 10317
rect 21550 9941 21556 10317
rect 21510 9929 21556 9941
rect 21628 10317 21674 10329
rect 21628 9941 21634 10317
rect 21668 9941 21674 10317
rect 21628 9929 21674 9941
rect 21746 10317 21792 10329
rect 21746 9941 21752 10317
rect 21786 9941 21792 10317
rect 21746 9929 21792 9941
rect 22158 9770 22192 10553
rect 21770 9769 21839 9770
rect 21885 9769 22192 9770
rect 20742 9764 21058 9769
rect 21770 9765 22192 9769
rect 20742 9753 21125 9764
rect 20742 9726 21074 9753
rect 20742 9597 20776 9726
rect 21058 9719 21074 9726
rect 21108 9719 21125 9753
rect 21058 9713 21125 9719
rect 21703 9754 22192 9765
rect 21703 9720 21720 9754
rect 21754 9726 22192 9754
rect 21754 9720 21770 9726
rect 21885 9725 22192 9726
rect 21703 9714 21770 9720
rect 20883 9686 20939 9698
rect 20883 9652 20889 9686
rect 20923 9685 20939 9686
rect 21996 9685 22052 9697
rect 20923 9669 21390 9685
rect 20923 9652 21340 9669
rect 20883 9636 21340 9652
rect 21324 9635 21340 9636
rect 21374 9635 21390 9669
rect 21324 9628 21390 9635
rect 21442 9670 22012 9685
rect 21442 9636 21458 9670
rect 21492 9651 22012 9670
rect 22046 9651 22052 9685
rect 21492 9636 22052 9651
rect 21442 9626 21509 9636
rect 21996 9635 22052 9636
rect 22158 9597 22192 9725
rect 22273 10375 22340 10399
rect 22273 10341 22290 10375
rect 22324 10341 22340 10375
rect 17957 9398 18346 9402
rect 17481 9386 17527 9398
rect 17481 9010 17487 9386
rect 17521 9010 17527 9386
rect 17481 8998 17527 9010
rect 17599 9386 17645 9398
rect 17599 9010 17605 9386
rect 17639 9010 17645 9386
rect 17599 8998 17645 9010
rect 17717 9386 17763 9398
rect 17717 9010 17723 9386
rect 17757 9034 17763 9386
rect 17834 9386 17880 9398
rect 17834 9210 17840 9386
rect 17874 9210 17880 9386
rect 17834 9198 17880 9210
rect 17952 9386 18346 9398
rect 18838 9585 18884 9597
rect 18838 9409 18844 9585
rect 18878 9409 18884 9585
rect 18838 9397 18884 9409
rect 18956 9585 19002 9597
rect 18956 9409 18962 9585
rect 18996 9409 19002 9585
rect 18956 9397 19002 9409
rect 19258 9585 19304 9597
rect 17952 9210 17958 9386
rect 17992 9373 18346 9386
rect 17992 9210 17998 9373
rect 18268 9370 18346 9373
rect 18268 9318 18278 9370
rect 18341 9318 18351 9370
rect 18273 9312 18346 9318
rect 17952 9198 17998 9210
rect 17840 9082 17875 9198
rect 18961 9103 18995 9397
rect 19258 9209 19264 9585
rect 19298 9209 19304 9585
rect 19258 9197 19304 9209
rect 19376 9585 19422 9597
rect 19376 9209 19382 9585
rect 19416 9209 19422 9585
rect 19376 9197 19422 9209
rect 19494 9585 19540 9597
rect 19494 9209 19500 9585
rect 19534 9209 19540 9585
rect 19494 9197 19540 9209
rect 19612 9585 19658 9597
rect 19612 9209 19618 9585
rect 19652 9209 19658 9585
rect 19612 9197 19658 9209
rect 19730 9585 19776 9597
rect 19730 9209 19736 9585
rect 19770 9209 19776 9585
rect 20136 9585 20182 9597
rect 20136 9409 20142 9585
rect 20176 9409 20182 9585
rect 20136 9397 20182 9409
rect 20254 9585 20300 9597
rect 20254 9409 20260 9585
rect 20294 9409 20300 9585
rect 20254 9397 20300 9409
rect 20736 9585 20782 9597
rect 20736 9409 20742 9585
rect 20776 9409 20782 9585
rect 20736 9397 20782 9409
rect 20854 9585 20900 9597
rect 20854 9409 20860 9585
rect 20894 9409 20900 9585
rect 20854 9397 20900 9409
rect 21156 9585 21202 9597
rect 19730 9197 19776 9209
rect 19618 9103 19652 9197
rect 20142 9103 20175 9397
rect 17971 9082 18079 9092
rect 17840 9034 17971 9082
rect 18961 9071 20175 9103
rect 20859 9103 20893 9397
rect 21156 9209 21162 9585
rect 21196 9209 21202 9585
rect 21156 9197 21202 9209
rect 21274 9585 21320 9597
rect 21274 9209 21280 9585
rect 21314 9209 21320 9585
rect 21274 9197 21320 9209
rect 21392 9585 21438 9597
rect 21392 9209 21398 9585
rect 21432 9209 21438 9585
rect 21392 9197 21438 9209
rect 21510 9585 21556 9597
rect 21510 9209 21516 9585
rect 21550 9209 21556 9585
rect 21510 9197 21556 9209
rect 21628 9585 21674 9597
rect 21628 9209 21634 9585
rect 21668 9209 21674 9585
rect 22034 9585 22080 9597
rect 22034 9409 22040 9585
rect 22074 9409 22080 9585
rect 22034 9397 22080 9409
rect 22152 9585 22198 9597
rect 22152 9409 22158 9585
rect 22192 9409 22198 9585
rect 22152 9397 22198 9409
rect 21628 9197 21674 9209
rect 21516 9103 21550 9197
rect 22040 9103 22073 9397
rect 20859 9071 22073 9103
rect 18079 9043 18230 9049
rect 17757 9010 17971 9034
rect 17717 8998 17971 9010
rect 16729 8994 17314 8996
rect 17723 8994 17971 8998
rect 16729 8966 17359 8994
rect 16729 8960 17596 8966
rect 16729 8926 17546 8960
rect 17580 8926 17596 8960
rect 16729 8910 17596 8926
rect 17648 8960 17714 8966
rect 17648 8926 17664 8960
rect 17698 8926 17714 8960
rect 17897 8950 17971 8994
rect 18218 8976 18230 9043
rect 19454 8986 19586 9071
rect 21352 8986 21484 9071
rect 18079 8970 18230 8976
rect 17971 8940 18079 8950
rect 16729 8894 17359 8910
rect 16729 8890 17314 8894
rect 16729 8889 16830 8890
rect 17259 8841 17359 8852
rect 17223 8735 17233 8841
rect 17345 8830 17359 8841
rect 17648 8830 17714 8926
rect 19444 8878 19454 8986
rect 19586 8878 19596 8986
rect 21342 8878 21352 8986
rect 21484 8878 21494 8986
rect 22273 8958 22340 10341
rect 17345 8782 17714 8830
rect 17345 8752 17359 8782
rect 17345 8735 17355 8752
rect 17647 8679 17713 8782
rect 19472 8742 19478 8878
rect 19545 8742 19551 8878
rect 19472 8730 19551 8742
rect 22273 8679 22339 8958
rect 17645 8599 22339 8679
rect 16387 8565 16550 8579
rect 16387 8497 16431 8565
rect 16501 8497 16550 8565
rect 16387 7778 16550 8497
rect 22395 8485 22405 8599
rect 22528 8485 22538 8599
rect 16387 7748 16551 7778
rect 16387 7680 16430 7748
rect 16500 7680 16551 7748
rect 20186 7747 20265 7759
rect 16387 7666 16551 7680
rect 17701 7687 17780 7699
rect 17701 7594 17707 7687
rect 17633 7574 17707 7594
rect 17774 7594 17780 7687
rect 20186 7628 20192 7747
rect 20259 7628 20265 7747
rect 21335 7744 21414 7756
rect 21335 7628 21341 7744
rect 21408 7628 21414 7744
rect 17774 7574 17853 7594
rect 17633 7466 17677 7574
rect 17809 7466 17853 7574
rect 19430 7532 19486 7540
rect 17633 7424 17853 7466
rect 18504 7524 19486 7532
rect 18504 7490 19446 7524
rect 19480 7490 19486 7524
rect 20149 7520 20159 7628
rect 20291 7565 20301 7628
rect 20291 7554 20303 7565
rect 20291 7520 20304 7554
rect 20560 7544 20616 7546
rect 18504 7474 19486 7490
rect 20159 7482 20304 7520
rect 18504 7473 19483 7474
rect 17237 7394 18214 7424
rect 17237 7288 17269 7394
rect 17473 7288 17505 7394
rect 17709 7288 17741 7394
rect 17945 7288 17977 7394
rect 18180 7288 18214 7394
rect 17230 7276 17276 7288
rect 17230 7100 17236 7276
rect 17270 7100 17276 7276
rect 17230 7088 17276 7100
rect 17348 7276 17394 7288
rect 17348 7100 17354 7276
rect 17388 7100 17394 7276
rect 17348 7088 17394 7100
rect 17466 7276 17512 7288
rect 17466 7100 17472 7276
rect 17506 7100 17512 7276
rect 17466 7088 17512 7100
rect 17584 7276 17630 7288
rect 17584 7100 17590 7276
rect 17624 7100 17630 7276
rect 17584 7088 17630 7100
rect 17702 7276 17748 7288
rect 17702 7100 17708 7276
rect 17742 7100 17748 7276
rect 17702 7088 17748 7100
rect 17820 7276 17866 7288
rect 17820 7100 17826 7276
rect 17860 7100 17866 7276
rect 17820 7088 17866 7100
rect 17938 7276 17984 7288
rect 17938 7100 17944 7276
rect 17978 7100 17984 7276
rect 17938 7088 17984 7100
rect 18056 7276 18102 7288
rect 18056 7100 18062 7276
rect 18096 7100 18102 7276
rect 18056 7088 18102 7100
rect 18174 7276 18220 7288
rect 18174 7100 18180 7276
rect 18214 7100 18220 7276
rect 18174 7088 18220 7100
rect 18292 7276 18338 7288
rect 18292 7100 18298 7276
rect 18332 7100 18338 7276
rect 18292 7088 18338 7100
rect 17353 6994 17389 7088
rect 17589 6994 17625 7088
rect 17825 6995 17861 7088
rect 17987 7040 18053 7047
rect 17987 7006 18003 7040
rect 18037 7006 18053 7040
rect 17987 6995 18053 7006
rect 17825 6994 18053 6995
rect 17353 6965 18053 6994
rect 17353 6964 17935 6965
rect 17473 6851 17507 6964
rect 17869 6923 17935 6964
rect 17869 6889 17885 6923
rect 17919 6889 17935 6923
rect 17869 6882 17935 6889
rect 18297 6883 18332 7088
rect 18504 6883 18571 7473
rect 20263 7450 20304 7482
rect 20550 7478 20560 7544
rect 20616 7478 20626 7544
rect 21296 7520 21306 7628
rect 21438 7565 21448 7628
rect 21438 7554 21450 7565
rect 21438 7520 21451 7554
rect 21306 7482 21451 7520
rect 21410 7454 21451 7482
rect 19679 7422 19949 7450
rect 19420 7356 19430 7422
rect 19496 7356 19506 7422
rect 19679 7360 19713 7422
rect 19915 7360 19949 7422
rect 20033 7422 20304 7450
rect 20821 7426 21091 7454
rect 20033 7360 20067 7422
rect 20269 7360 20304 7422
rect 20445 7410 20616 7426
rect 20445 7376 20576 7410
rect 20610 7376 20616 7410
rect 20445 7360 20616 7376
rect 20821 7364 20855 7426
rect 21057 7364 21091 7426
rect 21175 7426 21451 7454
rect 21175 7364 21209 7426
rect 21411 7364 21451 7426
rect 19555 7348 19601 7360
rect 19555 6972 19561 7348
rect 19595 6972 19601 7348
rect 19555 6960 19601 6972
rect 19673 7348 19719 7360
rect 19673 6972 19679 7348
rect 19713 6972 19719 7348
rect 19673 6960 19719 6972
rect 19791 7348 19837 7360
rect 19791 6972 19797 7348
rect 19831 6972 19837 7348
rect 19791 6960 19837 6972
rect 19909 7348 19955 7360
rect 19909 6972 19915 7348
rect 19949 6972 19955 7348
rect 19909 6960 19955 6972
rect 20027 7348 20073 7360
rect 20027 6972 20033 7348
rect 20067 6972 20073 7348
rect 20027 6960 20073 6972
rect 20145 7348 20191 7360
rect 20145 6972 20151 7348
rect 20185 6972 20191 7348
rect 20145 6960 20191 6972
rect 20263 7348 20309 7360
rect 20263 6972 20269 7348
rect 20303 6972 20309 7348
rect 20263 6960 20309 6972
rect 18297 6855 18571 6883
rect 17943 6851 18571 6855
rect 17467 6839 17513 6851
rect 17467 6463 17473 6839
rect 17507 6463 17513 6839
rect 17467 6451 17513 6463
rect 17585 6839 17631 6851
rect 17585 6463 17591 6839
rect 17625 6463 17631 6839
rect 17585 6451 17631 6463
rect 17703 6839 17749 6851
rect 17703 6463 17709 6839
rect 17743 6487 17749 6839
rect 17820 6839 17866 6851
rect 17820 6663 17826 6839
rect 17860 6663 17866 6839
rect 17820 6651 17866 6663
rect 17938 6839 18571 6851
rect 17938 6663 17944 6839
rect 17978 6826 18571 6839
rect 19561 6918 19595 6960
rect 19797 6918 19831 6960
rect 19561 6890 19831 6918
rect 19915 6919 19949 6960
rect 20151 6919 20185 6960
rect 19915 6890 20185 6919
rect 19561 6842 19595 6890
rect 17978 6663 17984 6826
rect 19561 6812 19624 6842
rect 17938 6651 17984 6663
rect 19589 6720 19624 6812
rect 19589 6684 19816 6720
rect 20086 6709 20096 6806
rect 20195 6709 20205 6806
rect 20269 6777 20303 6960
rect 20269 6723 20378 6777
rect 17826 6535 17861 6651
rect 19589 6577 19624 6684
rect 19750 6650 19816 6684
rect 19750 6616 19766 6650
rect 19800 6616 19816 6650
rect 20097 6708 20194 6709
rect 20097 6641 20154 6708
rect 19750 6610 19816 6616
rect 19991 6605 20260 6641
rect 19991 6577 20024 6605
rect 20227 6577 20260 6605
rect 20344 6577 20378 6723
rect 19465 6565 19511 6577
rect 17957 6535 18065 6545
rect 17826 6487 17957 6535
rect 18065 6499 18216 6505
rect 17743 6463 17957 6487
rect 17703 6451 17957 6463
rect 17709 6447 17957 6451
rect 16020 6446 16643 6447
rect 16020 6419 17345 6446
rect 16020 6413 17582 6419
rect 13958 6341 13992 6380
rect 14194 6341 14228 6380
rect 13958 6305 14228 6341
rect 14595 6342 14628 6380
rect 14831 6342 14864 6380
rect 14595 6306 14864 6342
rect 16020 6379 17532 6413
rect 17566 6379 17582 6413
rect 16020 6363 17582 6379
rect 17634 6413 17700 6419
rect 17634 6379 17650 6413
rect 17684 6379 17700 6413
rect 17883 6403 17957 6447
rect 18204 6432 18216 6499
rect 18065 6426 18216 6432
rect 17957 6393 18065 6403
rect 16020 6347 17345 6363
rect 16020 6346 17282 6347
rect 16020 6342 16817 6346
rect 16020 6341 16643 6342
rect 13958 6304 14124 6305
rect 13992 6225 14124 6304
rect 13982 6117 13992 6225
rect 14124 6117 14134 6225
rect 14014 5972 14020 6117
rect 14087 5972 14093 6117
rect 14014 5960 14093 5972
rect 16021 5954 16602 5962
rect 16020 5936 16602 5954
rect 16020 5823 16382 5936
rect 16586 5918 16602 5936
rect 16020 5822 16534 5823
rect 16586 5822 16603 5918
rect 16020 5812 16603 5822
rect 10596 5743 11573 5773
rect 13790 5771 13853 5788
rect 13715 5767 13853 5771
rect 10596 5637 10628 5743
rect 10832 5637 10864 5743
rect 11068 5637 11100 5743
rect 11304 5637 11336 5743
rect 11539 5637 11573 5743
rect 11883 5733 13853 5767
rect 11881 5704 13853 5733
rect 11881 5688 11927 5704
rect 13715 5702 13853 5704
rect 10589 5625 10635 5637
rect 10589 5449 10595 5625
rect 10629 5449 10635 5625
rect 10589 5437 10635 5449
rect 10707 5625 10753 5637
rect 10707 5449 10713 5625
rect 10747 5449 10753 5625
rect 10707 5437 10753 5449
rect 10825 5625 10871 5637
rect 10825 5449 10831 5625
rect 10865 5449 10871 5625
rect 10825 5437 10871 5449
rect 10943 5625 10989 5637
rect 10943 5449 10949 5625
rect 10983 5449 10989 5625
rect 10943 5437 10989 5449
rect 11061 5625 11107 5637
rect 11061 5449 11067 5625
rect 11101 5449 11107 5625
rect 11061 5437 11107 5449
rect 11179 5625 11225 5637
rect 11179 5449 11185 5625
rect 11219 5449 11225 5625
rect 11179 5437 11225 5449
rect 11297 5625 11343 5637
rect 11297 5449 11303 5625
rect 11337 5449 11343 5625
rect 11297 5437 11343 5449
rect 11415 5625 11461 5637
rect 11415 5449 11421 5625
rect 11455 5449 11461 5625
rect 11415 5437 11461 5449
rect 11533 5625 11579 5637
rect 11533 5449 11539 5625
rect 11573 5449 11579 5625
rect 11533 5437 11579 5449
rect 11651 5625 11697 5637
rect 11651 5449 11657 5625
rect 11691 5449 11697 5625
rect 11651 5437 11697 5449
rect 10712 5343 10748 5437
rect 10948 5343 10984 5437
rect 11184 5344 11220 5437
rect 11346 5389 11412 5396
rect 11346 5355 11362 5389
rect 11396 5355 11412 5389
rect 11346 5344 11412 5355
rect 11184 5343 11412 5344
rect 10712 5314 11412 5343
rect 10712 5313 11294 5314
rect 10832 5200 10866 5313
rect 11228 5272 11294 5313
rect 11228 5238 11244 5272
rect 11278 5238 11294 5272
rect 11228 5231 11294 5238
rect 11656 5219 11691 5437
rect 11880 5236 11927 5688
rect 14778 5697 14857 5709
rect 14778 5580 14784 5697
rect 14851 5580 14857 5697
rect 12839 5472 12849 5580
rect 12981 5472 12991 5580
rect 14737 5472 14747 5580
rect 14879 5472 14889 5580
rect 12849 5432 12981 5472
rect 14747 5432 14879 5472
rect 12848 5366 12981 5432
rect 14746 5366 14879 5432
rect 12177 5323 13650 5366
rect 11880 5220 11926 5236
rect 11845 5219 11926 5220
rect 11656 5204 11926 5219
rect 11302 5200 11926 5204
rect 10826 5188 10872 5200
rect 10561 4710 10571 4828
rect 10689 4796 10699 4828
rect 10826 4812 10832 5188
rect 10866 4812 10872 5188
rect 10826 4800 10872 4812
rect 10944 5188 10990 5200
rect 10944 4812 10950 5188
rect 10984 4812 10990 5188
rect 10944 4800 10990 4812
rect 11062 5188 11108 5200
rect 11062 4812 11068 5188
rect 11102 4836 11108 5188
rect 11179 5188 11225 5200
rect 11179 5012 11185 5188
rect 11219 5012 11225 5188
rect 11179 5000 11225 5012
rect 11297 5188 11926 5200
rect 11297 5012 11303 5188
rect 11337 5176 11926 5188
rect 11337 5175 11579 5176
rect 11337 5012 11343 5175
rect 11845 5174 11926 5176
rect 12177 5020 12211 5323
rect 12543 5220 12577 5323
rect 12779 5220 12813 5323
rect 13015 5220 13049 5323
rect 13251 5220 13285 5323
rect 12537 5208 12583 5220
rect 11297 5000 11343 5012
rect 12053 5008 12099 5020
rect 11185 4884 11220 5000
rect 11316 4884 11424 4894
rect 11185 4836 11316 4884
rect 11424 4845 11571 4851
rect 11102 4812 11316 4836
rect 11062 4800 11316 4812
rect 11068 4796 11316 4800
rect 10689 4768 10704 4796
rect 10689 4762 10941 4768
rect 10689 4728 10891 4762
rect 10925 4728 10941 4762
rect 10689 4712 10941 4728
rect 10993 4762 11059 4768
rect 10993 4728 11009 4762
rect 11043 4728 11059 4762
rect 11242 4752 11316 4796
rect 11559 4778 11571 4845
rect 12053 4832 12059 5008
rect 12093 4832 12099 5008
rect 12053 4820 12099 4832
rect 12171 5008 12217 5020
rect 12171 4832 12177 5008
rect 12211 4832 12217 5008
rect 12171 4820 12217 4832
rect 12289 5008 12335 5020
rect 12289 4832 12295 5008
rect 12329 4832 12335 5008
rect 12289 4820 12335 4832
rect 12407 5008 12453 5020
rect 12537 5008 12543 5208
rect 12407 4832 12413 5008
rect 12447 4832 12543 5008
rect 12577 4832 12583 5208
rect 12407 4820 12453 4832
rect 12537 4820 12583 4832
rect 12655 5208 12701 5220
rect 12655 4832 12661 5208
rect 12695 4832 12701 5208
rect 12655 4820 12701 4832
rect 12773 5208 12819 5220
rect 12773 4832 12779 5208
rect 12813 4832 12819 5208
rect 12773 4820 12819 4832
rect 12891 5208 12937 5220
rect 12891 4832 12897 5208
rect 12931 4832 12937 5208
rect 12891 4820 12937 4832
rect 13009 5208 13055 5220
rect 13009 4832 13015 5208
rect 13049 4832 13055 5208
rect 13009 4820 13055 4832
rect 13127 5208 13173 5220
rect 13127 4832 13133 5208
rect 13167 4832 13173 5208
rect 13127 4820 13173 4832
rect 13245 5208 13291 5220
rect 13245 4832 13251 5208
rect 13285 5008 13291 5208
rect 13616 5020 13650 5323
rect 14075 5323 15548 5366
rect 14075 5020 14109 5323
rect 14441 5220 14475 5323
rect 14677 5220 14711 5323
rect 14913 5220 14947 5323
rect 15149 5220 15183 5323
rect 14435 5208 14481 5220
rect 13374 5008 13420 5020
rect 13285 4832 13380 5008
rect 13414 4832 13420 5008
rect 13245 4820 13291 4832
rect 13374 4820 13420 4832
rect 13492 5008 13538 5020
rect 13492 4832 13498 5008
rect 13532 4832 13538 5008
rect 13492 4820 13538 4832
rect 13610 5008 13656 5020
rect 13610 4832 13616 5008
rect 13650 4832 13656 5008
rect 13610 4820 13656 4832
rect 13728 5008 13774 5020
rect 13728 4832 13734 5008
rect 13768 4832 13774 5008
rect 13728 4820 13774 4832
rect 13951 5008 13997 5020
rect 13951 4832 13957 5008
rect 13991 4832 13997 5008
rect 13951 4820 13997 4832
rect 14069 5008 14115 5020
rect 14069 4832 14075 5008
rect 14109 4832 14115 5008
rect 14069 4820 14115 4832
rect 14187 5008 14233 5020
rect 14187 4832 14193 5008
rect 14227 4832 14233 5008
rect 14187 4820 14233 4832
rect 14305 5008 14351 5020
rect 14435 5008 14441 5208
rect 14305 4832 14311 5008
rect 14345 4832 14441 5008
rect 14475 4832 14481 5208
rect 14305 4820 14351 4832
rect 14435 4820 14481 4832
rect 14553 5208 14599 5220
rect 14553 4832 14559 5208
rect 14593 4832 14599 5208
rect 14553 4820 14599 4832
rect 14671 5208 14717 5220
rect 14671 4832 14677 5208
rect 14711 4832 14717 5208
rect 14671 4820 14717 4832
rect 14789 5208 14835 5220
rect 14789 4832 14795 5208
rect 14829 4832 14835 5208
rect 14789 4820 14835 4832
rect 14907 5208 14953 5220
rect 14907 4832 14913 5208
rect 14947 4832 14953 5208
rect 14907 4820 14953 4832
rect 15025 5208 15071 5220
rect 15025 4832 15031 5208
rect 15065 4832 15071 5208
rect 15025 4820 15071 4832
rect 15143 5208 15189 5220
rect 15143 4832 15149 5208
rect 15183 5008 15189 5208
rect 15514 5020 15548 5323
rect 15272 5008 15318 5020
rect 15183 4832 15278 5008
rect 15312 4832 15318 5008
rect 15143 4820 15189 4832
rect 15272 4820 15318 4832
rect 15390 5008 15436 5020
rect 15390 4832 15396 5008
rect 15430 4832 15436 5008
rect 15390 4820 15436 4832
rect 15508 5008 15554 5020
rect 15508 4832 15514 5008
rect 15548 4832 15554 5008
rect 15508 4820 15554 4832
rect 15626 5008 15672 5020
rect 15626 4832 15632 5008
rect 15666 4832 15672 5008
rect 15626 4820 15672 4832
rect 11424 4772 11571 4778
rect 12059 4786 12093 4820
rect 12661 4786 12695 4820
rect 12897 4786 12931 4820
rect 11316 4742 11424 4752
rect 12059 4751 12218 4786
rect 12661 4751 12931 4786
rect 13498 4786 13532 4820
rect 13734 4786 13768 4820
rect 13498 4751 13768 4786
rect 13957 4786 13991 4820
rect 14559 4786 14593 4820
rect 14795 4786 14829 4820
rect 13957 4751 14116 4786
rect 14559 4751 14829 4786
rect 15396 4786 15430 4820
rect 15632 4786 15666 4820
rect 15396 4751 15666 4786
rect 10689 4710 10704 4712
rect 10604 4696 10704 4710
rect 10604 4653 10704 4654
rect 10225 4632 10704 4653
rect 10993 4632 11059 4728
rect 10225 4584 11059 4632
rect 10225 4555 10704 4584
rect 10225 4553 10330 4555
rect 10604 4554 10704 4555
rect 10058 4368 10068 4447
rect 10161 4368 10171 4447
rect 11061 4435 11140 4447
rect 10069 3194 10162 4368
rect 11061 4339 11067 4435
rect 10987 4319 11067 4339
rect 11134 4339 11140 4435
rect 11134 4319 11207 4339
rect 10987 4211 11031 4319
rect 11163 4211 11207 4319
rect 10987 4169 11207 4211
rect 10591 4139 11568 4169
rect 10591 4033 10623 4139
rect 10827 4033 10859 4139
rect 11063 4033 11095 4139
rect 11299 4033 11331 4139
rect 11534 4033 11568 4139
rect 10584 4021 10630 4033
rect 10584 3845 10590 4021
rect 10624 3845 10630 4021
rect 10584 3833 10630 3845
rect 10702 4021 10748 4033
rect 10702 3845 10708 4021
rect 10742 3845 10748 4021
rect 10702 3833 10748 3845
rect 10820 4021 10866 4033
rect 10820 3845 10826 4021
rect 10860 3845 10866 4021
rect 10820 3833 10866 3845
rect 10938 4021 10984 4033
rect 10938 3845 10944 4021
rect 10978 3845 10984 4021
rect 10938 3833 10984 3845
rect 11056 4021 11102 4033
rect 11056 3845 11062 4021
rect 11096 3845 11102 4021
rect 11056 3833 11102 3845
rect 11174 4021 11220 4033
rect 11174 3845 11180 4021
rect 11214 3845 11220 4021
rect 11174 3833 11220 3845
rect 11292 4021 11338 4033
rect 11292 3845 11298 4021
rect 11332 3845 11338 4021
rect 11292 3833 11338 3845
rect 11410 4021 11456 4033
rect 11410 3845 11416 4021
rect 11450 3845 11456 4021
rect 11410 3833 11456 3845
rect 11528 4021 11574 4033
rect 11528 3845 11534 4021
rect 11568 3845 11574 4021
rect 11528 3833 11574 3845
rect 11646 4021 11692 4033
rect 11646 3845 11652 4021
rect 11686 3845 11692 4021
rect 11646 3833 11692 3845
rect 12184 3967 12218 4751
rect 12897 4689 12931 4751
rect 12486 4651 13228 4689
rect 12486 4527 12520 4651
rect 12722 4527 12756 4651
rect 12958 4527 12992 4651
rect 13194 4527 13228 4651
rect 13484 4544 13494 4610
rect 13557 4544 13567 4610
rect 12480 4515 12526 4527
rect 12480 4139 12486 4515
rect 12520 4139 12526 4515
rect 12480 4127 12526 4139
rect 12598 4515 12644 4527
rect 12598 4139 12604 4515
rect 12638 4139 12644 4515
rect 12598 4127 12644 4139
rect 12716 4515 12762 4527
rect 12716 4139 12722 4515
rect 12756 4139 12762 4515
rect 12716 4127 12762 4139
rect 12834 4515 12880 4527
rect 12834 4139 12840 4515
rect 12874 4139 12880 4515
rect 12834 4127 12880 4139
rect 12952 4515 12998 4527
rect 12952 4139 12958 4515
rect 12992 4139 12998 4515
rect 12952 4127 12998 4139
rect 13070 4515 13116 4527
rect 13070 4139 13076 4515
rect 13110 4139 13116 4515
rect 13070 4127 13116 4139
rect 13188 4515 13234 4527
rect 13188 4139 13194 4515
rect 13228 4139 13234 4515
rect 13188 4127 13234 4139
rect 13600 3968 13634 4751
rect 13327 3967 13634 3968
rect 12184 3962 12500 3967
rect 13214 3962 13634 3967
rect 12184 3951 12567 3962
rect 12184 3924 12516 3951
rect 10707 3739 10743 3833
rect 10943 3739 10979 3833
rect 11179 3740 11215 3833
rect 11341 3785 11407 3792
rect 11341 3751 11357 3785
rect 11391 3751 11407 3785
rect 11341 3740 11407 3751
rect 11179 3739 11407 3740
rect 10707 3710 11407 3739
rect 10707 3709 11289 3710
rect 10827 3596 10861 3709
rect 11223 3668 11289 3709
rect 11223 3634 11239 3668
rect 11273 3634 11289 3668
rect 11223 3627 11289 3634
rect 11651 3600 11686 3833
rect 12184 3795 12218 3924
rect 12500 3917 12516 3924
rect 12550 3917 12567 3951
rect 12500 3911 12567 3917
rect 13147 3951 13634 3962
rect 13147 3917 13164 3951
rect 13198 3924 13634 3951
rect 13198 3917 13214 3924
rect 13327 3923 13634 3924
rect 13147 3911 13214 3917
rect 12325 3884 12381 3896
rect 12325 3850 12331 3884
rect 12365 3883 12381 3884
rect 13438 3883 13494 3895
rect 12365 3867 12832 3883
rect 12365 3850 12782 3867
rect 12325 3834 12782 3850
rect 12766 3833 12782 3834
rect 12816 3833 12832 3867
rect 12766 3826 12832 3833
rect 12884 3868 13454 3883
rect 12884 3834 12900 3868
rect 12934 3849 13454 3868
rect 13488 3849 13494 3883
rect 12934 3834 13494 3849
rect 12884 3824 12951 3834
rect 13438 3833 13494 3834
rect 13600 3795 13634 3923
rect 14082 3967 14116 4751
rect 14795 4689 14829 4751
rect 14384 4651 15126 4689
rect 14384 4527 14418 4651
rect 14620 4527 14654 4651
rect 14856 4527 14890 4651
rect 15092 4527 15126 4651
rect 14378 4515 14424 4527
rect 14378 4139 14384 4515
rect 14418 4139 14424 4515
rect 14378 4127 14424 4139
rect 14496 4515 14542 4527
rect 14496 4139 14502 4515
rect 14536 4139 14542 4515
rect 14496 4127 14542 4139
rect 14614 4515 14660 4527
rect 14614 4139 14620 4515
rect 14654 4139 14660 4515
rect 14614 4127 14660 4139
rect 14732 4515 14778 4527
rect 14732 4139 14738 4515
rect 14772 4139 14778 4515
rect 14732 4127 14778 4139
rect 14850 4515 14896 4527
rect 14850 4139 14856 4515
rect 14890 4139 14896 4515
rect 14850 4127 14896 4139
rect 14968 4515 15014 4527
rect 14968 4139 14974 4515
rect 15008 4139 15014 4515
rect 14968 4127 15014 4139
rect 15086 4515 15132 4527
rect 15086 4139 15092 4515
rect 15126 4139 15132 4515
rect 15086 4127 15132 4139
rect 15498 3968 15532 4751
rect 15110 3967 15179 3968
rect 15225 3967 15532 3968
rect 14082 3962 14398 3967
rect 15110 3963 15532 3967
rect 14082 3951 14465 3962
rect 14082 3924 14414 3951
rect 14082 3795 14116 3924
rect 14398 3917 14414 3924
rect 14448 3917 14465 3951
rect 14398 3911 14465 3917
rect 15043 3952 15532 3963
rect 15043 3918 15060 3952
rect 15094 3924 15532 3952
rect 15094 3918 15110 3924
rect 15225 3923 15532 3924
rect 15043 3912 15110 3918
rect 14223 3884 14279 3896
rect 14223 3850 14229 3884
rect 14263 3883 14279 3884
rect 15336 3883 15392 3895
rect 14263 3867 14730 3883
rect 14263 3850 14680 3867
rect 14223 3834 14680 3850
rect 14664 3833 14680 3834
rect 14714 3833 14730 3867
rect 14664 3826 14730 3833
rect 14782 3868 15352 3883
rect 14782 3834 14798 3868
rect 14832 3849 15352 3868
rect 15386 3849 15392 3883
rect 14832 3834 15392 3849
rect 14782 3824 14849 3834
rect 15336 3833 15392 3834
rect 15498 3795 15532 3923
rect 15613 4573 15680 4597
rect 15613 4539 15630 4573
rect 15664 4539 15680 4573
rect 11297 3596 11686 3600
rect 10821 3584 10867 3596
rect 10821 3208 10827 3584
rect 10861 3208 10867 3584
rect 10821 3196 10867 3208
rect 10939 3584 10985 3596
rect 10939 3208 10945 3584
rect 10979 3208 10985 3584
rect 10939 3196 10985 3208
rect 11057 3584 11103 3596
rect 11057 3208 11063 3584
rect 11097 3232 11103 3584
rect 11174 3584 11220 3596
rect 11174 3408 11180 3584
rect 11214 3408 11220 3584
rect 11174 3396 11220 3408
rect 11292 3584 11686 3596
rect 12178 3783 12224 3795
rect 12178 3607 12184 3783
rect 12218 3607 12224 3783
rect 12178 3595 12224 3607
rect 12296 3783 12342 3795
rect 12296 3607 12302 3783
rect 12336 3607 12342 3783
rect 12296 3595 12342 3607
rect 12598 3783 12644 3795
rect 11292 3408 11298 3584
rect 11332 3571 11686 3584
rect 11332 3408 11338 3571
rect 11608 3568 11686 3571
rect 11608 3516 11618 3568
rect 11681 3516 11691 3568
rect 11613 3510 11686 3516
rect 11292 3396 11338 3408
rect 11180 3280 11215 3396
rect 12301 3301 12335 3595
rect 12598 3407 12604 3783
rect 12638 3407 12644 3783
rect 12598 3395 12644 3407
rect 12716 3783 12762 3795
rect 12716 3407 12722 3783
rect 12756 3407 12762 3783
rect 12716 3395 12762 3407
rect 12834 3783 12880 3795
rect 12834 3407 12840 3783
rect 12874 3407 12880 3783
rect 12834 3395 12880 3407
rect 12952 3783 12998 3795
rect 12952 3407 12958 3783
rect 12992 3407 12998 3783
rect 12952 3395 12998 3407
rect 13070 3783 13116 3795
rect 13070 3407 13076 3783
rect 13110 3407 13116 3783
rect 13476 3783 13522 3795
rect 13476 3607 13482 3783
rect 13516 3607 13522 3783
rect 13476 3595 13522 3607
rect 13594 3783 13640 3795
rect 13594 3607 13600 3783
rect 13634 3607 13640 3783
rect 13594 3595 13640 3607
rect 14076 3783 14122 3795
rect 14076 3607 14082 3783
rect 14116 3607 14122 3783
rect 14076 3595 14122 3607
rect 14194 3783 14240 3795
rect 14194 3607 14200 3783
rect 14234 3607 14240 3783
rect 14194 3595 14240 3607
rect 14496 3783 14542 3795
rect 13070 3395 13116 3407
rect 12958 3301 12992 3395
rect 13482 3301 13515 3595
rect 11311 3280 11419 3290
rect 11180 3232 11311 3280
rect 12301 3269 13515 3301
rect 14199 3301 14233 3595
rect 14496 3407 14502 3783
rect 14536 3407 14542 3783
rect 14496 3395 14542 3407
rect 14614 3783 14660 3795
rect 14614 3407 14620 3783
rect 14654 3407 14660 3783
rect 14614 3395 14660 3407
rect 14732 3783 14778 3795
rect 14732 3407 14738 3783
rect 14772 3407 14778 3783
rect 14732 3395 14778 3407
rect 14850 3783 14896 3795
rect 14850 3407 14856 3783
rect 14890 3407 14896 3783
rect 14850 3395 14896 3407
rect 14968 3783 15014 3795
rect 14968 3407 14974 3783
rect 15008 3407 15014 3783
rect 15374 3783 15420 3795
rect 15374 3607 15380 3783
rect 15414 3607 15420 3783
rect 15374 3595 15420 3607
rect 15492 3783 15538 3795
rect 15492 3607 15498 3783
rect 15532 3607 15538 3783
rect 15492 3595 15538 3607
rect 14968 3395 15014 3407
rect 14856 3301 14890 3395
rect 15380 3301 15413 3595
rect 14199 3269 15413 3301
rect 11419 3245 11560 3251
rect 11097 3208 11311 3232
rect 11057 3196 11311 3208
rect 10069 3192 10654 3194
rect 11063 3192 11311 3196
rect 10069 3164 10699 3192
rect 10069 3158 10936 3164
rect 10069 3124 10886 3158
rect 10920 3124 10936 3158
rect 10069 3108 10936 3124
rect 10988 3158 11054 3164
rect 10988 3124 11004 3158
rect 11038 3124 11054 3158
rect 11237 3148 11311 3192
rect 11548 3178 11560 3245
rect 12794 3184 12926 3269
rect 14692 3184 14824 3269
rect 11419 3172 11560 3178
rect 11311 3138 11419 3148
rect 10069 3092 10699 3108
rect 10069 3088 10654 3092
rect 10069 3087 10170 3088
rect 10599 3039 10699 3050
rect 10563 2933 10573 3039
rect 10685 3028 10699 3039
rect 10988 3028 11054 3124
rect 12784 3076 12794 3184
rect 12926 3076 12936 3184
rect 14682 3076 14692 3184
rect 14824 3076 14834 3184
rect 15613 3156 15680 4539
rect 10685 2980 11054 3028
rect 10685 2950 10699 2980
rect 10685 2933 10695 2950
rect 10987 2877 11053 2980
rect 12815 2936 12821 3076
rect 12888 2936 12894 3076
rect 12815 2924 12894 2936
rect 15613 2877 15679 3156
rect 10985 2797 15679 2877
rect 14402 2299 14866 2331
rect 14954 2315 14964 2375
rect 15026 2315 15036 2375
rect 14402 2291 14865 2299
rect 14402 2142 14456 2291
rect 8839 1794 9568 1874
rect 8589 1781 9568 1794
rect 8549 1769 9568 1781
rect 8084 1656 8118 1769
rect 8554 1765 9568 1769
rect 14082 2042 14456 2142
rect 14516 2246 14747 2262
rect 14516 2212 14697 2246
rect 14731 2212 14747 2246
rect 14516 2206 14747 2212
rect 14799 2246 14865 2291
rect 14799 2212 14815 2246
rect 14849 2212 14865 2246
rect 14799 2206 14865 2212
rect 8480 1731 8546 1738
rect 8480 1697 8496 1731
rect 8530 1697 8546 1731
rect 8480 1656 8546 1697
rect 7964 1655 8546 1656
rect 7964 1626 8664 1655
rect 7964 1532 8000 1626
rect 8200 1532 8236 1626
rect 8436 1625 8664 1626
rect 8436 1532 8472 1625
rect 8598 1614 8664 1625
rect 8598 1580 8614 1614
rect 8648 1580 8664 1614
rect 8598 1573 8664 1580
rect 8908 1532 8943 1765
rect 7841 1520 7887 1532
rect 7841 1344 7847 1520
rect 7881 1344 7887 1520
rect 7841 1332 7887 1344
rect 7959 1520 8005 1532
rect 7959 1344 7965 1520
rect 7999 1344 8005 1520
rect 7959 1332 8005 1344
rect 8077 1520 8123 1532
rect 8077 1344 8083 1520
rect 8117 1344 8123 1520
rect 8077 1332 8123 1344
rect 8195 1520 8241 1532
rect 8195 1344 8201 1520
rect 8235 1344 8241 1520
rect 8195 1332 8241 1344
rect 8313 1520 8359 1532
rect 8313 1344 8319 1520
rect 8353 1344 8359 1520
rect 8313 1332 8359 1344
rect 8431 1520 8477 1532
rect 8431 1344 8437 1520
rect 8471 1344 8477 1520
rect 8431 1332 8477 1344
rect 8549 1520 8595 1532
rect 8549 1344 8555 1520
rect 8589 1344 8595 1520
rect 8549 1332 8595 1344
rect 8667 1520 8713 1532
rect 8667 1344 8673 1520
rect 8707 1344 8713 1520
rect 8667 1332 8713 1344
rect 8785 1520 8831 1532
rect 8785 1344 8791 1520
rect 8825 1344 8831 1520
rect 8785 1332 8831 1344
rect 8903 1520 8949 1532
rect 8903 1344 8909 1520
rect 8943 1344 8949 1520
rect 8903 1332 8949 1344
rect 7848 1226 7880 1332
rect 8084 1226 8116 1332
rect 8320 1226 8352 1332
rect 8556 1226 8588 1332
rect 8791 1226 8825 1332
rect 7848 1196 8825 1226
rect 8152 1168 8288 1196
rect 8152 1106 8188 1168
rect 8248 1106 8288 1168
rect 8152 1086 8288 1106
rect 772 1027 1545 1028
rect 14082 1027 14205 2042
rect 14516 2013 14570 2206
rect 14958 2178 15034 2315
rect 14874 2174 15034 2178
rect 772 928 14205 1027
rect 14243 1914 14570 2013
rect 14632 2162 14678 2174
rect 871 927 13806 928
rect -3115 877 -2715 883
rect -3277 843 -3103 877
rect -2727 843 -2715 877
rect -3808 820 -3408 826
rect -3954 786 -3796 820
rect -3420 786 -3408 820
rect -3954 584 -3911 786
rect -3808 780 -3408 786
rect -3808 702 -3408 708
rect -3808 668 -3796 702
rect -3420 668 -3408 702
rect -3808 662 -3408 668
rect -3277 641 -3239 843
rect -3115 837 -2715 843
rect -3115 759 -2715 765
rect -3115 725 -3103 759
rect -2727 725 -2715 759
rect -3115 719 -2715 725
rect -2550 671 -2499 688
rect -3115 641 -2715 647
rect -3277 607 -3103 641
rect -2727 607 -2715 641
rect -2550 637 -2539 671
rect -2505 637 -2499 671
rect -2550 621 -2499 637
rect -3115 601 -2715 607
rect -3808 584 -3408 590
rect -3954 550 -3796 584
rect -3420 550 -3408 584
rect -3954 219 -3911 550
rect -3808 544 -3408 550
rect -3596 461 -3420 544
rect -2555 508 -2512 621
rect -3608 455 -3408 461
rect -3608 421 -3596 455
rect -3420 421 -3408 455
rect -3608 415 -3408 421
rect -3257 369 -3191 381
rect -3608 337 -3408 343
rect -3608 303 -3596 337
rect -3420 303 -3339 337
rect -3257 315 -3251 369
rect -3197 315 -3191 369
rect -3257 303 -3191 315
rect -3608 297 -3408 303
rect -3374 235 -3339 303
rect -2556 235 -2511 508
rect -2471 397 -2422 884
rect -2383 877 -1983 883
rect -1889 877 -1857 909
rect 5 903 130 909
rect -2383 843 -2371 877
rect -1995 843 -1857 877
rect -2383 837 -1983 843
rect -2383 759 -1983 765
rect -2383 725 -2371 759
rect -1995 725 -1983 759
rect -2383 719 -1983 725
rect -2483 381 -2421 397
rect -2483 347 -2471 381
rect -2437 347 -2421 381
rect -2483 341 -2421 347
rect -2383 353 -2183 359
rect -1889 353 -1857 843
rect 3 898 130 903
rect 14243 898 14348 1914
rect 14632 1786 14638 2162
rect 14672 1786 14678 2162
rect 14632 1774 14678 1786
rect 14750 2162 14796 2174
rect 14750 1786 14756 2162
rect 14790 1786 14796 2162
rect 14750 1774 14796 1786
rect 14868 2162 15034 2174
rect 14868 1786 14874 2162
rect 14908 2135 15034 2162
rect 14908 1786 14914 2135
rect 14991 1974 15034 2135
rect 14868 1774 14914 1786
rect 14985 1969 15034 1974
rect 14985 1962 15031 1969
rect 14985 1786 14991 1962
rect 15025 1786 15031 1962
rect 14985 1774 15031 1786
rect 15103 1962 15149 1974
rect 15103 1786 15109 1962
rect 15143 1799 15149 1962
rect 16020 1879 16156 5812
rect 16724 4448 16817 6342
rect 16880 6283 17346 6305
rect 17634 6283 17700 6379
rect 19465 6389 19471 6565
rect 19505 6389 19511 6565
rect 19465 6377 19511 6389
rect 19583 6565 19629 6577
rect 19583 6389 19589 6565
rect 19623 6389 19629 6565
rect 19583 6377 19629 6389
rect 19701 6565 19747 6577
rect 19701 6389 19707 6565
rect 19741 6389 19747 6565
rect 19701 6377 19747 6389
rect 19819 6565 19865 6577
rect 19819 6389 19825 6565
rect 19859 6510 19865 6565
rect 19984 6565 20030 6577
rect 19984 6510 19990 6565
rect 19859 6422 19990 6510
rect 19859 6389 19865 6422
rect 19819 6377 19865 6389
rect 19984 6389 19990 6422
rect 20024 6389 20030 6565
rect 19984 6377 20030 6389
rect 20102 6565 20148 6577
rect 20102 6389 20108 6565
rect 20142 6389 20148 6565
rect 20102 6377 20148 6389
rect 20220 6565 20266 6577
rect 20220 6389 20226 6565
rect 20260 6389 20266 6565
rect 20220 6377 20266 6389
rect 20338 6565 20384 6577
rect 20338 6389 20344 6565
rect 20378 6389 20384 6565
rect 20338 6377 20384 6389
rect 19471 6338 19505 6377
rect 19707 6338 19741 6377
rect 19471 6303 19741 6338
rect 20108 6339 20141 6377
rect 20344 6339 20377 6377
rect 20108 6303 20377 6339
rect 16880 6235 17700 6283
rect 19505 6302 19741 6303
rect 16880 6204 17346 6235
rect 19505 6228 19637 6302
rect 16880 5948 16985 6204
rect 19495 6120 19505 6228
rect 19637 6120 19647 6228
rect 17721 6041 17800 6053
rect 16880 5842 16943 5948
rect 17055 5842 17065 5948
rect 17721 5944 17727 6041
rect 17647 5924 17727 5944
rect 17794 5944 17800 6041
rect 19525 5987 19531 6120
rect 19598 5987 19604 6120
rect 19525 5975 19604 5987
rect 17794 5924 17867 5944
rect 16880 5831 17029 5842
rect 16880 4654 16985 5831
rect 17647 5816 17691 5924
rect 17823 5816 17867 5924
rect 17647 5774 17867 5816
rect 20445 5789 20507 7360
rect 20697 7352 20743 7364
rect 20697 6976 20703 7352
rect 20737 6976 20743 7352
rect 20697 6964 20743 6976
rect 20815 7352 20861 7364
rect 20815 6976 20821 7352
rect 20855 6976 20861 7352
rect 20815 6964 20861 6976
rect 20933 7352 20979 7364
rect 20933 6976 20939 7352
rect 20973 6976 20979 7352
rect 20933 6964 20979 6976
rect 21051 7352 21097 7364
rect 21051 6976 21057 7352
rect 21091 6976 21097 7352
rect 21051 6964 21097 6976
rect 21169 7352 21215 7364
rect 21169 6976 21175 7352
rect 21209 6976 21215 7352
rect 21169 6964 21215 6976
rect 21287 7352 21333 7364
rect 21287 6976 21293 7352
rect 21327 6976 21333 7352
rect 21287 6964 21333 6976
rect 21405 7352 21451 7364
rect 21405 6976 21411 7352
rect 21445 6976 21451 7352
rect 21405 6964 21451 6976
rect 20703 6922 20737 6964
rect 20939 6922 20973 6964
rect 20703 6894 20973 6922
rect 21057 6923 21091 6964
rect 21293 6923 21327 6964
rect 21057 6894 21327 6923
rect 20703 6846 20737 6894
rect 20703 6816 20766 6846
rect 20731 6724 20766 6816
rect 21238 6786 21338 6807
rect 21238 6732 21252 6786
rect 21317 6732 21338 6786
rect 21238 6727 21338 6732
rect 21411 6781 21445 6964
rect 22626 6933 22778 11117
rect 23354 10317 23447 12211
rect 23510 12152 23976 12174
rect 24264 12152 24330 12248
rect 26095 12258 26101 12434
rect 26135 12258 26141 12434
rect 26095 12246 26141 12258
rect 26213 12434 26259 12446
rect 26213 12258 26219 12434
rect 26253 12258 26259 12434
rect 26213 12246 26259 12258
rect 26331 12434 26377 12446
rect 26331 12258 26337 12434
rect 26371 12258 26377 12434
rect 26331 12246 26377 12258
rect 26449 12434 26495 12446
rect 26449 12258 26455 12434
rect 26489 12379 26495 12434
rect 26614 12434 26660 12446
rect 26614 12379 26620 12434
rect 26489 12291 26620 12379
rect 26489 12258 26495 12291
rect 26449 12246 26495 12258
rect 26614 12258 26620 12291
rect 26654 12258 26660 12434
rect 26614 12246 26660 12258
rect 26732 12434 26778 12446
rect 26732 12258 26738 12434
rect 26772 12258 26778 12434
rect 26732 12246 26778 12258
rect 26850 12434 26896 12446
rect 26850 12258 26856 12434
rect 26890 12258 26896 12434
rect 26850 12246 26896 12258
rect 26968 12434 27014 12446
rect 26968 12258 26974 12434
rect 27008 12258 27014 12434
rect 26968 12246 27014 12258
rect 26101 12207 26135 12246
rect 26337 12207 26371 12246
rect 26101 12172 26371 12207
rect 26738 12208 26771 12246
rect 26974 12208 27007 12246
rect 26738 12172 27007 12208
rect 23510 12104 24330 12152
rect 26135 12171 26371 12172
rect 23510 12073 23976 12104
rect 26135 12097 26267 12171
rect 23510 11817 23615 12073
rect 26125 11989 26135 12097
rect 26267 11989 26277 12097
rect 24352 11908 24431 11920
rect 23510 11711 23573 11817
rect 23685 11711 23695 11817
rect 24352 11813 24358 11908
rect 24277 11793 24358 11813
rect 24425 11813 24431 11908
rect 26153 11846 26159 11989
rect 26226 11846 26232 11989
rect 26153 11834 26232 11846
rect 24425 11793 24497 11813
rect 23510 11700 23659 11711
rect 23510 10523 23615 11700
rect 24277 11685 24321 11793
rect 24453 11685 24497 11793
rect 24277 11643 24497 11685
rect 27075 11658 27137 13229
rect 27327 13221 27373 13233
rect 27327 12845 27333 13221
rect 27367 12845 27373 13221
rect 27327 12833 27373 12845
rect 27445 13221 27491 13233
rect 27445 12845 27451 13221
rect 27485 12845 27491 13221
rect 27445 12833 27491 12845
rect 27563 13221 27609 13233
rect 27563 12845 27569 13221
rect 27603 12845 27609 13221
rect 27563 12833 27609 12845
rect 27681 13221 27727 13233
rect 27681 12845 27687 13221
rect 27721 12845 27727 13221
rect 27681 12833 27727 12845
rect 27799 13221 27845 13233
rect 27799 12845 27805 13221
rect 27839 12845 27845 13221
rect 27799 12833 27845 12845
rect 27917 13221 27963 13233
rect 27917 12845 27923 13221
rect 27957 12845 27963 13221
rect 27917 12833 27963 12845
rect 28035 13221 28081 13233
rect 28035 12845 28041 13221
rect 28075 12845 28081 13221
rect 28035 12833 28081 12845
rect 27333 12791 27367 12833
rect 27569 12791 27603 12833
rect 27333 12763 27603 12791
rect 27687 12792 27721 12833
rect 27923 12792 27957 12833
rect 27687 12763 27957 12792
rect 27333 12715 27367 12763
rect 27333 12685 27396 12715
rect 27361 12593 27396 12685
rect 27868 12655 27968 12676
rect 27868 12601 27882 12655
rect 27947 12601 27968 12655
rect 27868 12596 27968 12601
rect 28041 12650 28075 12833
rect 28041 12596 28150 12650
rect 27361 12557 27588 12593
rect 27361 12450 27396 12557
rect 27522 12523 27588 12557
rect 27522 12489 27538 12523
rect 27572 12489 27588 12523
rect 27869 12581 27966 12596
rect 27869 12514 27926 12581
rect 27522 12483 27588 12489
rect 27763 12478 28032 12514
rect 27763 12450 27796 12478
rect 27999 12450 28032 12478
rect 28116 12450 28150 12596
rect 28850 12589 28860 12664
rect 28928 12589 29040 15532
rect 28877 12588 29040 12589
rect 28929 12578 29040 12588
rect 27237 12438 27283 12450
rect 27237 12262 27243 12438
rect 27277 12262 27283 12438
rect 27237 12250 27283 12262
rect 27355 12438 27401 12450
rect 27355 12262 27361 12438
rect 27395 12262 27401 12438
rect 27355 12250 27401 12262
rect 27473 12438 27519 12450
rect 27473 12262 27479 12438
rect 27513 12262 27519 12438
rect 27473 12250 27519 12262
rect 27591 12438 27637 12450
rect 27591 12262 27597 12438
rect 27631 12383 27637 12438
rect 27756 12438 27802 12450
rect 27756 12383 27762 12438
rect 27631 12295 27762 12383
rect 27631 12262 27637 12295
rect 27591 12250 27637 12262
rect 27756 12262 27762 12295
rect 27796 12262 27802 12438
rect 27756 12250 27802 12262
rect 27874 12438 27920 12450
rect 27874 12262 27880 12438
rect 27914 12262 27920 12438
rect 27874 12250 27920 12262
rect 27992 12438 28038 12450
rect 27992 12262 27998 12438
rect 28032 12262 28038 12438
rect 27992 12250 28038 12262
rect 28110 12438 28156 12450
rect 28110 12262 28116 12438
rect 28150 12262 28156 12438
rect 28110 12250 28156 12262
rect 27243 12211 27277 12250
rect 27479 12211 27513 12250
rect 27243 12175 27513 12211
rect 27880 12212 27913 12250
rect 28116 12212 28149 12250
rect 27880 12176 28149 12212
rect 27243 12174 27409 12175
rect 27277 12095 27409 12174
rect 27267 11987 27277 12095
rect 27409 11987 27419 12095
rect 27296 11848 27302 11987
rect 27369 11848 27375 11987
rect 27296 11836 27375 11848
rect 23881 11613 24858 11643
rect 27075 11641 27138 11658
rect 27000 11637 27138 11641
rect 23881 11507 23913 11613
rect 24117 11507 24149 11613
rect 24353 11507 24385 11613
rect 24589 11507 24621 11613
rect 24824 11507 24858 11613
rect 25168 11603 27138 11637
rect 25166 11574 27138 11603
rect 25166 11558 25212 11574
rect 27000 11572 27138 11574
rect 23874 11495 23920 11507
rect 23874 11319 23880 11495
rect 23914 11319 23920 11495
rect 23874 11307 23920 11319
rect 23992 11495 24038 11507
rect 23992 11319 23998 11495
rect 24032 11319 24038 11495
rect 23992 11307 24038 11319
rect 24110 11495 24156 11507
rect 24110 11319 24116 11495
rect 24150 11319 24156 11495
rect 24110 11307 24156 11319
rect 24228 11495 24274 11507
rect 24228 11319 24234 11495
rect 24268 11319 24274 11495
rect 24228 11307 24274 11319
rect 24346 11495 24392 11507
rect 24346 11319 24352 11495
rect 24386 11319 24392 11495
rect 24346 11307 24392 11319
rect 24464 11495 24510 11507
rect 24464 11319 24470 11495
rect 24504 11319 24510 11495
rect 24464 11307 24510 11319
rect 24582 11495 24628 11507
rect 24582 11319 24588 11495
rect 24622 11319 24628 11495
rect 24582 11307 24628 11319
rect 24700 11495 24746 11507
rect 24700 11319 24706 11495
rect 24740 11319 24746 11495
rect 24700 11307 24746 11319
rect 24818 11495 24864 11507
rect 24818 11319 24824 11495
rect 24858 11319 24864 11495
rect 24818 11307 24864 11319
rect 24936 11495 24982 11507
rect 24936 11319 24942 11495
rect 24976 11319 24982 11495
rect 24936 11307 24982 11319
rect 23997 11213 24033 11307
rect 24233 11213 24269 11307
rect 24469 11214 24505 11307
rect 24631 11259 24697 11266
rect 24631 11225 24647 11259
rect 24681 11225 24697 11259
rect 24631 11214 24697 11225
rect 24469 11213 24697 11214
rect 23997 11184 24697 11213
rect 23997 11183 24579 11184
rect 24117 11070 24151 11183
rect 24513 11142 24579 11183
rect 24513 11108 24529 11142
rect 24563 11108 24579 11142
rect 24513 11101 24579 11108
rect 24941 11089 24976 11307
rect 25165 11106 25212 11558
rect 28059 11563 28138 11575
rect 28059 11450 28065 11563
rect 28132 11450 28138 11563
rect 26124 11342 26134 11450
rect 26266 11342 26276 11450
rect 28022 11342 28032 11450
rect 28164 11342 28174 11450
rect 26134 11302 26266 11342
rect 28032 11302 28164 11342
rect 26133 11236 26266 11302
rect 28031 11236 28164 11302
rect 25462 11193 26935 11236
rect 25165 11090 25211 11106
rect 25130 11089 25211 11090
rect 24941 11074 25211 11089
rect 24587 11070 25211 11074
rect 24111 11058 24157 11070
rect 23846 10580 23856 10698
rect 23974 10666 23984 10698
rect 24111 10682 24117 11058
rect 24151 10682 24157 11058
rect 24111 10670 24157 10682
rect 24229 11058 24275 11070
rect 24229 10682 24235 11058
rect 24269 10682 24275 11058
rect 24229 10670 24275 10682
rect 24347 11058 24393 11070
rect 24347 10682 24353 11058
rect 24387 10706 24393 11058
rect 24464 11058 24510 11070
rect 24464 10882 24470 11058
rect 24504 10882 24510 11058
rect 24464 10870 24510 10882
rect 24582 11058 25211 11070
rect 24582 10882 24588 11058
rect 24622 11046 25211 11058
rect 24622 11045 24864 11046
rect 24622 10882 24628 11045
rect 25130 11044 25211 11046
rect 25462 10890 25496 11193
rect 25828 11090 25862 11193
rect 26064 11090 26098 11193
rect 26300 11090 26334 11193
rect 26536 11090 26570 11193
rect 25822 11078 25868 11090
rect 24582 10870 24628 10882
rect 25338 10878 25384 10890
rect 24470 10754 24505 10870
rect 24601 10754 24709 10764
rect 24470 10706 24601 10754
rect 24709 10714 24848 10720
rect 24387 10682 24601 10706
rect 24347 10670 24601 10682
rect 24353 10666 24601 10670
rect 23974 10638 23989 10666
rect 23974 10632 24226 10638
rect 23974 10598 24176 10632
rect 24210 10598 24226 10632
rect 23974 10582 24226 10598
rect 24278 10632 24344 10638
rect 24278 10598 24294 10632
rect 24328 10598 24344 10632
rect 24527 10622 24601 10666
rect 24836 10647 24848 10714
rect 25338 10702 25344 10878
rect 25378 10702 25384 10878
rect 25338 10690 25384 10702
rect 25456 10878 25502 10890
rect 25456 10702 25462 10878
rect 25496 10702 25502 10878
rect 25456 10690 25502 10702
rect 25574 10878 25620 10890
rect 25574 10702 25580 10878
rect 25614 10702 25620 10878
rect 25574 10690 25620 10702
rect 25692 10878 25738 10890
rect 25822 10878 25828 11078
rect 25692 10702 25698 10878
rect 25732 10702 25828 10878
rect 25862 10702 25868 11078
rect 25692 10690 25738 10702
rect 25822 10690 25868 10702
rect 25940 11078 25986 11090
rect 25940 10702 25946 11078
rect 25980 10702 25986 11078
rect 25940 10690 25986 10702
rect 26058 11078 26104 11090
rect 26058 10702 26064 11078
rect 26098 10702 26104 11078
rect 26058 10690 26104 10702
rect 26176 11078 26222 11090
rect 26176 10702 26182 11078
rect 26216 10702 26222 11078
rect 26176 10690 26222 10702
rect 26294 11078 26340 11090
rect 26294 10702 26300 11078
rect 26334 10702 26340 11078
rect 26294 10690 26340 10702
rect 26412 11078 26458 11090
rect 26412 10702 26418 11078
rect 26452 10702 26458 11078
rect 26412 10690 26458 10702
rect 26530 11078 26576 11090
rect 26530 10702 26536 11078
rect 26570 10878 26576 11078
rect 26901 10890 26935 11193
rect 27360 11193 28833 11236
rect 27360 10890 27394 11193
rect 27726 11090 27760 11193
rect 27962 11090 27996 11193
rect 28198 11090 28232 11193
rect 28434 11090 28468 11193
rect 27720 11078 27766 11090
rect 26659 10878 26705 10890
rect 26570 10702 26665 10878
rect 26699 10702 26705 10878
rect 26530 10690 26576 10702
rect 26659 10690 26705 10702
rect 26777 10878 26823 10890
rect 26777 10702 26783 10878
rect 26817 10702 26823 10878
rect 26777 10690 26823 10702
rect 26895 10878 26941 10890
rect 26895 10702 26901 10878
rect 26935 10702 26941 10878
rect 26895 10690 26941 10702
rect 27013 10878 27059 10890
rect 27013 10702 27019 10878
rect 27053 10702 27059 10878
rect 27013 10690 27059 10702
rect 27236 10878 27282 10890
rect 27236 10702 27242 10878
rect 27276 10702 27282 10878
rect 27236 10690 27282 10702
rect 27354 10878 27400 10890
rect 27354 10702 27360 10878
rect 27394 10702 27400 10878
rect 27354 10690 27400 10702
rect 27472 10878 27518 10890
rect 27472 10702 27478 10878
rect 27512 10702 27518 10878
rect 27472 10690 27518 10702
rect 27590 10878 27636 10890
rect 27720 10878 27726 11078
rect 27590 10702 27596 10878
rect 27630 10702 27726 10878
rect 27760 10702 27766 11078
rect 27590 10690 27636 10702
rect 27720 10690 27766 10702
rect 27838 11078 27884 11090
rect 27838 10702 27844 11078
rect 27878 10702 27884 11078
rect 27838 10690 27884 10702
rect 27956 11078 28002 11090
rect 27956 10702 27962 11078
rect 27996 10702 28002 11078
rect 27956 10690 28002 10702
rect 28074 11078 28120 11090
rect 28074 10702 28080 11078
rect 28114 10702 28120 11078
rect 28074 10690 28120 10702
rect 28192 11078 28238 11090
rect 28192 10702 28198 11078
rect 28232 10702 28238 11078
rect 28192 10690 28238 10702
rect 28310 11078 28356 11090
rect 28310 10702 28316 11078
rect 28350 10702 28356 11078
rect 28310 10690 28356 10702
rect 28428 11078 28474 11090
rect 28428 10702 28434 11078
rect 28468 10878 28474 11078
rect 28799 10890 28833 11193
rect 28557 10878 28603 10890
rect 28468 10702 28563 10878
rect 28597 10702 28603 10878
rect 28428 10690 28474 10702
rect 28557 10690 28603 10702
rect 28675 10878 28721 10890
rect 28675 10702 28681 10878
rect 28715 10702 28721 10878
rect 28675 10690 28721 10702
rect 28793 10878 28839 10890
rect 28793 10702 28799 10878
rect 28833 10702 28839 10878
rect 28793 10690 28839 10702
rect 28911 10878 28957 10890
rect 28911 10702 28917 10878
rect 28951 10702 28957 10878
rect 28911 10690 28957 10702
rect 24709 10641 24848 10647
rect 25344 10656 25378 10690
rect 25946 10656 25980 10690
rect 26182 10656 26216 10690
rect 24601 10612 24709 10622
rect 25344 10621 25503 10656
rect 25946 10621 26216 10656
rect 26783 10656 26817 10690
rect 27019 10656 27053 10690
rect 26783 10621 27053 10656
rect 27242 10656 27276 10690
rect 27844 10656 27878 10690
rect 28080 10656 28114 10690
rect 27242 10621 27401 10656
rect 27844 10621 28114 10656
rect 28681 10656 28715 10690
rect 28917 10656 28951 10690
rect 28681 10621 28951 10656
rect 23974 10580 23989 10582
rect 23889 10566 23989 10580
rect 23889 10523 23989 10524
rect 23510 10502 23989 10523
rect 24278 10502 24344 10598
rect 23510 10454 24344 10502
rect 23510 10425 23989 10454
rect 23510 10423 23615 10425
rect 23889 10424 23989 10425
rect 23343 10238 23353 10317
rect 23446 10238 23456 10317
rect 24344 10300 24423 10312
rect 22868 9911 22976 9923
rect 22864 9811 22874 9911
rect 22970 9811 22980 9911
rect 22868 9799 22976 9811
rect 23354 9064 23447 10238
rect 24344 10209 24350 10300
rect 24272 10189 24350 10209
rect 24417 10209 24423 10300
rect 24417 10189 24492 10209
rect 24272 10081 24316 10189
rect 24448 10081 24492 10189
rect 24272 10039 24492 10081
rect 23876 10009 24853 10039
rect 23876 9903 23908 10009
rect 24112 9903 24144 10009
rect 24348 9903 24380 10009
rect 24584 9903 24616 10009
rect 24819 9903 24853 10009
rect 23869 9891 23915 9903
rect 23869 9715 23875 9891
rect 23909 9715 23915 9891
rect 23869 9703 23915 9715
rect 23987 9891 24033 9903
rect 23987 9715 23993 9891
rect 24027 9715 24033 9891
rect 23987 9703 24033 9715
rect 24105 9891 24151 9903
rect 24105 9715 24111 9891
rect 24145 9715 24151 9891
rect 24105 9703 24151 9715
rect 24223 9891 24269 9903
rect 24223 9715 24229 9891
rect 24263 9715 24269 9891
rect 24223 9703 24269 9715
rect 24341 9891 24387 9903
rect 24341 9715 24347 9891
rect 24381 9715 24387 9891
rect 24341 9703 24387 9715
rect 24459 9891 24505 9903
rect 24459 9715 24465 9891
rect 24499 9715 24505 9891
rect 24459 9703 24505 9715
rect 24577 9891 24623 9903
rect 24577 9715 24583 9891
rect 24617 9715 24623 9891
rect 24577 9703 24623 9715
rect 24695 9891 24741 9903
rect 24695 9715 24701 9891
rect 24735 9715 24741 9891
rect 24695 9703 24741 9715
rect 24813 9891 24859 9903
rect 24813 9715 24819 9891
rect 24853 9715 24859 9891
rect 24813 9703 24859 9715
rect 24931 9891 24977 9903
rect 24931 9715 24937 9891
rect 24971 9715 24977 9891
rect 24931 9703 24977 9715
rect 25469 9837 25503 10621
rect 26182 10559 26216 10621
rect 25771 10521 26513 10559
rect 25771 10397 25805 10521
rect 26007 10397 26041 10521
rect 26243 10397 26277 10521
rect 26479 10397 26513 10521
rect 26769 10414 26779 10480
rect 26842 10414 26852 10480
rect 25765 10385 25811 10397
rect 25765 10009 25771 10385
rect 25805 10009 25811 10385
rect 25765 9997 25811 10009
rect 25883 10385 25929 10397
rect 25883 10009 25889 10385
rect 25923 10009 25929 10385
rect 25883 9997 25929 10009
rect 26001 10385 26047 10397
rect 26001 10009 26007 10385
rect 26041 10009 26047 10385
rect 26001 9997 26047 10009
rect 26119 10385 26165 10397
rect 26119 10009 26125 10385
rect 26159 10009 26165 10385
rect 26119 9997 26165 10009
rect 26237 10385 26283 10397
rect 26237 10009 26243 10385
rect 26277 10009 26283 10385
rect 26237 9997 26283 10009
rect 26355 10385 26401 10397
rect 26355 10009 26361 10385
rect 26395 10009 26401 10385
rect 26355 9997 26401 10009
rect 26473 10385 26519 10397
rect 26473 10009 26479 10385
rect 26513 10009 26519 10385
rect 26473 9997 26519 10009
rect 26885 9838 26919 10621
rect 26612 9837 26919 9838
rect 25469 9832 25785 9837
rect 26499 9832 26919 9837
rect 25469 9821 25852 9832
rect 25469 9794 25801 9821
rect 23992 9609 24028 9703
rect 24228 9609 24264 9703
rect 24464 9610 24500 9703
rect 24626 9655 24692 9662
rect 24626 9621 24642 9655
rect 24676 9621 24692 9655
rect 24626 9610 24692 9621
rect 24464 9609 24692 9610
rect 23992 9580 24692 9609
rect 23992 9579 24574 9580
rect 24112 9466 24146 9579
rect 24508 9538 24574 9579
rect 24508 9504 24524 9538
rect 24558 9504 24574 9538
rect 24508 9497 24574 9504
rect 24936 9470 24971 9703
rect 25469 9665 25503 9794
rect 25785 9787 25801 9794
rect 25835 9787 25852 9821
rect 25785 9781 25852 9787
rect 26432 9821 26919 9832
rect 26432 9787 26449 9821
rect 26483 9794 26919 9821
rect 26483 9787 26499 9794
rect 26612 9793 26919 9794
rect 26432 9781 26499 9787
rect 25610 9754 25666 9766
rect 25610 9720 25616 9754
rect 25650 9753 25666 9754
rect 26723 9753 26779 9765
rect 25650 9737 26117 9753
rect 25650 9720 26067 9737
rect 25610 9704 26067 9720
rect 26051 9703 26067 9704
rect 26101 9703 26117 9737
rect 26051 9696 26117 9703
rect 26169 9738 26739 9753
rect 26169 9704 26185 9738
rect 26219 9719 26739 9738
rect 26773 9719 26779 9753
rect 26219 9704 26779 9719
rect 26169 9694 26236 9704
rect 26723 9703 26779 9704
rect 26885 9665 26919 9793
rect 27367 9837 27401 10621
rect 28080 10559 28114 10621
rect 27669 10521 28411 10559
rect 27669 10397 27703 10521
rect 27905 10397 27939 10521
rect 28141 10397 28175 10521
rect 28377 10397 28411 10521
rect 27663 10385 27709 10397
rect 27663 10009 27669 10385
rect 27703 10009 27709 10385
rect 27663 9997 27709 10009
rect 27781 10385 27827 10397
rect 27781 10009 27787 10385
rect 27821 10009 27827 10385
rect 27781 9997 27827 10009
rect 27899 10385 27945 10397
rect 27899 10009 27905 10385
rect 27939 10009 27945 10385
rect 27899 9997 27945 10009
rect 28017 10385 28063 10397
rect 28017 10009 28023 10385
rect 28057 10009 28063 10385
rect 28017 9997 28063 10009
rect 28135 10385 28181 10397
rect 28135 10009 28141 10385
rect 28175 10009 28181 10385
rect 28135 9997 28181 10009
rect 28253 10385 28299 10397
rect 28253 10009 28259 10385
rect 28293 10009 28299 10385
rect 28253 9997 28299 10009
rect 28371 10385 28417 10397
rect 28371 10009 28377 10385
rect 28411 10009 28417 10385
rect 28371 9997 28417 10009
rect 28783 9838 28817 10621
rect 28395 9837 28464 9838
rect 28510 9837 28817 9838
rect 27367 9832 27683 9837
rect 28395 9833 28817 9837
rect 27367 9821 27750 9832
rect 27367 9794 27699 9821
rect 27367 9665 27401 9794
rect 27683 9787 27699 9794
rect 27733 9787 27750 9821
rect 27683 9781 27750 9787
rect 28328 9822 28817 9833
rect 28328 9788 28345 9822
rect 28379 9794 28817 9822
rect 28379 9788 28395 9794
rect 28510 9793 28817 9794
rect 28328 9782 28395 9788
rect 27508 9754 27564 9766
rect 27508 9720 27514 9754
rect 27548 9753 27564 9754
rect 28621 9753 28677 9765
rect 27548 9737 28015 9753
rect 27548 9720 27965 9737
rect 27508 9704 27965 9720
rect 27949 9703 27965 9704
rect 27999 9703 28015 9737
rect 27949 9696 28015 9703
rect 28067 9738 28637 9753
rect 28067 9704 28083 9738
rect 28117 9719 28637 9738
rect 28671 9719 28677 9753
rect 28117 9704 28677 9719
rect 28067 9694 28134 9704
rect 28621 9703 28677 9704
rect 28783 9665 28817 9793
rect 28898 10443 28965 10467
rect 28898 10409 28915 10443
rect 28949 10409 28965 10443
rect 24582 9466 24971 9470
rect 24106 9454 24152 9466
rect 24106 9078 24112 9454
rect 24146 9078 24152 9454
rect 24106 9066 24152 9078
rect 24224 9454 24270 9466
rect 24224 9078 24230 9454
rect 24264 9078 24270 9454
rect 24224 9066 24270 9078
rect 24342 9454 24388 9466
rect 24342 9078 24348 9454
rect 24382 9102 24388 9454
rect 24459 9454 24505 9466
rect 24459 9278 24465 9454
rect 24499 9278 24505 9454
rect 24459 9266 24505 9278
rect 24577 9454 24971 9466
rect 25463 9653 25509 9665
rect 25463 9477 25469 9653
rect 25503 9477 25509 9653
rect 25463 9465 25509 9477
rect 25581 9653 25627 9665
rect 25581 9477 25587 9653
rect 25621 9477 25627 9653
rect 25581 9465 25627 9477
rect 25883 9653 25929 9665
rect 24577 9278 24583 9454
rect 24617 9441 24971 9454
rect 24617 9278 24623 9441
rect 24893 9438 24971 9441
rect 24893 9386 24903 9438
rect 24966 9386 24976 9438
rect 24898 9380 24971 9386
rect 24577 9266 24623 9278
rect 24465 9150 24500 9266
rect 25586 9171 25620 9465
rect 25883 9277 25889 9653
rect 25923 9277 25929 9653
rect 25883 9265 25929 9277
rect 26001 9653 26047 9665
rect 26001 9277 26007 9653
rect 26041 9277 26047 9653
rect 26001 9265 26047 9277
rect 26119 9653 26165 9665
rect 26119 9277 26125 9653
rect 26159 9277 26165 9653
rect 26119 9265 26165 9277
rect 26237 9653 26283 9665
rect 26237 9277 26243 9653
rect 26277 9277 26283 9653
rect 26237 9265 26283 9277
rect 26355 9653 26401 9665
rect 26355 9277 26361 9653
rect 26395 9277 26401 9653
rect 26761 9653 26807 9665
rect 26761 9477 26767 9653
rect 26801 9477 26807 9653
rect 26761 9465 26807 9477
rect 26879 9653 26925 9665
rect 26879 9477 26885 9653
rect 26919 9477 26925 9653
rect 26879 9465 26925 9477
rect 27361 9653 27407 9665
rect 27361 9477 27367 9653
rect 27401 9477 27407 9653
rect 27361 9465 27407 9477
rect 27479 9653 27525 9665
rect 27479 9477 27485 9653
rect 27519 9477 27525 9653
rect 27479 9465 27525 9477
rect 27781 9653 27827 9665
rect 26355 9265 26401 9277
rect 26243 9171 26277 9265
rect 26767 9171 26800 9465
rect 24596 9150 24704 9160
rect 24465 9102 24596 9150
rect 25586 9139 26800 9171
rect 27484 9171 27518 9465
rect 27781 9277 27787 9653
rect 27821 9277 27827 9653
rect 27781 9265 27827 9277
rect 27899 9653 27945 9665
rect 27899 9277 27905 9653
rect 27939 9277 27945 9653
rect 27899 9265 27945 9277
rect 28017 9653 28063 9665
rect 28017 9277 28023 9653
rect 28057 9277 28063 9653
rect 28017 9265 28063 9277
rect 28135 9653 28181 9665
rect 28135 9277 28141 9653
rect 28175 9277 28181 9653
rect 28135 9265 28181 9277
rect 28253 9653 28299 9665
rect 28253 9277 28259 9653
rect 28293 9277 28299 9653
rect 28659 9653 28705 9665
rect 28659 9477 28665 9653
rect 28699 9477 28705 9653
rect 28659 9465 28705 9477
rect 28777 9653 28823 9665
rect 28777 9477 28783 9653
rect 28817 9477 28823 9653
rect 28777 9465 28823 9477
rect 28253 9265 28299 9277
rect 28141 9171 28175 9265
rect 28665 9171 28698 9465
rect 27484 9139 28698 9171
rect 24704 9109 24854 9115
rect 24382 9078 24596 9102
rect 24342 9066 24596 9078
rect 23354 9062 23939 9064
rect 24348 9062 24596 9066
rect 23354 9034 23984 9062
rect 23354 9028 24221 9034
rect 23354 8994 24171 9028
rect 24205 8994 24221 9028
rect 23354 8978 24221 8994
rect 24273 9028 24339 9034
rect 24273 8994 24289 9028
rect 24323 8994 24339 9028
rect 24522 9018 24596 9062
rect 24842 9042 24854 9109
rect 26079 9054 26211 9139
rect 27977 9054 28109 9139
rect 24704 9036 24854 9042
rect 24596 9008 24704 9018
rect 23354 8962 23984 8978
rect 23354 8958 23939 8962
rect 23354 8957 23455 8958
rect 23884 8909 23984 8920
rect 23848 8803 23858 8909
rect 23970 8898 23984 8909
rect 24273 8898 24339 8994
rect 26069 8946 26079 9054
rect 26211 8946 26221 9054
rect 27967 8946 27977 9054
rect 28109 8946 28119 9054
rect 28898 9026 28965 10409
rect 29111 9986 29211 15590
rect 30845 15458 30940 15461
rect 30840 15452 30942 15458
rect 30840 15380 30852 15452
rect 30930 15380 30942 15452
rect 30840 15374 30942 15380
rect 32098 15410 32543 15416
rect 29973 15315 30109 15335
rect 29973 15253 30009 15315
rect 30069 15253 30109 15315
rect 29973 15225 30109 15253
rect 29669 15195 30646 15225
rect 29669 15089 29701 15195
rect 29905 15089 29937 15195
rect 30141 15089 30173 15195
rect 30377 15089 30409 15195
rect 30612 15089 30646 15195
rect 29662 15077 29708 15089
rect 29662 14901 29668 15077
rect 29702 14901 29708 15077
rect 29662 14889 29708 14901
rect 29780 15077 29826 15089
rect 29780 14901 29786 15077
rect 29820 14901 29826 15077
rect 29780 14889 29826 14901
rect 29898 15077 29944 15089
rect 29898 14901 29904 15077
rect 29938 14901 29944 15077
rect 29898 14889 29944 14901
rect 30016 15077 30062 15089
rect 30016 14901 30022 15077
rect 30056 14901 30062 15077
rect 30016 14889 30062 14901
rect 30134 15077 30180 15089
rect 30134 14901 30140 15077
rect 30174 14901 30180 15077
rect 30134 14889 30180 14901
rect 30252 15077 30298 15089
rect 30252 14901 30258 15077
rect 30292 14901 30298 15077
rect 30252 14889 30298 14901
rect 30370 15077 30416 15089
rect 30370 14901 30376 15077
rect 30410 14901 30416 15077
rect 30370 14889 30416 14901
rect 30488 15077 30534 15089
rect 30488 14901 30494 15077
rect 30528 14901 30534 15077
rect 30488 14889 30534 14901
rect 30606 15077 30652 15089
rect 30606 14901 30612 15077
rect 30646 14901 30652 15077
rect 30606 14889 30652 14901
rect 30724 15077 30770 15089
rect 30724 14901 30730 15077
rect 30764 14901 30770 15077
rect 30724 14889 30770 14901
rect 29785 14795 29821 14889
rect 30021 14795 30057 14889
rect 30257 14796 30293 14889
rect 30419 14841 30485 14848
rect 30419 14807 30435 14841
rect 30469 14807 30485 14841
rect 30419 14796 30485 14807
rect 30257 14795 30485 14796
rect 29785 14766 30485 14795
rect 29785 14765 30367 14766
rect 29905 14652 29939 14765
rect 30301 14724 30367 14765
rect 30301 14690 30317 14724
rect 30351 14690 30367 14724
rect 30301 14683 30367 14690
rect 30729 14657 30764 14889
rect 30845 14657 30940 15374
rect 32098 15210 32110 15410
rect 32531 15210 32543 15410
rect 32098 15204 32266 15210
rect 32256 15136 32266 15204
rect 32398 15204 32543 15210
rect 32398 15136 32408 15204
rect 32266 15096 32398 15136
rect 32265 15030 32398 15096
rect 31594 14987 33067 15030
rect 31594 14684 31628 14987
rect 31960 14884 31994 14987
rect 32196 14884 32230 14987
rect 32432 14884 32466 14987
rect 32668 14884 32702 14987
rect 31954 14872 32000 14884
rect 30674 14656 30940 14657
rect 30375 14652 30940 14656
rect 29899 14640 29945 14652
rect 29899 14264 29905 14640
rect 29939 14264 29945 14640
rect 29899 14252 29945 14264
rect 30017 14640 30063 14652
rect 30017 14264 30023 14640
rect 30057 14264 30063 14640
rect 30017 14252 30063 14264
rect 30135 14640 30181 14652
rect 30135 14264 30141 14640
rect 30175 14291 30181 14640
rect 30252 14640 30298 14652
rect 30252 14464 30258 14640
rect 30292 14464 30298 14640
rect 30252 14457 30298 14464
rect 30370 14640 30940 14652
rect 30370 14464 30376 14640
rect 30410 14627 30940 14640
rect 30410 14464 30416 14627
rect 30660 14547 30940 14627
rect 30674 14546 30940 14547
rect 31470 14672 31516 14684
rect 31470 14496 31476 14672
rect 31510 14496 31516 14672
rect 31470 14484 31516 14496
rect 31588 14672 31634 14684
rect 31588 14496 31594 14672
rect 31628 14496 31634 14672
rect 31588 14484 31634 14496
rect 31706 14672 31752 14684
rect 31706 14496 31712 14672
rect 31746 14496 31752 14672
rect 31706 14484 31752 14496
rect 31824 14672 31870 14684
rect 31954 14672 31960 14872
rect 31824 14496 31830 14672
rect 31864 14496 31960 14672
rect 31994 14496 32000 14872
rect 31824 14484 31870 14496
rect 31954 14484 32000 14496
rect 32072 14872 32118 14884
rect 32072 14496 32078 14872
rect 32112 14496 32118 14872
rect 32072 14484 32118 14496
rect 32190 14872 32236 14884
rect 32190 14496 32196 14872
rect 32230 14496 32236 14872
rect 32190 14484 32236 14496
rect 32308 14872 32354 14884
rect 32308 14496 32314 14872
rect 32348 14496 32354 14872
rect 32308 14484 32354 14496
rect 32426 14872 32472 14884
rect 32426 14496 32432 14872
rect 32466 14496 32472 14872
rect 32426 14484 32472 14496
rect 32544 14872 32590 14884
rect 32544 14496 32550 14872
rect 32584 14496 32590 14872
rect 32544 14484 32590 14496
rect 32662 14872 32708 14884
rect 32662 14496 32668 14872
rect 32702 14672 32708 14872
rect 33033 14684 33067 14987
rect 33574 14907 33710 14927
rect 33574 14845 33610 14907
rect 33670 14845 33710 14907
rect 33574 14817 33710 14845
rect 33270 14787 34247 14817
rect 32791 14672 32837 14684
rect 32702 14496 32797 14672
rect 32831 14496 32837 14672
rect 32662 14484 32708 14496
rect 32791 14484 32837 14496
rect 32909 14672 32955 14684
rect 32909 14496 32915 14672
rect 32949 14496 32955 14672
rect 32909 14484 32955 14496
rect 33027 14672 33073 14684
rect 33027 14496 33033 14672
rect 33067 14496 33073 14672
rect 33027 14484 33073 14496
rect 33145 14672 33191 14684
rect 33270 14681 33302 14787
rect 33506 14681 33538 14787
rect 33742 14681 33774 14787
rect 33978 14681 34010 14787
rect 34213 14681 34247 14787
rect 33145 14496 33151 14672
rect 33185 14496 33191 14672
rect 33145 14484 33191 14496
rect 33263 14669 33309 14681
rect 33263 14493 33269 14669
rect 33303 14493 33309 14669
rect 30252 14452 30301 14457
rect 30370 14452 30416 14464
rect 30258 14291 30301 14452
rect 31476 14450 31510 14484
rect 32078 14450 32112 14484
rect 32314 14450 32348 14484
rect 31476 14415 31635 14450
rect 32078 14415 32348 14450
rect 32915 14450 32949 14484
rect 33151 14450 33185 14484
rect 33263 14481 33309 14493
rect 33381 14669 33427 14681
rect 33381 14493 33387 14669
rect 33421 14493 33427 14669
rect 33381 14481 33427 14493
rect 33499 14669 33545 14681
rect 33499 14493 33505 14669
rect 33539 14493 33545 14669
rect 33499 14481 33545 14493
rect 33617 14669 33663 14681
rect 33617 14493 33623 14669
rect 33657 14493 33663 14669
rect 33617 14481 33663 14493
rect 33735 14669 33781 14681
rect 33735 14493 33741 14669
rect 33775 14493 33781 14669
rect 33735 14481 33781 14493
rect 33853 14669 33899 14681
rect 33853 14493 33859 14669
rect 33893 14493 33899 14669
rect 33853 14481 33899 14493
rect 33971 14669 34017 14681
rect 33971 14493 33977 14669
rect 34011 14493 34017 14669
rect 33971 14481 34017 14493
rect 34089 14669 34135 14681
rect 34089 14493 34095 14669
rect 34129 14493 34135 14669
rect 34089 14481 34135 14493
rect 34207 14669 34253 14681
rect 34207 14493 34213 14669
rect 34247 14493 34253 14669
rect 34207 14481 34253 14493
rect 34325 14669 34371 14681
rect 34325 14493 34331 14669
rect 34365 14493 34371 14669
rect 34325 14481 34371 14493
rect 32915 14415 33185 14450
rect 31412 14333 31541 14334
rect 30175 14264 30301 14291
rect 30135 14252 30301 14264
rect 30141 14248 30301 14252
rect 29349 14246 29436 14247
rect 29349 14242 29732 14246
rect 29344 14168 29354 14242
rect 29433 14221 29732 14242
rect 29433 14220 29866 14221
rect 29433 14214 30014 14220
rect 29433 14180 29964 14214
rect 29998 14180 30014 14214
rect 29433 14168 30014 14180
rect 29026 9980 29211 9986
rect 29026 9882 29038 9980
rect 29170 9882 29211 9980
rect 29026 9876 29211 9882
rect 29111 9875 29211 9876
rect 29349 14164 30014 14168
rect 30066 14214 30132 14220
rect 30066 14180 30082 14214
rect 30116 14180 30132 14214
rect 23970 8850 24339 8898
rect 23970 8820 23984 8850
rect 23970 8803 23980 8820
rect 24272 8747 24338 8850
rect 26103 8808 26109 8946
rect 26176 8808 26182 8946
rect 26103 8796 26182 8808
rect 28898 8747 28964 9026
rect 24270 8667 28964 8747
rect 29349 8780 29439 14164
rect 30066 14135 30132 14180
rect 29499 14128 30132 14135
rect 29496 14032 29506 14128
rect 29587 14127 30132 14128
rect 29587 14095 30133 14127
rect 30225 14111 30301 14248
rect 31011 14330 31541 14333
rect 31011 14267 31463 14330
rect 31530 14267 31541 14330
rect 31011 14264 31541 14267
rect 29587 14032 29732 14095
rect 30221 14051 30231 14111
rect 30293 14051 30303 14111
rect 31011 14044 31153 14264
rect 31443 14208 31547 14214
rect 31443 14140 31455 14208
rect 31535 14140 31547 14208
rect 31443 14134 31547 14140
rect 29499 11941 29593 14032
rect 29968 12744 30104 12764
rect 29968 12682 30004 12744
rect 30064 12682 30104 12744
rect 29968 12654 30104 12682
rect 29664 12624 30641 12654
rect 29664 12518 29696 12624
rect 29900 12518 29932 12624
rect 30136 12518 30168 12624
rect 30372 12518 30404 12624
rect 30607 12518 30641 12624
rect 29657 12506 29703 12518
rect 29657 12330 29663 12506
rect 29697 12330 29703 12506
rect 29657 12318 29703 12330
rect 29775 12506 29821 12518
rect 29775 12330 29781 12506
rect 29815 12330 29821 12506
rect 29775 12318 29821 12330
rect 29893 12506 29939 12518
rect 29893 12330 29899 12506
rect 29933 12330 29939 12506
rect 29893 12318 29939 12330
rect 30011 12506 30057 12518
rect 30011 12330 30017 12506
rect 30051 12330 30057 12506
rect 30011 12318 30057 12330
rect 30129 12506 30175 12518
rect 30129 12330 30135 12506
rect 30169 12330 30175 12506
rect 30129 12318 30175 12330
rect 30247 12506 30293 12518
rect 30247 12330 30253 12506
rect 30287 12330 30293 12506
rect 30247 12318 30293 12330
rect 30365 12506 30411 12518
rect 30365 12330 30371 12506
rect 30405 12330 30411 12506
rect 30365 12318 30411 12330
rect 30483 12506 30529 12518
rect 30483 12330 30489 12506
rect 30523 12330 30529 12506
rect 30483 12318 30529 12330
rect 30601 12506 30647 12518
rect 30601 12330 30607 12506
rect 30641 12330 30647 12506
rect 30601 12318 30647 12330
rect 30719 12506 30765 12518
rect 30719 12330 30725 12506
rect 30759 12330 30765 12506
rect 30719 12318 30765 12330
rect 29780 12224 29816 12318
rect 30016 12224 30052 12318
rect 30252 12225 30288 12318
rect 30414 12270 30480 12277
rect 30414 12236 30430 12270
rect 30464 12236 30480 12270
rect 30414 12225 30480 12236
rect 30252 12224 30480 12225
rect 29780 12195 30480 12224
rect 29780 12194 30362 12195
rect 29900 12081 29934 12194
rect 30296 12153 30362 12194
rect 30296 12119 30312 12153
rect 30346 12119 30362 12153
rect 30296 12112 30362 12119
rect 30724 12085 30759 12318
rect 31011 12085 31152 14044
rect 31601 13631 31635 14415
rect 32314 14353 32348 14415
rect 31903 14315 32645 14353
rect 31713 14144 31723 14212
rect 31778 14144 31788 14212
rect 31903 14191 31937 14315
rect 32139 14191 32173 14315
rect 32375 14191 32409 14315
rect 32611 14191 32645 14315
rect 31897 14179 31943 14191
rect 31897 13803 31903 14179
rect 31937 13803 31943 14179
rect 31897 13791 31943 13803
rect 32015 14179 32061 14191
rect 32015 13803 32021 14179
rect 32055 13803 32061 14179
rect 32015 13791 32061 13803
rect 32133 14179 32179 14191
rect 32133 13803 32139 14179
rect 32173 13803 32179 14179
rect 32133 13791 32179 13803
rect 32251 14179 32297 14191
rect 32251 13803 32257 14179
rect 32291 13803 32297 14179
rect 32251 13791 32297 13803
rect 32369 14179 32415 14191
rect 32369 13803 32375 14179
rect 32409 13803 32415 14179
rect 32369 13791 32415 13803
rect 32487 14179 32533 14191
rect 32487 13803 32493 14179
rect 32527 13803 32533 14179
rect 32487 13791 32533 13803
rect 32605 14179 32651 14191
rect 32605 13803 32611 14179
rect 32645 13803 32651 14179
rect 32771 13974 32845 13986
rect 32767 13883 32777 13974
rect 32839 13883 32849 13974
rect 32771 13871 32845 13883
rect 32605 13791 32651 13803
rect 33017 13632 33051 14415
rect 33386 14387 33422 14481
rect 33622 14387 33658 14481
rect 33858 14388 33894 14481
rect 34020 14433 34086 14440
rect 34020 14399 34036 14433
rect 34070 14399 34086 14433
rect 34020 14388 34086 14399
rect 33858 14387 34086 14388
rect 33386 14358 34086 14387
rect 33386 14357 33968 14358
rect 33112 14325 33188 14330
rect 33109 14269 33119 14325
rect 33172 14324 33188 14325
rect 33172 14269 33438 14324
rect 33112 14264 33438 14269
rect 33233 14222 33324 14227
rect 33233 14133 33243 14222
rect 33316 14133 33324 14222
rect 33233 14121 33324 14133
rect 33270 13727 33324 14121
rect 33384 13812 33438 14264
rect 33506 14244 33540 14357
rect 33902 14316 33968 14357
rect 33902 14282 33918 14316
rect 33952 14282 33968 14316
rect 33902 14275 33968 14282
rect 34330 14248 34365 14481
rect 33976 14244 34365 14248
rect 33500 14232 33546 14244
rect 33500 13856 33506 14232
rect 33540 13856 33546 14232
rect 33500 13844 33546 13856
rect 33618 14232 33664 14244
rect 33618 13856 33624 14232
rect 33658 13856 33664 14232
rect 33618 13844 33664 13856
rect 33736 14232 33782 14244
rect 33736 13856 33742 14232
rect 33776 13883 33782 14232
rect 33853 14232 33899 14244
rect 33853 14056 33859 14232
rect 33893 14056 33899 14232
rect 33853 14049 33899 14056
rect 33971 14232 34365 14244
rect 33971 14056 33977 14232
rect 34011 14219 34365 14232
rect 34011 14056 34017 14219
rect 34190 14217 34365 14219
rect 34190 14159 34232 14217
rect 34344 14159 34365 14217
rect 34190 14130 34365 14159
rect 33853 14044 33902 14049
rect 33971 14044 34017 14056
rect 33859 13883 33902 14044
rect 33776 13856 33902 13883
rect 34000 13984 34328 13985
rect 34000 13977 34394 13984
rect 34000 13969 34254 13977
rect 34000 13888 34016 13969
rect 34124 13888 34254 13969
rect 34000 13883 34254 13888
rect 34377 13883 34394 13977
rect 34000 13871 34394 13883
rect 34244 13870 34394 13871
rect 33736 13844 33902 13856
rect 33742 13840 33902 13844
rect 33384 13806 33615 13812
rect 33384 13772 33565 13806
rect 33599 13772 33615 13806
rect 33384 13756 33615 13772
rect 33667 13806 33733 13812
rect 33667 13772 33683 13806
rect 33717 13772 33733 13806
rect 33667 13727 33733 13772
rect 33270 13719 33733 13727
rect 33270 13687 33734 13719
rect 33826 13703 33902 13840
rect 33822 13643 33832 13703
rect 33894 13643 33904 13703
rect 32744 13631 33051 13632
rect 31601 13626 31917 13631
rect 32631 13626 33051 13631
rect 31601 13615 31984 13626
rect 31601 13588 31933 13615
rect 31601 13459 31635 13588
rect 31917 13581 31933 13588
rect 31967 13581 31984 13615
rect 31917 13575 31984 13581
rect 32564 13615 33051 13626
rect 33830 13617 33900 13643
rect 32564 13581 32581 13615
rect 32615 13588 33051 13615
rect 32615 13581 32631 13588
rect 32744 13587 33051 13588
rect 32564 13575 32631 13581
rect 31742 13548 31798 13560
rect 31742 13514 31748 13548
rect 31782 13547 31798 13548
rect 32855 13547 32911 13559
rect 31782 13531 32249 13547
rect 31782 13514 32199 13531
rect 31742 13498 32199 13514
rect 32183 13497 32199 13498
rect 32233 13497 32249 13531
rect 32183 13490 32249 13497
rect 32301 13532 32871 13547
rect 32301 13498 32317 13532
rect 32351 13513 32871 13532
rect 32905 13513 32911 13547
rect 32351 13498 32911 13513
rect 32301 13488 32368 13498
rect 32855 13497 32911 13498
rect 33017 13459 33051 13587
rect 31595 13447 31641 13459
rect 31595 13271 31601 13447
rect 31635 13271 31641 13447
rect 31595 13259 31641 13271
rect 31713 13447 31759 13459
rect 31713 13271 31719 13447
rect 31753 13271 31759 13447
rect 31713 13259 31759 13271
rect 32015 13447 32061 13459
rect 31718 12965 31752 13259
rect 32015 13071 32021 13447
rect 32055 13071 32061 13447
rect 32015 13059 32061 13071
rect 32133 13447 32179 13459
rect 32133 13071 32139 13447
rect 32173 13071 32179 13447
rect 32133 13059 32179 13071
rect 32251 13447 32297 13459
rect 32251 13071 32257 13447
rect 32291 13071 32297 13447
rect 32251 13059 32297 13071
rect 32369 13447 32415 13459
rect 32369 13071 32375 13447
rect 32409 13071 32415 13447
rect 32369 13059 32415 13071
rect 32487 13447 32533 13459
rect 32487 13071 32493 13447
rect 32527 13071 32533 13447
rect 32893 13447 32939 13459
rect 32893 13271 32899 13447
rect 32933 13271 32939 13447
rect 32893 13259 32939 13271
rect 33011 13447 33057 13459
rect 33011 13271 33017 13447
rect 33051 13271 33057 13447
rect 33011 13259 33057 13271
rect 32487 13059 32533 13071
rect 32375 12965 32409 13059
rect 32899 12965 32932 13259
rect 31718 12933 32932 12965
rect 32084 12909 32490 12933
rect 32084 12786 32196 12909
rect 32370 12786 32490 12909
rect 32084 12742 32490 12786
rect 30370 12081 31152 12085
rect 29894 12069 29940 12081
rect 29499 11844 29832 11941
rect 29642 11801 29742 11813
rect 29642 11720 29653 11801
rect 29735 11720 29745 11801
rect 29642 11713 29742 11720
rect 29664 11564 29718 11713
rect 29778 11649 29832 11844
rect 29894 11693 29900 12069
rect 29934 11693 29940 12069
rect 29894 11681 29940 11693
rect 30012 12069 30058 12081
rect 30012 11693 30018 12069
rect 30052 11693 30058 12069
rect 30012 11681 30058 11693
rect 30130 12069 30176 12081
rect 30130 11693 30136 12069
rect 30170 11720 30176 12069
rect 30247 12069 30293 12081
rect 30247 11893 30253 12069
rect 30287 11893 30293 12069
rect 30247 11886 30293 11893
rect 30365 12069 31152 12081
rect 30365 11893 30371 12069
rect 30405 12056 31152 12069
rect 30405 11893 30411 12056
rect 30655 11974 31152 12056
rect 30247 11881 30296 11886
rect 30365 11881 30411 11893
rect 30253 11720 30296 11881
rect 30170 11693 30296 11720
rect 30130 11681 30296 11693
rect 30136 11677 30296 11681
rect 29778 11643 30009 11649
rect 29778 11609 29959 11643
rect 29993 11609 30009 11643
rect 29778 11593 30009 11609
rect 30061 11643 30127 11649
rect 30061 11609 30077 11643
rect 30111 11609 30127 11643
rect 30061 11564 30127 11609
rect 29664 11556 30127 11564
rect 29664 11524 30128 11556
rect 30220 11540 30296 11677
rect 30216 11480 30226 11540
rect 30288 11480 30298 11540
rect 32100 11319 32545 11325
rect 32100 11119 32112 11319
rect 32533 11119 32545 11319
rect 32100 11113 32268 11119
rect 32258 11045 32268 11113
rect 32400 11113 32545 11119
rect 32400 11045 32410 11113
rect 32268 11005 32400 11045
rect 32267 10939 32400 11005
rect 31596 10896 33069 10939
rect 31596 10593 31630 10896
rect 31962 10793 31996 10896
rect 32198 10793 32232 10896
rect 32434 10793 32468 10896
rect 32670 10793 32704 10896
rect 31956 10781 32002 10793
rect 31472 10581 31518 10593
rect 31472 10405 31478 10581
rect 31512 10405 31518 10581
rect 31472 10393 31518 10405
rect 31590 10581 31636 10593
rect 31590 10405 31596 10581
rect 31630 10405 31636 10581
rect 31590 10393 31636 10405
rect 31708 10581 31754 10593
rect 31708 10405 31714 10581
rect 31748 10405 31754 10581
rect 31708 10393 31754 10405
rect 31826 10581 31872 10593
rect 31956 10581 31962 10781
rect 31826 10405 31832 10581
rect 31866 10405 31962 10581
rect 31996 10405 32002 10781
rect 31826 10393 31872 10405
rect 31956 10393 32002 10405
rect 32074 10781 32120 10793
rect 32074 10405 32080 10781
rect 32114 10405 32120 10781
rect 32074 10393 32120 10405
rect 32192 10781 32238 10793
rect 32192 10405 32198 10781
rect 32232 10405 32238 10781
rect 32192 10393 32238 10405
rect 32310 10781 32356 10793
rect 32310 10405 32316 10781
rect 32350 10405 32356 10781
rect 32310 10393 32356 10405
rect 32428 10781 32474 10793
rect 32428 10405 32434 10781
rect 32468 10405 32474 10781
rect 32428 10393 32474 10405
rect 32546 10781 32592 10793
rect 32546 10405 32552 10781
rect 32586 10405 32592 10781
rect 32546 10393 32592 10405
rect 32664 10781 32710 10793
rect 32664 10405 32670 10781
rect 32704 10581 32710 10781
rect 33035 10593 33069 10896
rect 33576 10816 33712 10836
rect 33576 10754 33612 10816
rect 33672 10754 33712 10816
rect 33576 10726 33712 10754
rect 33272 10696 34249 10726
rect 32793 10581 32839 10593
rect 32704 10405 32799 10581
rect 32833 10405 32839 10581
rect 32664 10393 32710 10405
rect 32793 10393 32839 10405
rect 32911 10581 32957 10593
rect 32911 10405 32917 10581
rect 32951 10405 32957 10581
rect 32911 10393 32957 10405
rect 33029 10581 33075 10593
rect 33029 10405 33035 10581
rect 33069 10405 33075 10581
rect 33029 10393 33075 10405
rect 33147 10581 33193 10593
rect 33272 10590 33304 10696
rect 33508 10590 33540 10696
rect 33744 10590 33776 10696
rect 33980 10590 34012 10696
rect 34215 10590 34249 10696
rect 33147 10405 33153 10581
rect 33187 10405 33193 10581
rect 33147 10393 33193 10405
rect 33265 10578 33311 10590
rect 33265 10402 33271 10578
rect 33305 10402 33311 10578
rect 31478 10359 31512 10393
rect 32080 10359 32114 10393
rect 32316 10359 32350 10393
rect 31478 10324 31637 10359
rect 32080 10324 32350 10359
rect 32917 10359 32951 10393
rect 33153 10359 33187 10393
rect 33265 10390 33311 10402
rect 33383 10578 33429 10590
rect 33383 10402 33389 10578
rect 33423 10402 33429 10578
rect 33383 10390 33429 10402
rect 33501 10578 33547 10590
rect 33501 10402 33507 10578
rect 33541 10402 33547 10578
rect 33501 10390 33547 10402
rect 33619 10578 33665 10590
rect 33619 10402 33625 10578
rect 33659 10402 33665 10578
rect 33619 10390 33665 10402
rect 33737 10578 33783 10590
rect 33737 10402 33743 10578
rect 33777 10402 33783 10578
rect 33737 10390 33783 10402
rect 33855 10578 33901 10590
rect 33855 10402 33861 10578
rect 33895 10402 33901 10578
rect 33855 10390 33901 10402
rect 33973 10578 34019 10590
rect 33973 10402 33979 10578
rect 34013 10402 34019 10578
rect 33973 10390 34019 10402
rect 34091 10578 34137 10590
rect 34091 10402 34097 10578
rect 34131 10402 34137 10578
rect 34091 10390 34137 10402
rect 34209 10578 34255 10590
rect 34209 10402 34215 10578
rect 34249 10402 34255 10578
rect 34209 10390 34255 10402
rect 34327 10578 34373 10590
rect 34327 10402 34333 10578
rect 34367 10402 34373 10578
rect 34327 10390 34373 10402
rect 32917 10324 33187 10359
rect 30847 10176 31465 10239
rect 31532 10176 31542 10239
rect 30847 10175 31501 10176
rect 29968 9711 30104 9731
rect 29968 9649 30004 9711
rect 30064 9649 30104 9711
rect 29968 9621 30104 9649
rect 29664 9591 30641 9621
rect 29664 9485 29696 9591
rect 29900 9485 29932 9591
rect 30136 9485 30168 9591
rect 30372 9485 30404 9591
rect 30607 9485 30641 9591
rect 29657 9473 29703 9485
rect 29657 9297 29663 9473
rect 29697 9297 29703 9473
rect 29657 9285 29703 9297
rect 29775 9473 29821 9485
rect 29775 9297 29781 9473
rect 29815 9297 29821 9473
rect 29775 9285 29821 9297
rect 29893 9473 29939 9485
rect 29893 9297 29899 9473
rect 29933 9297 29939 9473
rect 29893 9285 29939 9297
rect 30011 9473 30057 9485
rect 30011 9297 30017 9473
rect 30051 9297 30057 9473
rect 30011 9285 30057 9297
rect 30129 9473 30175 9485
rect 30129 9297 30135 9473
rect 30169 9297 30175 9473
rect 30129 9285 30175 9297
rect 30247 9473 30293 9485
rect 30247 9297 30253 9473
rect 30287 9297 30293 9473
rect 30247 9285 30293 9297
rect 30365 9473 30411 9485
rect 30365 9297 30371 9473
rect 30405 9297 30411 9473
rect 30365 9285 30411 9297
rect 30483 9473 30529 9485
rect 30483 9297 30489 9473
rect 30523 9297 30529 9473
rect 30483 9285 30529 9297
rect 30601 9473 30647 9485
rect 30601 9297 30607 9473
rect 30641 9297 30647 9473
rect 30601 9285 30647 9297
rect 30719 9473 30765 9485
rect 30719 9297 30725 9473
rect 30759 9297 30765 9473
rect 30719 9285 30765 9297
rect 29780 9191 29816 9285
rect 30016 9191 30052 9285
rect 30252 9192 30288 9285
rect 30414 9237 30480 9244
rect 30414 9203 30430 9237
rect 30464 9203 30480 9237
rect 30414 9192 30480 9203
rect 30252 9191 30480 9192
rect 29780 9162 30480 9191
rect 29780 9161 30362 9162
rect 29900 9048 29934 9161
rect 30296 9120 30362 9161
rect 30296 9086 30312 9120
rect 30346 9086 30362 9120
rect 30296 9079 30362 9086
rect 30724 9052 30759 9285
rect 30847 9052 30938 10175
rect 30370 9048 30938 9052
rect 29894 9036 29940 9048
rect 29754 8900 29854 8908
rect 29748 8813 29758 8900
rect 29847 8813 29857 8900
rect 29754 8808 29854 8813
rect 29349 8680 29718 8780
rect 23504 8485 23514 8599
rect 23637 8485 23647 8599
rect 29664 8531 29718 8680
rect 29778 8616 29832 8808
rect 29894 8660 29900 9036
rect 29934 8660 29940 9036
rect 29894 8648 29940 8660
rect 30012 9036 30058 9048
rect 30012 8660 30018 9036
rect 30052 8660 30058 9036
rect 30012 8648 30058 8660
rect 30130 9036 30176 9048
rect 30130 8660 30136 9036
rect 30170 8687 30176 9036
rect 30247 9036 30293 9048
rect 30247 8860 30253 9036
rect 30287 8860 30293 9036
rect 30247 8853 30293 8860
rect 30365 9036 30938 9048
rect 30365 8860 30371 9036
rect 30405 9023 30938 9036
rect 30405 8860 30411 9023
rect 30655 8943 30938 9023
rect 31027 10050 31465 10113
rect 31532 10050 31542 10113
rect 30247 8848 30296 8853
rect 30365 8848 30411 8860
rect 30253 8687 30296 8848
rect 30170 8660 30296 8687
rect 30130 8648 30296 8660
rect 30136 8644 30296 8648
rect 29778 8610 30009 8616
rect 29778 8576 29959 8610
rect 29993 8576 30009 8610
rect 29778 8560 30009 8576
rect 30061 8610 30127 8616
rect 30061 8576 30077 8610
rect 30111 8576 30127 8610
rect 30061 8531 30127 8576
rect 29664 8523 30127 8531
rect 29664 8491 30128 8523
rect 30220 8507 30296 8644
rect 30216 8447 30226 8507
rect 30288 8447 30298 8507
rect 30039 7791 30175 7811
rect 26804 7740 26883 7752
rect 24325 7692 24404 7704
rect 24325 7595 24331 7692
rect 24255 7575 24331 7595
rect 24398 7595 24404 7692
rect 26804 7629 26810 7740
rect 26877 7629 26883 7740
rect 27952 7746 28031 7758
rect 27952 7629 27958 7746
rect 28025 7629 28031 7746
rect 30039 7729 30075 7791
rect 30135 7729 30175 7791
rect 30039 7701 30175 7729
rect 29735 7671 30712 7701
rect 24398 7575 24475 7595
rect 24255 7467 24299 7575
rect 24431 7467 24475 7575
rect 26052 7533 26108 7541
rect 24255 7425 24475 7467
rect 25126 7525 26108 7533
rect 25126 7491 26068 7525
rect 26102 7491 26108 7525
rect 26771 7521 26781 7629
rect 26913 7566 26923 7629
rect 26913 7555 26925 7566
rect 26913 7521 26926 7555
rect 27182 7545 27238 7547
rect 25126 7475 26108 7491
rect 26781 7483 26926 7521
rect 25126 7474 26105 7475
rect 23859 7395 24836 7425
rect 23859 7289 23891 7395
rect 24095 7289 24127 7395
rect 24331 7289 24363 7395
rect 24567 7289 24599 7395
rect 24802 7289 24836 7395
rect 23852 7277 23898 7289
rect 23852 7101 23858 7277
rect 23892 7101 23898 7277
rect 23852 7089 23898 7101
rect 23970 7277 24016 7289
rect 23970 7101 23976 7277
rect 24010 7101 24016 7277
rect 23970 7089 24016 7101
rect 24088 7277 24134 7289
rect 24088 7101 24094 7277
rect 24128 7101 24134 7277
rect 24088 7089 24134 7101
rect 24206 7277 24252 7289
rect 24206 7101 24212 7277
rect 24246 7101 24252 7277
rect 24206 7089 24252 7101
rect 24324 7277 24370 7289
rect 24324 7101 24330 7277
rect 24364 7101 24370 7277
rect 24324 7089 24370 7101
rect 24442 7277 24488 7289
rect 24442 7101 24448 7277
rect 24482 7101 24488 7277
rect 24442 7089 24488 7101
rect 24560 7277 24606 7289
rect 24560 7101 24566 7277
rect 24600 7101 24606 7277
rect 24560 7089 24606 7101
rect 24678 7277 24724 7289
rect 24678 7101 24684 7277
rect 24718 7101 24724 7277
rect 24678 7089 24724 7101
rect 24796 7277 24842 7289
rect 24796 7101 24802 7277
rect 24836 7101 24842 7277
rect 24796 7089 24842 7101
rect 24914 7277 24960 7289
rect 24914 7101 24920 7277
rect 24954 7101 24960 7277
rect 24914 7089 24960 7101
rect 23975 6995 24011 7089
rect 24211 6995 24247 7089
rect 24447 6996 24483 7089
rect 24609 7041 24675 7048
rect 24609 7007 24625 7041
rect 24659 7007 24675 7041
rect 24609 6996 24675 7007
rect 24447 6995 24675 6996
rect 23975 6966 24675 6995
rect 23975 6965 24557 6966
rect 22626 6795 22779 6933
rect 24095 6852 24129 6965
rect 24491 6924 24557 6965
rect 24491 6890 24507 6924
rect 24541 6890 24557 6924
rect 24491 6883 24557 6890
rect 24919 6884 24954 7089
rect 25126 6884 25193 7474
rect 26885 7451 26926 7483
rect 27172 7479 27182 7545
rect 27238 7479 27248 7545
rect 27918 7521 27928 7629
rect 28060 7566 28070 7629
rect 28060 7555 28072 7566
rect 29735 7565 29767 7671
rect 29971 7565 30003 7671
rect 30207 7565 30239 7671
rect 30443 7565 30475 7671
rect 30678 7565 30712 7671
rect 28060 7521 28073 7555
rect 27928 7483 28073 7521
rect 28032 7455 28073 7483
rect 26301 7423 26571 7451
rect 26042 7357 26052 7423
rect 26118 7357 26128 7423
rect 26301 7361 26335 7423
rect 26537 7361 26571 7423
rect 26655 7423 26926 7451
rect 27443 7427 27713 7455
rect 26655 7361 26689 7423
rect 26891 7361 26926 7423
rect 27067 7411 27238 7427
rect 27067 7377 27198 7411
rect 27232 7377 27238 7411
rect 27067 7361 27238 7377
rect 27443 7365 27477 7427
rect 27679 7365 27713 7427
rect 27797 7427 28073 7455
rect 27797 7365 27831 7427
rect 28033 7365 28073 7427
rect 29728 7553 29774 7565
rect 29728 7377 29734 7553
rect 29768 7377 29774 7553
rect 29728 7365 29774 7377
rect 29846 7553 29892 7565
rect 29846 7377 29852 7553
rect 29886 7377 29892 7553
rect 29846 7365 29892 7377
rect 29964 7553 30010 7565
rect 29964 7377 29970 7553
rect 30004 7377 30010 7553
rect 29964 7365 30010 7377
rect 30082 7553 30128 7565
rect 30082 7377 30088 7553
rect 30122 7377 30128 7553
rect 30082 7365 30128 7377
rect 30200 7553 30246 7565
rect 30200 7377 30206 7553
rect 30240 7377 30246 7553
rect 30200 7365 30246 7377
rect 30318 7553 30364 7565
rect 30318 7377 30324 7553
rect 30358 7377 30364 7553
rect 30318 7365 30364 7377
rect 30436 7553 30482 7565
rect 30436 7377 30442 7553
rect 30476 7377 30482 7553
rect 30436 7365 30482 7377
rect 30554 7553 30600 7565
rect 30554 7377 30560 7553
rect 30594 7377 30600 7553
rect 30554 7365 30600 7377
rect 30672 7553 30718 7565
rect 30672 7377 30678 7553
rect 30712 7377 30718 7553
rect 30672 7365 30718 7377
rect 30790 7553 30836 7565
rect 30790 7377 30796 7553
rect 30830 7377 30836 7553
rect 30790 7365 30836 7377
rect 26177 7349 26223 7361
rect 26177 6973 26183 7349
rect 26217 6973 26223 7349
rect 26177 6961 26223 6973
rect 26295 7349 26341 7361
rect 26295 6973 26301 7349
rect 26335 6973 26341 7349
rect 26295 6961 26341 6973
rect 26413 7349 26459 7361
rect 26413 6973 26419 7349
rect 26453 6973 26459 7349
rect 26413 6961 26459 6973
rect 26531 7349 26577 7361
rect 26531 6973 26537 7349
rect 26571 6973 26577 7349
rect 26531 6961 26577 6973
rect 26649 7349 26695 7361
rect 26649 6973 26655 7349
rect 26689 6973 26695 7349
rect 26649 6961 26695 6973
rect 26767 7349 26813 7361
rect 26767 6973 26773 7349
rect 26807 6973 26813 7349
rect 26767 6961 26813 6973
rect 26885 7349 26931 7361
rect 26885 6973 26891 7349
rect 26925 6973 26931 7349
rect 26885 6961 26931 6973
rect 24919 6856 25193 6884
rect 24565 6852 25193 6856
rect 21411 6727 21520 6781
rect 20731 6688 20958 6724
rect 20731 6581 20766 6688
rect 20892 6654 20958 6688
rect 20892 6620 20908 6654
rect 20942 6620 20958 6654
rect 21239 6712 21336 6727
rect 21239 6645 21296 6712
rect 20892 6614 20958 6620
rect 21133 6609 21402 6645
rect 21133 6581 21166 6609
rect 21369 6581 21402 6609
rect 21486 6581 21520 6727
rect 22337 6720 22347 6795
rect 22415 6720 22779 6795
rect 22364 6719 22779 6720
rect 24089 6840 24135 6852
rect 20607 6569 20653 6581
rect 20607 6393 20613 6569
rect 20647 6393 20653 6569
rect 20607 6381 20653 6393
rect 20725 6569 20771 6581
rect 20725 6393 20731 6569
rect 20765 6393 20771 6569
rect 20725 6381 20771 6393
rect 20843 6569 20889 6581
rect 20843 6393 20849 6569
rect 20883 6393 20889 6569
rect 20843 6381 20889 6393
rect 20961 6569 21007 6581
rect 20961 6393 20967 6569
rect 21001 6514 21007 6569
rect 21126 6569 21172 6581
rect 21126 6514 21132 6569
rect 21001 6426 21132 6514
rect 21001 6393 21007 6426
rect 20961 6381 21007 6393
rect 21126 6393 21132 6426
rect 21166 6393 21172 6569
rect 21126 6381 21172 6393
rect 21244 6569 21290 6581
rect 21244 6393 21250 6569
rect 21284 6393 21290 6569
rect 21244 6381 21290 6393
rect 21362 6569 21408 6581
rect 21362 6393 21368 6569
rect 21402 6393 21408 6569
rect 21362 6381 21408 6393
rect 21480 6569 21526 6581
rect 21480 6393 21486 6569
rect 21520 6393 21526 6569
rect 24089 6464 24095 6840
rect 24129 6464 24135 6840
rect 24089 6452 24135 6464
rect 24207 6840 24253 6852
rect 24207 6464 24213 6840
rect 24247 6464 24253 6840
rect 24207 6452 24253 6464
rect 24325 6840 24371 6852
rect 24325 6464 24331 6840
rect 24365 6488 24371 6840
rect 24442 6840 24488 6852
rect 24442 6664 24448 6840
rect 24482 6664 24488 6840
rect 24442 6652 24488 6664
rect 24560 6840 25193 6852
rect 24560 6664 24566 6840
rect 24600 6827 25193 6840
rect 26183 6919 26217 6961
rect 26419 6919 26453 6961
rect 26183 6891 26453 6919
rect 26537 6920 26571 6961
rect 26773 6920 26807 6961
rect 26537 6891 26807 6920
rect 26183 6843 26217 6891
rect 24600 6664 24606 6827
rect 26183 6813 26246 6843
rect 24560 6652 24606 6664
rect 26211 6721 26246 6813
rect 26211 6685 26438 6721
rect 26708 6710 26718 6807
rect 26817 6710 26827 6807
rect 26891 6778 26925 6961
rect 26891 6724 27000 6778
rect 24448 6536 24483 6652
rect 26211 6578 26246 6685
rect 26372 6651 26438 6685
rect 26372 6617 26388 6651
rect 26422 6617 26438 6651
rect 26719 6709 26816 6710
rect 26719 6642 26776 6709
rect 26372 6611 26438 6617
rect 26613 6606 26882 6642
rect 26613 6578 26646 6606
rect 26849 6578 26882 6606
rect 26966 6578 27000 6724
rect 26087 6566 26133 6578
rect 24579 6536 24687 6546
rect 24448 6488 24579 6536
rect 24687 6504 24832 6510
rect 24365 6464 24579 6488
rect 24325 6452 24579 6464
rect 24331 6448 24579 6452
rect 21480 6381 21526 6393
rect 22396 6447 23242 6448
rect 22396 6420 23967 6447
rect 22396 6414 24204 6420
rect 20613 6342 20647 6381
rect 20849 6342 20883 6381
rect 20613 6306 20883 6342
rect 21250 6343 21283 6381
rect 21486 6343 21519 6381
rect 21250 6307 21519 6343
rect 22396 6380 24154 6414
rect 24188 6380 24204 6414
rect 22396 6364 24204 6380
rect 24256 6414 24322 6420
rect 24256 6380 24272 6414
rect 24306 6380 24322 6414
rect 24505 6404 24579 6448
rect 24820 6437 24832 6504
rect 24687 6431 24832 6437
rect 24579 6394 24687 6404
rect 22396 6348 23967 6364
rect 22396 6347 23904 6348
rect 22396 6344 23439 6347
rect 20613 6305 20779 6306
rect 20647 6226 20779 6305
rect 20637 6118 20647 6226
rect 20779 6118 20789 6226
rect 20671 5990 20677 6118
rect 20744 5990 20750 6118
rect 20671 5978 20750 5990
rect 17251 5744 18228 5774
rect 20445 5772 20508 5789
rect 20370 5768 20508 5772
rect 17251 5638 17283 5744
rect 17487 5638 17519 5744
rect 17723 5638 17755 5744
rect 17959 5638 17991 5744
rect 18194 5638 18228 5744
rect 18538 5734 20508 5768
rect 18536 5705 20508 5734
rect 18536 5689 18582 5705
rect 20370 5703 20508 5705
rect 17244 5626 17290 5638
rect 17244 5450 17250 5626
rect 17284 5450 17290 5626
rect 17244 5438 17290 5450
rect 17362 5626 17408 5638
rect 17362 5450 17368 5626
rect 17402 5450 17408 5626
rect 17362 5438 17408 5450
rect 17480 5626 17526 5638
rect 17480 5450 17486 5626
rect 17520 5450 17526 5626
rect 17480 5438 17526 5450
rect 17598 5626 17644 5638
rect 17598 5450 17604 5626
rect 17638 5450 17644 5626
rect 17598 5438 17644 5450
rect 17716 5626 17762 5638
rect 17716 5450 17722 5626
rect 17756 5450 17762 5626
rect 17716 5438 17762 5450
rect 17834 5626 17880 5638
rect 17834 5450 17840 5626
rect 17874 5450 17880 5626
rect 17834 5438 17880 5450
rect 17952 5626 17998 5638
rect 17952 5450 17958 5626
rect 17992 5450 17998 5626
rect 17952 5438 17998 5450
rect 18070 5626 18116 5638
rect 18070 5450 18076 5626
rect 18110 5450 18116 5626
rect 18070 5438 18116 5450
rect 18188 5626 18234 5638
rect 18188 5450 18194 5626
rect 18228 5450 18234 5626
rect 18188 5438 18234 5450
rect 18306 5626 18352 5638
rect 18306 5450 18312 5626
rect 18346 5450 18352 5626
rect 18306 5438 18352 5450
rect 17367 5344 17403 5438
rect 17603 5344 17639 5438
rect 17839 5345 17875 5438
rect 18001 5390 18067 5397
rect 18001 5356 18017 5390
rect 18051 5356 18067 5390
rect 18001 5345 18067 5356
rect 17839 5344 18067 5345
rect 17367 5315 18067 5344
rect 17367 5314 17949 5315
rect 17487 5201 17521 5314
rect 17883 5273 17949 5314
rect 17883 5239 17899 5273
rect 17933 5239 17949 5273
rect 17883 5232 17949 5239
rect 18311 5220 18346 5438
rect 18535 5237 18582 5689
rect 21432 5699 21511 5711
rect 21432 5581 21438 5699
rect 21505 5581 21511 5699
rect 19494 5473 19504 5581
rect 19636 5473 19646 5581
rect 21392 5473 21402 5581
rect 21534 5473 21544 5581
rect 19504 5433 19636 5473
rect 21402 5433 21534 5473
rect 19503 5367 19636 5433
rect 21401 5367 21534 5433
rect 18832 5324 20305 5367
rect 18535 5221 18581 5237
rect 18500 5220 18581 5221
rect 18311 5205 18581 5220
rect 17957 5201 18581 5205
rect 17481 5189 17527 5201
rect 17216 4711 17226 4829
rect 17344 4797 17354 4829
rect 17481 4813 17487 5189
rect 17521 4813 17527 5189
rect 17481 4801 17527 4813
rect 17599 5189 17645 5201
rect 17599 4813 17605 5189
rect 17639 4813 17645 5189
rect 17599 4801 17645 4813
rect 17717 5189 17763 5201
rect 17717 4813 17723 5189
rect 17757 4837 17763 5189
rect 17834 5189 17880 5201
rect 17834 5013 17840 5189
rect 17874 5013 17880 5189
rect 17834 5001 17880 5013
rect 17952 5189 18581 5201
rect 17952 5013 17958 5189
rect 17992 5177 18581 5189
rect 17992 5176 18234 5177
rect 17992 5013 17998 5176
rect 18500 5175 18581 5177
rect 18832 5021 18866 5324
rect 19198 5221 19232 5324
rect 19434 5221 19468 5324
rect 19670 5221 19704 5324
rect 19906 5221 19940 5324
rect 19192 5209 19238 5221
rect 17952 5001 17998 5013
rect 18708 5009 18754 5021
rect 17840 4885 17875 5001
rect 17971 4885 18079 4895
rect 17840 4837 17971 4885
rect 18079 4848 18227 4854
rect 17757 4813 17971 4837
rect 17717 4801 17971 4813
rect 17723 4797 17971 4801
rect 17344 4769 17359 4797
rect 17344 4763 17596 4769
rect 17344 4729 17546 4763
rect 17580 4729 17596 4763
rect 17344 4713 17596 4729
rect 17648 4763 17714 4769
rect 17648 4729 17664 4763
rect 17698 4729 17714 4763
rect 17897 4753 17971 4797
rect 18215 4781 18227 4848
rect 18708 4833 18714 5009
rect 18748 4833 18754 5009
rect 18708 4821 18754 4833
rect 18826 5009 18872 5021
rect 18826 4833 18832 5009
rect 18866 4833 18872 5009
rect 18826 4821 18872 4833
rect 18944 5009 18990 5021
rect 18944 4833 18950 5009
rect 18984 4833 18990 5009
rect 18944 4821 18990 4833
rect 19062 5009 19108 5021
rect 19192 5009 19198 5209
rect 19062 4833 19068 5009
rect 19102 4833 19198 5009
rect 19232 4833 19238 5209
rect 19062 4821 19108 4833
rect 19192 4821 19238 4833
rect 19310 5209 19356 5221
rect 19310 4833 19316 5209
rect 19350 4833 19356 5209
rect 19310 4821 19356 4833
rect 19428 5209 19474 5221
rect 19428 4833 19434 5209
rect 19468 4833 19474 5209
rect 19428 4821 19474 4833
rect 19546 5209 19592 5221
rect 19546 4833 19552 5209
rect 19586 4833 19592 5209
rect 19546 4821 19592 4833
rect 19664 5209 19710 5221
rect 19664 4833 19670 5209
rect 19704 4833 19710 5209
rect 19664 4821 19710 4833
rect 19782 5209 19828 5221
rect 19782 4833 19788 5209
rect 19822 4833 19828 5209
rect 19782 4821 19828 4833
rect 19900 5209 19946 5221
rect 19900 4833 19906 5209
rect 19940 5009 19946 5209
rect 20271 5021 20305 5324
rect 20730 5324 22203 5367
rect 20730 5021 20764 5324
rect 21096 5221 21130 5324
rect 21332 5221 21366 5324
rect 21568 5221 21602 5324
rect 21804 5221 21838 5324
rect 21090 5209 21136 5221
rect 20029 5009 20075 5021
rect 19940 4833 20035 5009
rect 20069 4833 20075 5009
rect 19900 4821 19946 4833
rect 20029 4821 20075 4833
rect 20147 5009 20193 5021
rect 20147 4833 20153 5009
rect 20187 4833 20193 5009
rect 20147 4821 20193 4833
rect 20265 5009 20311 5021
rect 20265 4833 20271 5009
rect 20305 4833 20311 5009
rect 20265 4821 20311 4833
rect 20383 5009 20429 5021
rect 20383 4833 20389 5009
rect 20423 4833 20429 5009
rect 20383 4821 20429 4833
rect 20606 5009 20652 5021
rect 20606 4833 20612 5009
rect 20646 4833 20652 5009
rect 20606 4821 20652 4833
rect 20724 5009 20770 5021
rect 20724 4833 20730 5009
rect 20764 4833 20770 5009
rect 20724 4821 20770 4833
rect 20842 5009 20888 5021
rect 20842 4833 20848 5009
rect 20882 4833 20888 5009
rect 20842 4821 20888 4833
rect 20960 5009 21006 5021
rect 21090 5009 21096 5209
rect 20960 4833 20966 5009
rect 21000 4833 21096 5009
rect 21130 4833 21136 5209
rect 20960 4821 21006 4833
rect 21090 4821 21136 4833
rect 21208 5209 21254 5221
rect 21208 4833 21214 5209
rect 21248 4833 21254 5209
rect 21208 4821 21254 4833
rect 21326 5209 21372 5221
rect 21326 4833 21332 5209
rect 21366 4833 21372 5209
rect 21326 4821 21372 4833
rect 21444 5209 21490 5221
rect 21444 4833 21450 5209
rect 21484 4833 21490 5209
rect 21444 4821 21490 4833
rect 21562 5209 21608 5221
rect 21562 4833 21568 5209
rect 21602 4833 21608 5209
rect 21562 4821 21608 4833
rect 21680 5209 21726 5221
rect 21680 4833 21686 5209
rect 21720 4833 21726 5209
rect 21680 4821 21726 4833
rect 21798 5209 21844 5221
rect 21798 4833 21804 5209
rect 21838 5009 21844 5209
rect 22169 5021 22203 5324
rect 21927 5009 21973 5021
rect 21838 4833 21933 5009
rect 21967 4833 21973 5009
rect 21798 4821 21844 4833
rect 21927 4821 21973 4833
rect 22045 5009 22091 5021
rect 22045 4833 22051 5009
rect 22085 4833 22091 5009
rect 22045 4821 22091 4833
rect 22163 5009 22209 5021
rect 22163 4833 22169 5009
rect 22203 4833 22209 5009
rect 22163 4821 22209 4833
rect 22281 5009 22327 5021
rect 22281 4833 22287 5009
rect 22321 4833 22327 5009
rect 22281 4821 22327 4833
rect 18079 4775 18227 4781
rect 18714 4787 18748 4821
rect 19316 4787 19350 4821
rect 19552 4787 19586 4821
rect 17971 4743 18079 4753
rect 18714 4752 18873 4787
rect 19316 4752 19586 4787
rect 20153 4787 20187 4821
rect 20389 4787 20423 4821
rect 20153 4752 20423 4787
rect 20612 4787 20646 4821
rect 21214 4787 21248 4821
rect 21450 4787 21484 4821
rect 20612 4752 20771 4787
rect 21214 4752 21484 4787
rect 22051 4787 22085 4821
rect 22287 4787 22321 4821
rect 22051 4752 22321 4787
rect 17344 4711 17359 4713
rect 17259 4697 17359 4711
rect 17259 4654 17359 4655
rect 16880 4633 17359 4654
rect 17648 4633 17714 4729
rect 16880 4585 17714 4633
rect 16880 4556 17359 4585
rect 16880 4554 16985 4556
rect 17259 4555 17359 4556
rect 16713 4369 16723 4448
rect 16816 4369 16826 4448
rect 17716 4433 17795 4445
rect 16724 3195 16817 4369
rect 17716 4340 17722 4433
rect 17642 4320 17722 4340
rect 17789 4340 17795 4433
rect 17789 4320 17862 4340
rect 17642 4212 17686 4320
rect 17818 4212 17862 4320
rect 17642 4170 17862 4212
rect 17246 4140 18223 4170
rect 17246 4034 17278 4140
rect 17482 4034 17514 4140
rect 17718 4034 17750 4140
rect 17954 4034 17986 4140
rect 18189 4034 18223 4140
rect 17239 4022 17285 4034
rect 17239 3846 17245 4022
rect 17279 3846 17285 4022
rect 17239 3834 17285 3846
rect 17357 4022 17403 4034
rect 17357 3846 17363 4022
rect 17397 3846 17403 4022
rect 17357 3834 17403 3846
rect 17475 4022 17521 4034
rect 17475 3846 17481 4022
rect 17515 3846 17521 4022
rect 17475 3834 17521 3846
rect 17593 4022 17639 4034
rect 17593 3846 17599 4022
rect 17633 3846 17639 4022
rect 17593 3834 17639 3846
rect 17711 4022 17757 4034
rect 17711 3846 17717 4022
rect 17751 3846 17757 4022
rect 17711 3834 17757 3846
rect 17829 4022 17875 4034
rect 17829 3846 17835 4022
rect 17869 3846 17875 4022
rect 17829 3834 17875 3846
rect 17947 4022 17993 4034
rect 17947 3846 17953 4022
rect 17987 3846 17993 4022
rect 17947 3834 17993 3846
rect 18065 4022 18111 4034
rect 18065 3846 18071 4022
rect 18105 3846 18111 4022
rect 18065 3834 18111 3846
rect 18183 4022 18229 4034
rect 18183 3846 18189 4022
rect 18223 3846 18229 4022
rect 18183 3834 18229 3846
rect 18301 4022 18347 4034
rect 18301 3846 18307 4022
rect 18341 3846 18347 4022
rect 18301 3834 18347 3846
rect 18839 3968 18873 4752
rect 19552 4690 19586 4752
rect 19141 4652 19883 4690
rect 19141 4528 19175 4652
rect 19377 4528 19411 4652
rect 19613 4528 19647 4652
rect 19849 4528 19883 4652
rect 20139 4545 20149 4611
rect 20212 4545 20222 4611
rect 19135 4516 19181 4528
rect 19135 4140 19141 4516
rect 19175 4140 19181 4516
rect 19135 4128 19181 4140
rect 19253 4516 19299 4528
rect 19253 4140 19259 4516
rect 19293 4140 19299 4516
rect 19253 4128 19299 4140
rect 19371 4516 19417 4528
rect 19371 4140 19377 4516
rect 19411 4140 19417 4516
rect 19371 4128 19417 4140
rect 19489 4516 19535 4528
rect 19489 4140 19495 4516
rect 19529 4140 19535 4516
rect 19489 4128 19535 4140
rect 19607 4516 19653 4528
rect 19607 4140 19613 4516
rect 19647 4140 19653 4516
rect 19607 4128 19653 4140
rect 19725 4516 19771 4528
rect 19725 4140 19731 4516
rect 19765 4140 19771 4516
rect 19725 4128 19771 4140
rect 19843 4516 19889 4528
rect 19843 4140 19849 4516
rect 19883 4140 19889 4516
rect 19843 4128 19889 4140
rect 20255 3969 20289 4752
rect 19982 3968 20289 3969
rect 18839 3963 19155 3968
rect 19869 3963 20289 3968
rect 18839 3952 19222 3963
rect 18839 3925 19171 3952
rect 17362 3740 17398 3834
rect 17598 3740 17634 3834
rect 17834 3741 17870 3834
rect 17996 3786 18062 3793
rect 17996 3752 18012 3786
rect 18046 3752 18062 3786
rect 17996 3741 18062 3752
rect 17834 3740 18062 3741
rect 17362 3711 18062 3740
rect 17362 3710 17944 3711
rect 17482 3597 17516 3710
rect 17878 3669 17944 3710
rect 17878 3635 17894 3669
rect 17928 3635 17944 3669
rect 17878 3628 17944 3635
rect 18306 3601 18341 3834
rect 18839 3796 18873 3925
rect 19155 3918 19171 3925
rect 19205 3918 19222 3952
rect 19155 3912 19222 3918
rect 19802 3952 20289 3963
rect 19802 3918 19819 3952
rect 19853 3925 20289 3952
rect 19853 3918 19869 3925
rect 19982 3924 20289 3925
rect 19802 3912 19869 3918
rect 18980 3885 19036 3897
rect 18980 3851 18986 3885
rect 19020 3884 19036 3885
rect 20093 3884 20149 3896
rect 19020 3868 19487 3884
rect 19020 3851 19437 3868
rect 18980 3835 19437 3851
rect 19421 3834 19437 3835
rect 19471 3834 19487 3868
rect 19421 3827 19487 3834
rect 19539 3869 20109 3884
rect 19539 3835 19555 3869
rect 19589 3850 20109 3869
rect 20143 3850 20149 3884
rect 19589 3835 20149 3850
rect 19539 3825 19606 3835
rect 20093 3834 20149 3835
rect 20255 3796 20289 3924
rect 20737 3968 20771 4752
rect 21450 4690 21484 4752
rect 21039 4652 21781 4690
rect 21039 4528 21073 4652
rect 21275 4528 21309 4652
rect 21511 4528 21545 4652
rect 21747 4528 21781 4652
rect 21033 4516 21079 4528
rect 21033 4140 21039 4516
rect 21073 4140 21079 4516
rect 21033 4128 21079 4140
rect 21151 4516 21197 4528
rect 21151 4140 21157 4516
rect 21191 4140 21197 4516
rect 21151 4128 21197 4140
rect 21269 4516 21315 4528
rect 21269 4140 21275 4516
rect 21309 4140 21315 4516
rect 21269 4128 21315 4140
rect 21387 4516 21433 4528
rect 21387 4140 21393 4516
rect 21427 4140 21433 4516
rect 21387 4128 21433 4140
rect 21505 4516 21551 4528
rect 21505 4140 21511 4516
rect 21545 4140 21551 4516
rect 21505 4128 21551 4140
rect 21623 4516 21669 4528
rect 21623 4140 21629 4516
rect 21663 4140 21669 4516
rect 21623 4128 21669 4140
rect 21741 4516 21787 4528
rect 21741 4140 21747 4516
rect 21781 4140 21787 4516
rect 21741 4128 21787 4140
rect 22153 3969 22187 4752
rect 21765 3968 21834 3969
rect 21880 3968 22187 3969
rect 20737 3963 21053 3968
rect 21765 3964 22187 3968
rect 20737 3952 21120 3963
rect 20737 3925 21069 3952
rect 20737 3796 20771 3925
rect 21053 3918 21069 3925
rect 21103 3918 21120 3952
rect 21053 3912 21120 3918
rect 21698 3953 22187 3964
rect 21698 3919 21715 3953
rect 21749 3925 22187 3953
rect 21749 3919 21765 3925
rect 21880 3924 22187 3925
rect 21698 3913 21765 3919
rect 20878 3885 20934 3897
rect 20878 3851 20884 3885
rect 20918 3884 20934 3885
rect 21991 3884 22047 3896
rect 20918 3868 21385 3884
rect 20918 3851 21335 3868
rect 20878 3835 21335 3851
rect 21319 3834 21335 3835
rect 21369 3834 21385 3868
rect 21319 3827 21385 3834
rect 21437 3869 22007 3884
rect 21437 3835 21453 3869
rect 21487 3850 22007 3869
rect 22041 3850 22047 3884
rect 21487 3835 22047 3850
rect 21437 3825 21504 3835
rect 21991 3834 22047 3835
rect 22153 3796 22187 3924
rect 22268 4574 22335 4598
rect 22268 4540 22285 4574
rect 22319 4540 22335 4574
rect 17952 3597 18341 3601
rect 17476 3585 17522 3597
rect 17476 3209 17482 3585
rect 17516 3209 17522 3585
rect 17476 3197 17522 3209
rect 17594 3585 17640 3597
rect 17594 3209 17600 3585
rect 17634 3209 17640 3585
rect 17594 3197 17640 3209
rect 17712 3585 17758 3597
rect 17712 3209 17718 3585
rect 17752 3233 17758 3585
rect 17829 3585 17875 3597
rect 17829 3409 17835 3585
rect 17869 3409 17875 3585
rect 17829 3397 17875 3409
rect 17947 3585 18341 3597
rect 18833 3784 18879 3796
rect 18833 3608 18839 3784
rect 18873 3608 18879 3784
rect 18833 3596 18879 3608
rect 18951 3784 18997 3796
rect 18951 3608 18957 3784
rect 18991 3608 18997 3784
rect 18951 3596 18997 3608
rect 19253 3784 19299 3796
rect 17947 3409 17953 3585
rect 17987 3572 18341 3585
rect 17987 3409 17993 3572
rect 18263 3569 18341 3572
rect 18263 3517 18273 3569
rect 18336 3517 18346 3569
rect 18268 3511 18341 3517
rect 17947 3397 17993 3409
rect 17835 3281 17870 3397
rect 18956 3302 18990 3596
rect 19253 3408 19259 3784
rect 19293 3408 19299 3784
rect 19253 3396 19299 3408
rect 19371 3784 19417 3796
rect 19371 3408 19377 3784
rect 19411 3408 19417 3784
rect 19371 3396 19417 3408
rect 19489 3784 19535 3796
rect 19489 3408 19495 3784
rect 19529 3408 19535 3784
rect 19489 3396 19535 3408
rect 19607 3784 19653 3796
rect 19607 3408 19613 3784
rect 19647 3408 19653 3784
rect 19607 3396 19653 3408
rect 19725 3784 19771 3796
rect 19725 3408 19731 3784
rect 19765 3408 19771 3784
rect 20131 3784 20177 3796
rect 20131 3608 20137 3784
rect 20171 3608 20177 3784
rect 20131 3596 20177 3608
rect 20249 3784 20295 3796
rect 20249 3608 20255 3784
rect 20289 3608 20295 3784
rect 20249 3596 20295 3608
rect 20731 3784 20777 3796
rect 20731 3608 20737 3784
rect 20771 3608 20777 3784
rect 20731 3596 20777 3608
rect 20849 3784 20895 3796
rect 20849 3608 20855 3784
rect 20889 3608 20895 3784
rect 20849 3596 20895 3608
rect 21151 3784 21197 3796
rect 19725 3396 19771 3408
rect 19613 3302 19647 3396
rect 20137 3302 20170 3596
rect 17966 3281 18074 3291
rect 17835 3233 17966 3281
rect 18956 3270 20170 3302
rect 20854 3302 20888 3596
rect 21151 3408 21157 3784
rect 21191 3408 21197 3784
rect 21151 3396 21197 3408
rect 21269 3784 21315 3796
rect 21269 3408 21275 3784
rect 21309 3408 21315 3784
rect 21269 3396 21315 3408
rect 21387 3784 21433 3796
rect 21387 3408 21393 3784
rect 21427 3408 21433 3784
rect 21387 3396 21433 3408
rect 21505 3784 21551 3796
rect 21505 3408 21511 3784
rect 21545 3408 21551 3784
rect 21505 3396 21551 3408
rect 21623 3784 21669 3796
rect 21623 3408 21629 3784
rect 21663 3408 21669 3784
rect 22029 3784 22075 3796
rect 22029 3608 22035 3784
rect 22069 3608 22075 3784
rect 22029 3596 22075 3608
rect 22147 3784 22193 3796
rect 22147 3608 22153 3784
rect 22187 3608 22193 3784
rect 22147 3596 22193 3608
rect 21623 3396 21669 3408
rect 21511 3302 21545 3396
rect 22035 3302 22068 3596
rect 20854 3270 22068 3302
rect 18074 3239 18230 3245
rect 17752 3209 17966 3233
rect 17712 3197 17966 3209
rect 16724 3193 17309 3195
rect 17718 3193 17966 3197
rect 16724 3165 17354 3193
rect 16724 3159 17591 3165
rect 16724 3125 17541 3159
rect 17575 3125 17591 3159
rect 16724 3109 17591 3125
rect 17643 3159 17709 3165
rect 17643 3125 17659 3159
rect 17693 3125 17709 3159
rect 17892 3149 17966 3193
rect 18218 3172 18230 3239
rect 19449 3185 19581 3270
rect 21347 3185 21479 3270
rect 18074 3166 18230 3172
rect 17966 3139 18074 3149
rect 16724 3093 17354 3109
rect 16724 3089 17309 3093
rect 16724 3088 16825 3089
rect 17254 3040 17354 3051
rect 16384 3002 16552 3021
rect 16384 2915 16411 3002
rect 16513 2915 16552 3002
rect 17218 2934 17228 3040
rect 17340 3029 17354 3040
rect 17643 3029 17709 3125
rect 19439 3077 19449 3185
rect 19581 3077 19591 3185
rect 21337 3077 21347 3185
rect 21479 3077 21489 3185
rect 22268 3157 22335 4540
rect 22396 4111 22552 6344
rect 23237 6343 23439 6344
rect 22396 4013 22408 4111
rect 22540 4013 22552 4111
rect 22396 4007 22552 4013
rect 22679 5932 23223 5959
rect 22679 5826 23071 5932
rect 23183 5919 23223 5932
rect 23183 5826 23225 5919
rect 22679 5815 23225 5826
rect 22679 5814 23223 5815
rect 17340 2981 17709 3029
rect 17340 2951 17354 2981
rect 17340 2934 17350 2951
rect 16384 2909 16552 2915
rect 17642 2878 17708 2981
rect 19465 2937 19471 3077
rect 19538 2937 19544 3077
rect 19465 2925 19544 2937
rect 22268 2878 22334 3157
rect 17640 2798 22334 2878
rect 21051 2287 21515 2319
rect 21603 2303 21613 2363
rect 21675 2303 21685 2363
rect 21051 2279 21514 2287
rect 21051 2131 21105 2279
rect 15393 1799 16156 1879
rect 15143 1786 16156 1799
rect 15103 1774 16156 1786
rect 14638 1661 14672 1774
rect 15108 1770 16156 1774
rect 15458 1769 16156 1770
rect 20740 2030 21105 2131
rect 21165 2234 21396 2250
rect 21165 2200 21346 2234
rect 21380 2200 21396 2234
rect 21165 2194 21396 2200
rect 21448 2234 21514 2279
rect 21448 2200 21464 2234
rect 21498 2200 21514 2234
rect 21448 2194 21514 2200
rect 15034 1736 15100 1743
rect 15034 1702 15050 1736
rect 15084 1702 15100 1736
rect 15034 1661 15100 1702
rect 14518 1660 15100 1661
rect 14518 1631 15218 1660
rect 14518 1537 14554 1631
rect 14754 1537 14790 1631
rect 14990 1630 15218 1631
rect 14990 1537 15026 1630
rect 15152 1619 15218 1630
rect 15152 1585 15168 1619
rect 15202 1585 15218 1619
rect 15152 1578 15218 1585
rect 15462 1537 15497 1769
rect 14395 1525 14441 1537
rect 14395 1349 14401 1525
rect 14435 1349 14441 1525
rect 14395 1337 14441 1349
rect 14513 1525 14559 1537
rect 14513 1349 14519 1525
rect 14553 1349 14559 1525
rect 14513 1337 14559 1349
rect 14631 1525 14677 1537
rect 14631 1349 14637 1525
rect 14671 1349 14677 1525
rect 14631 1337 14677 1349
rect 14749 1525 14795 1537
rect 14749 1349 14755 1525
rect 14789 1349 14795 1525
rect 14749 1337 14795 1349
rect 14867 1525 14913 1537
rect 14867 1349 14873 1525
rect 14907 1349 14913 1525
rect 14867 1337 14913 1349
rect 14985 1525 15031 1537
rect 14985 1349 14991 1525
rect 15025 1349 15031 1525
rect 14985 1337 15031 1349
rect 15103 1525 15149 1537
rect 15103 1349 15109 1525
rect 15143 1349 15149 1525
rect 15103 1337 15149 1349
rect 15221 1525 15267 1537
rect 15221 1349 15227 1525
rect 15261 1349 15267 1525
rect 15221 1337 15267 1349
rect 15339 1525 15385 1537
rect 15339 1349 15345 1525
rect 15379 1349 15385 1525
rect 15339 1337 15385 1349
rect 15457 1525 15503 1537
rect 15457 1349 15463 1525
rect 15497 1349 15503 1525
rect 15457 1337 15503 1349
rect 14402 1231 14434 1337
rect 14638 1231 14670 1337
rect 14874 1231 14906 1337
rect 15110 1231 15142 1337
rect 15345 1231 15379 1337
rect 14402 1201 15379 1231
rect 14706 1173 14842 1201
rect 14706 1111 14742 1173
rect 14802 1111 14842 1173
rect 14706 1091 14842 1111
rect 20740 1001 20826 2030
rect 21165 2002 21219 2194
rect 21607 2166 21683 2303
rect 21523 2162 21683 2166
rect 20894 1995 21219 2002
rect 20889 1906 20899 1995
rect 20968 1906 21219 1995
rect 20894 1902 21219 1906
rect 21281 2150 21327 2162
rect 21281 1774 21287 2150
rect 21321 1774 21327 2150
rect 21281 1762 21327 1774
rect 21399 2150 21445 2162
rect 21399 1774 21405 2150
rect 21439 1774 21445 2150
rect 21399 1762 21445 1774
rect 21517 2150 21683 2162
rect 21517 1774 21523 2150
rect 21557 2123 21683 2150
rect 21557 1774 21563 2123
rect 21640 1962 21683 2123
rect 21517 1762 21563 1774
rect 21634 1957 21683 1962
rect 21634 1950 21680 1957
rect 21634 1774 21640 1950
rect 21674 1774 21680 1950
rect 21634 1762 21680 1774
rect 21752 1950 21798 1962
rect 21752 1774 21758 1950
rect 21792 1787 21798 1950
rect 22679 1867 22835 5814
rect 22935 4820 23222 4849
rect 22935 4714 23070 4820
rect 23182 4818 23222 4820
rect 23188 4807 23222 4818
rect 22935 4712 23076 4714
rect 23188 4712 23223 4807
rect 22935 4703 23223 4712
rect 22935 4702 23222 4703
rect 22935 4701 23190 4702
rect 22938 2364 23090 4701
rect 23346 4449 23439 6343
rect 23502 6284 23968 6306
rect 24256 6284 24322 6380
rect 26087 6390 26093 6566
rect 26127 6390 26133 6566
rect 26087 6378 26133 6390
rect 26205 6566 26251 6578
rect 26205 6390 26211 6566
rect 26245 6390 26251 6566
rect 26205 6378 26251 6390
rect 26323 6566 26369 6578
rect 26323 6390 26329 6566
rect 26363 6390 26369 6566
rect 26323 6378 26369 6390
rect 26441 6566 26487 6578
rect 26441 6390 26447 6566
rect 26481 6511 26487 6566
rect 26606 6566 26652 6578
rect 26606 6511 26612 6566
rect 26481 6423 26612 6511
rect 26481 6390 26487 6423
rect 26441 6378 26487 6390
rect 26606 6390 26612 6423
rect 26646 6390 26652 6566
rect 26606 6378 26652 6390
rect 26724 6566 26770 6578
rect 26724 6390 26730 6566
rect 26764 6390 26770 6566
rect 26724 6378 26770 6390
rect 26842 6566 26888 6578
rect 26842 6390 26848 6566
rect 26882 6390 26888 6566
rect 26842 6378 26888 6390
rect 26960 6566 27006 6578
rect 26960 6390 26966 6566
rect 27000 6390 27006 6566
rect 26960 6378 27006 6390
rect 26093 6339 26127 6378
rect 26329 6339 26363 6378
rect 26093 6304 26363 6339
rect 26730 6340 26763 6378
rect 26966 6340 26999 6378
rect 26730 6304 26999 6340
rect 23502 6236 24322 6284
rect 26127 6303 26363 6304
rect 23502 6205 23968 6236
rect 26127 6229 26259 6303
rect 23502 5949 23607 6205
rect 26117 6121 26127 6229
rect 26259 6121 26269 6229
rect 24340 6042 24419 6054
rect 23502 5843 23565 5949
rect 23677 5843 23687 5949
rect 24340 5945 24346 6042
rect 24269 5925 24346 5945
rect 24413 5945 24419 6042
rect 26156 5991 26162 6121
rect 26229 5991 26235 6121
rect 26156 5979 26235 5991
rect 24413 5925 24489 5945
rect 23502 5832 23651 5843
rect 23502 4655 23607 5832
rect 24269 5817 24313 5925
rect 24445 5817 24489 5925
rect 24269 5775 24489 5817
rect 27067 5790 27129 7361
rect 27319 7353 27365 7365
rect 27319 6977 27325 7353
rect 27359 6977 27365 7353
rect 27319 6965 27365 6977
rect 27437 7353 27483 7365
rect 27437 6977 27443 7353
rect 27477 6977 27483 7353
rect 27437 6965 27483 6977
rect 27555 7353 27601 7365
rect 27555 6977 27561 7353
rect 27595 6977 27601 7353
rect 27555 6965 27601 6977
rect 27673 7353 27719 7365
rect 27673 6977 27679 7353
rect 27713 6977 27719 7353
rect 27673 6965 27719 6977
rect 27791 7353 27837 7365
rect 27791 6977 27797 7353
rect 27831 6977 27837 7353
rect 27791 6965 27837 6977
rect 27909 7353 27955 7365
rect 27909 6977 27915 7353
rect 27949 6977 27955 7353
rect 27909 6965 27955 6977
rect 28027 7353 28073 7365
rect 28027 6977 28033 7353
rect 28067 6977 28073 7353
rect 29851 7271 29887 7365
rect 30087 7271 30123 7365
rect 30323 7272 30359 7365
rect 30485 7317 30551 7324
rect 30485 7283 30501 7317
rect 30535 7283 30551 7317
rect 30485 7272 30551 7283
rect 30323 7271 30551 7272
rect 29851 7242 30551 7271
rect 29851 7241 30433 7242
rect 29971 7128 30005 7241
rect 30367 7200 30433 7241
rect 30367 7166 30383 7200
rect 30417 7166 30433 7200
rect 30367 7159 30433 7166
rect 30795 7132 30830 7365
rect 30441 7131 30830 7132
rect 31027 7131 31118 10050
rect 31603 9540 31637 10324
rect 32316 10262 32350 10324
rect 31905 10224 32647 10262
rect 31715 10053 31725 10121
rect 31780 10053 31790 10121
rect 31905 10100 31939 10224
rect 32141 10100 32175 10224
rect 32377 10100 32411 10224
rect 32613 10100 32647 10224
rect 31899 10088 31945 10100
rect 31899 9712 31905 10088
rect 31939 9712 31945 10088
rect 31899 9700 31945 9712
rect 32017 10088 32063 10100
rect 32017 9712 32023 10088
rect 32057 9712 32063 10088
rect 32017 9700 32063 9712
rect 32135 10088 32181 10100
rect 32135 9712 32141 10088
rect 32175 9712 32181 10088
rect 32135 9700 32181 9712
rect 32253 10088 32299 10100
rect 32253 9712 32259 10088
rect 32293 9712 32299 10088
rect 32253 9700 32299 9712
rect 32371 10088 32417 10100
rect 32371 9712 32377 10088
rect 32411 9712 32417 10088
rect 32371 9700 32417 9712
rect 32489 10088 32535 10100
rect 32489 9712 32495 10088
rect 32529 9712 32535 10088
rect 32489 9700 32535 9712
rect 32607 10088 32653 10100
rect 32607 9712 32613 10088
rect 32647 9712 32653 10088
rect 32773 9883 32847 9895
rect 32769 9792 32779 9883
rect 32841 9792 32851 9883
rect 32773 9780 32847 9792
rect 32607 9700 32653 9712
rect 33019 9541 33053 10324
rect 33388 10296 33424 10390
rect 33624 10296 33660 10390
rect 33860 10297 33896 10390
rect 34022 10342 34088 10349
rect 34022 10308 34038 10342
rect 34072 10308 34088 10342
rect 34022 10297 34088 10308
rect 33860 10296 34088 10297
rect 33388 10267 34088 10296
rect 33388 10266 33970 10267
rect 33114 10234 33190 10239
rect 33111 10178 33121 10234
rect 33174 10233 33190 10234
rect 33174 10178 33440 10233
rect 33114 10173 33440 10178
rect 33235 10131 33326 10136
rect 33235 10042 33245 10131
rect 33318 10042 33326 10131
rect 33235 10030 33326 10042
rect 33272 9636 33326 10030
rect 33386 9721 33440 10173
rect 33508 10153 33542 10266
rect 33904 10225 33970 10266
rect 33904 10191 33920 10225
rect 33954 10191 33970 10225
rect 33904 10184 33970 10191
rect 34332 10157 34367 10390
rect 33978 10153 34367 10157
rect 33502 10141 33548 10153
rect 33502 9765 33508 10141
rect 33542 9765 33548 10141
rect 33502 9753 33548 9765
rect 33620 10141 33666 10153
rect 33620 9765 33626 10141
rect 33660 9765 33666 10141
rect 33620 9753 33666 9765
rect 33738 10141 33784 10153
rect 33738 9765 33744 10141
rect 33778 9792 33784 10141
rect 33855 10141 33901 10153
rect 33855 9965 33861 10141
rect 33895 9965 33901 10141
rect 33855 9958 33901 9965
rect 33973 10141 34367 10153
rect 33973 9965 33979 10141
rect 34013 10131 34367 10141
rect 34013 10128 34226 10131
rect 34013 9965 34019 10128
rect 34192 10060 34226 10128
rect 34353 10060 34367 10131
rect 34655 10089 34737 15590
rect 34192 10039 34367 10060
rect 33855 9953 33904 9958
rect 33973 9953 34019 9965
rect 33861 9792 33904 9953
rect 33778 9765 33904 9792
rect 33738 9753 33904 9765
rect 33744 9749 33904 9753
rect 33386 9715 33617 9721
rect 33386 9681 33567 9715
rect 33601 9681 33617 9715
rect 33386 9665 33617 9681
rect 33669 9715 33735 9721
rect 33669 9681 33685 9715
rect 33719 9681 33735 9715
rect 33669 9636 33735 9681
rect 33272 9628 33735 9636
rect 33272 9596 33736 9628
rect 33828 9612 33904 9749
rect 33824 9552 33834 9612
rect 33896 9552 33906 9612
rect 32746 9540 33053 9541
rect 31603 9535 31919 9540
rect 32633 9535 33053 9540
rect 31603 9524 31986 9535
rect 31603 9497 31935 9524
rect 31603 9368 31637 9497
rect 31919 9490 31935 9497
rect 31969 9490 31986 9524
rect 31919 9484 31986 9490
rect 32566 9524 33053 9535
rect 33832 9526 33902 9552
rect 32566 9490 32583 9524
rect 32617 9497 33053 9524
rect 32617 9490 32633 9497
rect 32746 9496 33053 9497
rect 32566 9484 32633 9490
rect 31744 9457 31800 9469
rect 31744 9423 31750 9457
rect 31784 9456 31800 9457
rect 32857 9456 32913 9468
rect 31784 9440 32251 9456
rect 31784 9423 32201 9440
rect 31744 9407 32201 9423
rect 32185 9406 32201 9407
rect 32235 9406 32251 9440
rect 32185 9399 32251 9406
rect 32303 9441 32873 9456
rect 32303 9407 32319 9441
rect 32353 9422 32873 9441
rect 32907 9422 32913 9456
rect 32353 9407 32913 9422
rect 32303 9397 32370 9407
rect 32857 9406 32913 9407
rect 33019 9368 33053 9496
rect 31597 9356 31643 9368
rect 31597 9180 31603 9356
rect 31637 9180 31643 9356
rect 31597 9168 31643 9180
rect 31715 9356 31761 9368
rect 31715 9180 31721 9356
rect 31755 9180 31761 9356
rect 31715 9168 31761 9180
rect 32017 9356 32063 9368
rect 31720 8874 31754 9168
rect 32017 8980 32023 9356
rect 32057 8980 32063 9356
rect 32017 8968 32063 8980
rect 32135 9356 32181 9368
rect 32135 8980 32141 9356
rect 32175 8980 32181 9356
rect 32135 8968 32181 8980
rect 32253 9356 32299 9368
rect 32253 8980 32259 9356
rect 32293 8980 32299 9356
rect 32253 8968 32299 8980
rect 32371 9356 32417 9368
rect 32371 8980 32377 9356
rect 32411 8980 32417 9356
rect 32371 8968 32417 8980
rect 32489 9356 32535 9368
rect 32489 8980 32495 9356
rect 32529 8980 32535 9356
rect 32895 9356 32941 9368
rect 32895 9180 32901 9356
rect 32935 9180 32941 9356
rect 32895 9168 32941 9180
rect 33013 9356 33059 9368
rect 33013 9180 33019 9356
rect 33053 9180 33059 9356
rect 33013 9168 33059 9180
rect 32489 8968 32535 8980
rect 32377 8874 32411 8968
rect 32901 8874 32934 9168
rect 31720 8842 32934 8874
rect 32086 8818 32492 8842
rect 32086 8695 32198 8818
rect 32372 8695 32492 8818
rect 32086 8651 32492 8695
rect 32100 7824 32545 7830
rect 32100 7624 32112 7824
rect 32533 7624 32545 7824
rect 32100 7618 32268 7624
rect 32258 7550 32268 7618
rect 32400 7618 32545 7624
rect 32400 7550 32410 7618
rect 32268 7510 32400 7550
rect 32267 7444 32400 7510
rect 30441 7128 31118 7131
rect 28027 6965 28073 6977
rect 29965 7116 30011 7128
rect 27325 6923 27359 6965
rect 27561 6923 27595 6965
rect 27325 6895 27595 6923
rect 27679 6924 27713 6965
rect 27915 6924 27949 6965
rect 27679 6895 27949 6924
rect 27325 6847 27359 6895
rect 27325 6817 27388 6847
rect 27353 6725 27388 6817
rect 27860 6787 27960 6808
rect 27860 6733 27874 6787
rect 27939 6733 27960 6787
rect 27860 6728 27960 6733
rect 28033 6782 28067 6965
rect 28033 6728 28142 6782
rect 27353 6689 27580 6725
rect 27353 6582 27388 6689
rect 27514 6655 27580 6689
rect 27514 6621 27530 6655
rect 27564 6621 27580 6655
rect 27861 6713 27958 6728
rect 27861 6646 27918 6713
rect 27514 6615 27580 6621
rect 27755 6610 28024 6646
rect 27755 6582 27788 6610
rect 27991 6582 28024 6610
rect 28108 6582 28142 6728
rect 29800 6779 29904 6787
rect 29800 6678 29810 6779
rect 29896 6696 29906 6779
rect 29965 6740 29971 7116
rect 30005 6740 30011 7116
rect 29965 6728 30011 6740
rect 30083 7116 30129 7128
rect 30083 6740 30089 7116
rect 30123 6740 30129 7116
rect 30083 6728 30129 6740
rect 30201 7116 30247 7128
rect 30201 6740 30207 7116
rect 30241 6767 30247 7116
rect 30318 7116 30364 7128
rect 30318 6940 30324 7116
rect 30358 6940 30364 7116
rect 30318 6933 30364 6940
rect 30436 7116 31118 7128
rect 30436 6940 30442 7116
rect 30476 7103 31118 7116
rect 30476 6940 30482 7103
rect 30726 7023 31118 7103
rect 31596 7401 33069 7444
rect 31596 7098 31630 7401
rect 31962 7298 31996 7401
rect 32198 7298 32232 7401
rect 32434 7298 32468 7401
rect 32670 7298 32704 7401
rect 31956 7286 32002 7298
rect 31472 7086 31518 7098
rect 30318 6928 30367 6933
rect 30436 6928 30482 6940
rect 30324 6767 30367 6928
rect 31472 6910 31478 7086
rect 31512 6910 31518 7086
rect 31472 6898 31518 6910
rect 31590 7086 31636 7098
rect 31590 6910 31596 7086
rect 31630 6910 31636 7086
rect 31590 6898 31636 6910
rect 31708 7086 31754 7098
rect 31708 6910 31714 7086
rect 31748 6910 31754 7086
rect 31708 6898 31754 6910
rect 31826 7086 31872 7098
rect 31956 7086 31962 7286
rect 31826 6910 31832 7086
rect 31866 6910 31962 7086
rect 31996 6910 32002 7286
rect 31826 6898 31872 6910
rect 31956 6898 32002 6910
rect 32074 7286 32120 7298
rect 32074 6910 32080 7286
rect 32114 6910 32120 7286
rect 32074 6898 32120 6910
rect 32192 7286 32238 7298
rect 32192 6910 32198 7286
rect 32232 6910 32238 7286
rect 32192 6898 32238 6910
rect 32310 7286 32356 7298
rect 32310 6910 32316 7286
rect 32350 6910 32356 7286
rect 32310 6898 32356 6910
rect 32428 7286 32474 7298
rect 32428 6910 32434 7286
rect 32468 6910 32474 7286
rect 32428 6898 32474 6910
rect 32546 7286 32592 7298
rect 32546 6910 32552 7286
rect 32586 6910 32592 7286
rect 32546 6898 32592 6910
rect 32664 7286 32710 7298
rect 32664 6910 32670 7286
rect 32704 7086 32710 7286
rect 33035 7098 33069 7401
rect 33576 7321 33712 7341
rect 33576 7259 33612 7321
rect 33672 7259 33712 7321
rect 33576 7231 33712 7259
rect 33272 7201 34249 7231
rect 32793 7086 32839 7098
rect 32704 6910 32799 7086
rect 32833 6910 32839 7086
rect 32664 6898 32710 6910
rect 32793 6898 32839 6910
rect 32911 7086 32957 7098
rect 32911 6910 32917 7086
rect 32951 6910 32957 7086
rect 32911 6898 32957 6910
rect 33029 7086 33075 7098
rect 33029 6910 33035 7086
rect 33069 6910 33075 7086
rect 33029 6898 33075 6910
rect 33147 7086 33193 7098
rect 33272 7095 33304 7201
rect 33508 7095 33540 7201
rect 33744 7095 33776 7201
rect 33980 7095 34012 7201
rect 34215 7095 34249 7201
rect 33147 6910 33153 7086
rect 33187 6910 33193 7086
rect 33147 6898 33193 6910
rect 33265 7083 33311 7095
rect 33265 6907 33271 7083
rect 33305 6907 33311 7083
rect 31478 6864 31512 6898
rect 32080 6864 32114 6898
rect 32316 6864 32350 6898
rect 31478 6829 31637 6864
rect 32080 6829 32350 6864
rect 32917 6864 32951 6898
rect 33153 6864 33187 6898
rect 33265 6895 33311 6907
rect 33383 7083 33429 7095
rect 33383 6907 33389 7083
rect 33423 6907 33429 7083
rect 33383 6895 33429 6907
rect 33501 7083 33547 7095
rect 33501 6907 33507 7083
rect 33541 6907 33547 7083
rect 33501 6895 33547 6907
rect 33619 7083 33665 7095
rect 33619 6907 33625 7083
rect 33659 6907 33665 7083
rect 33619 6895 33665 6907
rect 33737 7083 33783 7095
rect 33737 6907 33743 7083
rect 33777 6907 33783 7083
rect 33737 6895 33783 6907
rect 33855 7083 33901 7095
rect 33855 6907 33861 7083
rect 33895 6907 33901 7083
rect 33855 6895 33901 6907
rect 33973 7083 34019 7095
rect 33973 6907 33979 7083
rect 34013 6907 34019 7083
rect 33973 6895 34019 6907
rect 34091 7083 34137 7095
rect 34091 6907 34097 7083
rect 34131 6907 34137 7083
rect 34091 6895 34137 6907
rect 34209 7083 34255 7095
rect 34209 6907 34215 7083
rect 34249 6907 34255 7083
rect 34209 6895 34255 6907
rect 34327 7083 34373 7095
rect 34327 6907 34333 7083
rect 34367 6907 34373 7083
rect 34327 6895 34373 6907
rect 32917 6829 33187 6864
rect 30241 6740 30367 6767
rect 30201 6728 30367 6740
rect 30207 6724 30367 6728
rect 29896 6690 30080 6696
rect 29896 6678 30030 6690
rect 29800 6656 30030 6678
rect 30064 6656 30080 6690
rect 29800 6640 30080 6656
rect 30132 6690 30198 6696
rect 30132 6656 30148 6690
rect 30182 6656 30198 6690
rect 30132 6611 30198 6656
rect 29577 6605 30198 6611
rect 27229 6570 27275 6582
rect 27229 6394 27235 6570
rect 27269 6394 27275 6570
rect 27229 6382 27275 6394
rect 27347 6570 27393 6582
rect 27347 6394 27353 6570
rect 27387 6394 27393 6570
rect 27347 6382 27393 6394
rect 27465 6570 27511 6582
rect 27465 6394 27471 6570
rect 27505 6394 27511 6570
rect 27465 6382 27511 6394
rect 27583 6570 27629 6582
rect 27583 6394 27589 6570
rect 27623 6515 27629 6570
rect 27748 6570 27794 6582
rect 27748 6515 27754 6570
rect 27623 6427 27754 6515
rect 27623 6394 27629 6427
rect 27583 6382 27629 6394
rect 27748 6394 27754 6427
rect 27788 6394 27794 6570
rect 27748 6382 27794 6394
rect 27866 6570 27912 6582
rect 27866 6394 27872 6570
rect 27906 6394 27912 6570
rect 27866 6382 27912 6394
rect 27984 6570 28030 6582
rect 27984 6394 27990 6570
rect 28024 6394 28030 6570
rect 27984 6382 28030 6394
rect 28102 6570 28148 6582
rect 28102 6394 28108 6570
rect 28142 6394 28148 6570
rect 29572 6545 29582 6605
rect 29667 6603 30198 6605
rect 29667 6571 30199 6603
rect 30291 6587 30367 6724
rect 29667 6545 29677 6571
rect 29577 6538 29672 6545
rect 30287 6527 30297 6587
rect 30359 6527 30369 6587
rect 31024 6555 31465 6618
rect 31532 6555 31542 6618
rect 28102 6382 28148 6394
rect 27235 6343 27269 6382
rect 27471 6343 27505 6382
rect 27235 6307 27505 6343
rect 27872 6344 27905 6382
rect 28108 6344 28141 6382
rect 27872 6308 28141 6344
rect 27235 6306 27401 6307
rect 27269 6227 27401 6306
rect 27259 6119 27269 6227
rect 27401 6119 27411 6227
rect 27290 5982 27296 6119
rect 27363 5982 27369 6119
rect 27290 5970 27369 5982
rect 23873 5745 24850 5775
rect 27067 5773 27130 5790
rect 26992 5769 27130 5773
rect 23873 5639 23905 5745
rect 24109 5639 24141 5745
rect 24345 5639 24377 5745
rect 24581 5639 24613 5745
rect 24816 5639 24850 5745
rect 25160 5735 27130 5769
rect 25158 5706 27130 5735
rect 25158 5690 25204 5706
rect 26992 5704 27130 5706
rect 23866 5627 23912 5639
rect 23866 5451 23872 5627
rect 23906 5451 23912 5627
rect 23866 5439 23912 5451
rect 23984 5627 24030 5639
rect 23984 5451 23990 5627
rect 24024 5451 24030 5627
rect 23984 5439 24030 5451
rect 24102 5627 24148 5639
rect 24102 5451 24108 5627
rect 24142 5451 24148 5627
rect 24102 5439 24148 5451
rect 24220 5627 24266 5639
rect 24220 5451 24226 5627
rect 24260 5451 24266 5627
rect 24220 5439 24266 5451
rect 24338 5627 24384 5639
rect 24338 5451 24344 5627
rect 24378 5451 24384 5627
rect 24338 5439 24384 5451
rect 24456 5627 24502 5639
rect 24456 5451 24462 5627
rect 24496 5451 24502 5627
rect 24456 5439 24502 5451
rect 24574 5627 24620 5639
rect 24574 5451 24580 5627
rect 24614 5451 24620 5627
rect 24574 5439 24620 5451
rect 24692 5627 24738 5639
rect 24692 5451 24698 5627
rect 24732 5451 24738 5627
rect 24692 5439 24738 5451
rect 24810 5627 24856 5639
rect 24810 5451 24816 5627
rect 24850 5451 24856 5627
rect 24810 5439 24856 5451
rect 24928 5627 24974 5639
rect 24928 5451 24934 5627
rect 24968 5451 24974 5627
rect 24928 5439 24974 5451
rect 23989 5345 24025 5439
rect 24225 5345 24261 5439
rect 24461 5346 24497 5439
rect 24623 5391 24689 5398
rect 24623 5357 24639 5391
rect 24673 5357 24689 5391
rect 24623 5346 24689 5357
rect 24461 5345 24689 5346
rect 23989 5316 24689 5345
rect 23989 5315 24571 5316
rect 24109 5202 24143 5315
rect 24505 5274 24571 5315
rect 24505 5240 24521 5274
rect 24555 5240 24571 5274
rect 24505 5233 24571 5240
rect 24933 5221 24968 5439
rect 25157 5238 25204 5690
rect 28053 5697 28132 5709
rect 28053 5582 28059 5697
rect 28126 5582 28132 5697
rect 26116 5474 26126 5582
rect 26258 5474 26268 5582
rect 28014 5474 28024 5582
rect 28156 5474 28166 5582
rect 26126 5434 26258 5474
rect 28024 5434 28156 5474
rect 26125 5368 26258 5434
rect 28023 5368 28156 5434
rect 25454 5325 26927 5368
rect 25157 5222 25203 5238
rect 25122 5221 25203 5222
rect 24933 5206 25203 5221
rect 24579 5202 25203 5206
rect 24103 5190 24149 5202
rect 23838 4712 23848 4830
rect 23966 4798 23976 4830
rect 24103 4814 24109 5190
rect 24143 4814 24149 5190
rect 24103 4802 24149 4814
rect 24221 5190 24267 5202
rect 24221 4814 24227 5190
rect 24261 4814 24267 5190
rect 24221 4802 24267 4814
rect 24339 5190 24385 5202
rect 24339 4814 24345 5190
rect 24379 4838 24385 5190
rect 24456 5190 24502 5202
rect 24456 5014 24462 5190
rect 24496 5014 24502 5190
rect 24456 5002 24502 5014
rect 24574 5190 25203 5202
rect 24574 5014 24580 5190
rect 24614 5178 25203 5190
rect 24614 5177 24856 5178
rect 24614 5014 24620 5177
rect 25122 5176 25203 5178
rect 25454 5022 25488 5325
rect 25820 5222 25854 5325
rect 26056 5222 26090 5325
rect 26292 5222 26326 5325
rect 26528 5222 26562 5325
rect 25814 5210 25860 5222
rect 24574 5002 24620 5014
rect 25330 5010 25376 5022
rect 24462 4886 24497 5002
rect 24593 4886 24701 4896
rect 24462 4838 24593 4886
rect 24701 4855 24850 4861
rect 24379 4814 24593 4838
rect 24339 4802 24593 4814
rect 24345 4798 24593 4802
rect 23966 4770 23981 4798
rect 23966 4764 24218 4770
rect 23966 4730 24168 4764
rect 24202 4730 24218 4764
rect 23966 4714 24218 4730
rect 24270 4764 24336 4770
rect 24270 4730 24286 4764
rect 24320 4730 24336 4764
rect 24519 4754 24593 4798
rect 24838 4788 24850 4855
rect 25330 4834 25336 5010
rect 25370 4834 25376 5010
rect 25330 4822 25376 4834
rect 25448 5010 25494 5022
rect 25448 4834 25454 5010
rect 25488 4834 25494 5010
rect 25448 4822 25494 4834
rect 25566 5010 25612 5022
rect 25566 4834 25572 5010
rect 25606 4834 25612 5010
rect 25566 4822 25612 4834
rect 25684 5010 25730 5022
rect 25814 5010 25820 5210
rect 25684 4834 25690 5010
rect 25724 4834 25820 5010
rect 25854 4834 25860 5210
rect 25684 4822 25730 4834
rect 25814 4822 25860 4834
rect 25932 5210 25978 5222
rect 25932 4834 25938 5210
rect 25972 4834 25978 5210
rect 25932 4822 25978 4834
rect 26050 5210 26096 5222
rect 26050 4834 26056 5210
rect 26090 4834 26096 5210
rect 26050 4822 26096 4834
rect 26168 5210 26214 5222
rect 26168 4834 26174 5210
rect 26208 4834 26214 5210
rect 26168 4822 26214 4834
rect 26286 5210 26332 5222
rect 26286 4834 26292 5210
rect 26326 4834 26332 5210
rect 26286 4822 26332 4834
rect 26404 5210 26450 5222
rect 26404 4834 26410 5210
rect 26444 4834 26450 5210
rect 26404 4822 26450 4834
rect 26522 5210 26568 5222
rect 26522 4834 26528 5210
rect 26562 5010 26568 5210
rect 26893 5022 26927 5325
rect 27352 5325 28825 5368
rect 27352 5022 27386 5325
rect 27718 5222 27752 5325
rect 27954 5222 27988 5325
rect 28190 5222 28224 5325
rect 28426 5222 28460 5325
rect 27712 5210 27758 5222
rect 26651 5010 26697 5022
rect 26562 4834 26657 5010
rect 26691 4834 26697 5010
rect 26522 4822 26568 4834
rect 26651 4822 26697 4834
rect 26769 5010 26815 5022
rect 26769 4834 26775 5010
rect 26809 4834 26815 5010
rect 26769 4822 26815 4834
rect 26887 5010 26933 5022
rect 26887 4834 26893 5010
rect 26927 4834 26933 5010
rect 26887 4822 26933 4834
rect 27005 5010 27051 5022
rect 27005 4834 27011 5010
rect 27045 4834 27051 5010
rect 27005 4822 27051 4834
rect 27228 5010 27274 5022
rect 27228 4834 27234 5010
rect 27268 4834 27274 5010
rect 27228 4822 27274 4834
rect 27346 5010 27392 5022
rect 27346 4834 27352 5010
rect 27386 4834 27392 5010
rect 27346 4822 27392 4834
rect 27464 5010 27510 5022
rect 27464 4834 27470 5010
rect 27504 4834 27510 5010
rect 27464 4822 27510 4834
rect 27582 5010 27628 5022
rect 27712 5010 27718 5210
rect 27582 4834 27588 5010
rect 27622 4834 27718 5010
rect 27752 4834 27758 5210
rect 27582 4822 27628 4834
rect 27712 4822 27758 4834
rect 27830 5210 27876 5222
rect 27830 4834 27836 5210
rect 27870 4834 27876 5210
rect 27830 4822 27876 4834
rect 27948 5210 27994 5222
rect 27948 4834 27954 5210
rect 27988 4834 27994 5210
rect 27948 4822 27994 4834
rect 28066 5210 28112 5222
rect 28066 4834 28072 5210
rect 28106 4834 28112 5210
rect 28066 4822 28112 4834
rect 28184 5210 28230 5222
rect 28184 4834 28190 5210
rect 28224 4834 28230 5210
rect 28184 4822 28230 4834
rect 28302 5210 28348 5222
rect 28302 4834 28308 5210
rect 28342 4834 28348 5210
rect 28302 4822 28348 4834
rect 28420 5210 28466 5222
rect 28420 4834 28426 5210
rect 28460 5010 28466 5210
rect 28791 5022 28825 5325
rect 28549 5010 28595 5022
rect 28460 4834 28555 5010
rect 28589 4834 28595 5010
rect 28420 4822 28466 4834
rect 28549 4822 28595 4834
rect 28667 5010 28713 5022
rect 28667 4834 28673 5010
rect 28707 4834 28713 5010
rect 28667 4822 28713 4834
rect 28785 5010 28831 5022
rect 28785 4834 28791 5010
rect 28825 4834 28831 5010
rect 28785 4822 28831 4834
rect 28903 5010 28949 5022
rect 28903 4834 28909 5010
rect 28943 4834 28949 5010
rect 28903 4822 28949 4834
rect 24701 4782 24850 4788
rect 25336 4788 25370 4822
rect 25938 4788 25972 4822
rect 26174 4788 26208 4822
rect 24593 4744 24701 4754
rect 25336 4753 25495 4788
rect 25938 4753 26208 4788
rect 26775 4788 26809 4822
rect 27011 4788 27045 4822
rect 26775 4753 27045 4788
rect 27234 4788 27268 4822
rect 27836 4788 27870 4822
rect 28072 4788 28106 4822
rect 27234 4753 27393 4788
rect 27836 4753 28106 4788
rect 28673 4788 28707 4822
rect 28909 4788 28943 4822
rect 28673 4753 28943 4788
rect 23966 4712 23981 4714
rect 23881 4698 23981 4712
rect 23881 4655 23981 4656
rect 23502 4634 23981 4655
rect 24270 4634 24336 4730
rect 23502 4586 24336 4634
rect 23502 4557 23981 4586
rect 23502 4555 23607 4557
rect 23881 4556 23981 4557
rect 23335 4370 23345 4449
rect 23438 4370 23448 4449
rect 24337 4433 24416 4445
rect 23346 3196 23439 4370
rect 24337 4341 24343 4433
rect 24264 4321 24343 4341
rect 24410 4341 24416 4433
rect 24410 4321 24484 4341
rect 24264 4213 24308 4321
rect 24440 4213 24484 4321
rect 24264 4171 24484 4213
rect 23868 4141 24845 4171
rect 23868 4035 23900 4141
rect 24104 4035 24136 4141
rect 24340 4035 24372 4141
rect 24576 4035 24608 4141
rect 24811 4035 24845 4141
rect 23861 4023 23907 4035
rect 23861 3847 23867 4023
rect 23901 3847 23907 4023
rect 23861 3835 23907 3847
rect 23979 4023 24025 4035
rect 23979 3847 23985 4023
rect 24019 3847 24025 4023
rect 23979 3835 24025 3847
rect 24097 4023 24143 4035
rect 24097 3847 24103 4023
rect 24137 3847 24143 4023
rect 24097 3835 24143 3847
rect 24215 4023 24261 4035
rect 24215 3847 24221 4023
rect 24255 3847 24261 4023
rect 24215 3835 24261 3847
rect 24333 4023 24379 4035
rect 24333 3847 24339 4023
rect 24373 3847 24379 4023
rect 24333 3835 24379 3847
rect 24451 4023 24497 4035
rect 24451 3847 24457 4023
rect 24491 3847 24497 4023
rect 24451 3835 24497 3847
rect 24569 4023 24615 4035
rect 24569 3847 24575 4023
rect 24609 3847 24615 4023
rect 24569 3835 24615 3847
rect 24687 4023 24733 4035
rect 24687 3847 24693 4023
rect 24727 3847 24733 4023
rect 24687 3835 24733 3847
rect 24805 4023 24851 4035
rect 24805 3847 24811 4023
rect 24845 3847 24851 4023
rect 24805 3835 24851 3847
rect 24923 4023 24969 4035
rect 24923 3847 24929 4023
rect 24963 3847 24969 4023
rect 24923 3835 24969 3847
rect 25461 3969 25495 4753
rect 26174 4691 26208 4753
rect 25763 4653 26505 4691
rect 25763 4529 25797 4653
rect 25999 4529 26033 4653
rect 26235 4529 26269 4653
rect 26471 4529 26505 4653
rect 26761 4546 26771 4612
rect 26834 4546 26844 4612
rect 25757 4517 25803 4529
rect 25757 4141 25763 4517
rect 25797 4141 25803 4517
rect 25757 4129 25803 4141
rect 25875 4517 25921 4529
rect 25875 4141 25881 4517
rect 25915 4141 25921 4517
rect 25875 4129 25921 4141
rect 25993 4517 26039 4529
rect 25993 4141 25999 4517
rect 26033 4141 26039 4517
rect 25993 4129 26039 4141
rect 26111 4517 26157 4529
rect 26111 4141 26117 4517
rect 26151 4141 26157 4517
rect 26111 4129 26157 4141
rect 26229 4517 26275 4529
rect 26229 4141 26235 4517
rect 26269 4141 26275 4517
rect 26229 4129 26275 4141
rect 26347 4517 26393 4529
rect 26347 4141 26353 4517
rect 26387 4141 26393 4517
rect 26347 4129 26393 4141
rect 26465 4517 26511 4529
rect 26465 4141 26471 4517
rect 26505 4141 26511 4517
rect 26465 4129 26511 4141
rect 26877 3970 26911 4753
rect 26604 3969 26911 3970
rect 25461 3964 25777 3969
rect 26491 3964 26911 3969
rect 25461 3953 25844 3964
rect 25461 3926 25793 3953
rect 23984 3741 24020 3835
rect 24220 3741 24256 3835
rect 24456 3742 24492 3835
rect 24618 3787 24684 3794
rect 24618 3753 24634 3787
rect 24668 3753 24684 3787
rect 24618 3742 24684 3753
rect 24456 3741 24684 3742
rect 23984 3712 24684 3741
rect 23984 3711 24566 3712
rect 24104 3598 24138 3711
rect 24500 3670 24566 3711
rect 24500 3636 24516 3670
rect 24550 3636 24566 3670
rect 24500 3629 24566 3636
rect 24928 3602 24963 3835
rect 25461 3797 25495 3926
rect 25777 3919 25793 3926
rect 25827 3919 25844 3953
rect 25777 3913 25844 3919
rect 26424 3953 26911 3964
rect 26424 3919 26441 3953
rect 26475 3926 26911 3953
rect 26475 3919 26491 3926
rect 26604 3925 26911 3926
rect 26424 3913 26491 3919
rect 25602 3886 25658 3898
rect 25602 3852 25608 3886
rect 25642 3885 25658 3886
rect 26715 3885 26771 3897
rect 25642 3869 26109 3885
rect 25642 3852 26059 3869
rect 25602 3836 26059 3852
rect 26043 3835 26059 3836
rect 26093 3835 26109 3869
rect 26043 3828 26109 3835
rect 26161 3870 26731 3885
rect 26161 3836 26177 3870
rect 26211 3851 26731 3870
rect 26765 3851 26771 3885
rect 26211 3836 26771 3851
rect 26161 3826 26228 3836
rect 26715 3835 26771 3836
rect 26877 3797 26911 3925
rect 27359 3969 27393 4753
rect 28072 4691 28106 4753
rect 27661 4653 28403 4691
rect 27661 4529 27695 4653
rect 27897 4529 27931 4653
rect 28133 4529 28167 4653
rect 28369 4529 28403 4653
rect 27655 4517 27701 4529
rect 27655 4141 27661 4517
rect 27695 4141 27701 4517
rect 27655 4129 27701 4141
rect 27773 4517 27819 4529
rect 27773 4141 27779 4517
rect 27813 4141 27819 4517
rect 27773 4129 27819 4141
rect 27891 4517 27937 4529
rect 27891 4141 27897 4517
rect 27931 4141 27937 4517
rect 27891 4129 27937 4141
rect 28009 4517 28055 4529
rect 28009 4141 28015 4517
rect 28049 4141 28055 4517
rect 28009 4129 28055 4141
rect 28127 4517 28173 4529
rect 28127 4141 28133 4517
rect 28167 4141 28173 4517
rect 28127 4129 28173 4141
rect 28245 4517 28291 4529
rect 28245 4141 28251 4517
rect 28285 4141 28291 4517
rect 28245 4129 28291 4141
rect 28363 4517 28409 4529
rect 28363 4141 28369 4517
rect 28403 4141 28409 4517
rect 28363 4129 28409 4141
rect 28775 3970 28809 4753
rect 30036 4721 30172 4741
rect 30036 4659 30072 4721
rect 30132 4659 30172 4721
rect 30036 4631 30172 4659
rect 29732 4601 30709 4631
rect 28387 3969 28456 3970
rect 28502 3969 28809 3970
rect 27359 3964 27675 3969
rect 28387 3965 28809 3969
rect 27359 3953 27742 3964
rect 27359 3926 27691 3953
rect 27359 3797 27393 3926
rect 27675 3919 27691 3926
rect 27725 3919 27742 3953
rect 27675 3913 27742 3919
rect 28320 3954 28809 3965
rect 28320 3920 28337 3954
rect 28371 3926 28809 3954
rect 28371 3920 28387 3926
rect 28502 3925 28809 3926
rect 28320 3914 28387 3920
rect 27500 3886 27556 3898
rect 27500 3852 27506 3886
rect 27540 3885 27556 3886
rect 28613 3885 28669 3897
rect 27540 3869 28007 3885
rect 27540 3852 27957 3869
rect 27500 3836 27957 3852
rect 27941 3835 27957 3836
rect 27991 3835 28007 3869
rect 27941 3828 28007 3835
rect 28059 3870 28629 3885
rect 28059 3836 28075 3870
rect 28109 3851 28629 3870
rect 28663 3851 28669 3885
rect 28109 3836 28669 3851
rect 28059 3826 28126 3836
rect 28613 3835 28669 3836
rect 28775 3797 28809 3925
rect 28890 4575 28957 4599
rect 28890 4541 28907 4575
rect 28941 4541 28957 4575
rect 24574 3598 24963 3602
rect 24098 3586 24144 3598
rect 24098 3210 24104 3586
rect 24138 3210 24144 3586
rect 24098 3198 24144 3210
rect 24216 3586 24262 3598
rect 24216 3210 24222 3586
rect 24256 3210 24262 3586
rect 24216 3198 24262 3210
rect 24334 3586 24380 3598
rect 24334 3210 24340 3586
rect 24374 3234 24380 3586
rect 24451 3586 24497 3598
rect 24451 3410 24457 3586
rect 24491 3410 24497 3586
rect 24451 3398 24497 3410
rect 24569 3586 24963 3598
rect 25455 3785 25501 3797
rect 25455 3609 25461 3785
rect 25495 3609 25501 3785
rect 25455 3597 25501 3609
rect 25573 3785 25619 3797
rect 25573 3609 25579 3785
rect 25613 3609 25619 3785
rect 25573 3597 25619 3609
rect 25875 3785 25921 3797
rect 24569 3410 24575 3586
rect 24609 3573 24963 3586
rect 24609 3410 24615 3573
rect 24885 3570 24963 3573
rect 24885 3518 24895 3570
rect 24958 3518 24968 3570
rect 24890 3512 24963 3518
rect 24569 3398 24615 3410
rect 24457 3282 24492 3398
rect 25578 3303 25612 3597
rect 25875 3409 25881 3785
rect 25915 3409 25921 3785
rect 25875 3397 25921 3409
rect 25993 3785 26039 3797
rect 25993 3409 25999 3785
rect 26033 3409 26039 3785
rect 25993 3397 26039 3409
rect 26111 3785 26157 3797
rect 26111 3409 26117 3785
rect 26151 3409 26157 3785
rect 26111 3397 26157 3409
rect 26229 3785 26275 3797
rect 26229 3409 26235 3785
rect 26269 3409 26275 3785
rect 26229 3397 26275 3409
rect 26347 3785 26393 3797
rect 26347 3409 26353 3785
rect 26387 3409 26393 3785
rect 26753 3785 26799 3797
rect 26753 3609 26759 3785
rect 26793 3609 26799 3785
rect 26753 3597 26799 3609
rect 26871 3785 26917 3797
rect 26871 3609 26877 3785
rect 26911 3609 26917 3785
rect 26871 3597 26917 3609
rect 27353 3785 27399 3797
rect 27353 3609 27359 3785
rect 27393 3609 27399 3785
rect 27353 3597 27399 3609
rect 27471 3785 27517 3797
rect 27471 3609 27477 3785
rect 27511 3609 27517 3785
rect 27471 3597 27517 3609
rect 27773 3785 27819 3797
rect 26347 3397 26393 3409
rect 26235 3303 26269 3397
rect 26759 3303 26792 3597
rect 24588 3282 24696 3292
rect 24457 3234 24588 3282
rect 25578 3271 26792 3303
rect 27476 3303 27510 3597
rect 27773 3409 27779 3785
rect 27813 3409 27819 3785
rect 27773 3397 27819 3409
rect 27891 3785 27937 3797
rect 27891 3409 27897 3785
rect 27931 3409 27937 3785
rect 27891 3397 27937 3409
rect 28009 3785 28055 3797
rect 28009 3409 28015 3785
rect 28049 3409 28055 3785
rect 28009 3397 28055 3409
rect 28127 3785 28173 3797
rect 28127 3409 28133 3785
rect 28167 3409 28173 3785
rect 28127 3397 28173 3409
rect 28245 3785 28291 3797
rect 28245 3409 28251 3785
rect 28285 3409 28291 3785
rect 28651 3785 28697 3797
rect 28651 3609 28657 3785
rect 28691 3609 28697 3785
rect 28651 3597 28697 3609
rect 28769 3785 28815 3797
rect 28769 3609 28775 3785
rect 28809 3609 28815 3785
rect 28769 3597 28815 3609
rect 28245 3397 28291 3409
rect 28133 3303 28167 3397
rect 28657 3303 28690 3597
rect 27476 3271 28690 3303
rect 24696 3238 24841 3244
rect 24374 3210 24588 3234
rect 24334 3198 24588 3210
rect 23346 3194 23931 3196
rect 24340 3194 24588 3198
rect 23346 3166 23976 3194
rect 23346 3160 24213 3166
rect 23346 3126 24163 3160
rect 24197 3126 24213 3160
rect 23346 3110 24213 3126
rect 24265 3160 24331 3166
rect 24265 3126 24281 3160
rect 24315 3126 24331 3160
rect 24514 3150 24588 3194
rect 24829 3171 24841 3238
rect 26071 3186 26203 3271
rect 27969 3186 28101 3271
rect 24696 3165 24841 3171
rect 24588 3140 24696 3150
rect 23346 3094 23976 3110
rect 23346 3090 23931 3094
rect 23346 3089 23447 3090
rect 23876 3041 23976 3052
rect 23840 2935 23850 3041
rect 23962 3030 23976 3041
rect 24265 3030 24331 3126
rect 26061 3078 26071 3186
rect 26203 3078 26213 3186
rect 27959 3078 27969 3186
rect 28101 3078 28111 3186
rect 28890 3158 28957 4541
rect 29732 4495 29764 4601
rect 29968 4495 30000 4601
rect 30204 4495 30236 4601
rect 30440 4495 30472 4601
rect 30675 4495 30709 4601
rect 29725 4483 29771 4495
rect 29725 4307 29731 4483
rect 29765 4307 29771 4483
rect 29725 4295 29771 4307
rect 29843 4483 29889 4495
rect 29843 4307 29849 4483
rect 29883 4307 29889 4483
rect 29843 4295 29889 4307
rect 29961 4483 30007 4495
rect 29961 4307 29967 4483
rect 30001 4307 30007 4483
rect 29961 4295 30007 4307
rect 30079 4483 30125 4495
rect 30079 4307 30085 4483
rect 30119 4307 30125 4483
rect 30079 4295 30125 4307
rect 30197 4483 30243 4495
rect 30197 4307 30203 4483
rect 30237 4307 30243 4483
rect 30197 4295 30243 4307
rect 30315 4483 30361 4495
rect 30315 4307 30321 4483
rect 30355 4307 30361 4483
rect 30315 4295 30361 4307
rect 30433 4483 30479 4495
rect 30433 4307 30439 4483
rect 30473 4307 30479 4483
rect 30433 4295 30479 4307
rect 30551 4483 30597 4495
rect 30551 4307 30557 4483
rect 30591 4307 30597 4483
rect 30551 4295 30597 4307
rect 30669 4483 30715 4495
rect 30669 4307 30675 4483
rect 30709 4307 30715 4483
rect 30669 4295 30715 4307
rect 30787 4483 30833 4495
rect 30787 4307 30793 4483
rect 30827 4307 30833 4483
rect 30787 4295 30833 4307
rect 29848 4201 29884 4295
rect 30084 4201 30120 4295
rect 30320 4202 30356 4295
rect 30482 4247 30548 4254
rect 30482 4213 30498 4247
rect 30532 4213 30548 4247
rect 30482 4202 30548 4213
rect 30320 4201 30548 4202
rect 29848 4172 30548 4201
rect 29848 4171 30430 4172
rect 29018 4112 29174 4118
rect 29018 4014 29030 4112
rect 29162 4014 29174 4112
rect 29968 4058 30002 4171
rect 30364 4130 30430 4171
rect 30364 4096 30380 4130
rect 30414 4096 30430 4130
rect 30364 4089 30430 4096
rect 30792 4062 30827 4295
rect 30438 4061 30973 4062
rect 31024 4061 31119 6555
rect 31603 6045 31637 6829
rect 32316 6767 32350 6829
rect 31905 6729 32647 6767
rect 31715 6558 31725 6626
rect 31780 6558 31790 6626
rect 31905 6605 31939 6729
rect 32141 6605 32175 6729
rect 32377 6605 32411 6729
rect 32613 6605 32647 6729
rect 31899 6593 31945 6605
rect 31899 6217 31905 6593
rect 31939 6217 31945 6593
rect 31899 6205 31945 6217
rect 32017 6593 32063 6605
rect 32017 6217 32023 6593
rect 32057 6217 32063 6593
rect 32017 6205 32063 6217
rect 32135 6593 32181 6605
rect 32135 6217 32141 6593
rect 32175 6217 32181 6593
rect 32135 6205 32181 6217
rect 32253 6593 32299 6605
rect 32253 6217 32259 6593
rect 32293 6217 32299 6593
rect 32253 6205 32299 6217
rect 32371 6593 32417 6605
rect 32371 6217 32377 6593
rect 32411 6217 32417 6593
rect 32371 6205 32417 6217
rect 32489 6593 32535 6605
rect 32489 6217 32495 6593
rect 32529 6217 32535 6593
rect 32489 6205 32535 6217
rect 32607 6593 32653 6605
rect 32607 6217 32613 6593
rect 32647 6217 32653 6593
rect 32773 6388 32847 6400
rect 32769 6297 32779 6388
rect 32841 6297 32851 6388
rect 32773 6285 32847 6297
rect 32607 6205 32653 6217
rect 33019 6046 33053 6829
rect 33388 6801 33424 6895
rect 33624 6801 33660 6895
rect 33860 6802 33896 6895
rect 34022 6847 34088 6854
rect 34022 6813 34038 6847
rect 34072 6813 34088 6847
rect 34022 6802 34088 6813
rect 33860 6801 34088 6802
rect 33388 6772 34088 6801
rect 33388 6771 33970 6772
rect 33114 6739 33190 6744
rect 33111 6683 33121 6739
rect 33174 6738 33190 6739
rect 33174 6683 33440 6738
rect 33114 6678 33440 6683
rect 33235 6636 33326 6641
rect 33235 6547 33245 6636
rect 33318 6547 33326 6636
rect 33235 6535 33326 6547
rect 33272 6141 33326 6535
rect 33386 6226 33440 6678
rect 33508 6658 33542 6771
rect 33904 6730 33970 6771
rect 33904 6696 33920 6730
rect 33954 6696 33970 6730
rect 33904 6689 33970 6696
rect 34332 6662 34367 6895
rect 33978 6658 34367 6662
rect 33502 6646 33548 6658
rect 33502 6270 33508 6646
rect 33542 6270 33548 6646
rect 33502 6258 33548 6270
rect 33620 6646 33666 6658
rect 33620 6270 33626 6646
rect 33660 6270 33666 6646
rect 33620 6258 33666 6270
rect 33738 6646 33784 6658
rect 33738 6270 33744 6646
rect 33778 6297 33784 6646
rect 33855 6646 33901 6658
rect 33855 6470 33861 6646
rect 33895 6470 33901 6646
rect 33855 6463 33901 6470
rect 33973 6646 34367 6658
rect 33973 6470 33979 6646
rect 34013 6633 34367 6646
rect 34013 6470 34019 6633
rect 34192 6544 34367 6633
rect 34236 6543 34367 6544
rect 33855 6458 33904 6463
rect 33973 6458 34019 6470
rect 33861 6297 33904 6458
rect 33778 6270 33904 6297
rect 33738 6258 33904 6270
rect 33744 6254 33904 6258
rect 33386 6220 33617 6226
rect 33386 6186 33567 6220
rect 33601 6186 33617 6220
rect 33386 6170 33617 6186
rect 33669 6220 33735 6226
rect 33669 6186 33685 6220
rect 33719 6186 33735 6220
rect 33669 6141 33735 6186
rect 33272 6133 33735 6141
rect 33272 6101 33736 6133
rect 33828 6117 33904 6254
rect 33824 6057 33834 6117
rect 33896 6057 33906 6117
rect 32746 6045 33053 6046
rect 31603 6040 31919 6045
rect 32633 6040 33053 6045
rect 31603 6029 31986 6040
rect 31603 6002 31935 6029
rect 31603 5873 31637 6002
rect 31919 5995 31935 6002
rect 31969 5995 31986 6029
rect 31919 5989 31986 5995
rect 32566 6029 33053 6040
rect 33832 6031 33902 6057
rect 32566 5995 32583 6029
rect 32617 6002 33053 6029
rect 32617 5995 32633 6002
rect 32746 6001 33053 6002
rect 32566 5989 32633 5995
rect 31744 5962 31800 5974
rect 31744 5928 31750 5962
rect 31784 5961 31800 5962
rect 32857 5961 32913 5973
rect 31784 5945 32251 5961
rect 31784 5928 32201 5945
rect 31744 5912 32201 5928
rect 32185 5911 32201 5912
rect 32235 5911 32251 5945
rect 32185 5904 32251 5911
rect 32303 5946 32873 5961
rect 32303 5912 32319 5946
rect 32353 5927 32873 5946
rect 32907 5927 32913 5961
rect 32353 5912 32913 5927
rect 32303 5902 32370 5912
rect 32857 5911 32913 5912
rect 33019 5873 33053 6001
rect 31597 5861 31643 5873
rect 31597 5685 31603 5861
rect 31637 5685 31643 5861
rect 31597 5673 31643 5685
rect 31715 5861 31761 5873
rect 31715 5685 31721 5861
rect 31755 5685 31761 5861
rect 31715 5673 31761 5685
rect 32017 5861 32063 5873
rect 31720 5379 31754 5673
rect 32017 5485 32023 5861
rect 32057 5485 32063 5861
rect 32017 5473 32063 5485
rect 32135 5861 32181 5873
rect 32135 5485 32141 5861
rect 32175 5485 32181 5861
rect 32135 5473 32181 5485
rect 32253 5861 32299 5873
rect 32253 5485 32259 5861
rect 32293 5485 32299 5861
rect 32253 5473 32299 5485
rect 32371 5861 32417 5873
rect 32371 5485 32377 5861
rect 32411 5485 32417 5861
rect 32371 5473 32417 5485
rect 32489 5861 32535 5873
rect 32489 5485 32495 5861
rect 32529 5485 32535 5861
rect 32895 5861 32941 5873
rect 32895 5685 32901 5861
rect 32935 5685 32941 5861
rect 32895 5673 32941 5685
rect 33013 5861 33059 5873
rect 33013 5685 33019 5861
rect 33053 5685 33059 5861
rect 33013 5673 33059 5685
rect 32489 5473 32535 5485
rect 32377 5379 32411 5473
rect 32901 5379 32934 5673
rect 31720 5347 32934 5379
rect 32086 5323 32492 5347
rect 32086 5200 32198 5323
rect 32372 5200 32492 5323
rect 32086 5156 32492 5200
rect 30438 4058 31119 4061
rect 29018 4008 29174 4014
rect 29962 4046 30008 4058
rect 29410 3791 29520 3792
rect 29408 3790 29786 3791
rect 29408 3785 29787 3790
rect 29402 3695 29412 3785
rect 29496 3695 29787 3785
rect 29408 3691 29787 3695
rect 29410 3690 29520 3691
rect 29710 3690 29787 3691
rect 29732 3541 29786 3690
rect 29962 3670 29968 4046
rect 30002 3670 30008 4046
rect 29962 3658 30008 3670
rect 30080 4046 30126 4058
rect 30080 3670 30086 4046
rect 30120 3670 30126 4046
rect 30080 3658 30126 3670
rect 30198 4046 30244 4058
rect 30198 3670 30204 4046
rect 30238 3697 30244 4046
rect 30315 4046 30361 4058
rect 30315 3870 30321 4046
rect 30355 3870 30361 4046
rect 30315 3863 30361 3870
rect 30433 4046 31119 4058
rect 30433 3870 30439 4046
rect 30473 4033 31119 4046
rect 30473 3870 30479 4033
rect 30723 3953 31119 4033
rect 30315 3858 30364 3863
rect 30433 3858 30479 3870
rect 30321 3697 30364 3858
rect 34254 3835 34367 6543
rect 34652 6510 34740 10089
rect 34778 10046 34896 15675
rect 34778 10019 34898 10046
rect 34651 6486 34741 6510
rect 34651 6418 34662 6486
rect 34728 6418 34741 6486
rect 34651 6406 34741 6418
rect 34413 6387 34558 6400
rect 34413 6296 34428 6387
rect 34538 6296 34558 6387
rect 34413 6287 34558 6296
rect 30691 3831 34367 3835
rect 30238 3670 30364 3697
rect 30198 3658 30364 3670
rect 30204 3654 30364 3658
rect 29842 3638 29915 3643
rect 29836 3574 29846 3638
rect 29912 3626 29922 3638
rect 29912 3620 30077 3626
rect 29912 3586 30027 3620
rect 30061 3586 30077 3620
rect 29912 3574 30077 3586
rect 29842 3570 30077 3574
rect 30129 3620 30195 3626
rect 30129 3586 30145 3620
rect 30179 3586 30195 3620
rect 30129 3541 30195 3586
rect 29732 3533 30195 3541
rect 29732 3501 30196 3533
rect 30288 3517 30364 3654
rect 30688 3717 34367 3831
rect 30284 3457 30294 3517
rect 30356 3457 30366 3517
rect 23962 2982 24331 3030
rect 23962 2952 23976 2982
rect 23962 2935 23972 2952
rect 24264 2879 24330 2982
rect 26093 2943 26099 3078
rect 26166 2943 26172 3078
rect 26093 2931 26172 2943
rect 28890 2879 28956 3158
rect 24262 2799 28956 2879
rect 30688 2364 30853 3717
rect 32100 3476 32545 3482
rect 32100 3276 32112 3476
rect 32533 3276 32545 3476
rect 32100 3270 32268 3276
rect 32258 3202 32268 3270
rect 32400 3270 32545 3276
rect 34779 3347 34898 10019
rect 34779 3341 34902 3347
rect 34779 3275 34797 3341
rect 34890 3275 34902 3341
rect 32400 3202 32410 3270
rect 34779 3269 34902 3275
rect 34779 3267 34898 3269
rect 34956 3259 35046 16594
rect 35093 6405 35176 16769
rect 35218 9539 35298 16870
rect 35342 12681 35434 16988
rect 35755 15884 35897 18508
rect 36951 18518 37151 18524
rect 36951 18484 36963 18518
rect 37139 18484 37151 18518
rect 36951 18437 37151 18484
rect 36751 18431 37151 18437
rect 36607 18397 36763 18431
rect 37139 18397 37151 18431
rect 36607 17634 36664 18397
rect 36751 18391 37151 18397
rect 36751 18313 37151 18319
rect 36751 18279 36763 18313
rect 37139 18279 37151 18313
rect 36751 18273 37151 18279
rect 36751 18195 37151 18201
rect 36751 18161 36763 18195
rect 37139 18161 37151 18195
rect 36751 18155 37151 18161
rect 36751 18077 37151 18083
rect 36751 18043 36763 18077
rect 37139 18043 37151 18077
rect 36751 18037 37151 18043
rect 36751 17964 37151 17970
rect 36751 17930 36763 17964
rect 37139 17930 37277 17964
rect 36751 17924 37151 17930
rect 36751 17846 37151 17852
rect 36751 17812 36763 17846
rect 37139 17812 37151 17846
rect 36751 17806 37151 17812
rect 36751 17728 37151 17734
rect 36751 17694 36763 17728
rect 37139 17694 37151 17728
rect 36751 17688 37151 17694
rect 36507 17624 36664 17634
rect 36567 17544 36664 17624
rect 36751 17610 37151 17616
rect 36751 17576 36763 17610
rect 37139 17576 37151 17610
rect 36751 17570 37151 17576
rect 36507 17534 36664 17544
rect 36607 17256 36664 17534
rect 36751 17492 37151 17498
rect 36751 17458 36763 17492
rect 37139 17458 37151 17492
rect 36751 17452 37151 17458
rect 36751 17374 37151 17380
rect 36751 17340 36763 17374
rect 37139 17340 37151 17374
rect 36751 17334 37151 17340
rect 36751 17256 37151 17262
rect 36607 17222 36763 17256
rect 37139 17222 37151 17256
rect 36607 16665 36664 17222
rect 36751 17216 37151 17222
rect 36751 17137 37151 17143
rect 36751 17103 36763 17137
rect 37139 17103 37151 17137
rect 36751 17097 37151 17103
rect 36751 17019 37151 17025
rect 36751 16985 36763 17019
rect 37139 16985 37151 17019
rect 36751 16979 37151 16985
rect 36751 16901 37151 16907
rect 36751 16867 36763 16901
rect 37139 16867 37151 16901
rect 36751 16861 37151 16867
rect 36751 16783 37151 16789
rect 37235 16783 37277 17930
rect 37337 17786 37404 18838
rect 37437 18771 37522 18783
rect 37437 18700 37450 18771
rect 37513 18700 37522 18771
rect 37437 18691 37522 18700
rect 37914 18039 37961 18838
rect 38084 18039 38284 18044
rect 37914 18038 38284 18039
rect 37914 18005 38096 18038
rect 37337 17752 37354 17786
rect 37388 17752 37404 17786
rect 37337 17736 37404 17752
rect 37725 17804 37810 17816
rect 37725 17736 37733 17804
rect 37798 17736 37810 17804
rect 37725 17724 37810 17736
rect 37440 17686 37525 17698
rect 37440 17616 37450 17686
rect 37512 17616 37525 17686
rect 37440 17606 37525 17616
rect 37914 17567 37961 18005
rect 38084 18004 38096 18005
rect 38272 18004 38284 18038
rect 38084 17998 38284 18004
rect 38084 17920 38284 17926
rect 38084 17886 38096 17920
rect 38272 17886 38703 17920
rect 38084 17852 38284 17886
rect 38084 17846 38484 17852
rect 38084 17812 38096 17846
rect 38472 17812 38484 17846
rect 38084 17806 38484 17812
rect 38084 17728 38484 17734
rect 38084 17694 38096 17728
rect 38472 17694 38484 17728
rect 38084 17688 38484 17694
rect 38084 17610 38484 17616
rect 38557 17610 38623 17625
rect 38084 17576 38096 17610
rect 38472 17609 38623 17610
rect 38472 17576 38573 17609
rect 38084 17570 38484 17576
rect 38557 17575 38573 17576
rect 38607 17575 38623 17609
rect 37914 17551 38024 17567
rect 38557 17559 38623 17575
rect 38651 17622 38703 17886
rect 38651 17610 38781 17622
rect 37914 17517 37974 17551
rect 38008 17517 38024 17551
rect 37914 17501 38024 17517
rect 38651 17544 38725 17610
rect 38777 17544 38781 17610
rect 38651 17530 38781 17544
rect 38084 17492 38484 17498
rect 38084 17458 38096 17492
rect 38472 17458 38484 17492
rect 38084 17452 38484 17458
rect 37564 17445 37636 17451
rect 37564 17386 37570 17445
rect 37630 17386 37636 17445
rect 37567 17382 37634 17386
rect 37570 17376 37630 17382
rect 38084 17374 38484 17380
rect 38084 17340 38096 17374
rect 38472 17340 38484 17374
rect 38084 17334 38484 17340
rect 38084 17296 38284 17334
rect 38651 17296 38703 17530
rect 38084 17262 38096 17296
rect 38272 17262 38703 17296
rect 38084 17256 38284 17262
rect 37913 17178 37960 17179
rect 38084 17178 38284 17184
rect 37913 17144 38096 17178
rect 38272 17144 38284 17178
rect 36751 16749 36763 16783
rect 37139 16749 37363 16783
rect 36751 16743 37151 16749
rect 36951 16665 37151 16670
rect 36607 16664 37151 16665
rect 36607 16630 36963 16664
rect 37139 16630 37151 16664
rect 36607 16628 37151 16630
rect 36951 16624 37151 16628
rect 36951 16546 37151 16552
rect 36951 16512 36963 16546
rect 37139 16512 37151 16546
rect 36951 16506 37151 16512
rect 37297 16476 37363 16749
rect 37297 16442 37313 16476
rect 37347 16442 37363 16476
rect 36951 16428 37151 16434
rect 36951 16394 36963 16428
rect 37139 16394 37151 16428
rect 37297 16426 37363 16442
rect 36951 16388 37151 16394
rect 36951 16310 37151 16316
rect 37913 16310 37960 17144
rect 38084 17138 38284 17144
rect 36951 16276 36963 16310
rect 37139 16279 37960 16310
rect 37139 16278 38057 16279
rect 39202 16278 39594 16402
rect 37139 16276 39594 16278
rect 36951 16275 39594 16276
rect 36951 16270 37151 16275
rect 37505 16129 39594 16275
rect 37962 16128 39594 16129
rect 39202 16033 39594 16128
rect 35755 15873 37641 15884
rect 35753 15871 37641 15873
rect 35753 15814 37565 15871
rect 37633 15814 37641 15871
rect 35753 15803 37641 15814
rect 36951 15729 37151 15734
rect 36951 15728 37961 15729
rect 36951 15694 36963 15728
rect 37139 15694 37961 15728
rect 36951 15688 37151 15694
rect 36951 15610 37151 15616
rect 36951 15576 36963 15610
rect 37139 15576 37151 15610
rect 36951 15570 37151 15576
rect 36951 15492 37151 15498
rect 36951 15458 36963 15492
rect 37139 15458 37151 15492
rect 36951 15452 37151 15458
rect 36951 15374 37151 15380
rect 36951 15340 36963 15374
rect 37139 15340 37151 15374
rect 36951 15293 37151 15340
rect 36751 15287 37151 15293
rect 36607 15253 36763 15287
rect 37139 15253 37151 15287
rect 36607 14490 36664 15253
rect 36751 15247 37151 15253
rect 36751 15169 37151 15175
rect 36751 15135 36763 15169
rect 37139 15135 37151 15169
rect 36751 15129 37151 15135
rect 36751 15051 37151 15057
rect 36751 15017 36763 15051
rect 37139 15017 37151 15051
rect 36751 15011 37151 15017
rect 36751 14933 37151 14939
rect 36751 14899 36763 14933
rect 37139 14899 37151 14933
rect 36751 14893 37151 14899
rect 36751 14820 37151 14826
rect 36751 14786 36763 14820
rect 37139 14786 37277 14820
rect 36751 14780 37151 14786
rect 36751 14702 37151 14708
rect 36751 14668 36763 14702
rect 37139 14668 37151 14702
rect 36751 14662 37151 14668
rect 36751 14584 37151 14590
rect 36751 14550 36763 14584
rect 37139 14550 37151 14584
rect 36751 14544 37151 14550
rect 36507 14480 36664 14490
rect 36567 14400 36664 14480
rect 36751 14466 37151 14472
rect 36751 14432 36763 14466
rect 37139 14432 37151 14466
rect 36751 14426 37151 14432
rect 36507 14390 36664 14400
rect 36607 14112 36664 14390
rect 36751 14348 37151 14354
rect 36751 14314 36763 14348
rect 37139 14314 37151 14348
rect 36751 14308 37151 14314
rect 36751 14230 37151 14236
rect 36751 14196 36763 14230
rect 37139 14196 37151 14230
rect 36751 14190 37151 14196
rect 36751 14112 37151 14118
rect 36607 14078 36763 14112
rect 37139 14078 37151 14112
rect 36607 13521 36664 14078
rect 36751 14072 37151 14078
rect 36751 13993 37151 13999
rect 36751 13959 36763 13993
rect 37139 13959 37151 13993
rect 36751 13953 37151 13959
rect 36751 13875 37151 13881
rect 36751 13841 36763 13875
rect 37139 13841 37151 13875
rect 36751 13835 37151 13841
rect 36751 13757 37151 13763
rect 36751 13723 36763 13757
rect 37139 13723 37151 13757
rect 36751 13717 37151 13723
rect 36751 13639 37151 13645
rect 37235 13639 37277 14786
rect 37337 14642 37404 15694
rect 37437 15627 37522 15639
rect 37437 15556 37450 15627
rect 37513 15556 37522 15627
rect 37437 15547 37522 15556
rect 37914 14895 37961 15694
rect 38084 14895 38284 14900
rect 37914 14894 38284 14895
rect 37914 14861 38096 14894
rect 37337 14608 37354 14642
rect 37388 14608 37404 14642
rect 37337 14592 37404 14608
rect 37725 14660 37810 14672
rect 37725 14592 37733 14660
rect 37798 14592 37810 14660
rect 37725 14580 37810 14592
rect 37440 14542 37525 14554
rect 37440 14472 37450 14542
rect 37512 14472 37525 14542
rect 37440 14462 37525 14472
rect 37914 14423 37961 14861
rect 38084 14860 38096 14861
rect 38272 14860 38284 14894
rect 38084 14854 38284 14860
rect 38084 14776 38284 14782
rect 38084 14742 38096 14776
rect 38272 14742 38703 14776
rect 38084 14708 38284 14742
rect 38084 14702 38484 14708
rect 38084 14668 38096 14702
rect 38472 14668 38484 14702
rect 38084 14662 38484 14668
rect 38084 14584 38484 14590
rect 38084 14550 38096 14584
rect 38472 14550 38484 14584
rect 38084 14544 38484 14550
rect 38084 14466 38484 14472
rect 38557 14466 38623 14481
rect 38084 14432 38096 14466
rect 38472 14465 38623 14466
rect 38472 14432 38573 14465
rect 38084 14426 38484 14432
rect 38557 14431 38573 14432
rect 38607 14431 38623 14465
rect 37914 14407 38024 14423
rect 38557 14415 38623 14431
rect 38651 14478 38703 14742
rect 38651 14466 38781 14478
rect 37914 14373 37974 14407
rect 38008 14373 38024 14407
rect 37914 14357 38024 14373
rect 38651 14400 38725 14466
rect 38777 14400 38781 14466
rect 38651 14386 38781 14400
rect 38084 14348 38484 14354
rect 38084 14314 38096 14348
rect 38472 14314 38484 14348
rect 38084 14308 38484 14314
rect 37564 14301 37636 14307
rect 37564 14242 37570 14301
rect 37630 14242 37636 14301
rect 37567 14238 37634 14242
rect 37570 14232 37630 14238
rect 38084 14230 38484 14236
rect 38084 14196 38096 14230
rect 38472 14196 38484 14230
rect 38084 14190 38484 14196
rect 38084 14152 38284 14190
rect 38651 14152 38703 14386
rect 38084 14118 38096 14152
rect 38272 14118 38703 14152
rect 38084 14112 38284 14118
rect 37913 14034 37960 14035
rect 38084 14034 38284 14040
rect 37913 14000 38096 14034
rect 38272 14000 38284 14034
rect 36751 13605 36763 13639
rect 37139 13605 37363 13639
rect 36751 13599 37151 13605
rect 36951 13521 37151 13526
rect 36607 13520 37151 13521
rect 36607 13486 36963 13520
rect 37139 13486 37151 13520
rect 36607 13484 37151 13486
rect 36951 13480 37151 13484
rect 36951 13402 37151 13408
rect 36951 13368 36963 13402
rect 37139 13368 37151 13402
rect 36951 13362 37151 13368
rect 37297 13332 37363 13605
rect 37297 13298 37313 13332
rect 37347 13298 37363 13332
rect 36951 13284 37151 13290
rect 36951 13250 36963 13284
rect 37139 13250 37151 13284
rect 37297 13282 37363 13298
rect 36951 13244 37151 13250
rect 36951 13166 37151 13172
rect 37913 13166 37960 14000
rect 38084 13994 38284 14000
rect 36951 13132 36963 13166
rect 37139 13134 37960 13166
rect 39201 13134 39593 13258
rect 37139 13132 39593 13134
rect 36951 13131 39593 13132
rect 36951 13126 37151 13131
rect 37505 12985 39593 13131
rect 37641 12984 39593 12985
rect 39201 12889 39593 12984
rect 35342 12669 37646 12681
rect 35342 12612 37569 12669
rect 37637 12612 37646 12669
rect 35342 12600 37646 12612
rect 37729 12669 37813 12684
rect 37729 12612 37737 12669
rect 37805 12612 37813 12669
rect 37729 12610 37813 12612
rect 37737 12602 37805 12610
rect 36955 12527 37155 12532
rect 36955 12526 37965 12527
rect 36955 12492 36967 12526
rect 37143 12492 37965 12526
rect 36955 12486 37155 12492
rect 36955 12408 37155 12414
rect 36955 12374 36967 12408
rect 37143 12374 37155 12408
rect 36955 12368 37155 12374
rect 36955 12290 37155 12296
rect 36955 12256 36967 12290
rect 37143 12256 37155 12290
rect 36955 12250 37155 12256
rect 36955 12172 37155 12178
rect 36955 12138 36967 12172
rect 37143 12138 37155 12172
rect 36955 12091 37155 12138
rect 36755 12085 37155 12091
rect 36611 12051 36767 12085
rect 37143 12051 37155 12085
rect 36611 11288 36668 12051
rect 36755 12045 37155 12051
rect 36755 11967 37155 11973
rect 36755 11933 36767 11967
rect 37143 11933 37155 11967
rect 36755 11927 37155 11933
rect 36755 11849 37155 11855
rect 36755 11815 36767 11849
rect 37143 11815 37155 11849
rect 36755 11809 37155 11815
rect 36755 11731 37155 11737
rect 36755 11697 36767 11731
rect 37143 11697 37155 11731
rect 36755 11691 37155 11697
rect 36755 11618 37155 11624
rect 36755 11584 36767 11618
rect 37143 11584 37281 11618
rect 36755 11578 37155 11584
rect 36755 11500 37155 11506
rect 36755 11466 36767 11500
rect 37143 11466 37155 11500
rect 36755 11460 37155 11466
rect 36755 11382 37155 11388
rect 36755 11348 36767 11382
rect 37143 11348 37155 11382
rect 36755 11342 37155 11348
rect 36511 11278 36668 11288
rect 36571 11198 36668 11278
rect 36755 11264 37155 11270
rect 36755 11230 36767 11264
rect 37143 11230 37155 11264
rect 36755 11224 37155 11230
rect 36511 11188 36668 11198
rect 36611 10910 36668 11188
rect 36755 11146 37155 11152
rect 36755 11112 36767 11146
rect 37143 11112 37155 11146
rect 36755 11106 37155 11112
rect 36755 11028 37155 11034
rect 36755 10994 36767 11028
rect 37143 10994 37155 11028
rect 36755 10988 37155 10994
rect 36755 10910 37155 10916
rect 36611 10876 36767 10910
rect 37143 10876 37155 10910
rect 36611 10319 36668 10876
rect 36755 10870 37155 10876
rect 36755 10791 37155 10797
rect 36755 10757 36767 10791
rect 37143 10757 37155 10791
rect 36755 10751 37155 10757
rect 36755 10673 37155 10679
rect 36755 10639 36767 10673
rect 37143 10639 37155 10673
rect 36755 10633 37155 10639
rect 36755 10555 37155 10561
rect 36755 10521 36767 10555
rect 37143 10521 37155 10555
rect 36755 10515 37155 10521
rect 36755 10437 37155 10443
rect 37239 10437 37281 11584
rect 37341 11440 37408 12492
rect 37441 12425 37526 12437
rect 37441 12354 37454 12425
rect 37517 12354 37526 12425
rect 37441 12345 37526 12354
rect 37918 11693 37965 12492
rect 38088 11693 38288 11698
rect 37918 11692 38288 11693
rect 37918 11659 38100 11692
rect 37341 11406 37358 11440
rect 37392 11406 37408 11440
rect 37341 11390 37408 11406
rect 37729 11458 37814 11470
rect 37729 11390 37737 11458
rect 37802 11390 37814 11458
rect 37729 11378 37814 11390
rect 37444 11340 37529 11352
rect 37444 11270 37454 11340
rect 37516 11270 37529 11340
rect 37444 11260 37529 11270
rect 37918 11221 37965 11659
rect 38088 11658 38100 11659
rect 38276 11658 38288 11692
rect 38088 11652 38288 11658
rect 38088 11574 38288 11580
rect 38088 11540 38100 11574
rect 38276 11540 38707 11574
rect 38088 11506 38288 11540
rect 38088 11500 38488 11506
rect 38088 11466 38100 11500
rect 38476 11466 38488 11500
rect 38088 11460 38488 11466
rect 38088 11382 38488 11388
rect 38088 11348 38100 11382
rect 38476 11348 38488 11382
rect 38088 11342 38488 11348
rect 38088 11264 38488 11270
rect 38561 11264 38627 11279
rect 38088 11230 38100 11264
rect 38476 11263 38627 11264
rect 38476 11230 38577 11263
rect 38088 11224 38488 11230
rect 38561 11229 38577 11230
rect 38611 11229 38627 11263
rect 37918 11205 38028 11221
rect 38561 11213 38627 11229
rect 38655 11276 38707 11540
rect 38655 11264 38785 11276
rect 37918 11171 37978 11205
rect 38012 11171 38028 11205
rect 37918 11155 38028 11171
rect 38655 11198 38729 11264
rect 38781 11198 38785 11264
rect 38655 11184 38785 11198
rect 38088 11146 38488 11152
rect 38088 11112 38100 11146
rect 38476 11112 38488 11146
rect 38088 11106 38488 11112
rect 37568 11099 37640 11105
rect 37568 11040 37574 11099
rect 37634 11040 37640 11099
rect 37571 11036 37638 11040
rect 37574 11030 37634 11036
rect 38088 11028 38488 11034
rect 38088 10994 38100 11028
rect 38476 10994 38488 11028
rect 38088 10988 38488 10994
rect 38088 10950 38288 10988
rect 38655 10950 38707 11184
rect 38088 10916 38100 10950
rect 38276 10916 38707 10950
rect 38088 10910 38288 10916
rect 37917 10832 37964 10833
rect 38088 10832 38288 10838
rect 37917 10798 38100 10832
rect 38276 10798 38288 10832
rect 36755 10403 36767 10437
rect 37143 10403 37367 10437
rect 36755 10397 37155 10403
rect 36955 10319 37155 10324
rect 36611 10318 37155 10319
rect 36611 10284 36967 10318
rect 37143 10284 37155 10318
rect 36611 10282 37155 10284
rect 36955 10278 37155 10282
rect 36955 10200 37155 10206
rect 36955 10166 36967 10200
rect 37143 10166 37155 10200
rect 36955 10160 37155 10166
rect 37301 10130 37367 10403
rect 37301 10096 37317 10130
rect 37351 10096 37367 10130
rect 36955 10082 37155 10088
rect 36955 10048 36967 10082
rect 37143 10048 37155 10082
rect 37301 10080 37367 10096
rect 36955 10042 37155 10048
rect 36955 9964 37155 9970
rect 37917 9964 37964 10798
rect 38088 10792 38288 10798
rect 36955 9930 36967 9964
rect 37143 9934 37964 9964
rect 37143 9933 38033 9934
rect 39204 9933 39596 10057
rect 37143 9930 39596 9933
rect 36955 9929 39596 9930
rect 36955 9924 37155 9929
rect 37509 9784 39596 9929
rect 37509 9783 37655 9784
rect 37964 9783 39596 9784
rect 39204 9688 39596 9783
rect 35218 9538 37601 9539
rect 35218 9525 37645 9538
rect 35218 9468 37569 9525
rect 37637 9468 37645 9525
rect 35218 9466 37645 9468
rect 35218 9458 37637 9466
rect 36955 9383 37155 9388
rect 36955 9382 37965 9383
rect 36955 9348 36967 9382
rect 37143 9348 37965 9382
rect 36955 9342 37155 9348
rect 36955 9264 37155 9270
rect 36955 9230 36967 9264
rect 37143 9230 37155 9264
rect 36955 9224 37155 9230
rect 36955 9146 37155 9152
rect 36955 9112 36967 9146
rect 37143 9112 37155 9146
rect 36955 9106 37155 9112
rect 36955 9028 37155 9034
rect 36955 8994 36967 9028
rect 37143 8994 37155 9028
rect 36955 8947 37155 8994
rect 36755 8941 37155 8947
rect 36611 8907 36767 8941
rect 37143 8907 37155 8941
rect 36611 8144 36668 8907
rect 36755 8901 37155 8907
rect 36755 8823 37155 8829
rect 36755 8789 36767 8823
rect 37143 8789 37155 8823
rect 36755 8783 37155 8789
rect 36755 8705 37155 8711
rect 36755 8671 36767 8705
rect 37143 8671 37155 8705
rect 36755 8665 37155 8671
rect 36755 8587 37155 8593
rect 36755 8553 36767 8587
rect 37143 8553 37155 8587
rect 36755 8547 37155 8553
rect 36755 8474 37155 8480
rect 36755 8440 36767 8474
rect 37143 8440 37281 8474
rect 36755 8434 37155 8440
rect 36755 8356 37155 8362
rect 36755 8322 36767 8356
rect 37143 8322 37155 8356
rect 36755 8316 37155 8322
rect 36755 8238 37155 8244
rect 36755 8204 36767 8238
rect 37143 8204 37155 8238
rect 36755 8198 37155 8204
rect 36511 8134 36668 8144
rect 36571 8054 36668 8134
rect 36755 8120 37155 8126
rect 36755 8086 36767 8120
rect 37143 8086 37155 8120
rect 36755 8080 37155 8086
rect 36511 8044 36668 8054
rect 36611 7766 36668 8044
rect 36755 8002 37155 8008
rect 36755 7968 36767 8002
rect 37143 7968 37155 8002
rect 36755 7962 37155 7968
rect 36755 7884 37155 7890
rect 36755 7850 36767 7884
rect 37143 7850 37155 7884
rect 36755 7844 37155 7850
rect 36755 7766 37155 7772
rect 36611 7732 36767 7766
rect 37143 7732 37155 7766
rect 36611 7175 36668 7732
rect 36755 7726 37155 7732
rect 36755 7647 37155 7653
rect 36755 7613 36767 7647
rect 37143 7613 37155 7647
rect 36755 7607 37155 7613
rect 36755 7529 37155 7535
rect 36755 7495 36767 7529
rect 37143 7495 37155 7529
rect 36755 7489 37155 7495
rect 36755 7411 37155 7417
rect 36755 7377 36767 7411
rect 37143 7377 37155 7411
rect 36755 7371 37155 7377
rect 36755 7293 37155 7299
rect 37239 7293 37281 8440
rect 37341 8296 37408 9348
rect 37441 9281 37526 9293
rect 37441 9210 37454 9281
rect 37517 9210 37526 9281
rect 37441 9201 37526 9210
rect 37918 8549 37965 9348
rect 38088 8549 38288 8554
rect 37918 8548 38288 8549
rect 37918 8515 38100 8548
rect 37341 8262 37358 8296
rect 37392 8262 37408 8296
rect 37341 8246 37408 8262
rect 37729 8314 37814 8326
rect 37729 8246 37737 8314
rect 37802 8246 37814 8314
rect 37729 8234 37814 8246
rect 37444 8196 37529 8208
rect 37444 8126 37454 8196
rect 37516 8126 37529 8196
rect 37444 8116 37529 8126
rect 37918 8077 37965 8515
rect 38088 8514 38100 8515
rect 38276 8514 38288 8548
rect 38088 8508 38288 8514
rect 38088 8430 38288 8436
rect 38088 8396 38100 8430
rect 38276 8396 38707 8430
rect 38088 8362 38288 8396
rect 38088 8356 38488 8362
rect 38088 8322 38100 8356
rect 38476 8322 38488 8356
rect 38088 8316 38488 8322
rect 38088 8238 38488 8244
rect 38088 8204 38100 8238
rect 38476 8204 38488 8238
rect 38088 8198 38488 8204
rect 38088 8120 38488 8126
rect 38561 8120 38627 8135
rect 38088 8086 38100 8120
rect 38476 8119 38627 8120
rect 38476 8086 38577 8119
rect 38088 8080 38488 8086
rect 38561 8085 38577 8086
rect 38611 8085 38627 8119
rect 37918 8061 38028 8077
rect 38561 8069 38627 8085
rect 38655 8132 38707 8396
rect 38655 8120 38785 8132
rect 37918 8027 37978 8061
rect 38012 8027 38028 8061
rect 37918 8011 38028 8027
rect 38655 8054 38729 8120
rect 38781 8054 38785 8120
rect 38655 8040 38785 8054
rect 38088 8002 38488 8008
rect 38088 7968 38100 8002
rect 38476 7968 38488 8002
rect 38088 7962 38488 7968
rect 37568 7955 37640 7961
rect 37568 7896 37574 7955
rect 37634 7896 37640 7955
rect 37571 7892 37638 7896
rect 37574 7886 37634 7892
rect 38088 7884 38488 7890
rect 38088 7850 38100 7884
rect 38476 7850 38488 7884
rect 38088 7844 38488 7850
rect 38088 7806 38288 7844
rect 38655 7806 38707 8040
rect 38088 7772 38100 7806
rect 38276 7772 38707 7806
rect 38088 7766 38288 7772
rect 37917 7688 37964 7689
rect 38088 7688 38288 7694
rect 37917 7654 38100 7688
rect 38276 7654 38288 7688
rect 36755 7259 36767 7293
rect 37143 7259 37367 7293
rect 36755 7253 37155 7259
rect 36955 7175 37155 7180
rect 36611 7174 37155 7175
rect 36611 7140 36967 7174
rect 37143 7140 37155 7174
rect 36611 7138 37155 7140
rect 36955 7134 37155 7138
rect 36955 7056 37155 7062
rect 36955 7022 36967 7056
rect 37143 7022 37155 7056
rect 36955 7016 37155 7022
rect 37301 6986 37367 7259
rect 37301 6952 37317 6986
rect 37351 6952 37367 6986
rect 36955 6938 37155 6944
rect 36955 6904 36967 6938
rect 37143 6904 37155 6938
rect 37301 6936 37367 6952
rect 36955 6898 37155 6904
rect 36955 6820 37155 6826
rect 37917 6820 37964 7654
rect 38088 7648 38288 7654
rect 36955 6786 36967 6820
rect 37143 6789 37964 6820
rect 37143 6788 38057 6789
rect 39204 6788 39596 6912
rect 37143 6786 39596 6788
rect 36955 6785 39596 6786
rect 36955 6780 37155 6785
rect 37509 6639 39596 6785
rect 37964 6638 39596 6639
rect 39204 6543 39596 6638
rect 37557 6405 37641 6406
rect 35093 6393 37643 6405
rect 35093 6336 37565 6393
rect 37633 6336 37643 6393
rect 35093 6326 37643 6336
rect 37725 6393 37809 6408
rect 37725 6336 37733 6393
rect 37801 6336 37809 6393
rect 37725 6334 37809 6336
rect 37733 6326 37801 6334
rect 36951 6251 37151 6256
rect 36951 6250 37961 6251
rect 36951 6216 36963 6250
rect 37139 6216 37961 6250
rect 36951 6210 37151 6216
rect 36951 6132 37151 6138
rect 36951 6098 36963 6132
rect 37139 6098 37151 6132
rect 36951 6092 37151 6098
rect 36951 6014 37151 6020
rect 36951 5980 36963 6014
rect 37139 5980 37151 6014
rect 36951 5974 37151 5980
rect 36951 5896 37151 5902
rect 36951 5862 36963 5896
rect 37139 5862 37151 5896
rect 36951 5815 37151 5862
rect 36751 5809 37151 5815
rect 36607 5775 36763 5809
rect 37139 5775 37151 5809
rect 36607 5012 36664 5775
rect 36751 5769 37151 5775
rect 36751 5691 37151 5697
rect 36751 5657 36763 5691
rect 37139 5657 37151 5691
rect 36751 5651 37151 5657
rect 36751 5573 37151 5579
rect 36751 5539 36763 5573
rect 37139 5539 37151 5573
rect 36751 5533 37151 5539
rect 36751 5455 37151 5461
rect 36751 5421 36763 5455
rect 37139 5421 37151 5455
rect 36751 5415 37151 5421
rect 36751 5342 37151 5348
rect 36751 5308 36763 5342
rect 37139 5308 37277 5342
rect 36751 5302 37151 5308
rect 36751 5224 37151 5230
rect 36751 5190 36763 5224
rect 37139 5190 37151 5224
rect 36751 5184 37151 5190
rect 36751 5106 37151 5112
rect 36751 5072 36763 5106
rect 37139 5072 37151 5106
rect 36751 5066 37151 5072
rect 36507 5002 36664 5012
rect 36567 4922 36664 5002
rect 36751 4988 37151 4994
rect 36751 4954 36763 4988
rect 37139 4954 37151 4988
rect 36751 4948 37151 4954
rect 36507 4912 36664 4922
rect 36607 4634 36664 4912
rect 36751 4870 37151 4876
rect 36751 4836 36763 4870
rect 37139 4836 37151 4870
rect 36751 4830 37151 4836
rect 36751 4752 37151 4758
rect 36751 4718 36763 4752
rect 37139 4718 37151 4752
rect 36751 4712 37151 4718
rect 36751 4634 37151 4640
rect 36607 4600 36763 4634
rect 37139 4600 37151 4634
rect 36607 4043 36664 4600
rect 36751 4594 37151 4600
rect 36751 4515 37151 4521
rect 36751 4481 36763 4515
rect 37139 4481 37151 4515
rect 36751 4475 37151 4481
rect 36751 4397 37151 4403
rect 36751 4363 36763 4397
rect 37139 4363 37151 4397
rect 36751 4357 37151 4363
rect 36751 4279 37151 4285
rect 36751 4245 36763 4279
rect 37139 4245 37151 4279
rect 36751 4239 37151 4245
rect 36751 4161 37151 4167
rect 37235 4161 37277 5308
rect 37337 5164 37404 6216
rect 37437 6149 37522 6161
rect 37437 6078 37450 6149
rect 37513 6078 37522 6149
rect 37437 6069 37522 6078
rect 37914 5417 37961 6216
rect 38084 5417 38284 5422
rect 37914 5416 38284 5417
rect 37914 5383 38096 5416
rect 37337 5130 37354 5164
rect 37388 5130 37404 5164
rect 37337 5114 37404 5130
rect 37725 5182 37810 5194
rect 37725 5114 37733 5182
rect 37798 5114 37810 5182
rect 37725 5102 37810 5114
rect 37440 5064 37525 5076
rect 37440 4994 37450 5064
rect 37512 4994 37525 5064
rect 37440 4984 37525 4994
rect 37914 4945 37961 5383
rect 38084 5382 38096 5383
rect 38272 5382 38284 5416
rect 38084 5376 38284 5382
rect 38084 5298 38284 5304
rect 38084 5264 38096 5298
rect 38272 5264 38703 5298
rect 38084 5230 38284 5264
rect 38084 5224 38484 5230
rect 38084 5190 38096 5224
rect 38472 5190 38484 5224
rect 38084 5184 38484 5190
rect 38084 5106 38484 5112
rect 38084 5072 38096 5106
rect 38472 5072 38484 5106
rect 38084 5066 38484 5072
rect 38084 4988 38484 4994
rect 38557 4988 38623 5003
rect 38084 4954 38096 4988
rect 38472 4987 38623 4988
rect 38472 4954 38573 4987
rect 38084 4948 38484 4954
rect 38557 4953 38573 4954
rect 38607 4953 38623 4987
rect 37914 4929 38024 4945
rect 38557 4937 38623 4953
rect 38651 5000 38703 5264
rect 38651 4988 38781 5000
rect 37914 4895 37974 4929
rect 38008 4895 38024 4929
rect 37914 4879 38024 4895
rect 38651 4922 38725 4988
rect 38777 4922 38781 4988
rect 38651 4908 38781 4922
rect 38084 4870 38484 4876
rect 38084 4836 38096 4870
rect 38472 4836 38484 4870
rect 38084 4830 38484 4836
rect 37564 4823 37636 4829
rect 37564 4764 37570 4823
rect 37630 4764 37636 4823
rect 37567 4760 37634 4764
rect 37570 4754 37630 4760
rect 38084 4752 38484 4758
rect 38084 4718 38096 4752
rect 38472 4718 38484 4752
rect 38084 4712 38484 4718
rect 38084 4674 38284 4712
rect 38651 4674 38703 4908
rect 38084 4640 38096 4674
rect 38272 4640 38703 4674
rect 38084 4634 38284 4640
rect 37913 4556 37960 4557
rect 38084 4556 38284 4562
rect 37913 4522 38096 4556
rect 38272 4522 38284 4556
rect 36751 4127 36763 4161
rect 37139 4127 37363 4161
rect 36751 4121 37151 4127
rect 36951 4043 37151 4048
rect 36607 4042 37151 4043
rect 36607 4008 36963 4042
rect 37139 4008 37151 4042
rect 36607 4006 37151 4008
rect 36951 4002 37151 4006
rect 36951 3924 37151 3930
rect 36951 3890 36963 3924
rect 37139 3890 37151 3924
rect 36951 3884 37151 3890
rect 37297 3854 37363 4127
rect 37297 3820 37313 3854
rect 37347 3820 37363 3854
rect 36951 3806 37151 3812
rect 36951 3772 36963 3806
rect 37139 3772 37151 3806
rect 37297 3804 37363 3820
rect 36951 3766 37151 3772
rect 36951 3688 37151 3694
rect 37913 3688 37960 4522
rect 38084 4516 38284 4522
rect 36951 3654 36963 3688
rect 37139 3658 37960 3688
rect 39200 3658 39592 3784
rect 37139 3654 39592 3658
rect 36951 3653 39592 3654
rect 36951 3648 37151 3653
rect 37505 3508 39592 3653
rect 39200 3413 39592 3508
rect 37557 3259 37641 3262
rect 34956 3249 37643 3259
rect 32268 3162 32400 3202
rect 34956 3192 37565 3249
rect 37633 3192 37643 3249
rect 34956 3182 37643 3192
rect 37725 3249 37809 3259
rect 37725 3192 37733 3249
rect 37801 3192 37809 3249
rect 37725 3190 37809 3192
rect 37733 3182 37801 3190
rect 34956 3181 35046 3182
rect 32267 3096 32400 3162
rect 36951 3107 37151 3112
rect 36951 3106 37961 3107
rect 31596 3053 33069 3096
rect 36951 3072 36963 3106
rect 37139 3072 37961 3106
rect 36951 3066 37151 3072
rect 31596 2750 31630 3053
rect 31962 2950 31996 3053
rect 32198 2950 32232 3053
rect 32434 2950 32468 3053
rect 32670 2950 32704 3053
rect 31956 2938 32002 2950
rect 31472 2738 31518 2750
rect 31472 2562 31478 2738
rect 31512 2562 31518 2738
rect 31472 2550 31518 2562
rect 31590 2738 31636 2750
rect 31590 2562 31596 2738
rect 31630 2562 31636 2738
rect 31590 2550 31636 2562
rect 31708 2738 31754 2750
rect 31708 2562 31714 2738
rect 31748 2562 31754 2738
rect 31708 2550 31754 2562
rect 31826 2738 31872 2750
rect 31956 2738 31962 2938
rect 31826 2562 31832 2738
rect 31866 2562 31962 2738
rect 31996 2562 32002 2938
rect 31826 2550 31872 2562
rect 31956 2550 32002 2562
rect 32074 2938 32120 2950
rect 32074 2562 32080 2938
rect 32114 2562 32120 2938
rect 32074 2550 32120 2562
rect 32192 2938 32238 2950
rect 32192 2562 32198 2938
rect 32232 2562 32238 2938
rect 32192 2550 32238 2562
rect 32310 2938 32356 2950
rect 32310 2562 32316 2938
rect 32350 2562 32356 2938
rect 32310 2550 32356 2562
rect 32428 2938 32474 2950
rect 32428 2562 32434 2938
rect 32468 2562 32474 2938
rect 32428 2550 32474 2562
rect 32546 2938 32592 2950
rect 32546 2562 32552 2938
rect 32586 2562 32592 2938
rect 32546 2550 32592 2562
rect 32664 2938 32710 2950
rect 32664 2562 32670 2938
rect 32704 2738 32710 2938
rect 33035 2750 33069 3053
rect 33576 2973 33712 2993
rect 33576 2911 33612 2973
rect 33672 2911 33712 2973
rect 36951 2988 37151 2994
rect 36951 2954 36963 2988
rect 37139 2954 37151 2988
rect 36951 2948 37151 2954
rect 33576 2883 33712 2911
rect 33272 2853 34249 2883
rect 32793 2738 32839 2750
rect 32704 2562 32799 2738
rect 32833 2562 32839 2738
rect 32664 2550 32710 2562
rect 32793 2550 32839 2562
rect 32911 2738 32957 2750
rect 32911 2562 32917 2738
rect 32951 2562 32957 2738
rect 32911 2550 32957 2562
rect 33029 2738 33075 2750
rect 33029 2562 33035 2738
rect 33069 2562 33075 2738
rect 33029 2550 33075 2562
rect 33147 2738 33193 2750
rect 33272 2747 33304 2853
rect 33508 2747 33540 2853
rect 33744 2747 33776 2853
rect 33980 2747 34012 2853
rect 34215 2747 34249 2853
rect 36951 2870 37151 2876
rect 36951 2836 36963 2870
rect 37139 2836 37151 2870
rect 36951 2830 37151 2836
rect 36951 2752 37151 2758
rect 33147 2562 33153 2738
rect 33187 2562 33193 2738
rect 33147 2550 33193 2562
rect 33265 2735 33311 2747
rect 33265 2559 33271 2735
rect 33305 2559 33311 2735
rect 31478 2516 31512 2550
rect 32080 2516 32114 2550
rect 32316 2516 32350 2550
rect 31478 2481 31637 2516
rect 32080 2481 32350 2516
rect 32917 2516 32951 2550
rect 33153 2516 33187 2550
rect 33265 2547 33311 2559
rect 33383 2735 33429 2747
rect 33383 2559 33389 2735
rect 33423 2559 33429 2735
rect 33383 2547 33429 2559
rect 33501 2735 33547 2747
rect 33501 2559 33507 2735
rect 33541 2559 33547 2735
rect 33501 2547 33547 2559
rect 33619 2735 33665 2747
rect 33619 2559 33625 2735
rect 33659 2559 33665 2735
rect 33619 2547 33665 2559
rect 33737 2735 33783 2747
rect 33737 2559 33743 2735
rect 33777 2559 33783 2735
rect 33737 2547 33783 2559
rect 33855 2735 33901 2747
rect 33855 2559 33861 2735
rect 33895 2559 33901 2735
rect 33855 2547 33901 2559
rect 33973 2735 34019 2747
rect 33973 2559 33979 2735
rect 34013 2559 34019 2735
rect 33973 2547 34019 2559
rect 34091 2735 34137 2747
rect 34091 2559 34097 2735
rect 34131 2559 34137 2735
rect 34091 2547 34137 2559
rect 34209 2735 34255 2747
rect 34209 2559 34215 2735
rect 34249 2559 34255 2735
rect 34209 2547 34255 2559
rect 34327 2735 34373 2747
rect 34327 2559 34333 2735
rect 34367 2559 34373 2735
rect 36951 2718 36963 2752
rect 37139 2718 37151 2752
rect 36951 2671 37151 2718
rect 36751 2665 37151 2671
rect 34327 2547 34373 2559
rect 36607 2631 36763 2665
rect 37139 2631 37151 2665
rect 32917 2481 33187 2516
rect 22938 2213 30853 2364
rect 31446 2400 31543 2406
rect 31446 2329 31458 2400
rect 31531 2396 31543 2400
rect 31532 2333 31543 2396
rect 31531 2329 31543 2333
rect 31446 2323 31543 2329
rect 23017 2211 30853 2213
rect 31024 2270 31488 2271
rect 31024 2207 31465 2270
rect 31532 2207 31542 2270
rect 31024 2204 31488 2207
rect 28510 2135 29798 2136
rect 22042 1787 22835 1867
rect 21792 1774 22835 1787
rect 21752 1762 22835 1774
rect 21287 1649 21321 1762
rect 21757 1758 22835 1762
rect 25436 2134 29922 2135
rect 25436 2125 29923 2134
rect 25436 2035 29826 2125
rect 29910 2035 29923 2125
rect 25436 2029 29923 2035
rect 25436 2028 29922 2029
rect 21683 1724 21749 1731
rect 21683 1690 21699 1724
rect 21733 1690 21749 1724
rect 21683 1649 21749 1690
rect 21167 1648 21749 1649
rect 21167 1619 21867 1648
rect 21167 1525 21203 1619
rect 21403 1525 21439 1619
rect 21639 1618 21867 1619
rect 21639 1525 21675 1618
rect 21801 1607 21867 1618
rect 21801 1573 21817 1607
rect 21851 1573 21867 1607
rect 21801 1566 21867 1573
rect 22111 1525 22146 1758
rect 21044 1513 21090 1525
rect 21044 1337 21050 1513
rect 21084 1337 21090 1513
rect 21044 1325 21090 1337
rect 21162 1513 21208 1525
rect 21162 1337 21168 1513
rect 21202 1337 21208 1513
rect 21162 1325 21208 1337
rect 21280 1513 21326 1525
rect 21280 1337 21286 1513
rect 21320 1337 21326 1513
rect 21280 1325 21326 1337
rect 21398 1513 21444 1525
rect 21398 1337 21404 1513
rect 21438 1337 21444 1513
rect 21398 1325 21444 1337
rect 21516 1513 21562 1525
rect 21516 1337 21522 1513
rect 21556 1337 21562 1513
rect 21516 1325 21562 1337
rect 21634 1513 21680 1525
rect 21634 1337 21640 1513
rect 21674 1337 21680 1513
rect 21634 1325 21680 1337
rect 21752 1513 21798 1525
rect 21752 1337 21758 1513
rect 21792 1337 21798 1513
rect 21752 1325 21798 1337
rect 21870 1513 21916 1525
rect 21870 1337 21876 1513
rect 21910 1337 21916 1513
rect 21870 1325 21916 1337
rect 21988 1513 22034 1525
rect 21988 1337 21994 1513
rect 22028 1337 22034 1513
rect 21988 1325 22034 1337
rect 22106 1513 22152 1525
rect 22106 1337 22112 1513
rect 22146 1337 22152 1513
rect 22106 1325 22152 1337
rect 21051 1219 21083 1325
rect 21287 1219 21319 1325
rect 21523 1219 21555 1325
rect 21759 1219 21791 1325
rect 21994 1219 22028 1325
rect 21051 1189 22028 1219
rect 21355 1161 21491 1189
rect 21355 1099 21391 1161
rect 21451 1099 21491 1161
rect 21355 1079 21491 1099
rect 3 897 1545 898
rect 13924 897 14348 898
rect 3 821 15 897
rect 109 892 14348 897
rect 109 888 7656 892
rect 109 821 2616 888
rect 3 819 2616 821
rect 2712 819 7656 888
rect 3 818 7656 819
rect 7756 818 14348 892
rect 3 815 14348 818
rect 5 813 14348 815
rect 14862 926 20826 1001
rect 871 812 13970 813
rect 491 782 14037 784
rect 14862 782 14943 926
rect 25436 887 25592 2028
rect 30043 1876 30179 1896
rect 30043 1814 30079 1876
rect 30139 1814 30179 1876
rect 30043 1786 30179 1814
rect 29739 1756 30716 1786
rect 29739 1650 29771 1756
rect 29975 1650 30007 1756
rect 30211 1650 30243 1756
rect 30447 1650 30479 1756
rect 30682 1650 30716 1756
rect 29732 1638 29778 1650
rect 29732 1462 29738 1638
rect 29772 1462 29778 1638
rect 29732 1450 29778 1462
rect 29850 1638 29896 1650
rect 29850 1462 29856 1638
rect 29890 1462 29896 1638
rect 29850 1450 29896 1462
rect 29968 1638 30014 1650
rect 29968 1462 29974 1638
rect 30008 1462 30014 1638
rect 29968 1450 30014 1462
rect 30086 1638 30132 1650
rect 30086 1462 30092 1638
rect 30126 1462 30132 1638
rect 30086 1450 30132 1462
rect 30204 1638 30250 1650
rect 30204 1462 30210 1638
rect 30244 1462 30250 1638
rect 30204 1450 30250 1462
rect 30322 1638 30368 1650
rect 30322 1462 30328 1638
rect 30362 1462 30368 1638
rect 30322 1450 30368 1462
rect 30440 1638 30486 1650
rect 30440 1462 30446 1638
rect 30480 1462 30486 1638
rect 30440 1450 30486 1462
rect 30558 1638 30604 1650
rect 30558 1462 30564 1638
rect 30598 1462 30604 1638
rect 30558 1450 30604 1462
rect 30676 1638 30722 1650
rect 30676 1462 30682 1638
rect 30716 1462 30722 1638
rect 30676 1450 30722 1462
rect 30794 1638 30840 1650
rect 30794 1462 30800 1638
rect 30834 1462 30840 1638
rect 30794 1450 30840 1462
rect 28753 1391 29337 1392
rect 491 776 14943 782
rect 491 690 502 776
rect 601 690 14943 776
rect 491 682 14943 690
rect 871 681 14943 682
rect 14971 806 25592 887
rect 25630 1382 29338 1391
rect 25630 1292 29241 1382
rect 29325 1292 29338 1382
rect 29855 1356 29891 1450
rect 30091 1356 30127 1450
rect 30327 1357 30363 1450
rect 30489 1402 30555 1409
rect 30489 1368 30505 1402
rect 30539 1368 30555 1402
rect 30489 1357 30555 1368
rect 30327 1356 30555 1357
rect 29855 1327 30555 1356
rect 29855 1326 30437 1327
rect 25630 1286 29338 1292
rect 25630 1285 29337 1286
rect 25630 1284 27815 1285
rect 14971 805 20661 806
rect 594 642 1545 643
rect 594 641 13986 642
rect 14971 641 15055 805
rect 25630 764 25786 1284
rect 29975 1213 30009 1326
rect 30371 1285 30437 1326
rect 30371 1251 30387 1285
rect 30421 1251 30437 1285
rect 30371 1244 30437 1251
rect 30799 1217 30834 1450
rect 31024 1217 31119 2204
rect 31603 1697 31637 2481
rect 32316 2419 32350 2481
rect 31905 2381 32647 2419
rect 31715 2210 31725 2278
rect 31780 2210 31790 2278
rect 31905 2257 31939 2381
rect 32141 2257 32175 2381
rect 32377 2257 32411 2381
rect 32613 2257 32647 2381
rect 31899 2245 31945 2257
rect 31899 1869 31905 2245
rect 31939 1869 31945 2245
rect 31899 1857 31945 1869
rect 32017 2245 32063 2257
rect 32017 1869 32023 2245
rect 32057 1869 32063 2245
rect 32017 1857 32063 1869
rect 32135 2245 32181 2257
rect 32135 1869 32141 2245
rect 32175 1869 32181 2245
rect 32135 1857 32181 1869
rect 32253 2245 32299 2257
rect 32253 1869 32259 2245
rect 32293 1869 32299 2245
rect 32253 1857 32299 1869
rect 32371 2245 32417 2257
rect 32371 1869 32377 2245
rect 32411 1869 32417 2245
rect 32371 1857 32417 1869
rect 32489 2245 32535 2257
rect 32489 1869 32495 2245
rect 32529 1869 32535 2245
rect 32489 1857 32535 1869
rect 32607 2245 32653 2257
rect 32607 1869 32613 2245
rect 32647 1869 32653 2245
rect 32773 2040 32847 2052
rect 32769 1949 32779 2040
rect 32841 1949 32851 2040
rect 32773 1937 32847 1949
rect 32607 1857 32653 1869
rect 33019 1698 33053 2481
rect 33388 2453 33424 2547
rect 33624 2453 33660 2547
rect 33860 2454 33896 2547
rect 34022 2499 34088 2506
rect 34022 2465 34038 2499
rect 34072 2465 34088 2499
rect 34022 2454 34088 2465
rect 33860 2453 34088 2454
rect 33388 2424 34088 2453
rect 33388 2423 33970 2424
rect 33114 2391 33190 2396
rect 33111 2335 33121 2391
rect 33174 2390 33190 2391
rect 33174 2335 33440 2390
rect 33114 2330 33440 2335
rect 33235 2288 33326 2293
rect 33235 2199 33245 2288
rect 33318 2199 33326 2288
rect 33235 2187 33326 2199
rect 33272 1793 33326 2187
rect 33386 1878 33440 2330
rect 33508 2310 33542 2423
rect 33904 2382 33970 2423
rect 33904 2348 33920 2382
rect 33954 2348 33970 2382
rect 33904 2341 33970 2348
rect 34332 2314 34367 2547
rect 33978 2310 34367 2314
rect 33502 2298 33548 2310
rect 33502 1922 33508 2298
rect 33542 1922 33548 2298
rect 33502 1910 33548 1922
rect 33620 2298 33666 2310
rect 33620 1922 33626 2298
rect 33660 1922 33666 2298
rect 33620 1910 33666 1922
rect 33738 2298 33784 2310
rect 33738 1922 33744 2298
rect 33778 1949 33784 2298
rect 33855 2298 33901 2310
rect 33855 2122 33861 2298
rect 33895 2122 33901 2298
rect 33855 2115 33901 2122
rect 33973 2299 34367 2310
rect 33973 2298 34210 2299
rect 33973 2122 33979 2298
rect 34013 2285 34210 2298
rect 34013 2122 34019 2285
rect 34192 2211 34210 2285
rect 34352 2211 34367 2299
rect 34192 2196 34367 2211
rect 33855 2110 33904 2115
rect 33973 2110 34019 2122
rect 33861 1949 33904 2110
rect 33778 1922 33904 1949
rect 33738 1910 33904 1922
rect 33744 1906 33904 1910
rect 33386 1872 33617 1878
rect 33386 1838 33567 1872
rect 33601 1838 33617 1872
rect 33386 1822 33617 1838
rect 33669 1872 33735 1878
rect 33669 1838 33685 1872
rect 33719 1838 33735 1872
rect 33669 1793 33735 1838
rect 33272 1785 33735 1793
rect 33272 1753 33736 1785
rect 33828 1769 33904 1906
rect 36607 1868 36664 2631
rect 36751 2625 37151 2631
rect 36751 2547 37151 2553
rect 36751 2513 36763 2547
rect 37139 2513 37151 2547
rect 36751 2507 37151 2513
rect 36751 2429 37151 2435
rect 36751 2395 36763 2429
rect 37139 2395 37151 2429
rect 36751 2389 37151 2395
rect 36751 2311 37151 2317
rect 36751 2277 36763 2311
rect 37139 2277 37151 2311
rect 36751 2271 37151 2277
rect 36751 2198 37151 2204
rect 36751 2164 36763 2198
rect 37139 2164 37277 2198
rect 36751 2158 37151 2164
rect 36751 2080 37151 2086
rect 36751 2046 36763 2080
rect 37139 2046 37151 2080
rect 36751 2040 37151 2046
rect 36751 1962 37151 1968
rect 36751 1928 36763 1962
rect 37139 1928 37151 1962
rect 36751 1922 37151 1928
rect 36507 1858 36664 1868
rect 36567 1778 36664 1858
rect 36751 1844 37151 1850
rect 36751 1810 36763 1844
rect 37139 1810 37151 1844
rect 36751 1804 37151 1810
rect 33824 1709 33834 1769
rect 33896 1709 33906 1769
rect 36507 1768 36664 1778
rect 32746 1697 33053 1698
rect 31603 1692 31919 1697
rect 32633 1692 33053 1697
rect 31603 1681 31986 1692
rect 31603 1654 31935 1681
rect 31603 1525 31637 1654
rect 31919 1647 31935 1654
rect 31969 1647 31986 1681
rect 31919 1641 31986 1647
rect 32566 1681 33053 1692
rect 33832 1683 33902 1709
rect 32566 1647 32583 1681
rect 32617 1654 33053 1681
rect 32617 1647 32633 1654
rect 32746 1653 33053 1654
rect 32566 1641 32633 1647
rect 31744 1614 31800 1626
rect 31744 1580 31750 1614
rect 31784 1613 31800 1614
rect 32857 1613 32913 1625
rect 31784 1597 32251 1613
rect 31784 1580 32201 1597
rect 31744 1564 32201 1580
rect 32185 1563 32201 1564
rect 32235 1563 32251 1597
rect 32185 1556 32251 1563
rect 32303 1598 32873 1613
rect 32303 1564 32319 1598
rect 32353 1579 32873 1598
rect 32907 1579 32913 1613
rect 32353 1564 32913 1579
rect 32303 1554 32370 1564
rect 32857 1563 32913 1564
rect 33019 1525 33053 1653
rect 31597 1513 31643 1525
rect 31597 1337 31603 1513
rect 31637 1337 31643 1513
rect 31597 1325 31643 1337
rect 31715 1513 31761 1525
rect 31715 1337 31721 1513
rect 31755 1337 31761 1513
rect 31715 1325 31761 1337
rect 32017 1513 32063 1525
rect 30445 1213 31119 1217
rect 29969 1201 30015 1213
rect 594 639 15055 641
rect 594 633 7464 639
rect 594 567 619 633
rect 763 567 7464 633
rect 7556 567 15055 639
rect 594 558 15055 567
rect 871 557 15055 558
rect 13963 556 15055 557
rect 15083 682 25786 764
rect 191 508 1545 509
rect 15083 508 15161 682
rect 25630 681 25786 682
rect 25835 1075 26240 1077
rect 25835 1073 29533 1075
rect 25835 1066 29907 1073
rect 25835 976 29410 1066
rect 29494 976 29907 1066
rect 25835 971 29907 976
rect 25835 970 29533 971
rect 25835 969 26240 970
rect 25835 641 25991 969
rect 29853 781 29907 971
rect 29969 825 29975 1201
rect 30009 825 30015 1201
rect 29969 813 30015 825
rect 30087 1201 30133 1213
rect 30087 825 30093 1201
rect 30127 825 30133 1201
rect 30087 813 30133 825
rect 30205 1201 30251 1213
rect 30205 825 30211 1201
rect 30245 852 30251 1201
rect 30322 1201 30368 1213
rect 30322 1025 30328 1201
rect 30362 1025 30368 1201
rect 30322 1018 30368 1025
rect 30440 1201 31119 1213
rect 30440 1025 30446 1201
rect 30480 1188 31119 1201
rect 30480 1025 30486 1188
rect 30730 1108 31119 1188
rect 30322 1013 30371 1018
rect 30440 1013 30486 1025
rect 31720 1031 31754 1325
rect 32017 1137 32023 1513
rect 32057 1137 32063 1513
rect 32017 1125 32063 1137
rect 32135 1513 32181 1525
rect 32135 1137 32141 1513
rect 32175 1137 32181 1513
rect 32135 1125 32181 1137
rect 32253 1513 32299 1525
rect 32253 1137 32259 1513
rect 32293 1137 32299 1513
rect 32253 1125 32299 1137
rect 32371 1513 32417 1525
rect 32371 1137 32377 1513
rect 32411 1137 32417 1513
rect 32371 1125 32417 1137
rect 32489 1513 32535 1525
rect 32489 1137 32495 1513
rect 32529 1137 32535 1513
rect 32895 1513 32941 1525
rect 32895 1337 32901 1513
rect 32935 1337 32941 1513
rect 32895 1325 32941 1337
rect 33013 1513 33059 1525
rect 33013 1337 33019 1513
rect 33053 1337 33059 1513
rect 33013 1325 33059 1337
rect 36607 1490 36664 1768
rect 36751 1726 37151 1732
rect 36751 1692 36763 1726
rect 37139 1692 37151 1726
rect 36751 1686 37151 1692
rect 36751 1608 37151 1614
rect 36751 1574 36763 1608
rect 37139 1574 37151 1608
rect 36751 1568 37151 1574
rect 36751 1490 37151 1496
rect 36607 1456 36763 1490
rect 37139 1456 37151 1490
rect 32489 1125 32535 1137
rect 32377 1031 32411 1125
rect 32901 1031 32934 1325
rect 30328 852 30371 1013
rect 31720 999 32934 1031
rect 30245 825 30371 852
rect 30205 813 30371 825
rect 30211 809 30371 813
rect 29853 775 30084 781
rect 29853 741 30034 775
rect 30068 741 30084 775
rect 29853 725 30084 741
rect 30136 775 30202 781
rect 30136 741 30152 775
rect 30186 741 30202 775
rect 191 493 15161 508
rect 191 422 204 493
rect 318 422 15161 493
rect 191 407 15161 422
rect 15189 632 25991 641
rect 15189 564 20896 632
rect 20965 564 25991 632
rect 15189 557 25991 564
rect 26038 720 26194 722
rect 29722 720 29785 721
rect 26038 717 29797 720
rect 26038 642 29723 717
rect 29784 696 29797 717
rect 30136 696 30202 741
rect 29784 688 30202 696
rect 29784 656 30203 688
rect 30295 672 30371 809
rect 32086 975 32492 999
rect 32086 852 32198 975
rect 32372 852 32492 975
rect 36607 899 36664 1456
rect 36751 1450 37151 1456
rect 36751 1371 37151 1377
rect 36751 1337 36763 1371
rect 37139 1337 37151 1371
rect 36751 1331 37151 1337
rect 36751 1253 37151 1259
rect 36751 1219 36763 1253
rect 37139 1219 37151 1253
rect 36751 1213 37151 1219
rect 36751 1135 37151 1141
rect 36751 1101 36763 1135
rect 37139 1101 37151 1135
rect 36751 1095 37151 1101
rect 36751 1017 37151 1023
rect 37235 1017 37277 2164
rect 37337 2020 37404 3072
rect 37437 3005 37522 3017
rect 37437 2934 37450 3005
rect 37513 2934 37522 3005
rect 37437 2925 37522 2934
rect 37914 2273 37961 3072
rect 38084 2273 38284 2278
rect 37914 2272 38284 2273
rect 37914 2239 38096 2272
rect 37337 1986 37354 2020
rect 37388 1986 37404 2020
rect 37337 1970 37404 1986
rect 37725 2038 37810 2050
rect 37725 1970 37733 2038
rect 37798 1970 37810 2038
rect 37725 1958 37810 1970
rect 37440 1920 37525 1932
rect 37440 1850 37450 1920
rect 37512 1850 37525 1920
rect 37440 1840 37525 1850
rect 37914 1801 37961 2239
rect 38084 2238 38096 2239
rect 38272 2238 38284 2272
rect 38084 2232 38284 2238
rect 38084 2154 38284 2160
rect 38084 2120 38096 2154
rect 38272 2120 38703 2154
rect 38084 2086 38284 2120
rect 38084 2080 38484 2086
rect 38084 2046 38096 2080
rect 38472 2046 38484 2080
rect 38084 2040 38484 2046
rect 38084 1962 38484 1968
rect 38084 1928 38096 1962
rect 38472 1928 38484 1962
rect 38084 1922 38484 1928
rect 38084 1844 38484 1850
rect 38557 1844 38623 1859
rect 38084 1810 38096 1844
rect 38472 1843 38623 1844
rect 38472 1810 38573 1843
rect 38084 1804 38484 1810
rect 38557 1809 38573 1810
rect 38607 1809 38623 1843
rect 37914 1785 38024 1801
rect 38557 1793 38623 1809
rect 38651 1856 38703 2120
rect 38651 1844 38781 1856
rect 37914 1751 37974 1785
rect 38008 1751 38024 1785
rect 37914 1735 38024 1751
rect 38651 1778 38725 1844
rect 38777 1778 38781 1844
rect 38651 1764 38781 1778
rect 38084 1726 38484 1732
rect 38084 1692 38096 1726
rect 38472 1692 38484 1726
rect 38084 1686 38484 1692
rect 37564 1679 37636 1685
rect 37564 1620 37570 1679
rect 37630 1620 37636 1679
rect 37567 1616 37634 1620
rect 37570 1610 37630 1616
rect 38084 1608 38484 1614
rect 38084 1574 38096 1608
rect 38472 1574 38484 1608
rect 38084 1568 38484 1574
rect 38084 1530 38284 1568
rect 38651 1530 38703 1764
rect 38084 1496 38096 1530
rect 38272 1496 38703 1530
rect 38084 1490 38284 1496
rect 37913 1412 37960 1413
rect 38084 1412 38284 1418
rect 37913 1378 38096 1412
rect 38272 1378 38284 1412
rect 36751 983 36763 1017
rect 37139 983 37363 1017
rect 36751 977 37151 983
rect 36951 899 37151 904
rect 36607 898 37151 899
rect 36607 864 36963 898
rect 37139 864 37151 898
rect 36607 862 37151 864
rect 36951 858 37151 862
rect 32086 808 32492 852
rect 36951 780 37151 786
rect 36951 746 36963 780
rect 37139 746 37151 780
rect 36951 740 37151 746
rect 37297 710 37363 983
rect 37297 676 37313 710
rect 37347 676 37363 710
rect 29784 642 29797 656
rect 26038 632 29797 642
rect 191 406 14045 407
rect 871 405 14045 406
rect 6 370 146 371
rect 6 369 1545 370
rect 2717 369 2923 371
rect 15189 369 15284 557
rect 6 367 15284 369
rect -2383 319 -2371 353
rect -2195 320 -1857 353
rect 3 361 15284 367
rect -2195 319 -2183 320
rect -2383 313 -2183 319
rect 3 278 15 361
rect 122 355 15284 361
rect 122 289 2748 355
rect 2892 289 15284 355
rect 122 278 15284 289
rect 3 272 15284 278
rect 6 268 15284 272
rect 15312 507 20168 508
rect 26038 507 26194 632
rect 30291 612 30301 672
rect 30363 612 30373 672
rect 36951 662 37151 668
rect 36951 628 36963 662
rect 37139 628 37151 662
rect 37297 660 37363 676
rect 36951 622 37151 628
rect 15312 407 26194 507
rect 36951 544 37151 550
rect 37913 544 37960 1378
rect 38084 1372 38284 1378
rect 36951 510 36963 544
rect 37139 510 37960 544
rect 39197 510 39589 640
rect 36951 509 39589 510
rect 36951 504 37151 509
rect 6 267 146 268
rect 871 267 13814 268
rect -2383 235 -2183 241
rect -3608 219 -3408 225
rect -3954 185 -3596 219
rect -3420 185 -3408 219
rect -3608 179 -3408 185
rect -3374 201 -2371 235
rect -2195 201 -2183 235
rect 15312 230 15402 407
rect 37505 390 39589 509
rect 39197 269 39589 390
rect -3608 101 -3408 107
rect -3374 101 -3339 201
rect -2383 195 -2183 201
rect 2454 210 15402 230
rect 2454 156 2462 210
rect 2557 156 15402 210
rect 2454 149 15402 156
rect -3608 67 -3596 101
rect -3420 67 -3339 101
rect -2705 137 -2591 149
rect -3608 61 -3408 67
rect -2705 35 -2699 137
rect -2597 35 -2591 137
rect -2705 23 -2591 35
<< via1 >>
rect 4391 28180 4522 28302
rect 6283 27798 6415 27906
rect 8765 27852 8897 27960
rect 9166 27862 9222 27876
rect 9166 27828 9182 27862
rect 9182 27828 9216 27862
rect 9216 27828 9222 27862
rect 9166 27810 9222 27828
rect 9912 27852 10044 27960
rect 8036 27738 8102 27754
rect 8036 27704 8052 27738
rect 8052 27704 8086 27738
rect 8086 27704 8102 27738
rect 8036 27688 8102 27704
rect 12796 27795 12928 27903
rect 15278 27849 15410 27957
rect 8702 27041 8801 27138
rect 6563 26735 6671 26867
rect -832 23256 -674 23393
rect -3253 16170 -3187 16236
rect -3057 16184 -2997 16248
rect -2997 16184 -2996 16248
rect -4055 15418 -4001 15428
rect -4055 15380 -4047 15418
rect -4047 15380 -4009 15418
rect -4009 15380 -4001 15418
rect -4055 15374 -4001 15380
rect -1831 15480 -1773 15486
rect -1831 15430 -1825 15480
rect -1825 15430 -1783 15480
rect -1783 15430 -1773 15480
rect -1831 15424 -1773 15430
rect -3247 14794 -3193 14848
rect -2684 14528 -2605 14605
rect -3255 14102 -3189 14168
rect -3059 14115 -2999 14177
rect -4057 13350 -4003 13360
rect -4057 13312 -4049 13350
rect -4049 13312 -4011 13350
rect -4011 13312 -4003 13350
rect -4057 13306 -4003 13312
rect -1833 13412 -1775 13418
rect -1833 13362 -1827 13412
rect -1827 13362 -1785 13412
rect -1785 13362 -1775 13412
rect -1833 13356 -1775 13362
rect -3249 12726 -3195 12780
rect -2681 12462 -2610 12536
rect -3253 12033 -3187 12099
rect -3056 12048 -2997 12108
rect -2997 12048 -2996 12108
rect -4055 11281 -4001 11291
rect -4055 11243 -4047 11281
rect -4047 11243 -4009 11281
rect -4009 11243 -4001 11281
rect -4055 11237 -4001 11243
rect -1831 11343 -1773 11349
rect -1831 11293 -1825 11343
rect -1825 11293 -1783 11343
rect -1783 11293 -1773 11343
rect -1831 11287 -1773 11293
rect -3247 10657 -3193 10711
rect -2674 10394 -2611 10459
rect -1209 12315 -1143 12389
rect -1342 10230 -1280 10294
rect -3255 9965 -3189 10031
rect -3057 9979 -3002 10040
rect -4057 9213 -4003 9223
rect -4057 9175 -4049 9213
rect -4049 9175 -4011 9213
rect -4011 9175 -4003 9213
rect -4057 9169 -4003 9175
rect -1833 9275 -1775 9281
rect -1833 9225 -1827 9275
rect -1827 9225 -1785 9275
rect -1785 9225 -1775 9275
rect -1833 9219 -1775 9225
rect -3249 8589 -3195 8643
rect -2682 8327 -2609 8391
rect -3255 7896 -3189 7962
rect -3058 7910 -3002 7971
rect -4057 7144 -4003 7154
rect -4057 7106 -4049 7144
rect -4049 7106 -4011 7144
rect -4011 7106 -4003 7144
rect -4057 7100 -4003 7106
rect -1833 7206 -1775 7212
rect -1833 7156 -1827 7206
rect -1827 7156 -1785 7206
rect -1785 7156 -1775 7206
rect -1833 7150 -1775 7156
rect -3249 6520 -3195 6574
rect -2679 6259 -2614 6325
rect -3257 5828 -3191 5894
rect -3059 5842 -3003 5904
rect -4059 5076 -4005 5086
rect -4059 5038 -4051 5076
rect -4051 5038 -4013 5076
rect -4013 5038 -4005 5076
rect -4059 5032 -4005 5038
rect -1835 5138 -1777 5144
rect -1835 5088 -1829 5138
rect -1829 5088 -1787 5138
rect -1787 5088 -1777 5138
rect -1835 5082 -1777 5088
rect -3251 4452 -3197 4506
rect -2679 4188 -2614 4258
rect -3255 3759 -3189 3825
rect -3055 3774 -3003 3834
rect -4057 3007 -4003 3017
rect -4057 2969 -4049 3007
rect -4049 2969 -4011 3007
rect -4011 2969 -4003 3007
rect -4057 2963 -4003 2969
rect -1833 3069 -1775 3075
rect -1833 3019 -1827 3069
rect -1827 3019 -1785 3069
rect -1785 3019 -1775 3069
rect -1833 3013 -1775 3019
rect -3249 2383 -3195 2437
rect -2682 2119 -2609 2189
rect -651 16282 -590 16334
rect 8111 26452 8243 26560
rect 5549 26174 5661 26280
rect 6297 26148 6429 26256
rect 9858 27064 9923 27118
rect 15679 27859 15735 27873
rect 15679 27825 15695 27859
rect 15695 27825 15729 27859
rect 15729 27825 15735 27859
rect 15679 27807 15735 27825
rect 16425 27849 16557 27957
rect 14549 27735 14615 27751
rect 14549 27701 14565 27735
rect 14565 27701 14599 27735
rect 14599 27701 14615 27735
rect 14549 27685 14615 27701
rect 19330 27790 19462 27898
rect 21812 27844 21944 27952
rect 10953 27052 11021 27127
rect 9253 26450 9385 26558
rect 8110 25805 8242 25913
rect 10008 25805 10140 25913
rect 5832 25043 5950 25161
rect 6577 25085 6685 25217
rect 11432 26694 11668 26838
rect 15215 27038 15314 27135
rect 13076 26732 13184 26864
rect 5329 24701 5422 24780
rect 6292 24544 6424 24652
rect 8755 24927 8818 24943
rect 8755 24893 8784 24927
rect 8784 24893 8818 24927
rect 8755 24877 8818 24893
rect 11567 25146 11679 25148
rect 11567 25042 11685 25146
rect 11573 25040 11685 25042
rect 6879 23849 6942 23901
rect 6572 23481 6680 23613
rect 5834 23266 5946 23372
rect 8055 23409 8187 23517
rect 9953 23409 10085 23517
rect 14624 26449 14756 26557
rect 12062 26171 12174 26277
rect 12810 26145 12942 26253
rect 16371 27061 16436 27115
rect 22213 27854 22269 27868
rect 22213 27820 22229 27854
rect 22229 27820 22263 27854
rect 22263 27820 22269 27854
rect 22213 27802 22269 27820
rect 22959 27844 23091 27952
rect 21083 27730 21149 27746
rect 21083 27696 21099 27730
rect 21099 27696 21133 27730
rect 21133 27696 21149 27730
rect 21083 27680 21149 27696
rect 25888 27794 26020 27902
rect 28370 27848 28502 27956
rect 17466 27049 17534 27124
rect 15766 26447 15898 26555
rect 14623 25802 14755 25910
rect 16521 25802 16653 25910
rect 12345 25040 12463 25158
rect 13090 25082 13198 25214
rect 17969 26688 18202 26845
rect 21749 27033 21848 27130
rect 19610 26727 19718 26859
rect 11842 24698 11935 24777
rect 12805 24541 12937 24649
rect 15268 24924 15331 24940
rect 15268 24890 15297 24924
rect 15297 24890 15331 24924
rect 15268 24874 15331 24890
rect 18101 25141 18213 25143
rect 18101 25037 18219 25141
rect 18107 25035 18219 25037
rect 13392 23846 13455 23898
rect 13085 23478 13193 23610
rect 12347 23263 12459 23369
rect 14568 23406 14700 23514
rect 16466 23406 16598 23514
rect 21158 26444 21290 26552
rect 18596 26166 18708 26272
rect 19344 26140 19476 26248
rect 22905 27056 22970 27110
rect 28771 27858 28827 27872
rect 28771 27824 28787 27858
rect 28787 27824 28821 27858
rect 28821 27824 28827 27858
rect 28771 27806 28827 27824
rect 29517 27848 29649 27956
rect 27641 27734 27707 27750
rect 27641 27700 27657 27734
rect 27657 27700 27691 27734
rect 27691 27700 27707 27734
rect 27641 27684 27707 27700
rect 24000 27044 24068 27119
rect 22300 26442 22432 26550
rect 21157 25797 21289 25905
rect 23055 25797 23187 25905
rect 18879 25035 18997 25153
rect 19624 25077 19732 25209
rect 24529 26683 24776 26846
rect 28307 27037 28406 27134
rect 26168 26731 26276 26863
rect 18376 24693 18469 24772
rect 19339 24536 19471 24644
rect 21802 24919 21865 24935
rect 21802 24885 21831 24919
rect 21831 24885 21865 24919
rect 21802 24869 21865 24885
rect 24659 25145 24771 25147
rect 24659 25041 24777 25145
rect 24665 25039 24777 25041
rect 19926 23841 19989 23893
rect 19619 23473 19727 23605
rect 18881 23258 18993 23364
rect 21102 23401 21234 23509
rect 23000 23401 23132 23509
rect 27716 26448 27848 26556
rect 25154 26170 25266 26276
rect 25902 26144 26034 26252
rect 29463 27060 29528 27114
rect 30558 27048 30626 27123
rect 28858 26446 28990 26554
rect 27715 25801 27847 25909
rect 29613 25801 29745 25909
rect 25437 25039 25555 25157
rect 26182 25081 26290 25213
rect 24934 24697 25027 24776
rect 25897 24540 26029 24648
rect 28360 24923 28423 24939
rect 28360 24889 28389 24923
rect 28389 24889 28423 24923
rect 28360 24873 28423 24889
rect 26484 23845 26547 23897
rect 26177 23477 26285 23609
rect 25439 23262 25551 23368
rect 27660 23405 27792 23513
rect 29558 23405 29690 23513
rect 11268 22994 11396 23072
rect 17781 22810 17892 22921
rect 24369 22620 24503 22738
rect 5860 22244 5992 22352
rect 6682 22254 6738 22268
rect 6682 22220 6688 22254
rect 6688 22220 6722 22254
rect 6722 22220 6738 22254
rect 6682 22202 6738 22220
rect 7007 22244 7139 22352
rect 5981 21456 6046 21510
rect 6519 20842 6651 20950
rect 7802 22130 7868 22146
rect 7802 22096 7818 22130
rect 7818 22096 7852 22130
rect 7852 22096 7868 22130
rect 7802 22080 7868 22096
rect 9489 22190 9621 22298
rect 12418 22240 12550 22348
rect 13240 22250 13296 22264
rect 13240 22216 13246 22250
rect 13246 22216 13280 22250
rect 13280 22216 13296 22250
rect 13240 22198 13296 22216
rect 13565 22240 13697 22348
rect 7103 21433 7202 21530
rect 9233 21127 9341 21259
rect 11441 21440 11509 21515
rect 12539 21452 12604 21506
rect 10755 21083 10979 21219
rect 7661 20844 7793 20952
rect 9475 20540 9607 20648
rect 10243 20566 10355 20672
rect 5764 20197 5896 20305
rect 7662 20197 7794 20305
rect 9219 19477 9327 19609
rect 7086 19319 7149 19335
rect 7086 19285 7120 19319
rect 7120 19285 7149 19319
rect 7086 19269 7149 19285
rect 9954 19435 10072 19553
rect 10737 20549 10738 20655
rect 10738 20549 10849 20655
rect 13077 20838 13209 20946
rect 14360 22126 14426 22142
rect 14360 22092 14376 22126
rect 14376 22092 14410 22126
rect 14410 22092 14426 22126
rect 14360 22076 14426 22092
rect 16047 22186 16179 22294
rect 18952 22245 19084 22353
rect 19774 22255 19830 22269
rect 19774 22221 19780 22255
rect 19780 22221 19814 22255
rect 19814 22221 19830 22255
rect 19774 22203 19830 22221
rect 20099 22245 20231 22353
rect 13661 21429 13760 21526
rect 15791 21123 15899 21255
rect 17975 21445 18043 21520
rect 19073 21457 19138 21511
rect 17298 21077 17548 21233
rect 14219 20840 14351 20948
rect 16033 20536 16165 20644
rect 16801 20562 16913 20668
rect 12322 20193 12454 20301
rect 14220 20193 14352 20301
rect 10738 19541 10850 19543
rect 10732 19437 10850 19541
rect 15777 19473 15885 19605
rect 10732 19435 10844 19437
rect 10482 19093 10575 19172
rect 9480 18936 9612 19044
rect 8962 18241 9025 18293
rect 5819 17801 5951 17909
rect 7717 17801 7849 17909
rect 9224 17873 9332 18005
rect 9958 17658 10070 17764
rect 13644 19315 13707 19331
rect 13644 19281 13678 19315
rect 13678 19281 13707 19315
rect 13644 19265 13707 19281
rect 16512 19431 16630 19549
rect 17295 20646 17407 20651
rect 17295 20549 17301 20646
rect 17301 20549 17404 20646
rect 17404 20549 17407 20646
rect 17295 20545 17407 20549
rect 19611 20843 19743 20951
rect 20894 22131 20960 22147
rect 20894 22097 20910 22131
rect 20910 22097 20944 22131
rect 20944 22097 20960 22131
rect 20894 22081 20960 22097
rect 22581 22191 22713 22299
rect 25465 22248 25597 22356
rect 26287 22258 26343 22272
rect 26287 22224 26293 22258
rect 26293 22224 26327 22258
rect 26327 22224 26343 22258
rect 26287 22206 26343 22224
rect 26612 22248 26744 22356
rect 20195 21434 20294 21531
rect 22325 21128 22433 21260
rect 24488 21448 24556 21523
rect 25586 21460 25651 21514
rect 23847 21085 24075 21222
rect 20753 20845 20885 20953
rect 22567 20541 22699 20649
rect 23335 20567 23447 20673
rect 18856 20198 18988 20306
rect 20754 20198 20886 20306
rect 17296 19537 17408 19539
rect 17290 19433 17408 19537
rect 22311 19478 22419 19610
rect 17290 19431 17402 19433
rect 17040 19089 17133 19168
rect 16038 18932 16170 19040
rect 15520 18237 15583 18289
rect 12377 17797 12509 17905
rect 14275 17797 14407 17905
rect 15782 17869 15890 18001
rect 16516 17654 16628 17760
rect 20178 19320 20241 19336
rect 20178 19286 20212 19320
rect 20212 19286 20241 19320
rect 20178 19270 20241 19286
rect 23046 19436 23164 19554
rect 23829 20650 23941 20656
rect 23829 20558 23837 20650
rect 23837 20558 23935 20650
rect 23935 20558 23941 20650
rect 23829 20550 23941 20558
rect 26124 20846 26256 20954
rect 27407 22134 27473 22150
rect 27407 22100 27423 22134
rect 27423 22100 27457 22134
rect 27457 22100 27473 22134
rect 27407 22084 27473 22100
rect 29094 22194 29226 22302
rect 26708 21437 26807 21534
rect 28838 21131 28946 21263
rect 30360 21085 30592 21216
rect 27266 20848 27398 20956
rect 29080 20544 29212 20652
rect 29848 20570 29960 20676
rect 25369 20201 25501 20309
rect 27267 20201 27399 20309
rect 23830 19542 23942 19544
rect 23824 19438 23942 19542
rect 28824 19481 28932 19613
rect 23824 19436 23936 19438
rect 23574 19094 23667 19173
rect 22572 18937 22704 19045
rect 22054 18242 22117 18294
rect 18911 17802 19043 17910
rect 20809 17802 20941 17910
rect 22316 17874 22424 18006
rect 23050 17659 23162 17765
rect 26691 19323 26754 19339
rect 26691 19289 26725 19323
rect 26725 19289 26754 19323
rect 26691 19273 26754 19289
rect 29559 19439 29677 19557
rect 37569 25234 37637 25291
rect 37737 25287 37805 25291
rect 37737 25238 37741 25287
rect 37741 25238 37801 25287
rect 37801 25238 37805 25287
rect 37737 25234 37805 25238
rect 30343 19545 30455 19547
rect 30337 19441 30455 19545
rect 30337 19439 30449 19441
rect 30087 19097 30180 19176
rect 29085 18940 29217 19048
rect 28567 18245 28630 18297
rect 25424 17805 25556 17913
rect 27322 17805 27454 17913
rect 28829 17877 28937 18009
rect 36511 23896 36571 23900
rect 36511 23824 36517 23896
rect 36517 23824 36571 23896
rect 36511 23820 36571 23824
rect 37454 25043 37517 25047
rect 37454 24983 37458 25043
rect 37458 24983 37513 25043
rect 37513 24983 37517 25043
rect 37454 24976 37517 24983
rect 37737 24076 37802 24080
rect 37737 24016 37742 24076
rect 37742 24016 37797 24076
rect 37797 24016 37802 24076
rect 37737 24012 37802 24016
rect 37454 23958 37516 23962
rect 37454 23898 37457 23958
rect 37457 23898 37512 23958
rect 37512 23898 37516 23958
rect 37454 23892 37516 23898
rect 38729 23882 38781 23886
rect 38729 23824 38775 23882
rect 38775 23824 38781 23882
rect 38729 23820 38781 23824
rect 37574 23708 37634 23721
rect 37574 23674 37588 23708
rect 37588 23674 37622 23708
rect 37622 23674 37634 23708
rect 37574 23662 37634 23674
rect 34490 22236 34558 22246
rect 34490 22173 34502 22236
rect 34502 22173 34551 22236
rect 34551 22173 34558 22236
rect 34490 22163 34558 22173
rect 37569 22090 37637 22147
rect 37737 22143 37805 22147
rect 37737 22094 37741 22143
rect 37741 22094 37801 22143
rect 37801 22094 37805 22143
rect 37737 22090 37805 22094
rect 36511 20752 36571 20756
rect 36511 20680 36517 20752
rect 36517 20680 36571 20752
rect 36511 20676 36571 20680
rect 37454 21899 37517 21903
rect 37454 21839 37458 21899
rect 37458 21839 37513 21899
rect 37513 21839 37517 21899
rect 37454 21832 37517 21839
rect 37737 20932 37802 20936
rect 37737 20872 37742 20932
rect 37742 20872 37797 20932
rect 37797 20872 37802 20932
rect 37737 20868 37802 20872
rect 37454 20814 37516 20818
rect 37454 20754 37457 20814
rect 37457 20754 37512 20814
rect 37512 20754 37516 20814
rect 37454 20748 37516 20754
rect 38729 20738 38781 20742
rect 38729 20680 38775 20738
rect 38775 20680 38781 20738
rect 38729 20676 38781 20680
rect 37574 20564 37634 20577
rect 37574 20530 37588 20564
rect 37588 20530 37622 20564
rect 37622 20530 37634 20564
rect 37574 20518 37634 20530
rect 37565 18958 37633 19015
rect 37733 19011 37801 19015
rect 37733 18962 37737 19011
rect 37737 18962 37797 19011
rect 37797 18962 37801 19011
rect 37733 18958 37801 18962
rect 29563 17662 29675 17768
rect 30617 16591 30768 16592
rect 30607 16502 30768 16591
rect 30617 16501 30768 16502
rect 24097 16345 24246 16433
rect 17570 16198 17726 16286
rect 23973 16242 24059 16251
rect 23973 16184 23984 16242
rect 23984 16184 24052 16242
rect 24052 16184 24059 16242
rect 23973 16176 24059 16184
rect 11000 16029 11129 16126
rect 17450 16123 17537 16130
rect 17450 16067 17459 16123
rect 17459 16067 17530 16123
rect 17530 16067 17537 16123
rect 17450 16060 17537 16067
rect 34744 15871 34888 15952
rect 10875 15790 10968 15797
rect 10875 15745 10883 15790
rect 10883 15745 10962 15790
rect 10962 15745 10968 15790
rect 10875 15736 10968 15745
rect 8153 15400 8213 15462
rect 14702 15399 14762 15461
rect 21356 15420 21416 15482
rect -651 14192 -594 14246
rect 8375 14250 8437 14258
rect 8375 14204 8381 14250
rect 8381 14204 8433 14250
rect 8433 14204 8437 14250
rect 8375 14198 8437 14204
rect 135 13866 219 13924
rect 373 13536 441 13539
rect 373 13491 380 13536
rect 380 13491 437 13536
rect 437 13491 441 13536
rect 373 13487 441 13491
rect 1489 13500 1549 13562
rect 4479 13323 4513 13355
rect 4513 13323 4580 13355
rect 4580 13323 4611 13355
rect 4479 13247 4611 13323
rect 6961 13373 6995 13409
rect 6995 13373 7062 13409
rect 7062 13373 7093 13409
rect 6961 13301 7093 13373
rect 17 12313 107 12405
rect 1711 12350 1773 12358
rect 1711 12304 1717 12350
rect 1717 12304 1769 12350
rect 1769 12304 1773 12350
rect 1711 12298 1773 12304
rect 7362 13311 7418 13325
rect 7362 13277 7378 13311
rect 7378 13277 7412 13311
rect 7412 13277 7418 13311
rect 7362 13259 7418 13277
rect 8108 13375 8137 13409
rect 8137 13375 8204 13409
rect 8204 13375 8240 13409
rect 8108 13301 8240 13375
rect 6232 13187 6298 13203
rect 6232 13153 6248 13187
rect 6248 13153 6282 13187
rect 6282 13153 6298 13187
rect 6232 13137 6298 13153
rect 6898 12490 6997 12587
rect 4759 12283 4867 12316
rect -655 12129 -592 12190
rect 4759 12216 4854 12283
rect 4854 12216 4867 12283
rect 4759 12184 4867 12216
rect 3251 11606 3363 11712
rect 1481 10915 1541 10977
rect 3250 10598 3362 10600
rect 3250 10494 3368 10598
rect 3256 10492 3368 10494
rect -655 10065 -592 10126
rect 6307 11912 6439 12009
rect 6307 11901 6340 11912
rect 6340 11901 6407 11912
rect 6407 11901 6439 11912
rect 3745 11623 3857 11729
rect 4493 11672 4525 11705
rect 4525 11672 4592 11705
rect 4592 11672 4625 11705
rect 4493 11597 4625 11672
rect 8054 12513 8119 12567
rect 14924 14249 14986 14257
rect 14924 14203 14930 14249
rect 14930 14203 14982 14249
rect 14982 14203 14986 14249
rect 14924 14197 14986 14203
rect 14358 13768 14415 13822
rect 21578 14270 21640 14278
rect 21578 14224 21584 14270
rect 21584 14224 21636 14270
rect 21636 14224 21640 14270
rect 21578 14218 21640 14224
rect 11028 13411 11062 13443
rect 11062 13411 11129 13443
rect 11129 13411 11160 13443
rect 11028 13335 11160 13411
rect 13510 13462 13545 13497
rect 13545 13462 13612 13497
rect 13612 13462 13642 13497
rect 13510 13389 13642 13462
rect 13911 13399 13967 13413
rect 13911 13365 13927 13399
rect 13927 13365 13961 13399
rect 13961 13365 13967 13399
rect 13911 13347 13967 13365
rect 14657 13464 14689 13497
rect 14689 13464 14756 13497
rect 14756 13464 14789 13497
rect 14657 13389 14789 13464
rect 12781 13275 12847 13291
rect 12781 13241 12797 13275
rect 12797 13241 12831 13275
rect 12831 13241 12847 13275
rect 12781 13225 12847 13241
rect 13447 12578 13546 12675
rect 11308 12365 11416 12404
rect 11308 12298 11400 12365
rect 11400 12298 11416 12365
rect 11308 12272 11416 12298
rect 7449 11914 7581 12007
rect 7449 11899 7478 11914
rect 7478 11899 7545 11914
rect 7545 11899 7581 11914
rect 9800 11694 9912 11800
rect 6306 11254 6438 11362
rect 8204 11330 8237 11362
rect 8237 11330 8304 11362
rect 8304 11330 8336 11362
rect 8204 11254 8336 11330
rect 4028 10492 4146 10610
rect 4773 10633 4881 10666
rect 4773 10566 4869 10633
rect 4869 10566 4881 10633
rect 4773 10534 4881 10566
rect 3525 10150 3618 10229
rect 174 9684 261 9788
rect -656 7994 -589 8061
rect -650 5933 -594 5987
rect 971 9687 1048 9783
rect 1703 9765 1765 9773
rect 1703 9719 1709 9765
rect 1709 9719 1761 9765
rect 1761 9719 1765 9765
rect 1703 9713 1765 9719
rect 4488 10066 4523 10101
rect 4523 10066 4590 10101
rect 4590 10066 4620 10101
rect 4488 9993 4620 10066
rect 6951 10376 7014 10392
rect 6951 10342 6980 10376
rect 6980 10342 7014 10376
rect 6951 10326 7014 10342
rect 5075 9298 5138 9350
rect 4768 9025 4876 9062
rect 4768 8958 4867 9025
rect 4867 8958 4876 9025
rect 4768 8930 4876 8958
rect 4030 8715 4142 8821
rect 6251 8872 6383 8966
rect 6251 8858 6280 8872
rect 6280 8858 6347 8872
rect 6347 8858 6383 8872
rect 8149 8858 8281 8966
rect 1462 7637 1522 7699
rect 4471 7543 4501 7575
rect 4501 7543 4568 7575
rect 4568 7543 4603 7575
rect 4471 7467 4603 7543
rect 6953 7598 6981 7629
rect 6981 7598 7048 7629
rect 7048 7598 7085 7629
rect 6953 7521 7085 7598
rect 7354 7531 7410 7545
rect 7354 7497 7370 7531
rect 7370 7497 7404 7531
rect 7404 7497 7410 7531
rect 7354 7479 7410 7497
rect 8100 7595 8137 7629
rect 8137 7595 8204 7629
rect 8204 7595 8232 7629
rect 8100 7521 8232 7595
rect 6224 7407 6290 7423
rect 6224 7373 6240 7407
rect 6240 7373 6274 7407
rect 6274 7373 6290 7407
rect 6224 7357 6290 7373
rect 1684 6487 1746 6495
rect 1684 6441 1690 6487
rect 1690 6441 1742 6487
rect 1742 6441 1746 6487
rect 1684 6435 1746 6441
rect 6890 6710 6989 6807
rect 4751 6496 4859 6536
rect 4751 6429 4844 6496
rect 4844 6429 4859 6496
rect 4751 6404 4859 6429
rect 3243 5826 3355 5932
rect 1478 4877 1538 4939
rect 6299 6135 6431 6229
rect 6299 6121 6321 6135
rect 6321 6121 6388 6135
rect 6388 6121 6431 6135
rect 3737 5843 3849 5949
rect 4485 5890 4522 5925
rect 4522 5890 4589 5925
rect 4589 5890 4617 5925
rect 4485 5817 4617 5890
rect 8046 6733 8111 6787
rect 12856 12008 12988 12097
rect 12856 11989 12885 12008
rect 12885 11989 12952 12008
rect 12952 11989 12988 12008
rect 10294 11711 10406 11817
rect 11042 11759 11076 11793
rect 11076 11759 11143 11793
rect 11143 11759 11174 11793
rect 11042 11685 11174 11759
rect 14603 12601 14668 12655
rect 15698 12589 15766 12664
rect 13998 12000 14130 12095
rect 13998 11987 14024 12000
rect 14024 11987 14091 12000
rect 14091 11987 14130 12000
rect 12855 11342 12987 11450
rect 14753 11417 14791 11450
rect 14791 11417 14858 11450
rect 14858 11417 14885 11450
rect 14753 11342 14885 11417
rect 10577 10580 10695 10698
rect 11322 10715 11430 10754
rect 11322 10648 11418 10715
rect 11418 10648 11430 10715
rect 11322 10622 11430 10648
rect 10074 10238 10167 10317
rect 11037 10159 11068 10189
rect 11068 10159 11135 10189
rect 11135 10159 11169 10189
rect 11037 10081 11169 10159
rect 13500 10464 13563 10480
rect 13500 10430 13529 10464
rect 13529 10430 13563 10464
rect 13500 10414 13563 10430
rect 11624 9386 11687 9438
rect 11317 9114 11425 9150
rect 11317 9047 11415 9114
rect 11415 9047 11425 9114
rect 11317 9018 11425 9047
rect 10579 8803 10691 8909
rect 12800 8957 12932 9054
rect 12800 8946 12829 8957
rect 12829 8946 12896 8957
rect 12896 8946 12932 8957
rect 14698 8946 14830 9054
rect 15767 9888 15887 9977
rect 11022 7541 11056 7573
rect 11056 7541 11123 7573
rect 11123 7541 11154 7573
rect 11022 7465 11154 7541
rect 13504 7594 13537 7627
rect 13537 7594 13604 7627
rect 13604 7594 13636 7627
rect 13504 7519 13636 7594
rect 13905 7529 13961 7543
rect 13905 7495 13921 7529
rect 13921 7495 13955 7529
rect 13955 7495 13961 7529
rect 13905 7477 13961 7495
rect 14651 7594 14685 7627
rect 14685 7594 14752 7627
rect 14752 7594 14783 7627
rect 14651 7519 14783 7594
rect 12775 7405 12841 7421
rect 12775 7371 12791 7405
rect 12791 7371 12825 7405
rect 12825 7371 12841 7405
rect 12775 7355 12841 7371
rect 9141 6721 9209 6796
rect 13441 6708 13540 6805
rect 11302 6490 11410 6534
rect 11302 6423 11394 6490
rect 11394 6423 11410 6490
rect 11302 6402 11410 6423
rect 7441 6130 7573 6227
rect 7441 6119 7474 6130
rect 7474 6119 7541 6130
rect 7541 6119 7573 6130
rect 6298 5474 6430 5582
rect 8196 5549 8228 5582
rect 8228 5549 8295 5582
rect 8295 5549 8328 5582
rect 8196 5474 8328 5549
rect 4020 4712 4138 4830
rect 4765 4846 4873 4886
rect 4765 4779 4852 4846
rect 4852 4779 4873 4846
rect 4765 4754 4873 4779
rect 3517 4370 3610 4449
rect 16 4044 103 4125
rect 369 4056 450 4119
rect -650 3865 -594 3919
rect -650 1803 -594 1857
rect -3257 1691 -3191 1757
rect -3060 1704 -3001 1769
rect -4059 939 -4005 949
rect -4059 901 -4051 939
rect -4051 901 -4013 939
rect -4013 901 -4005 939
rect -4059 895 -4005 901
rect -1835 1001 -1777 1007
rect -1835 951 -1829 1001
rect -1829 951 -1787 1001
rect -1787 951 -1777 1001
rect -1835 945 -1777 951
rect 1700 3727 1762 3735
rect 1700 3681 1706 3727
rect 1706 3681 1758 3727
rect 1758 3681 1762 3727
rect 1700 3675 1762 3681
rect 4480 4291 4511 4321
rect 4511 4291 4578 4321
rect 4578 4291 4612 4321
rect 4480 4213 4612 4291
rect 6943 4596 7006 4612
rect 6943 4562 6972 4596
rect 6972 4562 7006 4596
rect 6943 4546 7006 4562
rect 5067 3518 5130 3570
rect 4760 3254 4868 3282
rect 4760 3187 4852 3254
rect 4852 3187 4868 3254
rect 4760 3150 4868 3187
rect 4022 2935 4134 3041
rect 6243 3086 6375 3186
rect 6243 3078 6273 3086
rect 6273 3078 6340 3086
rect 6340 3078 6375 3086
rect 8141 3078 8273 3186
rect 9794 5824 9906 5930
rect 8410 2364 8472 2370
rect 8410 2318 8416 2364
rect 8416 2318 8468 2364
rect 8468 2318 8472 2364
rect 8410 2310 8472 2318
rect 7471 2045 7547 2131
rect 7702 1913 7831 2004
rect 12850 6132 12982 6227
rect 12850 6119 12879 6132
rect 12879 6119 12946 6132
rect 12946 6119 12982 6132
rect 10288 5841 10400 5947
rect 11036 5897 11067 5923
rect 11067 5897 11134 5923
rect 11134 5897 11168 5923
rect 11036 5815 11168 5897
rect 14597 6731 14662 6785
rect 17682 13341 17715 13375
rect 17715 13341 17782 13375
rect 17782 13341 17814 13375
rect 17682 13267 17814 13341
rect 20164 13397 20196 13429
rect 20196 13397 20263 13429
rect 20263 13397 20296 13429
rect 20164 13321 20296 13397
rect 20565 13331 20621 13345
rect 20565 13297 20581 13331
rect 20581 13297 20615 13331
rect 20615 13297 20621 13331
rect 20565 13279 20621 13297
rect 21311 13396 21343 13429
rect 21343 13396 21410 13429
rect 21410 13396 21443 13429
rect 21311 13321 21443 13396
rect 19435 13207 19501 13223
rect 19435 13173 19451 13207
rect 19451 13173 19485 13207
rect 19485 13173 19501 13207
rect 19435 13157 19501 13173
rect 20101 12510 20200 12607
rect 17962 12299 18070 12336
rect 17962 12232 18050 12299
rect 18050 12232 18070 12299
rect 17962 12204 18070 12232
rect 16453 10618 16565 10620
rect 16453 10514 16571 10618
rect 16459 10513 16571 10514
rect 16459 10512 16571 10513
rect 19510 11936 19642 12029
rect 19510 11921 19538 11936
rect 19538 11921 19605 11936
rect 19605 11921 19642 11936
rect 16948 11643 17060 11749
rect 17696 11693 17730 11725
rect 17730 11693 17797 11725
rect 17797 11693 17828 11725
rect 17696 11617 17828 11693
rect 21257 12533 21322 12587
rect 24307 13410 24335 13443
rect 24335 13410 24402 13443
rect 24402 13410 24439 13443
rect 24307 13335 24439 13410
rect 26789 13462 26819 13497
rect 26819 13462 26886 13497
rect 26886 13462 26921 13497
rect 26789 13389 26921 13462
rect 27190 13399 27246 13413
rect 27190 13365 27206 13399
rect 27206 13365 27240 13399
rect 27240 13365 27246 13399
rect 27190 13347 27246 13365
rect 27936 13468 27968 13497
rect 27968 13468 28035 13497
rect 28035 13468 28068 13497
rect 27936 13389 28068 13468
rect 26060 13275 26126 13291
rect 26060 13241 26076 13275
rect 26076 13241 26110 13275
rect 26110 13241 26126 13275
rect 26060 13225 26126 13241
rect 26726 12578 26825 12675
rect 24587 12375 24695 12404
rect 24587 12308 24682 12375
rect 24682 12308 24695 12375
rect 24587 12272 24695 12308
rect 20652 11939 20784 12027
rect 20652 11919 20684 11939
rect 20684 11919 20751 11939
rect 20751 11919 20784 11939
rect 23079 11694 23191 11800
rect 19509 11274 19641 11382
rect 21407 11345 21437 11382
rect 21437 11345 21504 11382
rect 21504 11345 21539 11382
rect 21407 11274 21539 11345
rect 17231 10512 17349 10630
rect 17976 10648 18084 10686
rect 17976 10581 18067 10648
rect 18067 10581 18084 10648
rect 17976 10554 18084 10581
rect 16728 10170 16821 10249
rect 17691 10090 17725 10121
rect 17725 10090 17792 10121
rect 17792 10090 17823 10121
rect 17691 10013 17823 10090
rect 20154 10396 20217 10412
rect 20154 10362 20183 10396
rect 20183 10362 20217 10396
rect 20154 10346 20217 10362
rect 18278 9318 18341 9370
rect 17971 9043 18079 9082
rect 17971 8976 18069 9043
rect 18069 8976 18079 9043
rect 17971 8950 18079 8976
rect 17233 8735 17345 8841
rect 19454 8891 19586 8986
rect 19454 8878 19478 8891
rect 19478 8878 19545 8891
rect 19545 8878 19586 8891
rect 21352 8878 21484 8986
rect 22405 8590 22528 8599
rect 22405 8491 22414 8590
rect 22414 8491 22520 8590
rect 22520 8491 22528 8590
rect 22405 8485 22528 8491
rect 17677 7538 17707 7574
rect 17707 7538 17774 7574
rect 17774 7538 17809 7574
rect 17677 7466 17809 7538
rect 20159 7598 20192 7628
rect 20192 7598 20259 7628
rect 20259 7598 20291 7628
rect 20159 7520 20291 7598
rect 20560 7530 20616 7544
rect 20560 7496 20576 7530
rect 20576 7496 20610 7530
rect 20610 7496 20616 7530
rect 20560 7478 20616 7496
rect 21306 7595 21341 7628
rect 21341 7595 21408 7628
rect 21408 7595 21438 7628
rect 21306 7520 21438 7595
rect 19430 7406 19496 7422
rect 19430 7372 19446 7406
rect 19446 7372 19480 7406
rect 19480 7372 19496 7406
rect 19430 7356 19496 7372
rect 20096 6709 20195 6806
rect 17957 6499 18065 6535
rect 17957 6432 18055 6499
rect 18055 6432 18065 6499
rect 17957 6403 18065 6432
rect 13992 6121 14124 6225
rect 13992 6117 14020 6121
rect 14020 6117 14087 6121
rect 14087 6117 14124 6121
rect 16382 5823 16586 5936
rect 16534 5822 16586 5823
rect 12849 5472 12981 5580
rect 14747 5548 14784 5580
rect 14784 5548 14851 5580
rect 14851 5548 14879 5580
rect 14747 5472 14879 5548
rect 10571 4710 10689 4828
rect 11316 4845 11424 4884
rect 11316 4778 11410 4845
rect 11410 4778 11424 4845
rect 11316 4752 11424 4778
rect 10068 4368 10161 4447
rect 11031 4286 11067 4319
rect 11067 4286 11134 4319
rect 11134 4286 11163 4319
rect 11031 4211 11163 4286
rect 13494 4594 13557 4610
rect 13494 4560 13523 4594
rect 13523 4560 13557 4594
rect 13494 4544 13557 4560
rect 11618 3516 11681 3568
rect 11311 3245 11419 3280
rect 11311 3178 11399 3245
rect 11399 3178 11419 3245
rect 11311 3148 11419 3178
rect 10573 2933 10685 3039
rect 12794 3085 12926 3184
rect 12794 3076 12821 3085
rect 12821 3076 12888 3085
rect 12888 3076 12926 3085
rect 14692 3076 14824 3184
rect 14964 2369 15026 2375
rect 14964 2323 14970 2369
rect 14970 2323 15022 2369
rect 15022 2323 15026 2369
rect 14964 2315 15026 2323
rect 8188 1106 8248 1168
rect -3251 315 -3197 369
rect 19505 6136 19637 6228
rect 19505 6120 19531 6136
rect 19531 6120 19598 6136
rect 19598 6120 19637 6136
rect 16943 5842 17055 5948
rect 17691 5892 17727 5924
rect 17727 5892 17794 5924
rect 17794 5892 17823 5924
rect 17691 5816 17823 5892
rect 21252 6732 21317 6786
rect 26135 11995 26267 12097
rect 26135 11989 26159 11995
rect 26159 11989 26226 11995
rect 26226 11989 26267 11995
rect 23573 11711 23685 11817
rect 24321 11759 24358 11793
rect 24358 11759 24425 11793
rect 24425 11759 24453 11793
rect 24321 11685 24453 11759
rect 27882 12601 27947 12655
rect 28860 12589 28928 12664
rect 27277 11997 27409 12095
rect 27277 11987 27302 11997
rect 27302 11987 27369 11997
rect 27369 11987 27409 11997
rect 26134 11342 26266 11450
rect 28032 11414 28065 11450
rect 28065 11414 28132 11450
rect 28132 11414 28164 11450
rect 28032 11342 28164 11414
rect 23856 10580 23974 10698
rect 24601 10714 24709 10754
rect 24601 10647 24687 10714
rect 24687 10647 24709 10714
rect 24601 10622 24709 10647
rect 23353 10238 23446 10317
rect 22874 9811 22970 9911
rect 24316 10151 24350 10189
rect 24350 10151 24417 10189
rect 24417 10151 24448 10189
rect 24316 10081 24448 10151
rect 26779 10464 26842 10480
rect 26779 10430 26808 10464
rect 26808 10430 26842 10464
rect 26779 10414 26842 10430
rect 24903 9386 24966 9438
rect 24596 9109 24704 9150
rect 24596 9042 24693 9109
rect 24693 9042 24704 9109
rect 24596 9018 24704 9042
rect 23858 8803 23970 8909
rect 26079 8957 26211 9054
rect 26079 8946 26109 8957
rect 26109 8946 26176 8957
rect 26176 8946 26211 8957
rect 27977 8946 28109 9054
rect 30009 15253 30069 15315
rect 32266 15210 32398 15244
rect 32266 15136 32398 15210
rect 33610 14845 33670 14907
rect 29354 14168 29433 14242
rect 29506 14032 29587 14128
rect 31463 14267 31530 14330
rect 30231 14103 30293 14111
rect 30231 14057 30237 14103
rect 30237 14057 30289 14103
rect 30289 14057 30293 14103
rect 30231 14051 30293 14057
rect 31463 14141 31530 14204
rect 30004 12682 30064 12744
rect 31723 14195 31778 14212
rect 31723 14161 31728 14195
rect 31728 14161 31762 14195
rect 31762 14161 31778 14195
rect 31723 14144 31778 14161
rect 32777 13883 32839 13974
rect 33119 14314 33172 14325
rect 33119 14280 33128 14314
rect 33128 14280 33162 14314
rect 33162 14280 33172 14314
rect 33119 14269 33172 14280
rect 33243 14133 33316 14222
rect 34232 14159 34344 14217
rect 34016 13888 34124 13969
rect 33832 13695 33894 13703
rect 33832 13649 33838 13695
rect 33838 13649 33890 13695
rect 33890 13649 33894 13695
rect 33832 13643 33894 13649
rect 32196 12900 32370 12909
rect 32196 12798 32215 12900
rect 32215 12798 32350 12900
rect 32350 12798 32370 12900
rect 32196 12786 32370 12798
rect 29653 11720 29735 11801
rect 30226 11532 30288 11540
rect 30226 11486 30232 11532
rect 30232 11486 30284 11532
rect 30284 11486 30288 11532
rect 30226 11480 30288 11486
rect 32268 11119 32400 11153
rect 32268 11045 32400 11119
rect 33612 10754 33672 10816
rect 31465 10176 31532 10239
rect 30004 9649 30064 9711
rect 29758 8813 29847 8900
rect 23514 8590 23637 8599
rect 23514 8491 23523 8590
rect 23523 8491 23629 8590
rect 23629 8491 23637 8590
rect 23514 8485 23637 8491
rect 31465 10050 31532 10113
rect 30226 8499 30288 8507
rect 30226 8453 30232 8499
rect 30232 8453 30284 8499
rect 30284 8453 30288 8499
rect 30226 8447 30288 8453
rect 30075 7729 30135 7791
rect 24299 7543 24331 7575
rect 24331 7543 24398 7575
rect 24398 7543 24431 7575
rect 24299 7467 24431 7543
rect 26781 7591 26810 7629
rect 26810 7591 26877 7629
rect 26877 7591 26913 7629
rect 26781 7521 26913 7591
rect 27182 7531 27238 7545
rect 27182 7497 27198 7531
rect 27198 7497 27232 7531
rect 27232 7497 27238 7531
rect 27182 7479 27238 7497
rect 27928 7597 27958 7629
rect 27958 7597 28025 7629
rect 28025 7597 28060 7629
rect 27928 7521 28060 7597
rect 26052 7407 26118 7423
rect 26052 7373 26068 7407
rect 26068 7373 26102 7407
rect 26102 7373 26118 7407
rect 26052 7357 26118 7373
rect 22347 6720 22415 6795
rect 26718 6710 26817 6807
rect 24579 6504 24687 6536
rect 24579 6437 24671 6504
rect 24671 6437 24687 6504
rect 24579 6404 24687 6437
rect 20647 6139 20779 6226
rect 20647 6118 20677 6139
rect 20677 6118 20744 6139
rect 20744 6118 20779 6139
rect 19504 5473 19636 5581
rect 21402 5550 21438 5581
rect 21438 5550 21505 5581
rect 21505 5550 21534 5581
rect 21402 5473 21534 5550
rect 17226 4711 17344 4829
rect 17971 4848 18079 4885
rect 17971 4781 18066 4848
rect 18066 4781 18079 4848
rect 17971 4753 18079 4781
rect 16723 4369 16816 4448
rect 17686 4284 17722 4320
rect 17722 4284 17789 4320
rect 17789 4284 17818 4320
rect 17686 4212 17818 4284
rect 20149 4595 20212 4611
rect 20149 4561 20178 4595
rect 20178 4561 20212 4595
rect 20149 4545 20212 4561
rect 18273 3517 18336 3569
rect 17966 3239 18074 3281
rect 17966 3172 18069 3239
rect 18069 3172 18074 3239
rect 17966 3149 18074 3172
rect 16411 2990 16513 3002
rect 16411 2922 16430 2990
rect 16430 2922 16500 2990
rect 16500 2922 16513 2990
rect 16411 2915 16513 2922
rect 17228 2934 17340 3040
rect 19449 3086 19581 3185
rect 19449 3077 19471 3086
rect 19471 3077 19538 3086
rect 19538 3077 19581 3086
rect 21347 3077 21479 3185
rect 23071 5826 23183 5932
rect 21613 2357 21675 2363
rect 21613 2311 21619 2357
rect 21619 2311 21671 2357
rect 21671 2311 21675 2357
rect 21613 2303 21675 2311
rect 14742 1111 14802 1173
rect 20899 1906 20968 1995
rect 23070 4818 23182 4820
rect 23070 4714 23188 4818
rect 23076 4712 23188 4714
rect 26127 6140 26259 6229
rect 26127 6121 26162 6140
rect 26162 6121 26229 6140
rect 26229 6121 26259 6140
rect 23565 5843 23677 5949
rect 24313 5893 24346 5925
rect 24346 5893 24413 5925
rect 24413 5893 24445 5925
rect 24313 5817 24445 5893
rect 31725 10104 31780 10121
rect 31725 10070 31730 10104
rect 31730 10070 31764 10104
rect 31764 10070 31780 10104
rect 31725 10053 31780 10070
rect 32779 9792 32841 9883
rect 33121 10223 33174 10234
rect 33121 10189 33130 10223
rect 33130 10189 33164 10223
rect 33164 10189 33174 10223
rect 33121 10178 33174 10189
rect 33245 10042 33318 10131
rect 33834 9604 33896 9612
rect 33834 9558 33840 9604
rect 33840 9558 33892 9604
rect 33892 9558 33896 9604
rect 33834 9552 33896 9558
rect 32198 8809 32372 8818
rect 32198 8707 32217 8809
rect 32217 8707 32352 8809
rect 32352 8707 32372 8809
rect 32198 8695 32372 8707
rect 32268 7624 32400 7658
rect 32268 7550 32400 7624
rect 27874 6733 27939 6787
rect 29810 6678 29896 6779
rect 33612 7259 33672 7321
rect 29582 6545 29667 6605
rect 30297 6579 30359 6587
rect 30297 6533 30303 6579
rect 30303 6533 30355 6579
rect 30355 6533 30359 6579
rect 30297 6527 30359 6533
rect 31465 6555 31532 6618
rect 27269 6131 27401 6227
rect 27269 6119 27296 6131
rect 27296 6119 27363 6131
rect 27363 6119 27401 6131
rect 26126 5474 26258 5582
rect 28024 5548 28059 5582
rect 28059 5548 28126 5582
rect 28126 5548 28156 5582
rect 28024 5474 28156 5548
rect 23848 4712 23966 4830
rect 24593 4855 24701 4886
rect 24593 4788 24689 4855
rect 24689 4788 24701 4855
rect 24593 4754 24701 4788
rect 23345 4370 23438 4449
rect 24308 4284 24343 4321
rect 24343 4284 24410 4321
rect 24410 4284 24440 4321
rect 24308 4213 24440 4284
rect 26771 4596 26834 4612
rect 26771 4562 26800 4596
rect 26800 4562 26834 4596
rect 26771 4546 26834 4562
rect 30072 4659 30132 4721
rect 24895 3518 24958 3570
rect 24588 3238 24696 3282
rect 24588 3171 24680 3238
rect 24680 3171 24696 3238
rect 24588 3150 24696 3171
rect 23850 2935 23962 3041
rect 26071 3092 26203 3186
rect 26071 3078 26099 3092
rect 26099 3078 26166 3092
rect 26166 3078 26203 3092
rect 27969 3078 28101 3186
rect 29037 4023 29154 4104
rect 31725 6609 31780 6626
rect 31725 6575 31730 6609
rect 31730 6575 31764 6609
rect 31764 6575 31780 6609
rect 31725 6558 31780 6575
rect 32779 6297 32841 6388
rect 33121 6728 33174 6739
rect 33121 6694 33130 6728
rect 33130 6694 33164 6728
rect 33164 6694 33174 6728
rect 33121 6683 33174 6694
rect 33245 6547 33318 6636
rect 33834 6109 33896 6117
rect 33834 6063 33840 6109
rect 33840 6063 33892 6109
rect 33892 6063 33896 6109
rect 33834 6057 33896 6063
rect 32198 5314 32372 5323
rect 32198 5212 32217 5314
rect 32217 5212 32352 5314
rect 32352 5212 32372 5314
rect 32198 5200 32372 5212
rect 29412 3695 29496 3785
rect 34428 6375 34538 6387
rect 34428 6303 34434 6375
rect 34434 6303 34529 6375
rect 34529 6303 34538 6375
rect 34428 6296 34538 6303
rect 29846 3574 29912 3638
rect 30294 3509 30356 3517
rect 30294 3463 30300 3509
rect 30300 3463 30352 3509
rect 30352 3463 30356 3509
rect 30294 3457 30356 3463
rect 32268 3276 32400 3310
rect 32268 3202 32400 3276
rect 36507 17620 36567 17624
rect 36507 17548 36513 17620
rect 36513 17548 36567 17620
rect 36507 17544 36567 17548
rect 37450 18767 37513 18771
rect 37450 18707 37454 18767
rect 37454 18707 37509 18767
rect 37509 18707 37513 18767
rect 37450 18700 37513 18707
rect 37733 17800 37798 17804
rect 37733 17740 37738 17800
rect 37738 17740 37793 17800
rect 37793 17740 37798 17800
rect 37733 17736 37798 17740
rect 37450 17682 37512 17686
rect 37450 17622 37453 17682
rect 37453 17622 37508 17682
rect 37508 17622 37512 17682
rect 37450 17616 37512 17622
rect 38725 17606 38777 17610
rect 38725 17548 38771 17606
rect 38771 17548 38777 17606
rect 38725 17544 38777 17548
rect 37570 17432 37630 17445
rect 37570 17398 37584 17432
rect 37584 17398 37618 17432
rect 37618 17398 37630 17432
rect 37570 17386 37630 17398
rect 37565 15814 37633 15871
rect 36507 14476 36567 14480
rect 36507 14404 36513 14476
rect 36513 14404 36567 14476
rect 36507 14400 36567 14404
rect 37450 15623 37513 15627
rect 37450 15563 37454 15623
rect 37454 15563 37509 15623
rect 37509 15563 37513 15623
rect 37450 15556 37513 15563
rect 37733 14656 37798 14660
rect 37733 14596 37738 14656
rect 37738 14596 37793 14656
rect 37793 14596 37798 14656
rect 37733 14592 37798 14596
rect 37450 14538 37512 14542
rect 37450 14478 37453 14538
rect 37453 14478 37508 14538
rect 37508 14478 37512 14538
rect 37450 14472 37512 14478
rect 38725 14462 38777 14466
rect 38725 14404 38771 14462
rect 38771 14404 38777 14462
rect 38725 14400 38777 14404
rect 37570 14288 37630 14301
rect 37570 14254 37584 14288
rect 37584 14254 37618 14288
rect 37618 14254 37630 14288
rect 37570 14242 37630 14254
rect 37569 12612 37637 12669
rect 37737 12665 37805 12669
rect 37737 12616 37741 12665
rect 37741 12616 37801 12665
rect 37801 12616 37805 12665
rect 37737 12612 37805 12616
rect 36511 11274 36571 11278
rect 36511 11202 36517 11274
rect 36517 11202 36571 11274
rect 36511 11198 36571 11202
rect 37454 12421 37517 12425
rect 37454 12361 37458 12421
rect 37458 12361 37513 12421
rect 37513 12361 37517 12421
rect 37454 12354 37517 12361
rect 37737 11454 37802 11458
rect 37737 11394 37742 11454
rect 37742 11394 37797 11454
rect 37797 11394 37802 11454
rect 37737 11390 37802 11394
rect 37454 11336 37516 11340
rect 37454 11276 37457 11336
rect 37457 11276 37512 11336
rect 37512 11276 37516 11336
rect 37454 11270 37516 11276
rect 38729 11260 38781 11264
rect 38729 11202 38775 11260
rect 38775 11202 38781 11260
rect 38729 11198 38781 11202
rect 37574 11086 37634 11099
rect 37574 11052 37588 11086
rect 37588 11052 37622 11086
rect 37622 11052 37634 11086
rect 37574 11040 37634 11052
rect 37569 9468 37637 9525
rect 36511 8130 36571 8134
rect 36511 8058 36517 8130
rect 36517 8058 36571 8130
rect 36511 8054 36571 8058
rect 37454 9277 37517 9281
rect 37454 9217 37458 9277
rect 37458 9217 37513 9277
rect 37513 9217 37517 9277
rect 37454 9210 37517 9217
rect 37737 8310 37802 8314
rect 37737 8250 37742 8310
rect 37742 8250 37797 8310
rect 37797 8250 37802 8310
rect 37737 8246 37802 8250
rect 37454 8192 37516 8196
rect 37454 8132 37457 8192
rect 37457 8132 37512 8192
rect 37512 8132 37516 8192
rect 37454 8126 37516 8132
rect 38729 8116 38781 8120
rect 38729 8058 38775 8116
rect 38775 8058 38781 8116
rect 38729 8054 38781 8058
rect 37574 7942 37634 7955
rect 37574 7908 37588 7942
rect 37588 7908 37622 7942
rect 37622 7908 37634 7942
rect 37574 7896 37634 7908
rect 37565 6336 37633 6393
rect 37733 6389 37801 6393
rect 37733 6340 37737 6389
rect 37737 6340 37797 6389
rect 37797 6340 37801 6389
rect 37733 6336 37801 6340
rect 36507 4998 36567 5002
rect 36507 4926 36513 4998
rect 36513 4926 36567 4998
rect 36507 4922 36567 4926
rect 37450 6145 37513 6149
rect 37450 6085 37454 6145
rect 37454 6085 37509 6145
rect 37509 6085 37513 6145
rect 37450 6078 37513 6085
rect 37733 5178 37798 5182
rect 37733 5118 37738 5178
rect 37738 5118 37793 5178
rect 37793 5118 37798 5178
rect 37733 5114 37798 5118
rect 37450 5060 37512 5064
rect 37450 5000 37453 5060
rect 37453 5000 37508 5060
rect 37508 5000 37512 5060
rect 37450 4994 37512 5000
rect 38725 4984 38777 4988
rect 38725 4926 38771 4984
rect 38771 4926 38777 4984
rect 38725 4922 38777 4926
rect 37570 4810 37630 4823
rect 37570 4776 37584 4810
rect 37584 4776 37618 4810
rect 37618 4776 37630 4810
rect 37570 4764 37630 4776
rect 37565 3192 37633 3249
rect 37733 3245 37801 3249
rect 37733 3196 37737 3245
rect 37737 3196 37797 3245
rect 37797 3196 37801 3245
rect 37733 3192 37801 3196
rect 33612 2911 33672 2973
rect 31465 2333 31531 2396
rect 31531 2333 31532 2396
rect 31465 2207 31532 2270
rect 29826 2035 29910 2125
rect 21391 1099 21451 1161
rect 2616 819 2712 888
rect 7656 818 7756 892
rect 30079 1814 30139 1876
rect 502 690 601 776
rect 29241 1292 29325 1382
rect 31725 2261 31780 2278
rect 31725 2227 31730 2261
rect 31730 2227 31764 2261
rect 31764 2227 31780 2261
rect 31725 2210 31780 2227
rect 32779 1949 32841 2040
rect 33121 2380 33174 2391
rect 33121 2346 33130 2380
rect 33130 2346 33164 2380
rect 33164 2346 33174 2380
rect 33121 2335 33174 2346
rect 33245 2199 33318 2288
rect 34210 2211 34352 2299
rect 36507 1854 36567 1858
rect 36507 1782 36513 1854
rect 36513 1782 36567 1854
rect 36507 1778 36567 1782
rect 33834 1761 33896 1769
rect 33834 1715 33840 1761
rect 33840 1715 33892 1761
rect 33892 1715 33896 1761
rect 33834 1709 33896 1715
rect 7464 567 7556 639
rect 29410 976 29494 1066
rect 20896 564 20965 632
rect 29723 642 29784 717
rect 32198 966 32372 975
rect 32198 864 32217 966
rect 32217 864 32352 966
rect 32352 864 32372 966
rect 32198 852 32372 864
rect 37450 3001 37513 3005
rect 37450 2941 37454 3001
rect 37454 2941 37509 3001
rect 37509 2941 37513 3001
rect 37450 2934 37513 2941
rect 37733 2034 37798 2038
rect 37733 1974 37738 2034
rect 37738 1974 37793 2034
rect 37793 1974 37798 2034
rect 37733 1970 37798 1974
rect 37450 1916 37512 1920
rect 37450 1856 37453 1916
rect 37453 1856 37508 1916
rect 37508 1856 37512 1916
rect 37450 1850 37512 1856
rect 38725 1840 38777 1844
rect 38725 1782 38771 1840
rect 38771 1782 38777 1840
rect 38725 1778 38777 1782
rect 37570 1666 37630 1679
rect 37570 1632 37584 1666
rect 37584 1632 37618 1666
rect 37618 1632 37630 1666
rect 37570 1620 37630 1632
rect 30301 664 30363 672
rect 30301 618 30307 664
rect 30307 618 30359 664
rect 30359 618 30363 664
rect 30301 612 30363 618
rect 2462 156 2557 210
rect -2680 54 -2616 119
<< metal2 >>
rect 4376 28302 4535 28322
rect 4376 28180 4391 28302
rect 4522 28180 4535 28302
rect -845 23405 -661 23415
rect -845 23234 -661 23244
rect 4376 21521 4535 28180
rect 8754 27971 8907 27981
rect 6272 27917 6425 27927
rect 9901 27971 10054 27981
rect 9166 27876 9222 27886
rect 8754 27832 8907 27842
rect 6272 27778 6425 27788
rect 9041 27810 9166 27872
rect 9222 27810 9223 27872
rect 15267 27968 15420 27978
rect 9901 27832 10054 27842
rect 12785 27914 12938 27924
rect 8036 27761 8102 27764
rect 7110 27754 8102 27761
rect 7110 27688 8036 27754
rect 6543 26725 6553 26878
rect 6682 26725 6692 26878
rect 5069 26290 5282 26291
rect 5550 26290 5666 26291
rect 5069 26280 5666 26290
rect 5069 26268 5549 26280
rect 5069 26165 5091 26268
rect 5233 26174 5549 26268
rect 5661 26174 5666 26280
rect 5233 26165 5666 26174
rect 5069 26148 5666 26165
rect 6286 26267 6439 26277
rect 5069 26147 5282 26148
rect 6286 26128 6439 26138
rect 5051 25169 5189 25173
rect 5045 25168 5294 25169
rect 5832 25168 5950 25171
rect 5045 25163 5950 25168
rect 5045 25037 5051 25163
rect 5189 25161 5950 25163
rect 5189 25043 5832 25161
rect 6557 25075 6567 25228
rect 6696 25075 6706 25228
rect 5189 25037 5950 25043
rect 5045 25033 5950 25037
rect 5051 25027 5189 25033
rect 5319 24789 5434 24799
rect 5319 24682 5434 24692
rect 5829 23382 5945 25033
rect 6281 24663 6434 24673
rect 6281 24524 6434 24534
rect 6879 23905 6942 23911
rect 7110 23905 7178 27688
rect 8036 27678 8102 27688
rect 9041 27149 9101 27810
rect 9166 27800 9222 27810
rect 16414 27968 16567 27978
rect 15679 27873 15735 27883
rect 15267 27829 15420 27839
rect 12785 27775 12938 27785
rect 15554 27807 15679 27869
rect 15735 27807 15736 27869
rect 21801 27963 21954 27973
rect 16414 27829 16567 27839
rect 19319 27909 19472 27919
rect 14549 27758 14615 27761
rect 8963 27148 9101 27149
rect 8701 27138 9101 27148
rect 8701 27041 8702 27138
rect 8801 27041 9101 27138
rect 13623 27751 14615 27758
rect 13623 27685 14549 27751
rect 9858 27127 9923 27128
rect 10953 27127 11021 27137
rect 9857 27118 10953 27127
rect 9857 27064 9858 27118
rect 9923 27064 10953 27118
rect 9857 27053 10953 27064
rect 10953 27042 11021 27052
rect 8701 27033 9101 27041
rect 8701 27029 9010 27033
rect 11249 26864 11382 26865
rect 11249 26838 11692 26864
rect 11249 26694 11432 26838
rect 11668 26694 11692 26838
rect 13056 26722 13066 26875
rect 13195 26722 13205 26875
rect 11249 26670 11692 26694
rect 8101 26570 8254 26580
rect 8101 26431 8254 26441
rect 9243 26568 9396 26578
rect 9243 26429 9396 26439
rect 8099 25924 8252 25934
rect 8099 25785 8252 25795
rect 9997 25924 10150 25934
rect 9997 25785 10150 25795
rect 8740 24953 8818 24963
rect 8740 24857 8818 24867
rect 6874 23901 7178 23905
rect 6874 23849 6879 23901
rect 6942 23849 7178 23901
rect 6874 23843 7178 23849
rect 6879 23839 6942 23843
rect 6552 23471 6562 23624
rect 6691 23471 6701 23624
rect 8045 23527 8198 23537
rect 8045 23388 8198 23398
rect 9943 23527 10096 23537
rect 9943 23388 10096 23398
rect 5829 23372 5946 23382
rect 5829 23266 5834 23372
rect 5829 23256 5946 23266
rect 5829 23255 5945 23256
rect 11249 23072 11413 26670
rect 11495 26294 11775 26317
rect 11495 26170 11523 26294
rect 11752 26287 11775 26294
rect 12063 26287 12179 26288
rect 11752 26277 12179 26287
rect 11752 26171 12062 26277
rect 12174 26171 12179 26277
rect 11752 26170 12179 26171
rect 11495 26145 12179 26170
rect 12799 26264 12952 26274
rect 11495 26144 11775 26145
rect 12799 26125 12952 26135
rect 11555 25166 11720 25176
rect 11555 25165 11723 25166
rect 12345 25165 12463 25168
rect 11555 25158 12463 25165
rect 11555 25148 12345 25158
rect 11555 25042 11567 25148
rect 11679 25146 12345 25148
rect 11555 25040 11573 25042
rect 11685 25040 12345 25146
rect 13070 25072 13080 25225
rect 13209 25072 13219 25225
rect 11555 25033 12463 25040
rect 11561 25031 12463 25033
rect 11598 25030 12463 25031
rect 11832 24786 11947 24796
rect 11832 24679 11947 24689
rect 12342 23379 12458 25030
rect 12794 24660 12947 24670
rect 12794 24521 12947 24531
rect 13392 23902 13455 23908
rect 13623 23902 13691 27685
rect 14549 27675 14615 27685
rect 15554 27146 15614 27807
rect 15679 27797 15735 27807
rect 22948 27963 23101 27973
rect 22213 27868 22269 27878
rect 21801 27824 21954 27834
rect 19319 27770 19472 27780
rect 22088 27802 22213 27864
rect 22269 27802 22270 27864
rect 28359 27967 28512 27977
rect 22948 27824 23101 27834
rect 25877 27913 26030 27923
rect 21083 27753 21149 27756
rect 15476 27145 15614 27146
rect 15214 27135 15614 27145
rect 15214 27038 15215 27135
rect 15314 27038 15614 27135
rect 20157 27746 21149 27753
rect 20157 27680 21083 27746
rect 16371 27124 16436 27125
rect 17466 27124 17534 27134
rect 16370 27115 17466 27124
rect 16370 27061 16371 27115
rect 16436 27061 17466 27115
rect 16370 27050 17466 27061
rect 17466 27039 17534 27049
rect 15214 27030 15614 27038
rect 15214 27026 15523 27030
rect 17766 26845 18221 26864
rect 17766 26688 17969 26845
rect 18202 26688 18221 26845
rect 19590 26717 19600 26870
rect 19729 26717 19739 26870
rect 17766 26665 18221 26688
rect 14614 26567 14767 26577
rect 14614 26428 14767 26438
rect 15756 26565 15909 26575
rect 15756 26426 15909 26436
rect 14612 25921 14765 25931
rect 14612 25782 14765 25792
rect 16510 25921 16663 25931
rect 16510 25782 16663 25792
rect 15253 24950 15331 24960
rect 15253 24854 15331 24864
rect 13387 23898 13691 23902
rect 13387 23846 13392 23898
rect 13455 23846 13691 23898
rect 13387 23840 13691 23846
rect 13392 23836 13455 23840
rect 13065 23468 13075 23621
rect 13204 23468 13214 23621
rect 14558 23524 14711 23534
rect 14558 23385 14711 23395
rect 16456 23524 16609 23534
rect 16456 23385 16609 23395
rect 12342 23369 12459 23379
rect 12342 23263 12347 23369
rect 12342 23253 12459 23263
rect 12342 23252 12458 23253
rect 11249 22994 11268 23072
rect 11396 22994 11413 23072
rect 11249 22982 11413 22994
rect 17766 22921 17913 26665
rect 18149 26664 18221 26665
rect 18105 26317 18331 26318
rect 18056 26300 18331 26317
rect 18056 26160 18082 26300
rect 18300 26282 18331 26300
rect 18597 26282 18713 26283
rect 18300 26272 18713 26282
rect 18300 26166 18596 26272
rect 18708 26166 18713 26272
rect 18300 26160 18713 26166
rect 18056 26140 18713 26160
rect 19333 26259 19486 26269
rect 18056 26139 18315 26140
rect 19333 26120 19486 26130
rect 18089 25161 18254 25171
rect 18089 25160 18257 25161
rect 18879 25160 18997 25163
rect 18089 25153 18997 25160
rect 18089 25143 18879 25153
rect 18089 25037 18101 25143
rect 18213 25141 18879 25143
rect 18089 25035 18107 25037
rect 18219 25035 18879 25141
rect 19604 25067 19614 25220
rect 19743 25067 19753 25220
rect 18089 25028 18997 25035
rect 18095 25026 18997 25028
rect 18132 25025 18997 25026
rect 18366 24781 18481 24791
rect 18366 24674 18481 24684
rect 18876 23374 18992 25025
rect 19328 24655 19481 24665
rect 19328 24516 19481 24526
rect 19926 23897 19989 23903
rect 20157 23897 20225 27680
rect 21083 27670 21149 27680
rect 22088 27141 22148 27802
rect 22213 27792 22269 27802
rect 29506 27967 29659 27977
rect 28771 27872 28827 27882
rect 28359 27828 28512 27838
rect 25877 27774 26030 27784
rect 28646 27806 28771 27868
rect 28827 27806 28828 27868
rect 29506 27828 29659 27838
rect 27641 27757 27707 27760
rect 22010 27140 22148 27141
rect 21748 27130 22148 27140
rect 21748 27033 21749 27130
rect 21848 27033 22148 27130
rect 26715 27750 27707 27757
rect 26715 27684 27641 27750
rect 22905 27119 22970 27120
rect 24000 27119 24068 27129
rect 22904 27110 24000 27119
rect 22904 27056 22905 27110
rect 22970 27056 24000 27110
rect 22904 27045 24000 27056
rect 24000 27034 24068 27044
rect 21748 27025 22148 27033
rect 21748 27021 22057 27025
rect 24692 26865 24786 26866
rect 24354 26846 24786 26865
rect 24354 26683 24529 26846
rect 24776 26683 24786 26846
rect 26148 26721 26158 26874
rect 26287 26721 26297 26874
rect 24354 26669 24786 26683
rect 24354 26668 24768 26669
rect 21148 26562 21301 26572
rect 21148 26423 21301 26433
rect 22290 26560 22443 26570
rect 22290 26421 22443 26431
rect 21146 25916 21299 25926
rect 21146 25777 21299 25787
rect 23044 25916 23197 25926
rect 23044 25777 23197 25787
rect 21787 24945 21865 24955
rect 21787 24849 21865 24859
rect 19921 23893 20225 23897
rect 19921 23841 19926 23893
rect 19989 23841 20225 23893
rect 19921 23835 20225 23841
rect 19926 23831 19989 23835
rect 19599 23463 19609 23616
rect 19738 23463 19748 23616
rect 21092 23519 21245 23529
rect 21092 23380 21245 23390
rect 22990 23519 23143 23529
rect 22990 23380 23143 23390
rect 18876 23364 18993 23374
rect 18876 23258 18881 23364
rect 18876 23248 18993 23258
rect 18876 23247 18992 23248
rect 17766 22810 17781 22921
rect 17892 22810 17913 22921
rect 17766 22797 17913 22810
rect 24354 22738 24513 26668
rect 24588 26302 24884 26322
rect 24588 26157 24606 26302
rect 24858 26286 24884 26302
rect 25155 26286 25271 26287
rect 24858 26276 25271 26286
rect 24858 26170 25154 26276
rect 25266 26170 25271 26276
rect 24858 26157 25271 26170
rect 24588 26144 25271 26157
rect 25891 26263 26044 26273
rect 25891 26124 26044 26134
rect 24647 25165 24812 25175
rect 24647 25164 24815 25165
rect 25437 25164 25555 25167
rect 24647 25157 25555 25164
rect 24647 25147 25437 25157
rect 24647 25041 24659 25147
rect 24771 25145 25437 25147
rect 24647 25039 24665 25041
rect 24777 25039 25437 25145
rect 26162 25071 26172 25224
rect 26301 25071 26311 25224
rect 24647 25032 25555 25039
rect 24653 25030 25555 25032
rect 24690 25029 25555 25030
rect 24924 24785 25039 24795
rect 24924 24678 25039 24688
rect 25434 23378 25550 25029
rect 25886 24659 26039 24669
rect 25886 24520 26039 24530
rect 26484 23901 26547 23907
rect 26715 23901 26783 27684
rect 27641 27674 27707 27684
rect 28646 27145 28706 27806
rect 28771 27796 28827 27806
rect 28568 27144 28706 27145
rect 28306 27134 28706 27144
rect 28306 27037 28307 27134
rect 28406 27037 28706 27134
rect 29463 27123 29528 27124
rect 30558 27123 30626 27133
rect 29462 27114 30558 27123
rect 29462 27060 29463 27114
rect 29528 27060 30558 27114
rect 29462 27049 30558 27060
rect 30558 27038 30626 27048
rect 28306 27029 28706 27037
rect 28306 27025 28615 27029
rect 27706 26566 27859 26576
rect 27706 26427 27859 26437
rect 28848 26564 29001 26574
rect 28848 26425 29001 26435
rect 27704 25920 27857 25930
rect 27704 25781 27857 25791
rect 29602 25920 29755 25930
rect 29602 25781 29755 25791
rect 35009 25294 37482 25295
rect 35009 25207 37528 25294
rect 37561 25291 37646 25302
rect 37728 25291 37813 25302
rect 37559 25234 37569 25291
rect 37637 25234 37647 25291
rect 37727 25234 37737 25291
rect 37805 25234 37815 25291
rect 28345 24949 28423 24959
rect 28345 24853 28423 24863
rect 26479 23897 26783 23901
rect 26479 23845 26484 23897
rect 26547 23845 26783 23897
rect 26479 23839 26783 23845
rect 26484 23835 26547 23839
rect 26157 23467 26167 23620
rect 26296 23467 26306 23620
rect 27650 23523 27803 23533
rect 27650 23384 27803 23394
rect 29548 23523 29701 23533
rect 29548 23384 29701 23394
rect 25434 23368 25551 23378
rect 25434 23262 25439 23368
rect 25434 23252 25551 23262
rect 25434 23251 25550 23252
rect 24354 22620 24369 22738
rect 24503 22620 24513 22738
rect 24354 22606 24513 22620
rect 5850 22363 6003 22373
rect 6997 22363 7150 22373
rect 6682 22268 6738 22278
rect 5850 22224 6003 22234
rect 6681 22202 6682 22264
rect 6738 22202 6863 22264
rect 12408 22359 12561 22369
rect 6997 22224 7150 22234
rect 9479 22309 9632 22319
rect 6682 22192 6738 22202
rect 6803 21541 6863 22202
rect 13555 22359 13708 22369
rect 13240 22264 13296 22274
rect 12408 22220 12561 22230
rect 13239 22198 13240 22260
rect 13296 22198 13421 22260
rect 18942 22364 19095 22374
rect 13555 22220 13708 22230
rect 16037 22305 16190 22315
rect 13240 22188 13296 22198
rect 9479 22170 9632 22180
rect 7802 22153 7868 22156
rect 7802 22146 8794 22153
rect 7868 22080 8794 22146
rect 7802 22070 7868 22080
rect 6803 21540 6941 21541
rect 6803 21530 7203 21540
rect 4376 21519 5127 21521
rect 5981 21519 6046 21520
rect 4376 21510 6047 21519
rect 4376 21466 5981 21510
rect 4375 21456 5981 21466
rect 6046 21456 6047 21510
rect 4375 21445 6047 21456
rect 4375 21357 5409 21445
rect 6803 21433 7103 21530
rect 7202 21433 7203 21530
rect 6803 21425 7203 21433
rect 6894 21421 7203 21425
rect 6508 20960 6661 20970
rect 6508 20821 6661 20831
rect 7650 20962 7803 20972
rect 7650 20823 7803 20833
rect 5754 20316 5907 20326
rect 5754 20177 5907 20187
rect 7652 20316 7805 20326
rect 7652 20177 7805 20187
rect 7086 19345 7164 19355
rect 7086 19249 7164 19259
rect 8726 18297 8794 22080
rect 13361 21537 13421 22198
rect 20089 22364 20242 22374
rect 19774 22269 19830 22279
rect 18942 22225 19095 22235
rect 19773 22203 19774 22265
rect 19830 22203 19955 22265
rect 25455 22367 25608 22377
rect 20089 22225 20242 22235
rect 22571 22310 22724 22320
rect 19774 22193 19830 22203
rect 16037 22166 16190 22176
rect 14360 22149 14426 22152
rect 14360 22142 15352 22149
rect 14426 22076 15352 22142
rect 14360 22066 14426 22076
rect 13361 21536 13499 21537
rect 13361 21526 13761 21536
rect 11441 21515 11509 21525
rect 12539 21515 12604 21516
rect 11509 21506 12605 21515
rect 11509 21452 12539 21506
rect 12604 21452 12605 21506
rect 11509 21441 12605 21452
rect 11441 21430 11509 21440
rect 13361 21429 13661 21526
rect 13760 21429 13761 21526
rect 13361 21421 13761 21429
rect 13452 21417 13761 21421
rect 9212 21117 9222 21270
rect 9351 21117 9361 21270
rect 10731 21219 11142 21238
rect 10731 21083 10755 21219
rect 10979 21083 11142 21219
rect 10731 21065 11142 21083
rect 10238 20682 10354 20683
rect 10694 20682 10861 20683
rect 10238 20672 10861 20682
rect 9465 20659 9618 20669
rect 10238 20566 10243 20672
rect 10355 20655 10861 20672
rect 10355 20566 10737 20655
rect 10238 20549 10737 20566
rect 10849 20549 10861 20655
rect 10238 20540 10861 20549
rect 9465 20520 9618 20530
rect 9198 19467 9208 19620
rect 9337 19467 9347 19620
rect 9954 19560 10072 19563
rect 10697 19561 10862 19571
rect 10694 19560 10862 19561
rect 9954 19553 10862 19560
rect 10072 19543 10862 19553
rect 10072 19541 10738 19543
rect 10072 19435 10732 19541
rect 10850 19437 10862 19543
rect 10844 19435 10862 19437
rect 9954 19428 10862 19435
rect 9954 19426 10856 19428
rect 9954 19425 10819 19426
rect 9470 19055 9623 19065
rect 9470 18916 9623 18926
rect 8962 18297 9025 18303
rect 8726 18293 9030 18297
rect 8726 18241 8962 18293
rect 9025 18241 9030 18293
rect 8726 18235 9030 18241
rect 8962 18231 9025 18235
rect 5808 17919 5961 17929
rect 5808 17780 5961 17790
rect 7706 17919 7859 17929
rect 9203 17863 9213 18016
rect 9342 17863 9352 18016
rect 7706 17780 7859 17790
rect 9959 17774 10075 19425
rect 10470 19181 10585 19191
rect 10470 19074 10585 19084
rect 9958 17764 10075 17774
rect 10070 17658 10075 17764
rect 9958 17648 10075 17658
rect 9959 17647 10075 17648
rect -651 16339 -590 16344
rect -3062 16334 -586 16339
rect -3062 16282 -651 16334
rect -590 16282 -586 16334
rect -3062 16281 -586 16282
rect -3062 16248 -2991 16281
rect -651 16272 -590 16281
rect -3253 16236 -3187 16242
rect -3062 16184 -3057 16248
rect -2996 16184 -2991 16248
rect -3062 16172 -2991 16184
rect 10988 16186 11142 21065
rect 13066 20956 13219 20966
rect 13066 20817 13219 20827
rect 14208 20958 14361 20968
rect 14208 20819 14361 20829
rect 12312 20312 12465 20322
rect 12312 20173 12465 20183
rect 14210 20312 14363 20322
rect 14210 20173 14363 20183
rect 13644 19341 13722 19351
rect 13644 19245 13722 19255
rect 15284 18293 15352 22076
rect 19895 21542 19955 22203
rect 26602 22367 26755 22377
rect 26287 22272 26343 22282
rect 25455 22228 25608 22238
rect 26286 22206 26287 22268
rect 26343 22206 26468 22268
rect 26602 22228 26755 22238
rect 29084 22313 29237 22323
rect 26287 22196 26343 22206
rect 22571 22171 22724 22181
rect 20894 22154 20960 22157
rect 20894 22147 21886 22154
rect 20960 22081 21886 22147
rect 20894 22071 20960 22081
rect 19895 21541 20033 21542
rect 19895 21531 20295 21541
rect 17975 21520 18043 21530
rect 19073 21520 19138 21521
rect 18043 21511 19139 21520
rect 18043 21457 19073 21511
rect 19138 21457 19139 21511
rect 18043 21446 19139 21457
rect 17975 21435 18043 21445
rect 19895 21434 20195 21531
rect 20294 21434 20295 21531
rect 19895 21426 20295 21434
rect 19986 21422 20295 21426
rect 15770 21113 15780 21266
rect 15909 21113 15919 21266
rect 17283 21233 17738 21245
rect 17283 21077 17298 21233
rect 17548 21077 17738 21233
rect 17283 21060 17738 21077
rect 17553 20835 17738 21060
rect 17554 20704 17738 20835
rect 19600 20961 19753 20971
rect 19600 20822 19753 20832
rect 20742 20963 20895 20973
rect 20742 20824 20895 20834
rect 16796 20678 16912 20679
rect 17252 20678 17419 20679
rect 16796 20668 17419 20678
rect 16023 20655 16176 20665
rect 16796 20562 16801 20668
rect 16913 20651 17419 20668
rect 16913 20562 17295 20651
rect 16796 20545 17295 20562
rect 17407 20545 17419 20651
rect 16796 20536 17419 20545
rect 16023 20516 16176 20526
rect 15756 19463 15766 19616
rect 15895 19463 15905 19616
rect 16512 19556 16630 19559
rect 17255 19557 17420 19567
rect 17252 19556 17420 19557
rect 16512 19549 17420 19556
rect 16630 19539 17420 19549
rect 16630 19537 17296 19539
rect 16630 19431 17290 19537
rect 17408 19433 17420 19539
rect 17402 19431 17420 19433
rect 16512 19424 17420 19431
rect 16512 19422 17414 19424
rect 16512 19421 17377 19422
rect 16028 19051 16181 19061
rect 16028 18912 16181 18922
rect 15520 18293 15583 18299
rect 15284 18289 15588 18293
rect 15284 18237 15520 18289
rect 15583 18237 15588 18289
rect 15284 18231 15588 18237
rect 15520 18227 15583 18231
rect 12366 17915 12519 17925
rect 12366 17776 12519 17786
rect 14264 17915 14417 17925
rect 15761 17859 15771 18012
rect 15900 17859 15910 18012
rect 14264 17776 14417 17786
rect 16517 17770 16633 19421
rect 17028 19177 17143 19187
rect 17028 19070 17143 19080
rect 16516 17760 16633 17770
rect 16628 17654 16633 17760
rect 16516 17644 16633 17654
rect 16517 17643 16633 17644
rect 17553 16375 17738 20704
rect 18846 20317 18999 20327
rect 18846 20178 18999 20188
rect 20744 20317 20897 20327
rect 20744 20178 20897 20188
rect 20178 19346 20256 19356
rect 20178 19250 20256 19260
rect 21818 18298 21886 22081
rect 26408 21545 26468 22206
rect 29084 22174 29237 22184
rect 34475 22246 34575 22258
rect 34475 22163 34490 22246
rect 34558 22163 34575 22246
rect 27407 22157 27473 22160
rect 27407 22150 28399 22157
rect 27473 22084 28399 22150
rect 27407 22074 27473 22084
rect 26408 21544 26546 21545
rect 26408 21534 26808 21544
rect 24488 21523 24556 21533
rect 25586 21523 25651 21524
rect 24556 21514 25652 21523
rect 24556 21460 25586 21514
rect 25651 21460 25652 21514
rect 24556 21449 25652 21460
rect 24488 21438 24556 21448
rect 26408 21437 26708 21534
rect 26807 21437 26808 21534
rect 26408 21429 26808 21437
rect 26499 21425 26808 21429
rect 22304 21118 22314 21271
rect 22443 21118 22453 21271
rect 23826 21222 24263 21239
rect 23826 21085 23847 21222
rect 24075 21085 24263 21222
rect 23826 21065 24263 21085
rect 23330 20683 23446 20684
rect 23786 20683 23953 20684
rect 23330 20673 23953 20683
rect 22557 20660 22710 20670
rect 23330 20567 23335 20673
rect 23447 20656 23953 20673
rect 23447 20567 23829 20656
rect 23330 20550 23829 20567
rect 23941 20550 23953 20656
rect 23330 20541 23953 20550
rect 22557 20521 22710 20531
rect 22290 19468 22300 19621
rect 22429 19468 22439 19621
rect 23046 19561 23164 19564
rect 23789 19562 23954 19572
rect 23786 19561 23954 19562
rect 23046 19554 23954 19561
rect 23164 19544 23954 19554
rect 23164 19542 23830 19544
rect 23164 19436 23824 19542
rect 23942 19438 23954 19544
rect 23936 19436 23954 19438
rect 23046 19429 23954 19436
rect 23046 19427 23948 19429
rect 23046 19426 23911 19427
rect 22562 19056 22715 19066
rect 22562 18917 22715 18927
rect 22054 18298 22117 18304
rect 21818 18294 22122 18298
rect 21818 18242 22054 18294
rect 22117 18242 22122 18294
rect 21818 18236 22122 18242
rect 22054 18232 22117 18236
rect 18900 17920 19053 17930
rect 18900 17781 19053 17791
rect 20798 17920 20951 17930
rect 22295 17864 22305 18017
rect 22434 17864 22444 18017
rect 20798 17781 20951 17791
rect 23051 17775 23167 19426
rect 23562 19182 23677 19192
rect 23562 19075 23677 19085
rect 23050 17765 23167 17775
rect 23162 17659 23167 17765
rect 23050 17649 23167 17659
rect 23051 17648 23167 17649
rect 24082 16433 24261 21065
rect 26113 20964 26266 20974
rect 26113 20825 26266 20835
rect 27255 20966 27408 20976
rect 27255 20827 27408 20837
rect 25359 20320 25512 20330
rect 25359 20181 25512 20191
rect 27257 20320 27410 20330
rect 27257 20181 27410 20191
rect 26691 19349 26769 19359
rect 26691 19253 26769 19263
rect 28331 18301 28399 22084
rect 28817 21121 28827 21274
rect 28956 21121 28966 21274
rect 30707 21237 30780 21240
rect 30336 21216 30780 21237
rect 30336 21085 30360 21216
rect 30592 21085 30780 21216
rect 30336 21071 30780 21085
rect 30593 20982 30780 21071
rect 30239 20724 30501 20746
rect 29843 20686 29959 20687
rect 30239 20686 30262 20724
rect 29843 20676 30262 20686
rect 29070 20663 29223 20673
rect 29843 20570 29848 20676
rect 29960 20570 30262 20676
rect 29843 20568 30262 20570
rect 30480 20568 30501 20724
rect 29843 20544 30501 20568
rect 29070 20524 29223 20534
rect 28803 19471 28813 19624
rect 28942 19471 28952 19624
rect 29559 19564 29677 19567
rect 30302 19565 30467 19575
rect 30299 19564 30467 19565
rect 29559 19557 30467 19564
rect 29677 19547 30467 19557
rect 29677 19545 30343 19547
rect 29677 19439 30337 19545
rect 30455 19441 30467 19547
rect 30449 19439 30467 19441
rect 29559 19432 30467 19439
rect 29559 19430 30461 19432
rect 29559 19429 30424 19430
rect 29075 19059 29228 19069
rect 29075 18920 29228 18930
rect 28567 18301 28630 18307
rect 28331 18297 28635 18301
rect 28331 18245 28567 18297
rect 28630 18245 28635 18297
rect 28331 18239 28635 18245
rect 28567 18235 28630 18239
rect 25413 17923 25566 17933
rect 25413 17784 25566 17794
rect 27311 17923 27464 17933
rect 28808 17867 28818 18020
rect 28947 17867 28957 18020
rect 27311 17784 27464 17794
rect 29564 17778 29680 19429
rect 30075 19185 30190 19195
rect 30075 19078 30190 19088
rect 29563 17768 29680 17778
rect 29675 17662 29680 17768
rect 29563 17652 29680 17662
rect 29564 17651 29680 17652
rect 30594 16592 30780 20982
rect 30594 16591 30617 16592
rect 30594 16502 30607 16591
rect 30594 16501 30617 16502
rect 30768 16501 30780 16592
rect 30594 16488 30780 16501
rect 30707 16486 30780 16488
rect 17553 16286 17739 16375
rect 24082 16345 24097 16433
rect 24246 16345 24261 16433
rect 24082 16332 24261 16345
rect 17553 16198 17570 16286
rect 17726 16198 17739 16286
rect -4073 15362 -4063 15440
rect -3993 15362 -3983 15440
rect -3253 14848 -3187 16170
rect 10988 16126 11143 16186
rect 17553 16185 17739 16198
rect 23966 16267 24065 16277
rect 23966 16155 24065 16165
rect 10988 16029 11000 16126
rect 11129 16082 11143 16126
rect 17441 16137 17541 16147
rect 11129 16029 11142 16082
rect 17441 16042 17541 16052
rect 10988 16019 11142 16029
rect 10861 15801 10979 15811
rect 10861 15723 10979 15733
rect -1843 15420 -1833 15492
rect -1763 15420 -1753 15492
rect 21356 15482 21416 15492
rect 8153 15462 8213 15472
rect 8153 15390 8213 15400
rect 14702 15461 14762 15471
rect 21356 15410 21416 15420
rect 14702 15389 14762 15399
rect 30009 15315 30069 15325
rect 30009 15243 30069 15253
rect 32255 15255 32408 15265
rect 32255 15116 32408 15126
rect -3253 14794 -3247 14848
rect -3193 14794 -3187 14848
rect 33610 14907 33670 14917
rect 33610 14835 33670 14845
rect -2694 14613 -2598 14623
rect -2694 14506 -2598 14516
rect 31463 14335 31530 14340
rect 31456 14330 33172 14335
rect 21578 14286 21640 14288
rect 21578 14278 21642 14286
rect 21640 14276 21642 14278
rect 8375 14266 8437 14268
rect 8375 14258 8439 14266
rect 8437 14256 8439 14258
rect -651 14253 -594 14256
rect -3068 14246 -586 14253
rect -3068 14192 -651 14246
rect -594 14192 -586 14246
rect -3068 14182 -586 14192
rect 8375 14184 8439 14194
rect 14924 14265 14986 14267
rect 14924 14257 14988 14265
rect 14986 14255 14988 14257
rect 31456 14267 31463 14330
rect 31530 14325 33172 14330
rect 31530 14269 33119 14325
rect 31530 14267 33172 14269
rect 31456 14259 33172 14267
rect 31463 14257 31530 14259
rect 29354 14243 29433 14252
rect 21578 14204 21642 14214
rect 25405 14242 29433 14243
rect 14924 14183 14988 14193
rect -3068 14177 -2992 14182
rect -3255 14168 -3189 14174
rect -3068 14115 -3059 14177
rect -2999 14115 -2992 14177
rect -3068 14104 -2992 14115
rect 25405 14168 29354 14242
rect 33243 14222 33316 14232
rect 31463 14213 31530 14214
rect 31723 14213 33243 14222
rect 25405 14167 29433 14168
rect -4075 13294 -4065 13372
rect -3995 13294 -3985 13372
rect -3255 12780 -3189 14102
rect 349 14038 465 14048
rect 339 13982 349 14028
rect 465 14027 17242 14028
rect 25405 14027 25474 14167
rect 29354 14158 29433 14167
rect 31455 14212 33243 14213
rect 31455 14204 31723 14212
rect 31455 14141 31463 14204
rect 31530 14144 31723 14204
rect 31778 14144 33243 14212
rect 31530 14141 33243 14144
rect 29506 14128 29587 14138
rect 31455 14134 33243 14141
rect 31456 14133 31545 14134
rect 34219 14229 34357 14239
rect 34219 14137 34357 14147
rect 31463 14131 31530 14133
rect 465 13982 25474 14027
rect 339 13968 25474 13982
rect 25528 14120 25602 14121
rect 25528 14119 27862 14120
rect 25528 14038 29506 14119
rect 25528 13940 25602 14038
rect 27676 14037 29506 14038
rect 33243 14123 33316 14133
rect 30231 14119 30293 14121
rect 30231 14111 30295 14119
rect 30293 14109 30295 14111
rect 30231 14037 30295 14047
rect 29506 14022 29587 14032
rect 129 13924 25602 13940
rect 129 13866 135 13924
rect 219 13874 25602 13924
rect 32777 13974 34134 13984
rect 32839 13969 34134 13974
rect 32839 13888 34016 13969
rect 34124 13888 34134 13969
rect 32839 13883 34134 13888
rect 219 13866 230 13874
rect 129 13855 230 13866
rect 1489 13562 1549 13572
rect 373 13543 441 13549
rect 362 13539 453 13543
rect 362 13487 373 13539
rect 441 13487 453 13539
rect 1489 13490 1549 13500
rect -1845 13352 -1835 13424
rect -1765 13352 -1755 13424
rect -3255 12726 -3249 12780
rect -3195 12726 -3189 12780
rect -2692 12543 -2600 12553
rect -2692 12441 -2600 12451
rect -1216 12405 117 12417
rect -1216 12389 17 12405
rect -1216 12315 -1209 12389
rect -1143 12315 17 12389
rect -1216 12313 17 12315
rect 107 12313 117 12405
rect -1216 12305 117 12313
rect 17 12303 107 12305
rect -655 12198 -592 12200
rect -3069 12190 -584 12198
rect -3069 12129 -655 12190
rect -592 12129 -584 12190
rect -3069 12124 -584 12129
rect -3068 12108 -2991 12124
rect -655 12119 -592 12124
rect -3253 12099 -3187 12105
rect -3068 12048 -3056 12108
rect -2996 12048 -2991 12108
rect -3068 12036 -2991 12048
rect -4073 11225 -4063 11303
rect -3993 11225 -3983 11303
rect -3253 10711 -3187 12033
rect -1843 11283 -1833 11355
rect -1763 11283 -1753 11355
rect -3253 10657 -3247 10711
rect -3193 10657 -3187 10711
rect -2686 10471 -2601 10481
rect -2686 10375 -2601 10385
rect -1351 10294 -472 10304
rect -1351 10230 -1342 10294
rect -1280 10230 -472 10294
rect -1351 10218 -472 10230
rect -655 10133 -592 10136
rect -3070 10126 -585 10133
rect -3070 10065 -655 10126
rect -592 10065 -585 10126
rect -3070 10058 -585 10065
rect -3069 10040 -2990 10058
rect -655 10055 -592 10058
rect -3255 10031 -3189 10037
rect -3069 9979 -3057 10040
rect -3002 9979 -2990 10040
rect -3069 9969 -2990 9979
rect -4075 9157 -4065 9235
rect -3995 9157 -3985 9235
rect -3255 8643 -3189 9965
rect -1845 9215 -1835 9287
rect -1765 9215 -1755 9287
rect -3255 8589 -3249 8643
rect -3195 8589 -3189 8643
rect -2691 8401 -2602 8411
rect -2691 8306 -2602 8316
rect -656 8065 -589 8071
rect -3068 8061 -585 8065
rect -3068 7994 -656 8061
rect -589 7994 -585 8061
rect -3068 7990 -585 7994
rect -3068 7971 -2988 7990
rect -656 7984 -589 7990
rect -3255 7962 -3189 7968
rect -3068 7910 -3058 7971
rect -3002 7910 -2988 7971
rect -3068 7900 -2988 7910
rect -4075 7088 -4065 7166
rect -3995 7088 -3985 7166
rect -3255 6574 -3189 7896
rect -1845 7146 -1835 7218
rect -1765 7146 -1755 7218
rect -3255 6520 -3249 6574
rect -3195 6520 -3189 6574
rect -2688 6332 -2604 6342
rect -2688 6239 -2604 6249
rect -3069 5987 -585 5998
rect -3069 5933 -650 5987
rect -594 5933 -585 5987
rect -3069 5923 -585 5933
rect -3069 5904 -2989 5923
rect -3257 5894 -3191 5900
rect -3069 5842 -3059 5904
rect -3003 5842 -2989 5904
rect -3069 5832 -2989 5842
rect -4077 5020 -4067 5098
rect -3997 5020 -3987 5098
rect -3257 4506 -3191 5828
rect -1847 5078 -1837 5150
rect -1767 5078 -1757 5150
rect -3257 4452 -3251 4506
rect -3197 4452 -3191 4506
rect -2689 4265 -2606 4275
rect -2689 4171 -2606 4181
rect -540 4136 -472 10218
rect 174 9794 261 9798
rect 362 9794 453 13487
rect 1711 12366 1773 12368
rect 1711 12358 1775 12366
rect 1773 12356 1775 12358
rect 1711 12284 1775 12294
rect 1481 10977 1541 10987
rect 1481 10905 1541 10915
rect 165 9788 1049 9794
rect 165 9684 174 9788
rect 261 9783 1049 9788
rect 261 9687 971 9783
rect 1048 9687 1049 9783
rect 1703 9781 1765 9783
rect 1703 9773 1767 9781
rect 1765 9771 1767 9773
rect 1703 9699 1767 9709
rect 261 9684 1049 9687
rect 165 9677 1049 9684
rect 174 9674 261 9677
rect -540 4135 94 4136
rect -540 4125 103 4135
rect -540 4044 16 4125
rect -540 4034 103 4044
rect 356 4127 459 4137
rect 356 4038 459 4048
rect -540 4033 94 4034
rect -3069 3919 -585 3929
rect -3069 3865 -650 3919
rect -594 3865 -585 3919
rect -3069 3854 -585 3865
rect -3069 3834 -2989 3854
rect -3255 3825 -3189 3831
rect -3069 3774 -3055 3834
rect -3003 3774 -2989 3834
rect -3069 3763 -2989 3774
rect -4075 2951 -4065 3029
rect -3995 2951 -3985 3029
rect -3255 2437 -3189 3759
rect -1845 3009 -1835 3081
rect -1765 3009 -1755 3081
rect -3255 2383 -3249 2437
rect -3195 2383 -3189 2437
rect -2691 2196 -2601 2206
rect -2691 2099 -2601 2109
rect -650 1866 -594 1867
rect -3070 1857 -585 1866
rect -3070 1803 -650 1857
rect -594 1803 -585 1857
rect -3070 1791 -585 1803
rect -3070 1769 -2989 1791
rect -3257 1757 -3191 1763
rect -3070 1704 -3060 1769
rect -3001 1704 -2989 1769
rect -3070 1699 -2989 1704
rect -3060 1694 -3001 1699
rect -4077 883 -4067 961
rect -3997 883 -3987 961
rect -3257 369 -3191 1691
rect -1847 941 -1837 1013
rect -1767 941 -1757 1013
rect 492 776 610 9677
rect 1462 7699 1522 7709
rect 1462 7627 1522 7637
rect 1684 6503 1746 6505
rect 1684 6495 1748 6503
rect 1746 6493 1748 6495
rect 1684 6421 1748 6431
rect 1478 4939 1538 4949
rect 1478 4867 1538 4877
rect 1700 3743 1762 3745
rect 1700 3735 1764 3743
rect 1762 3733 1764 3735
rect 1700 3661 1764 3671
rect 492 690 502 776
rect 601 690 610 776
rect 492 682 610 690
rect 502 680 601 682
rect -3257 315 -3251 369
rect -3197 315 -3191 369
rect 2455 210 2562 13874
rect 32777 13873 34134 13883
rect 2603 13842 18762 13844
rect 29236 13842 29297 13843
rect 2603 13822 29328 13842
rect 2603 13768 14358 13822
rect 14415 13768 29328 13822
rect 2603 13749 29328 13768
rect 2603 13748 25587 13749
rect 2604 888 2722 13748
rect 29236 13622 29328 13749
rect 33832 13711 33894 13713
rect 33832 13703 33896 13711
rect 33894 13701 33896 13703
rect 33832 13629 33896 13639
rect 13499 13508 13652 13518
rect 11017 13454 11170 13464
rect 6950 13420 7103 13430
rect 4468 13366 4621 13376
rect 8097 13420 8250 13430
rect 7362 13325 7418 13335
rect 6950 13281 7103 13291
rect 4468 13227 4621 13237
rect 7237 13259 7362 13321
rect 7418 13259 7419 13321
rect 14646 13508 14799 13518
rect 13911 13413 13967 13423
rect 13499 13369 13652 13379
rect 11017 13315 11170 13325
rect 13786 13347 13911 13409
rect 13967 13347 13968 13409
rect 26778 13508 26931 13518
rect 24296 13454 24449 13464
rect 20153 13440 20306 13450
rect 14646 13369 14799 13379
rect 17671 13386 17824 13396
rect 12781 13298 12847 13301
rect 8097 13281 8250 13291
rect 11855 13291 12847 13298
rect 6232 13210 6298 13213
rect 5306 13203 6298 13210
rect 5306 13137 6232 13203
rect 4739 12174 4749 12327
rect 4878 12174 4888 12327
rect 3239 11739 3406 11740
rect 3746 11739 3862 11740
rect 3239 11729 3862 11739
rect 3239 11712 3745 11729
rect 3239 11606 3251 11712
rect 3363 11623 3745 11712
rect 3857 11623 3862 11729
rect 3363 11606 3862 11623
rect 3239 11597 3862 11606
rect 4482 11716 4635 11726
rect 4482 11577 4635 11587
rect 3238 10618 3403 10628
rect 3238 10617 3406 10618
rect 4028 10617 4146 10620
rect 3238 10610 4146 10617
rect 3238 10600 4028 10610
rect 3238 10494 3250 10600
rect 3362 10598 4028 10600
rect 3238 10492 3256 10494
rect 3368 10492 4028 10598
rect 4753 10524 4763 10677
rect 4892 10524 4902 10677
rect 3238 10485 4146 10492
rect 3244 10483 4146 10485
rect 3281 10482 4146 10483
rect 3515 10238 3630 10248
rect 3515 10131 3630 10141
rect 4025 8831 4141 10482
rect 4477 10112 4630 10122
rect 4477 9973 4630 9983
rect 5075 9354 5138 9360
rect 5306 9354 5374 13137
rect 6232 13127 6298 13137
rect 7237 12598 7297 13259
rect 7362 13249 7418 13259
rect 7159 12597 7297 12598
rect 6897 12587 7297 12597
rect 6897 12490 6898 12587
rect 6997 12490 7297 12587
rect 11855 13225 12781 13291
rect 8054 12576 8119 12577
rect 9149 12576 9363 12586
rect 8053 12567 9187 12576
rect 8053 12513 8054 12567
rect 8119 12513 9187 12567
rect 8053 12502 9187 12513
rect 6897 12482 7297 12490
rect 9149 12501 9187 12502
rect 9332 12501 9363 12576
rect 9149 12488 9363 12501
rect 6897 12478 7206 12482
rect 11288 12262 11298 12415
rect 11427 12262 11437 12415
rect 6297 12019 6450 12029
rect 6297 11880 6450 11890
rect 7439 12017 7592 12027
rect 7439 11878 7592 11888
rect 9788 11827 9955 11828
rect 10295 11827 10411 11828
rect 9788 11817 10411 11827
rect 9788 11800 10294 11817
rect 9788 11694 9800 11800
rect 9912 11711 10294 11800
rect 10406 11711 10411 11817
rect 9912 11694 10411 11711
rect 9788 11685 10411 11694
rect 11031 11804 11184 11814
rect 11031 11665 11184 11675
rect 6295 11373 6448 11383
rect 6295 11234 6448 11244
rect 8193 11373 8346 11383
rect 8193 11234 8346 11244
rect 10577 10705 10695 10708
rect 9785 10698 10695 10705
rect 9785 10580 10577 10698
rect 11302 10612 11312 10765
rect 11441 10612 11451 10765
rect 9785 10570 10695 10580
rect 6936 10402 7014 10412
rect 6936 10306 7014 10316
rect 5070 9350 5374 9354
rect 5070 9298 5075 9350
rect 5138 9298 5374 9350
rect 5070 9292 5374 9298
rect 5075 9288 5138 9292
rect 4748 8920 4758 9073
rect 4887 8920 4897 9073
rect 6241 8976 6394 8986
rect 6241 8837 6394 8847
rect 8139 8976 8292 8986
rect 8139 8837 8292 8847
rect 4025 8821 4142 8831
rect 4025 8715 4030 8821
rect 4025 8705 4142 8715
rect 4025 8704 4141 8705
rect 9785 8386 9951 10570
rect 10064 10326 10179 10336
rect 10064 10219 10179 10229
rect 10574 8919 10690 10570
rect 11026 10200 11179 10210
rect 11026 10061 11179 10071
rect 11624 9442 11687 9448
rect 11855 9442 11923 13225
rect 12781 13215 12847 13225
rect 13786 12686 13846 13347
rect 13911 13337 13967 13347
rect 21300 13440 21453 13450
rect 20565 13345 20621 13355
rect 20153 13301 20306 13311
rect 17671 13247 17824 13257
rect 20440 13279 20565 13341
rect 20621 13279 20622 13341
rect 27925 13508 28078 13518
rect 27190 13413 27246 13423
rect 26778 13369 26931 13379
rect 24296 13315 24449 13325
rect 27065 13347 27190 13409
rect 27246 13347 27247 13409
rect 27925 13369 28078 13379
rect 21300 13301 21453 13311
rect 26060 13298 26126 13301
rect 25134 13291 26126 13298
rect 19435 13230 19501 13233
rect 13708 12685 13846 12686
rect 13446 12675 13846 12685
rect 13446 12578 13447 12675
rect 13546 12578 13846 12675
rect 18509 13223 19501 13230
rect 18509 13157 19435 13223
rect 14603 12664 14668 12665
rect 15698 12664 15766 12674
rect 14602 12655 15698 12664
rect 14602 12601 14603 12655
rect 14668 12601 15698 12655
rect 14602 12590 15698 12601
rect 15698 12579 15766 12589
rect 13446 12570 13846 12578
rect 13446 12566 13755 12570
rect 17942 12194 17952 12347
rect 18081 12194 18091 12347
rect 12846 12107 12999 12117
rect 12846 11968 12999 11978
rect 13988 12105 14141 12115
rect 13988 11966 14141 11976
rect 15767 11759 16711 11762
rect 16949 11759 17065 11760
rect 15767 11749 17065 11759
rect 15767 11643 16948 11749
rect 17060 11643 17065 11749
rect 15767 11617 17065 11643
rect 17685 11736 17838 11746
rect 12844 11461 12997 11471
rect 12844 11322 12997 11332
rect 14742 11461 14895 11471
rect 14742 11322 14895 11332
rect 13485 10490 13563 10500
rect 13485 10394 13563 10404
rect 15767 9977 15887 11617
rect 17685 11597 17838 11607
rect 16441 10638 16606 10648
rect 16441 10637 16609 10638
rect 17231 10637 17349 10640
rect 16441 10630 17349 10637
rect 16441 10620 17231 10630
rect 16441 10514 16453 10620
rect 16565 10618 17231 10620
rect 16441 10512 16459 10514
rect 16571 10512 17231 10618
rect 17956 10544 17966 10697
rect 18095 10544 18105 10697
rect 16441 10505 17349 10512
rect 16447 10503 17349 10505
rect 16484 10502 17349 10503
rect 16718 10258 16833 10268
rect 16718 10151 16833 10161
rect 15767 9878 15887 9888
rect 11619 9438 11923 9442
rect 11619 9386 11624 9438
rect 11687 9386 11923 9438
rect 11619 9380 11923 9386
rect 11624 9376 11687 9380
rect 11297 9008 11307 9161
rect 11436 9008 11446 9161
rect 12790 9064 12943 9074
rect 12790 8925 12943 8935
rect 14688 9064 14841 9074
rect 14688 8925 14841 8935
rect 10574 8909 10691 8919
rect 10574 8803 10579 8909
rect 10574 8793 10691 8803
rect 17228 8851 17344 10502
rect 17680 10132 17833 10142
rect 17680 9993 17833 10003
rect 18278 9374 18341 9380
rect 18509 9374 18577 13157
rect 19435 13147 19501 13157
rect 20440 12618 20500 13279
rect 20565 13269 20621 13279
rect 20362 12617 20500 12618
rect 20100 12607 20500 12617
rect 20100 12510 20101 12607
rect 20200 12510 20500 12607
rect 25134 13225 26060 13291
rect 21257 12596 21322 12597
rect 22321 12596 22418 12606
rect 21256 12587 22321 12596
rect 21256 12533 21257 12587
rect 21322 12533 22321 12587
rect 21256 12522 22321 12533
rect 22418 12522 22419 12596
rect 22321 12512 22418 12522
rect 20100 12502 20500 12510
rect 20100 12498 20409 12502
rect 24567 12262 24577 12415
rect 24706 12262 24716 12415
rect 19500 12039 19653 12049
rect 19500 11900 19653 11910
rect 20642 12037 20795 12047
rect 20642 11898 20795 11908
rect 23067 11827 23234 11828
rect 23574 11827 23690 11828
rect 23067 11817 23690 11827
rect 23067 11800 23573 11817
rect 23067 11694 23079 11800
rect 23191 11711 23573 11800
rect 23685 11711 23690 11817
rect 23191 11694 23690 11711
rect 23067 11685 23690 11694
rect 24310 11804 24463 11814
rect 24310 11665 24463 11675
rect 19498 11393 19651 11403
rect 19498 11254 19651 11264
rect 21396 11393 21549 11403
rect 21396 11254 21549 11264
rect 23856 10705 23974 10708
rect 23093 10698 23974 10705
rect 23093 10580 23856 10698
rect 24581 10612 24591 10765
rect 24720 10612 24730 10765
rect 23093 10571 23974 10580
rect 20139 10422 20217 10432
rect 20139 10326 20217 10336
rect 22874 9911 22970 9921
rect 22874 9801 22970 9811
rect 18273 9370 18577 9374
rect 18273 9318 18278 9370
rect 18341 9318 18577 9370
rect 18273 9312 18577 9318
rect 18278 9308 18341 9312
rect 17951 8940 17961 9093
rect 18090 8940 18100 9093
rect 19444 8996 19597 9006
rect 19444 8857 19597 8867
rect 21342 8996 21495 9006
rect 21342 8857 21495 8867
rect 17228 8841 17345 8851
rect 10574 8792 10690 8793
rect 17228 8735 17233 8841
rect 17228 8725 17345 8735
rect 17228 8724 17344 8725
rect 22394 8607 22536 8617
rect 22394 8464 22536 8473
rect 9785 8240 15699 8386
rect 9874 8235 15699 8240
rect 23094 8364 23204 10571
rect 23235 10570 23974 10571
rect 23343 10326 23458 10336
rect 23343 10219 23458 10229
rect 23853 8919 23969 10570
rect 24305 10200 24458 10210
rect 24305 10061 24458 10071
rect 24903 9442 24966 9448
rect 25134 9442 25202 13225
rect 26060 13215 26126 13225
rect 27065 12686 27125 13347
rect 27190 13337 27246 13347
rect 26987 12685 27125 12686
rect 26725 12675 27125 12685
rect 26725 12578 26726 12675
rect 26825 12578 27125 12675
rect 27882 12664 27947 12665
rect 28860 12664 28928 12674
rect 27881 12655 28860 12664
rect 27881 12601 27882 12655
rect 27947 12601 28860 12655
rect 27881 12590 28860 12601
rect 28860 12579 28928 12589
rect 26725 12570 27125 12578
rect 26725 12566 27034 12570
rect 26125 12107 26278 12117
rect 26125 11968 26278 11978
rect 27267 12105 27420 12115
rect 27267 11966 27420 11976
rect 29236 11812 29327 13622
rect 32177 12925 32388 12935
rect 32177 12758 32388 12768
rect 30004 12744 30064 12754
rect 30004 12672 30064 12682
rect 29236 11801 29735 11812
rect 29236 11720 29653 11801
rect 29236 11711 29735 11720
rect 29653 11710 29735 11711
rect 30226 11548 30288 11550
rect 30226 11540 30290 11548
rect 30288 11538 30290 11540
rect 26123 11461 26276 11471
rect 26123 11322 26276 11332
rect 28021 11461 28174 11471
rect 30226 11466 30290 11476
rect 28021 11322 28174 11332
rect 32257 11164 32410 11174
rect 32257 11025 32410 11035
rect 33612 10816 33672 10826
rect 33612 10744 33672 10754
rect 26764 10490 26842 10500
rect 26764 10394 26842 10404
rect 31465 10244 31532 10249
rect 31458 10239 33174 10244
rect 31458 10176 31465 10239
rect 31532 10234 33174 10239
rect 31532 10178 33121 10234
rect 31532 10176 33174 10178
rect 31458 10168 33174 10176
rect 31465 10166 31532 10168
rect 33245 10131 33318 10141
rect 31465 10122 31532 10123
rect 31725 10122 33245 10131
rect 31457 10121 33245 10122
rect 31457 10113 31725 10121
rect 31457 10050 31465 10113
rect 31532 10053 31725 10113
rect 31780 10053 33245 10121
rect 31532 10050 33245 10053
rect 31457 10043 33245 10050
rect 31458 10042 31547 10043
rect 31465 10040 31532 10042
rect 33245 10032 33318 10042
rect 34475 9894 34575 22163
rect 35009 22158 35115 25207
rect 37444 25058 37528 25207
rect 37561 25206 37646 25234
rect 37728 25206 37813 25234
rect 37442 25047 37528 25058
rect 37442 24976 37454 25047
rect 37517 24976 37528 25047
rect 37442 24965 37528 24976
rect 37444 23962 37528 24965
rect 36473 23812 36483 23912
rect 36575 23812 36585 23912
rect 37444 23892 37454 23962
rect 37516 23892 37528 23962
rect 37444 23883 37528 23892
rect 37564 23721 37643 25206
rect 37729 24080 37813 25206
rect 37729 24012 37737 24080
rect 37802 24012 37813 24080
rect 37729 24001 37813 24012
rect 38717 23816 38727 23892
rect 38785 23816 38795 23892
rect 37564 23662 37574 23721
rect 37634 23662 37644 23721
rect 35009 22079 37529 22158
rect 37561 22147 37646 22158
rect 37728 22147 37813 22158
rect 37559 22090 37569 22147
rect 37637 22090 37647 22147
rect 37727 22090 37737 22147
rect 37805 22090 37815 22147
rect 35009 19026 35115 22079
rect 37444 22035 37529 22079
rect 37561 22062 37646 22090
rect 37728 22062 37813 22090
rect 37444 21914 37528 22035
rect 37442 21903 37528 21914
rect 37442 21832 37454 21903
rect 37517 21832 37528 21903
rect 37442 21821 37528 21832
rect 37444 20818 37528 21821
rect 36473 20668 36483 20768
rect 36575 20668 36585 20768
rect 37444 20748 37454 20818
rect 37516 20748 37528 20818
rect 37444 20739 37528 20748
rect 37564 20577 37643 22062
rect 37729 20936 37813 22062
rect 37729 20868 37737 20936
rect 37802 20868 37813 20936
rect 37729 20857 37813 20868
rect 38717 20672 38727 20748
rect 38785 20672 38795 20748
rect 37564 20518 37574 20577
rect 37634 20518 37644 20577
rect 35009 18947 37524 19026
rect 37557 19015 37642 19026
rect 37724 19015 37809 19026
rect 37555 18958 37565 19015
rect 37633 18958 37643 19015
rect 37723 18958 37733 19015
rect 37801 18958 37811 19015
rect 35009 15964 35115 18947
rect 37440 18782 37524 18947
rect 37557 18930 37642 18958
rect 37724 18930 37809 18958
rect 37438 18771 37524 18782
rect 37438 18700 37450 18771
rect 37513 18700 37524 18771
rect 37438 18689 37524 18700
rect 37440 17686 37524 18689
rect 36469 17536 36479 17636
rect 36571 17536 36581 17636
rect 37440 17616 37450 17686
rect 37512 17616 37524 17686
rect 37440 17607 37524 17616
rect 37560 17445 37639 18930
rect 37725 17804 37809 18930
rect 37725 17736 37733 17804
rect 37798 17736 37809 17804
rect 37725 17725 37809 17736
rect 38713 17540 38723 17616
rect 38781 17540 38791 17616
rect 37560 17386 37570 17445
rect 37630 17386 37640 17445
rect 34720 15952 35115 15964
rect 34720 15871 34744 15952
rect 34888 15884 35115 15952
rect 34888 15871 37525 15884
rect 37557 15871 37642 15882
rect 37725 15875 37809 15885
rect 34720 15861 37525 15871
rect 34720 15860 34970 15861
rect 33958 9893 34575 9894
rect 32779 9883 34575 9893
rect 32841 9792 34575 9883
rect 32779 9782 34575 9792
rect 34357 9781 34575 9782
rect 35009 15804 37525 15861
rect 37555 15814 37565 15871
rect 37633 15814 37643 15871
rect 35009 12680 35115 15804
rect 37439 15769 37525 15804
rect 37557 15786 37642 15814
rect 37440 15638 37524 15769
rect 37438 15627 37524 15638
rect 37438 15556 37450 15627
rect 37513 15556 37524 15627
rect 37438 15545 37524 15556
rect 37440 14542 37524 15545
rect 36469 14392 36479 14492
rect 36571 14392 36581 14492
rect 37440 14472 37450 14542
rect 37512 14472 37524 14542
rect 37440 14463 37524 14472
rect 37560 14301 37639 15786
rect 37725 15778 37736 15875
rect 37799 15778 37809 15875
rect 37725 14660 37809 15778
rect 37725 14592 37733 14660
rect 37798 14592 37809 14660
rect 37725 14581 37809 14592
rect 38713 14396 38723 14472
rect 38781 14396 38791 14472
rect 37560 14242 37570 14301
rect 37630 14242 37640 14301
rect 35009 12602 37528 12680
rect 37561 12669 37646 12680
rect 37728 12669 37813 12680
rect 37559 12612 37569 12669
rect 37637 12612 37647 12669
rect 37727 12612 37737 12669
rect 37805 12612 37815 12669
rect 30004 9711 30064 9721
rect 30004 9639 30064 9649
rect 33834 9620 33896 9622
rect 33834 9612 33898 9620
rect 33896 9610 33898 9612
rect 33834 9538 33898 9548
rect 24898 9438 25202 9442
rect 24898 9386 24903 9438
rect 24966 9386 25202 9438
rect 24898 9380 25202 9386
rect 35009 9536 35115 12602
rect 37444 12436 37528 12602
rect 37561 12584 37646 12612
rect 37728 12584 37813 12612
rect 37442 12425 37528 12436
rect 37442 12354 37454 12425
rect 37517 12354 37528 12425
rect 37442 12343 37528 12354
rect 37444 11340 37528 12343
rect 36473 11190 36483 11290
rect 36575 11190 36585 11290
rect 37444 11270 37454 11340
rect 37516 11270 37528 11340
rect 37444 11261 37528 11270
rect 37564 11099 37643 12584
rect 37729 11458 37813 12584
rect 37729 11390 37737 11458
rect 37802 11390 37813 11458
rect 37729 11379 37813 11390
rect 38717 11194 38727 11270
rect 38785 11194 38795 11270
rect 37564 11040 37574 11099
rect 37634 11040 37644 11099
rect 35009 9458 37529 9536
rect 37561 9525 37646 9536
rect 37728 9528 37814 9539
rect 37559 9468 37569 9525
rect 37637 9468 37647 9525
rect 24903 9376 24966 9380
rect 24576 9008 24586 9161
rect 24715 9008 24725 9161
rect 26069 9064 26222 9074
rect 26069 8925 26222 8935
rect 27967 9064 28120 9074
rect 27967 8925 28120 8935
rect 23853 8909 23970 8919
rect 23853 8803 23858 8909
rect 29758 8901 29847 8910
rect 23853 8793 23970 8803
rect 29242 8900 29847 8901
rect 29242 8813 29758 8900
rect 29242 8809 29847 8813
rect 23853 8792 23969 8793
rect 23503 8607 23645 8617
rect 23503 8463 23645 8473
rect 6942 7640 7095 7650
rect 4460 7586 4613 7596
rect 8089 7640 8242 7650
rect 7354 7545 7410 7555
rect 6942 7501 7095 7511
rect 4460 7447 4613 7457
rect 7229 7479 7354 7541
rect 7410 7479 7411 7541
rect 13493 7638 13646 7648
rect 8089 7501 8242 7511
rect 11011 7584 11164 7594
rect 6224 7430 6290 7433
rect 5298 7423 6290 7430
rect 5298 7357 6224 7423
rect 4731 6394 4741 6547
rect 4870 6394 4880 6547
rect 3231 5959 3398 5960
rect 3738 5959 3854 5960
rect 3231 5949 3854 5959
rect 3231 5932 3737 5949
rect 3231 5826 3243 5932
rect 3355 5843 3737 5932
rect 3849 5843 3854 5949
rect 3355 5826 3854 5843
rect 3231 5817 3854 5826
rect 4474 5936 4627 5946
rect 4474 5797 4627 5807
rect 3127 4848 3361 4853
rect 3127 4843 3395 4848
rect 3361 4838 3395 4843
rect 3361 4837 3398 4838
rect 4020 4837 4138 4840
rect 3361 4830 4138 4837
rect 3361 4712 4020 4830
rect 4745 4744 4755 4897
rect 4884 4744 4894 4897
rect 3361 4706 4138 4712
rect 3127 4702 4138 4706
rect 3127 4696 3361 4702
rect 3507 4458 3622 4468
rect 3507 4351 3622 4361
rect 4017 3051 4133 4702
rect 4469 4332 4622 4342
rect 4469 4193 4622 4203
rect 5067 3574 5130 3580
rect 5298 3574 5366 7357
rect 6224 7347 6290 7357
rect 7229 6818 7289 7479
rect 7354 7469 7410 7479
rect 14640 7638 14793 7648
rect 13905 7543 13961 7553
rect 13493 7499 13646 7509
rect 11011 7445 11164 7455
rect 13780 7477 13905 7539
rect 13961 7477 13962 7539
rect 14640 7499 14793 7509
rect 12775 7428 12841 7431
rect 7151 6817 7289 6818
rect 6889 6807 7289 6817
rect 6889 6710 6890 6807
rect 6989 6710 7289 6807
rect 11849 7421 12841 7428
rect 11849 7355 12775 7421
rect 8046 6796 8111 6797
rect 9141 6796 9209 6806
rect 8045 6787 9141 6796
rect 8045 6733 8046 6787
rect 8111 6733 9141 6787
rect 8045 6722 9141 6733
rect 9141 6711 9209 6721
rect 6889 6702 7289 6710
rect 6889 6698 7198 6702
rect 11282 6392 11292 6545
rect 11421 6392 11431 6545
rect 6289 6239 6442 6249
rect 6289 6100 6442 6110
rect 7431 6237 7584 6247
rect 7431 6098 7584 6108
rect 10289 5957 10405 5958
rect 10028 5954 10405 5957
rect 9782 5947 10405 5954
rect 9782 5930 10288 5947
rect 9782 5824 9794 5930
rect 9906 5841 10288 5930
rect 10400 5841 10405 5947
rect 9906 5824 10405 5841
rect 9782 5815 10405 5824
rect 11025 5934 11178 5944
rect 11025 5795 11178 5805
rect 6287 5593 6440 5603
rect 6287 5454 6440 5464
rect 8185 5593 8338 5603
rect 8185 5454 8338 5464
rect 9762 4836 9985 4846
rect 10571 4835 10689 4838
rect 9985 4828 10689 4835
rect 9985 4710 10571 4828
rect 11296 4742 11306 4895
rect 11435 4742 11445 4895
rect 9985 4700 10689 4710
rect 9762 4690 9985 4700
rect 6928 4622 7006 4632
rect 6928 4526 7006 4536
rect 10058 4456 10173 4466
rect 10058 4349 10173 4359
rect 5062 3570 5366 3574
rect 5062 3518 5067 3570
rect 5130 3518 5366 3570
rect 5062 3512 5366 3518
rect 5067 3508 5130 3512
rect 4740 3140 4750 3293
rect 4879 3140 4889 3293
rect 6233 3196 6386 3206
rect 6233 3057 6386 3067
rect 8131 3196 8284 3206
rect 8131 3057 8284 3067
rect 4017 3041 4134 3051
rect 4017 2935 4022 3041
rect 4017 2925 4134 2935
rect 10568 3049 10684 4700
rect 11020 4330 11173 4340
rect 11020 4191 11173 4201
rect 11618 3572 11681 3578
rect 11849 3572 11917 7355
rect 12775 7345 12841 7355
rect 13780 6816 13840 7477
rect 13905 7467 13961 7477
rect 13702 6815 13840 6816
rect 13440 6805 13840 6815
rect 13440 6708 13441 6805
rect 13540 6708 13840 6805
rect 14597 6794 14662 6795
rect 15565 6794 15695 8235
rect 23094 8232 29003 8364
rect 23094 8231 23198 8232
rect 28874 8208 29003 8232
rect 28874 8119 29004 8208
rect 20148 7639 20301 7649
rect 17666 7585 17819 7595
rect 21295 7639 21448 7649
rect 20560 7544 20616 7554
rect 20148 7500 20301 7510
rect 17666 7446 17819 7456
rect 20435 7478 20560 7540
rect 20616 7478 20617 7540
rect 26770 7640 26923 7650
rect 21295 7500 21448 7510
rect 24288 7586 24441 7596
rect 19430 7429 19496 7432
rect 14596 6785 15695 6794
rect 14596 6731 14597 6785
rect 14662 6731 15695 6785
rect 14596 6720 15695 6731
rect 15565 6717 15695 6720
rect 18504 7422 19496 7429
rect 18504 7356 19430 7422
rect 13440 6700 13840 6708
rect 13440 6696 13749 6700
rect 17937 6393 17947 6546
rect 18076 6393 18086 6546
rect 12840 6237 12993 6247
rect 12840 6098 12993 6108
rect 13982 6235 14135 6245
rect 13982 6096 14135 6106
rect 16370 5959 16536 5961
rect 16370 5958 16604 5959
rect 16944 5958 17060 5959
rect 16370 5948 17060 5958
rect 16370 5936 16943 5948
rect 16370 5823 16382 5936
rect 16586 5842 16943 5936
rect 17055 5842 17060 5948
rect 16370 5822 16534 5823
rect 16586 5822 17060 5842
rect 16370 5816 17060 5822
rect 17680 5935 17833 5945
rect 16370 5815 16594 5816
rect 17680 5796 17833 5806
rect 12838 5591 12991 5601
rect 12838 5452 12991 5462
rect 14736 5591 14889 5601
rect 14736 5452 14889 5462
rect 16436 4837 16601 4847
rect 16436 4836 16604 4837
rect 17226 4836 17344 4839
rect 16436 4829 17344 4836
rect 16436 4821 17226 4829
rect 16436 4709 16443 4821
rect 16587 4711 17226 4821
rect 17951 4743 17961 4896
rect 18090 4743 18100 4896
rect 16587 4709 17344 4711
rect 16436 4704 17344 4709
rect 16442 4702 17344 4704
rect 16443 4701 17344 4702
rect 16443 4699 16587 4701
rect 13479 4620 13557 4630
rect 13479 4524 13557 4534
rect 16713 4457 16828 4467
rect 16713 4350 16828 4360
rect 11613 3568 11917 3572
rect 11613 3516 11618 3568
rect 11681 3516 11917 3568
rect 11613 3510 11917 3516
rect 11618 3506 11681 3510
rect 11291 3138 11301 3291
rect 11430 3138 11440 3291
rect 12784 3194 12937 3204
rect 12784 3055 12937 3065
rect 14682 3194 14835 3204
rect 14682 3055 14835 3065
rect 17223 3050 17339 4701
rect 17675 4331 17828 4341
rect 17675 4192 17828 4202
rect 18273 3573 18336 3579
rect 18504 3573 18572 7356
rect 19430 7346 19496 7356
rect 20435 6817 20495 7478
rect 20560 7468 20616 7478
rect 27917 7640 28070 7650
rect 27182 7545 27238 7555
rect 26770 7501 26923 7511
rect 24288 7447 24441 7457
rect 27057 7479 27182 7541
rect 27238 7479 27239 7541
rect 27917 7501 28070 7511
rect 26052 7430 26118 7433
rect 20357 6816 20495 6817
rect 20095 6806 20495 6816
rect 20095 6709 20096 6806
rect 20195 6709 20495 6806
rect 25126 7423 26118 7430
rect 25126 7357 26052 7423
rect 21252 6795 21317 6796
rect 22347 6795 22415 6805
rect 21251 6786 22347 6795
rect 21251 6732 21252 6786
rect 21317 6732 22347 6786
rect 21251 6721 22347 6732
rect 22347 6710 22415 6720
rect 20095 6701 20495 6709
rect 20095 6697 20404 6701
rect 24559 6394 24569 6547
rect 24698 6394 24708 6547
rect 19495 6238 19648 6248
rect 19495 6099 19648 6109
rect 20637 6236 20790 6246
rect 20637 6097 20790 6107
rect 23566 5959 23682 5960
rect 23059 5949 23682 5959
rect 23059 5932 23565 5949
rect 23059 5826 23071 5932
rect 23183 5843 23565 5932
rect 23677 5843 23682 5949
rect 23183 5826 23682 5843
rect 23059 5817 23682 5826
rect 24302 5936 24455 5946
rect 24302 5797 24455 5807
rect 19493 5592 19646 5602
rect 19493 5453 19646 5463
rect 21391 5592 21544 5602
rect 21391 5453 21544 5463
rect 23058 4838 23223 4848
rect 23058 4837 23226 4838
rect 23848 4837 23966 4840
rect 23058 4830 23966 4837
rect 23058 4820 23848 4830
rect 23058 4714 23070 4820
rect 23182 4818 23848 4820
rect 23058 4712 23076 4714
rect 23188 4712 23848 4818
rect 24573 4744 24583 4897
rect 24712 4744 24722 4897
rect 23058 4705 23966 4712
rect 23064 4703 23966 4705
rect 23101 4702 23966 4703
rect 20134 4621 20212 4631
rect 20134 4525 20212 4535
rect 23335 4458 23450 4468
rect 23335 4351 23450 4361
rect 18268 3569 18572 3573
rect 18268 3517 18273 3569
rect 18336 3517 18572 3569
rect 18268 3511 18572 3517
rect 18273 3507 18336 3511
rect 17946 3139 17956 3292
rect 18085 3139 18095 3292
rect 19439 3195 19592 3205
rect 19439 3056 19592 3066
rect 21337 3195 21490 3205
rect 21337 3056 21490 3066
rect 23845 3051 23961 4702
rect 24297 4332 24450 4342
rect 24297 4193 24450 4203
rect 24895 3574 24958 3580
rect 25126 3574 25194 7357
rect 26052 7347 26118 7357
rect 27057 6818 27117 7479
rect 27182 7469 27238 7479
rect 26979 6817 27117 6818
rect 26717 6807 27117 6817
rect 26717 6710 26718 6807
rect 26817 6710 27117 6807
rect 27874 6796 27939 6797
rect 28874 6796 29005 8119
rect 27873 6787 29005 6796
rect 27873 6733 27874 6787
rect 27939 6733 29005 6787
rect 27873 6722 29005 6733
rect 28874 6720 29005 6722
rect 28969 6719 29005 6720
rect 26717 6702 27117 6710
rect 26717 6698 27026 6702
rect 26117 6239 26270 6249
rect 26117 6100 26270 6110
rect 27259 6237 27412 6247
rect 27259 6098 27412 6108
rect 26115 5593 26268 5603
rect 26115 5454 26268 5464
rect 28013 5593 28166 5603
rect 28013 5454 28166 5464
rect 26756 4622 26834 4632
rect 26756 4526 26834 4536
rect 29029 4110 29161 4120
rect 29029 4004 29161 4014
rect 24890 3570 25194 3574
rect 24890 3518 24895 3570
rect 24958 3518 25194 3570
rect 29242 3651 29339 8809
rect 29758 8803 29847 8809
rect 32179 8834 32390 8844
rect 32179 8667 32390 8677
rect 30226 8515 30288 8517
rect 30226 8507 30290 8515
rect 30288 8505 30290 8507
rect 30226 8433 30290 8443
rect 30075 7791 30135 7801
rect 30075 7719 30135 7729
rect 32257 7669 32410 7679
rect 32257 7530 32410 7540
rect 33612 7321 33672 7331
rect 33612 7249 33672 7259
rect 29810 6779 29896 6789
rect 31458 6756 31551 6760
rect 29810 6668 29896 6678
rect 31428 6750 31565 6756
rect 31428 6673 31458 6750
rect 31551 6749 31565 6750
rect 31551 6739 33174 6749
rect 31551 6683 33121 6739
rect 31551 6673 33174 6683
rect 31428 6666 31565 6673
rect 31458 6663 31551 6666
rect 33245 6636 33318 6646
rect 31465 6627 31532 6628
rect 31725 6627 33245 6636
rect 31457 6626 33245 6627
rect 31457 6618 31725 6626
rect 29582 6605 29667 6615
rect 29582 6535 29667 6545
rect 30297 6595 30359 6597
rect 30297 6587 30361 6595
rect 30359 6585 30361 6587
rect 31457 6555 31465 6618
rect 31532 6558 31725 6618
rect 31780 6558 33245 6626
rect 31532 6555 33245 6558
rect 31457 6548 33245 6555
rect 31458 6547 31547 6548
rect 31465 6545 31532 6547
rect 33245 6537 33318 6547
rect 30297 6513 30361 6523
rect 35009 6405 35115 9458
rect 37444 9418 37529 9458
rect 37561 9440 37646 9468
rect 37728 9455 37737 9528
rect 37807 9455 37814 9528
rect 37444 9292 37528 9418
rect 37442 9281 37528 9292
rect 37442 9210 37454 9281
rect 37517 9210 37528 9281
rect 37442 9199 37528 9210
rect 37444 8196 37528 9199
rect 36473 8046 36483 8146
rect 36575 8046 36585 8146
rect 37444 8126 37454 8196
rect 37516 8126 37528 8196
rect 37444 8117 37528 8126
rect 37564 7955 37643 9440
rect 37728 9422 37814 9455
rect 37729 8314 37813 9422
rect 37729 8246 37737 8314
rect 37802 8246 37813 8314
rect 37729 8235 37813 8246
rect 38717 8050 38727 8126
rect 38785 8050 38795 8126
rect 37564 7896 37574 7955
rect 37634 7896 37644 7955
rect 35009 6404 37509 6405
rect 34072 6398 34554 6399
rect 32779 6388 34554 6398
rect 32841 6387 34554 6388
rect 32841 6297 34428 6387
rect 32779 6296 34428 6297
rect 34538 6296 34554 6387
rect 32779 6287 34554 6296
rect 35009 6326 37524 6404
rect 37557 6393 37642 6404
rect 37724 6393 37809 6404
rect 37555 6336 37565 6393
rect 37633 6336 37643 6393
rect 37723 6336 37733 6393
rect 37801 6336 37811 6393
rect 34428 6286 34538 6287
rect 33834 6125 33896 6127
rect 33834 6117 33898 6125
rect 33896 6115 33898 6117
rect 33834 6043 33898 6053
rect 32179 5339 32390 5349
rect 32179 5172 32390 5182
rect 30072 4721 30132 4731
rect 30072 4649 30132 4659
rect 29412 3785 29496 3795
rect 29412 3686 29496 3695
rect 29242 3649 29880 3651
rect 29242 3648 29905 3649
rect 29242 3638 29912 3648
rect 29242 3574 29846 3638
rect 29242 3564 29912 3574
rect 31023 3621 34559 3709
rect 29242 3562 29837 3564
rect 24890 3512 25194 3518
rect 30294 3525 30356 3527
rect 30294 3517 30358 3525
rect 30356 3515 30358 3517
rect 24895 3508 24958 3512
rect 30294 3443 30358 3453
rect 24568 3140 24578 3293
rect 24707 3140 24717 3293
rect 26061 3196 26214 3206
rect 26061 3057 26214 3067
rect 27959 3196 28112 3206
rect 27959 3057 28112 3067
rect 10568 3039 10685 3049
rect 10568 2933 10573 3039
rect 17223 3040 17340 3050
rect 4017 2924 4133 2925
rect 10568 2923 10685 2933
rect 16384 3002 16552 3012
rect 10568 2922 10684 2923
rect 16384 2915 16411 3002
rect 16513 2915 16552 3002
rect 17223 2934 17228 3040
rect 17223 2924 17340 2934
rect 23845 3041 23962 3051
rect 23845 2935 23850 3041
rect 23845 2925 23962 2935
rect 23845 2924 23961 2925
rect 17223 2923 17339 2924
rect 16384 2667 16552 2915
rect 31023 2667 31117 3621
rect 32257 3321 32410 3331
rect 32257 3182 32410 3192
rect 33612 2973 33672 2983
rect 33612 2901 33672 2911
rect 16384 2493 31117 2667
rect 16483 2492 31117 2493
rect 31465 2401 31532 2406
rect 31458 2396 33174 2401
rect 8410 2374 8474 2384
rect 8472 2310 8474 2312
rect 8410 2302 8474 2310
rect 14964 2379 15028 2389
rect 15026 2315 15028 2317
rect 14964 2307 15028 2315
rect 21613 2367 21677 2377
rect 14964 2305 15026 2307
rect 31458 2333 31465 2396
rect 31532 2391 33174 2396
rect 31532 2335 33121 2391
rect 31532 2333 33174 2335
rect 31458 2325 33174 2333
rect 31465 2323 31532 2325
rect 34210 2308 34352 2309
rect 34445 2308 34559 3621
rect 35009 3260 35115 6326
rect 37440 6160 37524 6326
rect 37557 6308 37642 6336
rect 37724 6308 37809 6336
rect 37438 6149 37524 6160
rect 37438 6078 37450 6149
rect 37513 6078 37524 6149
rect 37438 6067 37524 6078
rect 37440 5064 37524 6067
rect 36469 4914 36479 5014
rect 36571 4914 36581 5014
rect 37440 4994 37450 5064
rect 37512 4994 37524 5064
rect 37440 4985 37524 4994
rect 37560 4823 37639 6308
rect 37725 5182 37809 6308
rect 37725 5114 37733 5182
rect 37798 5114 37809 5182
rect 37725 5103 37809 5114
rect 38713 4918 38723 4994
rect 38781 4918 38791 4994
rect 37560 4764 37570 4823
rect 37630 4764 37640 4823
rect 35009 3182 37524 3260
rect 37557 3249 37642 3260
rect 37724 3249 37809 3259
rect 37555 3192 37565 3249
rect 37633 3192 37643 3249
rect 37723 3192 37733 3249
rect 37801 3192 37811 3249
rect 37440 3016 37524 3182
rect 37557 3164 37642 3192
rect 37724 3164 37809 3192
rect 37438 3005 37524 3016
rect 37438 2934 37450 3005
rect 37513 2934 37524 3005
rect 37438 2923 37524 2934
rect 21675 2303 21677 2305
rect 8410 2300 8472 2302
rect 21613 2295 21677 2303
rect 34197 2299 34559 2308
rect 21613 2293 21675 2295
rect 33245 2288 33318 2298
rect 31465 2279 31532 2280
rect 31725 2279 33245 2288
rect 31457 2278 33245 2279
rect 31457 2270 31725 2278
rect 31457 2207 31465 2270
rect 31532 2210 31725 2270
rect 31780 2210 33245 2278
rect 31532 2207 33245 2210
rect 31457 2200 33245 2207
rect 31458 2199 31547 2200
rect 34197 2211 34210 2299
rect 34352 2211 34559 2299
rect 34197 2200 34559 2211
rect 31465 2197 31532 2199
rect 33245 2189 33318 2199
rect 7471 2139 7547 2141
rect 2604 819 2616 888
rect 2712 819 2722 888
rect 2604 813 2722 819
rect 7464 2131 7556 2139
rect 7464 2045 7471 2131
rect 7547 2045 7556 2131
rect 2616 809 2712 813
rect 7464 639 7556 2045
rect 29826 2125 29910 2135
rect 34961 2051 35087 2052
rect 34151 2050 35087 2051
rect 29826 2025 29910 2035
rect 32779 2040 35087 2050
rect 7651 2004 7831 2014
rect 7651 1913 7702 2004
rect 20899 1995 20968 2005
rect 7651 1903 7831 1913
rect 20891 1906 20899 1995
rect 20968 1906 20969 1995
rect 32841 2034 35087 2040
rect 32841 1961 34981 2034
rect 35068 1961 35087 2034
rect 32841 1949 35087 1961
rect 32779 1942 35087 1949
rect 32779 1939 34968 1942
rect 7651 892 7760 1903
rect 8188 1168 8248 1178
rect 8188 1096 8248 1106
rect 14742 1173 14802 1183
rect 14742 1101 14802 1111
rect 7651 818 7656 892
rect 7756 818 7760 892
rect 7651 812 7760 818
rect 7656 808 7756 812
rect 7464 557 7556 567
rect 20891 747 20969 1906
rect 37440 1920 37524 2923
rect 30079 1876 30139 1886
rect 30079 1804 30139 1814
rect 33834 1777 33896 1779
rect 33834 1769 33898 1777
rect 36469 1770 36479 1870
rect 36571 1770 36581 1870
rect 37440 1850 37450 1920
rect 37512 1850 37524 1920
rect 37440 1841 37524 1850
rect 33896 1767 33898 1769
rect 33834 1695 33898 1705
rect 37560 1679 37639 3164
rect 37725 2038 37809 3164
rect 37725 1970 37733 2038
rect 37798 1970 37809 2038
rect 37725 1959 37809 1970
rect 38713 1774 38723 1850
rect 38781 1774 38791 1850
rect 37560 1620 37570 1679
rect 37630 1620 37640 1679
rect 29241 1382 29325 1392
rect 29241 1282 29325 1292
rect 21391 1161 21451 1171
rect 21391 1089 21451 1099
rect 29410 1066 29494 1076
rect 29410 966 29494 976
rect 32179 991 32390 1001
rect 32179 824 32390 834
rect 20891 632 20970 747
rect 29723 717 29784 727
rect 29723 632 29784 642
rect 30301 680 30363 682
rect 30301 672 30365 680
rect 30363 670 30365 672
rect 20891 564 20896 632
rect 20965 564 20970 632
rect 30301 598 30365 608
rect 20891 561 20970 564
rect 20896 554 20965 561
rect 2455 156 2462 210
rect 2557 204 2562 210
rect 2557 156 2561 204
rect 2455 145 2561 156
rect -2690 128 -2604 138
rect -2690 33 -2604 43
<< via2 >>
rect -845 23393 -661 23405
rect -845 23256 -832 23393
rect -832 23256 -674 23393
rect -674 23256 -661 23393
rect -845 23244 -661 23256
rect 8754 27960 8907 27971
rect 6272 27906 6425 27917
rect 6272 27798 6283 27906
rect 6283 27798 6415 27906
rect 6415 27798 6425 27906
rect 8754 27852 8765 27960
rect 8765 27852 8897 27960
rect 8897 27852 8907 27960
rect 9901 27960 10054 27971
rect 8754 27842 8907 27852
rect 6272 27788 6425 27798
rect 9901 27852 9912 27960
rect 9912 27852 10044 27960
rect 10044 27852 10054 27960
rect 15267 27957 15420 27968
rect 9901 27842 10054 27852
rect 12785 27903 12938 27914
rect 6553 26867 6682 26878
rect 6553 26735 6563 26867
rect 6563 26735 6671 26867
rect 6671 26735 6682 26867
rect 6553 26725 6682 26735
rect 5091 26165 5233 26268
rect 6286 26256 6439 26267
rect 6286 26148 6297 26256
rect 6297 26148 6429 26256
rect 6429 26148 6439 26256
rect 6286 26138 6439 26148
rect 5051 25037 5189 25163
rect 6567 25217 6696 25228
rect 6567 25085 6577 25217
rect 6577 25085 6685 25217
rect 6685 25085 6696 25217
rect 6567 25075 6696 25085
rect 5319 24780 5434 24789
rect 5319 24701 5329 24780
rect 5329 24701 5422 24780
rect 5422 24701 5434 24780
rect 5319 24692 5434 24701
rect 6281 24652 6434 24663
rect 6281 24544 6292 24652
rect 6292 24544 6424 24652
rect 6424 24544 6434 24652
rect 6281 24534 6434 24544
rect 12785 27795 12796 27903
rect 12796 27795 12928 27903
rect 12928 27795 12938 27903
rect 15267 27849 15278 27957
rect 15278 27849 15410 27957
rect 15410 27849 15420 27957
rect 16414 27957 16567 27968
rect 15267 27839 15420 27849
rect 12785 27785 12938 27795
rect 16414 27849 16425 27957
rect 16425 27849 16557 27957
rect 16557 27849 16567 27957
rect 21801 27952 21954 27963
rect 16414 27839 16567 27849
rect 19319 27898 19472 27909
rect 13066 26864 13195 26875
rect 13066 26732 13076 26864
rect 13076 26732 13184 26864
rect 13184 26732 13195 26864
rect 13066 26722 13195 26732
rect 8101 26560 8254 26570
rect 8101 26452 8111 26560
rect 8111 26452 8243 26560
rect 8243 26452 8254 26560
rect 8101 26441 8254 26452
rect 9243 26558 9396 26568
rect 9243 26450 9253 26558
rect 9253 26450 9385 26558
rect 9385 26450 9396 26558
rect 9243 26439 9396 26450
rect 8099 25913 8252 25924
rect 8099 25805 8110 25913
rect 8110 25805 8242 25913
rect 8242 25805 8252 25913
rect 8099 25795 8252 25805
rect 9997 25913 10150 25924
rect 9997 25805 10008 25913
rect 10008 25805 10140 25913
rect 10140 25805 10150 25913
rect 9997 25795 10150 25805
rect 8740 24943 8818 24953
rect 8740 24877 8755 24943
rect 8755 24877 8818 24943
rect 8740 24867 8818 24877
rect 6562 23613 6691 23624
rect 6562 23481 6572 23613
rect 6572 23481 6680 23613
rect 6680 23481 6691 23613
rect 6562 23471 6691 23481
rect 8045 23517 8198 23527
rect 8045 23409 8055 23517
rect 8055 23409 8187 23517
rect 8187 23409 8198 23517
rect 8045 23398 8198 23409
rect 9943 23517 10096 23527
rect 9943 23409 9953 23517
rect 9953 23409 10085 23517
rect 10085 23409 10096 23517
rect 9943 23398 10096 23409
rect 11523 26170 11752 26294
rect 12799 26253 12952 26264
rect 12799 26145 12810 26253
rect 12810 26145 12942 26253
rect 12942 26145 12952 26253
rect 12799 26135 12952 26145
rect 13080 25214 13209 25225
rect 13080 25082 13090 25214
rect 13090 25082 13198 25214
rect 13198 25082 13209 25214
rect 13080 25072 13209 25082
rect 11832 24777 11947 24786
rect 11832 24698 11842 24777
rect 11842 24698 11935 24777
rect 11935 24698 11947 24777
rect 11832 24689 11947 24698
rect 12794 24649 12947 24660
rect 12794 24541 12805 24649
rect 12805 24541 12937 24649
rect 12937 24541 12947 24649
rect 12794 24531 12947 24541
rect 19319 27790 19330 27898
rect 19330 27790 19462 27898
rect 19462 27790 19472 27898
rect 21801 27844 21812 27952
rect 21812 27844 21944 27952
rect 21944 27844 21954 27952
rect 22948 27952 23101 27963
rect 21801 27834 21954 27844
rect 19319 27780 19472 27790
rect 22948 27844 22959 27952
rect 22959 27844 23091 27952
rect 23091 27844 23101 27952
rect 28359 27956 28512 27967
rect 22948 27834 23101 27844
rect 25877 27902 26030 27913
rect 19600 26859 19729 26870
rect 19600 26727 19610 26859
rect 19610 26727 19718 26859
rect 19718 26727 19729 26859
rect 19600 26717 19729 26727
rect 14614 26557 14767 26567
rect 14614 26449 14624 26557
rect 14624 26449 14756 26557
rect 14756 26449 14767 26557
rect 14614 26438 14767 26449
rect 15756 26555 15909 26565
rect 15756 26447 15766 26555
rect 15766 26447 15898 26555
rect 15898 26447 15909 26555
rect 15756 26436 15909 26447
rect 14612 25910 14765 25921
rect 14612 25802 14623 25910
rect 14623 25802 14755 25910
rect 14755 25802 14765 25910
rect 14612 25792 14765 25802
rect 16510 25910 16663 25921
rect 16510 25802 16521 25910
rect 16521 25802 16653 25910
rect 16653 25802 16663 25910
rect 16510 25792 16663 25802
rect 15253 24940 15331 24950
rect 15253 24874 15268 24940
rect 15268 24874 15331 24940
rect 15253 24864 15331 24874
rect 13075 23610 13204 23621
rect 13075 23478 13085 23610
rect 13085 23478 13193 23610
rect 13193 23478 13204 23610
rect 13075 23468 13204 23478
rect 14558 23514 14711 23524
rect 14558 23406 14568 23514
rect 14568 23406 14700 23514
rect 14700 23406 14711 23514
rect 14558 23395 14711 23406
rect 16456 23514 16609 23524
rect 16456 23406 16466 23514
rect 16466 23406 16598 23514
rect 16598 23406 16609 23514
rect 16456 23395 16609 23406
rect 18082 26160 18300 26300
rect 19333 26248 19486 26259
rect 19333 26140 19344 26248
rect 19344 26140 19476 26248
rect 19476 26140 19486 26248
rect 19333 26130 19486 26140
rect 19614 25209 19743 25220
rect 19614 25077 19624 25209
rect 19624 25077 19732 25209
rect 19732 25077 19743 25209
rect 19614 25067 19743 25077
rect 18366 24772 18481 24781
rect 18366 24693 18376 24772
rect 18376 24693 18469 24772
rect 18469 24693 18481 24772
rect 18366 24684 18481 24693
rect 19328 24644 19481 24655
rect 19328 24536 19339 24644
rect 19339 24536 19471 24644
rect 19471 24536 19481 24644
rect 19328 24526 19481 24536
rect 25877 27794 25888 27902
rect 25888 27794 26020 27902
rect 26020 27794 26030 27902
rect 28359 27848 28370 27956
rect 28370 27848 28502 27956
rect 28502 27848 28512 27956
rect 29506 27956 29659 27967
rect 28359 27838 28512 27848
rect 25877 27784 26030 27794
rect 29506 27848 29517 27956
rect 29517 27848 29649 27956
rect 29649 27848 29659 27956
rect 29506 27838 29659 27848
rect 26158 26863 26287 26874
rect 26158 26731 26168 26863
rect 26168 26731 26276 26863
rect 26276 26731 26287 26863
rect 26158 26721 26287 26731
rect 21148 26552 21301 26562
rect 21148 26444 21158 26552
rect 21158 26444 21290 26552
rect 21290 26444 21301 26552
rect 21148 26433 21301 26444
rect 22290 26550 22443 26560
rect 22290 26442 22300 26550
rect 22300 26442 22432 26550
rect 22432 26442 22443 26550
rect 22290 26431 22443 26442
rect 21146 25905 21299 25916
rect 21146 25797 21157 25905
rect 21157 25797 21289 25905
rect 21289 25797 21299 25905
rect 21146 25787 21299 25797
rect 23044 25905 23197 25916
rect 23044 25797 23055 25905
rect 23055 25797 23187 25905
rect 23187 25797 23197 25905
rect 23044 25787 23197 25797
rect 21787 24935 21865 24945
rect 21787 24869 21802 24935
rect 21802 24869 21865 24935
rect 21787 24859 21865 24869
rect 19609 23605 19738 23616
rect 19609 23473 19619 23605
rect 19619 23473 19727 23605
rect 19727 23473 19738 23605
rect 19609 23463 19738 23473
rect 21092 23509 21245 23519
rect 21092 23401 21102 23509
rect 21102 23401 21234 23509
rect 21234 23401 21245 23509
rect 21092 23390 21245 23401
rect 22990 23509 23143 23519
rect 22990 23401 23000 23509
rect 23000 23401 23132 23509
rect 23132 23401 23143 23509
rect 22990 23390 23143 23401
rect 24606 26157 24858 26302
rect 25891 26252 26044 26263
rect 25891 26144 25902 26252
rect 25902 26144 26034 26252
rect 26034 26144 26044 26252
rect 25891 26134 26044 26144
rect 26172 25213 26301 25224
rect 26172 25081 26182 25213
rect 26182 25081 26290 25213
rect 26290 25081 26301 25213
rect 26172 25071 26301 25081
rect 24924 24776 25039 24785
rect 24924 24697 24934 24776
rect 24934 24697 25027 24776
rect 25027 24697 25039 24776
rect 24924 24688 25039 24697
rect 25886 24648 26039 24659
rect 25886 24540 25897 24648
rect 25897 24540 26029 24648
rect 26029 24540 26039 24648
rect 25886 24530 26039 24540
rect 27706 26556 27859 26566
rect 27706 26448 27716 26556
rect 27716 26448 27848 26556
rect 27848 26448 27859 26556
rect 27706 26437 27859 26448
rect 28848 26554 29001 26564
rect 28848 26446 28858 26554
rect 28858 26446 28990 26554
rect 28990 26446 29001 26554
rect 28848 26435 29001 26446
rect 27704 25909 27857 25920
rect 27704 25801 27715 25909
rect 27715 25801 27847 25909
rect 27847 25801 27857 25909
rect 27704 25791 27857 25801
rect 29602 25909 29755 25920
rect 29602 25801 29613 25909
rect 29613 25801 29745 25909
rect 29745 25801 29755 25909
rect 29602 25791 29755 25801
rect 28345 24939 28423 24949
rect 28345 24873 28360 24939
rect 28360 24873 28423 24939
rect 28345 24863 28423 24873
rect 26167 23609 26296 23620
rect 26167 23477 26177 23609
rect 26177 23477 26285 23609
rect 26285 23477 26296 23609
rect 26167 23467 26296 23477
rect 27650 23513 27803 23523
rect 27650 23405 27660 23513
rect 27660 23405 27792 23513
rect 27792 23405 27803 23513
rect 27650 23394 27803 23405
rect 29548 23513 29701 23523
rect 29548 23405 29558 23513
rect 29558 23405 29690 23513
rect 29690 23405 29701 23513
rect 29548 23394 29701 23405
rect 5850 22352 6003 22363
rect 5850 22244 5860 22352
rect 5860 22244 5992 22352
rect 5992 22244 6003 22352
rect 6997 22352 7150 22363
rect 5850 22234 6003 22244
rect 6997 22244 7007 22352
rect 7007 22244 7139 22352
rect 7139 22244 7150 22352
rect 12408 22348 12561 22359
rect 6997 22234 7150 22244
rect 9479 22298 9632 22309
rect 9479 22190 9489 22298
rect 9489 22190 9621 22298
rect 9621 22190 9632 22298
rect 12408 22240 12418 22348
rect 12418 22240 12550 22348
rect 12550 22240 12561 22348
rect 13555 22348 13708 22359
rect 12408 22230 12561 22240
rect 13555 22240 13565 22348
rect 13565 22240 13697 22348
rect 13697 22240 13708 22348
rect 18942 22353 19095 22364
rect 13555 22230 13708 22240
rect 16037 22294 16190 22305
rect 9479 22180 9632 22190
rect 6508 20950 6661 20960
rect 6508 20842 6519 20950
rect 6519 20842 6651 20950
rect 6651 20842 6661 20950
rect 6508 20831 6661 20842
rect 7650 20952 7803 20962
rect 7650 20844 7661 20952
rect 7661 20844 7793 20952
rect 7793 20844 7803 20952
rect 7650 20833 7803 20844
rect 5754 20305 5907 20316
rect 5754 20197 5764 20305
rect 5764 20197 5896 20305
rect 5896 20197 5907 20305
rect 5754 20187 5907 20197
rect 7652 20305 7805 20316
rect 7652 20197 7662 20305
rect 7662 20197 7794 20305
rect 7794 20197 7805 20305
rect 7652 20187 7805 20197
rect 7086 19335 7164 19345
rect 7086 19269 7149 19335
rect 7149 19269 7164 19335
rect 7086 19259 7164 19269
rect 16037 22186 16047 22294
rect 16047 22186 16179 22294
rect 16179 22186 16190 22294
rect 18942 22245 18952 22353
rect 18952 22245 19084 22353
rect 19084 22245 19095 22353
rect 20089 22353 20242 22364
rect 18942 22235 19095 22245
rect 20089 22245 20099 22353
rect 20099 22245 20231 22353
rect 20231 22245 20242 22353
rect 25455 22356 25608 22367
rect 20089 22235 20242 22245
rect 22571 22299 22724 22310
rect 16037 22176 16190 22186
rect 9222 21259 9351 21270
rect 9222 21127 9233 21259
rect 9233 21127 9341 21259
rect 9341 21127 9351 21259
rect 9222 21117 9351 21127
rect 9465 20648 9618 20659
rect 9465 20540 9475 20648
rect 9475 20540 9607 20648
rect 9607 20540 9618 20648
rect 9465 20530 9618 20540
rect 9208 19609 9337 19620
rect 9208 19477 9219 19609
rect 9219 19477 9327 19609
rect 9327 19477 9337 19609
rect 9208 19467 9337 19477
rect 9470 19044 9623 19055
rect 9470 18936 9480 19044
rect 9480 18936 9612 19044
rect 9612 18936 9623 19044
rect 9470 18926 9623 18936
rect 5808 17909 5961 17919
rect 5808 17801 5819 17909
rect 5819 17801 5951 17909
rect 5951 17801 5961 17909
rect 5808 17790 5961 17801
rect 7706 17909 7859 17919
rect 7706 17801 7717 17909
rect 7717 17801 7849 17909
rect 7849 17801 7859 17909
rect 9213 18005 9342 18016
rect 9213 17873 9224 18005
rect 9224 17873 9332 18005
rect 9332 17873 9342 18005
rect 9213 17863 9342 17873
rect 7706 17790 7859 17801
rect 10470 19172 10585 19181
rect 10470 19093 10482 19172
rect 10482 19093 10575 19172
rect 10575 19093 10585 19172
rect 10470 19084 10585 19093
rect 13066 20946 13219 20956
rect 13066 20838 13077 20946
rect 13077 20838 13209 20946
rect 13209 20838 13219 20946
rect 13066 20827 13219 20838
rect 14208 20948 14361 20958
rect 14208 20840 14219 20948
rect 14219 20840 14351 20948
rect 14351 20840 14361 20948
rect 14208 20829 14361 20840
rect 12312 20301 12465 20312
rect 12312 20193 12322 20301
rect 12322 20193 12454 20301
rect 12454 20193 12465 20301
rect 12312 20183 12465 20193
rect 14210 20301 14363 20312
rect 14210 20193 14220 20301
rect 14220 20193 14352 20301
rect 14352 20193 14363 20301
rect 14210 20183 14363 20193
rect 13644 19331 13722 19341
rect 13644 19265 13707 19331
rect 13707 19265 13722 19331
rect 13644 19255 13722 19265
rect 22571 22191 22581 22299
rect 22581 22191 22713 22299
rect 22713 22191 22724 22299
rect 25455 22248 25465 22356
rect 25465 22248 25597 22356
rect 25597 22248 25608 22356
rect 26602 22356 26755 22367
rect 25455 22238 25608 22248
rect 26602 22248 26612 22356
rect 26612 22248 26744 22356
rect 26744 22248 26755 22356
rect 26602 22238 26755 22248
rect 29084 22302 29237 22313
rect 22571 22181 22724 22191
rect 15780 21255 15909 21266
rect 15780 21123 15791 21255
rect 15791 21123 15899 21255
rect 15899 21123 15909 21255
rect 15780 21113 15909 21123
rect 19600 20951 19753 20961
rect 19600 20843 19611 20951
rect 19611 20843 19743 20951
rect 19743 20843 19753 20951
rect 19600 20832 19753 20843
rect 20742 20953 20895 20963
rect 20742 20845 20753 20953
rect 20753 20845 20885 20953
rect 20885 20845 20895 20953
rect 20742 20834 20895 20845
rect 16023 20644 16176 20655
rect 16023 20536 16033 20644
rect 16033 20536 16165 20644
rect 16165 20536 16176 20644
rect 16023 20526 16176 20536
rect 15766 19605 15895 19616
rect 15766 19473 15777 19605
rect 15777 19473 15885 19605
rect 15885 19473 15895 19605
rect 15766 19463 15895 19473
rect 16028 19040 16181 19051
rect 16028 18932 16038 19040
rect 16038 18932 16170 19040
rect 16170 18932 16181 19040
rect 16028 18922 16181 18932
rect 12366 17905 12519 17915
rect 12366 17797 12377 17905
rect 12377 17797 12509 17905
rect 12509 17797 12519 17905
rect 12366 17786 12519 17797
rect 14264 17905 14417 17915
rect 14264 17797 14275 17905
rect 14275 17797 14407 17905
rect 14407 17797 14417 17905
rect 15771 18001 15900 18012
rect 15771 17869 15782 18001
rect 15782 17869 15890 18001
rect 15890 17869 15900 18001
rect 15771 17859 15900 17869
rect 14264 17786 14417 17797
rect 17028 19168 17143 19177
rect 17028 19089 17040 19168
rect 17040 19089 17133 19168
rect 17133 19089 17143 19168
rect 17028 19080 17143 19089
rect 18846 20306 18999 20317
rect 18846 20198 18856 20306
rect 18856 20198 18988 20306
rect 18988 20198 18999 20306
rect 18846 20188 18999 20198
rect 20744 20306 20897 20317
rect 20744 20198 20754 20306
rect 20754 20198 20886 20306
rect 20886 20198 20897 20306
rect 20744 20188 20897 20198
rect 20178 19336 20256 19346
rect 20178 19270 20241 19336
rect 20241 19270 20256 19336
rect 20178 19260 20256 19270
rect 29084 22194 29094 22302
rect 29094 22194 29226 22302
rect 29226 22194 29237 22302
rect 29084 22184 29237 22194
rect 22314 21260 22443 21271
rect 22314 21128 22325 21260
rect 22325 21128 22433 21260
rect 22433 21128 22443 21260
rect 22314 21118 22443 21128
rect 22557 20649 22710 20660
rect 22557 20541 22567 20649
rect 22567 20541 22699 20649
rect 22699 20541 22710 20649
rect 22557 20531 22710 20541
rect 22300 19610 22429 19621
rect 22300 19478 22311 19610
rect 22311 19478 22419 19610
rect 22419 19478 22429 19610
rect 22300 19468 22429 19478
rect 22562 19045 22715 19056
rect 22562 18937 22572 19045
rect 22572 18937 22704 19045
rect 22704 18937 22715 19045
rect 22562 18927 22715 18937
rect 18900 17910 19053 17920
rect 18900 17802 18911 17910
rect 18911 17802 19043 17910
rect 19043 17802 19053 17910
rect 18900 17791 19053 17802
rect 20798 17910 20951 17920
rect 20798 17802 20809 17910
rect 20809 17802 20941 17910
rect 20941 17802 20951 17910
rect 22305 18006 22434 18017
rect 22305 17874 22316 18006
rect 22316 17874 22424 18006
rect 22424 17874 22434 18006
rect 22305 17864 22434 17874
rect 20798 17791 20951 17802
rect 23562 19173 23677 19182
rect 23562 19094 23574 19173
rect 23574 19094 23667 19173
rect 23667 19094 23677 19173
rect 23562 19085 23677 19094
rect 26113 20954 26266 20964
rect 26113 20846 26124 20954
rect 26124 20846 26256 20954
rect 26256 20846 26266 20954
rect 26113 20835 26266 20846
rect 27255 20956 27408 20966
rect 27255 20848 27266 20956
rect 27266 20848 27398 20956
rect 27398 20848 27408 20956
rect 27255 20837 27408 20848
rect 25359 20309 25512 20320
rect 25359 20201 25369 20309
rect 25369 20201 25501 20309
rect 25501 20201 25512 20309
rect 25359 20191 25512 20201
rect 27257 20309 27410 20320
rect 27257 20201 27267 20309
rect 27267 20201 27399 20309
rect 27399 20201 27410 20309
rect 27257 20191 27410 20201
rect 26691 19339 26769 19349
rect 26691 19273 26754 19339
rect 26754 19273 26769 19339
rect 26691 19263 26769 19273
rect 28827 21263 28956 21274
rect 28827 21131 28838 21263
rect 28838 21131 28946 21263
rect 28946 21131 28956 21263
rect 28827 21121 28956 21131
rect 29070 20652 29223 20663
rect 29070 20544 29080 20652
rect 29080 20544 29212 20652
rect 29212 20544 29223 20652
rect 30262 20568 30480 20724
rect 29070 20534 29223 20544
rect 28813 19613 28942 19624
rect 28813 19481 28824 19613
rect 28824 19481 28932 19613
rect 28932 19481 28942 19613
rect 28813 19471 28942 19481
rect 29075 19048 29228 19059
rect 29075 18940 29085 19048
rect 29085 18940 29217 19048
rect 29217 18940 29228 19048
rect 29075 18930 29228 18940
rect 25413 17913 25566 17923
rect 25413 17805 25424 17913
rect 25424 17805 25556 17913
rect 25556 17805 25566 17913
rect 25413 17794 25566 17805
rect 27311 17913 27464 17923
rect 27311 17805 27322 17913
rect 27322 17805 27454 17913
rect 27454 17805 27464 17913
rect 28818 18009 28947 18020
rect 28818 17877 28829 18009
rect 28829 17877 28937 18009
rect 28937 17877 28947 18009
rect 28818 17867 28947 17877
rect 27311 17794 27464 17805
rect 30075 19176 30190 19185
rect 30075 19097 30087 19176
rect 30087 19097 30180 19176
rect 30180 19097 30190 19176
rect 30075 19088 30190 19097
rect -4063 15428 -3993 15440
rect -4063 15374 -4055 15428
rect -4055 15374 -4001 15428
rect -4001 15374 -3993 15428
rect -4063 15362 -3993 15374
rect 23966 16251 24065 16267
rect 23966 16176 23973 16251
rect 23973 16176 24059 16251
rect 24059 16176 24065 16251
rect 23966 16165 24065 16176
rect 17441 16130 17541 16137
rect 17441 16060 17450 16130
rect 17450 16060 17537 16130
rect 17537 16060 17541 16130
rect 17441 16052 17541 16060
rect 10861 15797 10979 15801
rect 10861 15736 10875 15797
rect 10875 15736 10968 15797
rect 10968 15736 10979 15797
rect 10861 15733 10979 15736
rect -1833 15486 -1763 15492
rect -1833 15424 -1831 15486
rect -1831 15424 -1773 15486
rect -1773 15424 -1763 15486
rect -1833 15420 -1763 15424
rect 8153 15400 8213 15462
rect 14702 15399 14762 15461
rect 21356 15420 21416 15482
rect 30009 15253 30069 15315
rect 32255 15244 32408 15255
rect 32255 15136 32266 15244
rect 32266 15136 32398 15244
rect 32398 15136 32408 15244
rect 32255 15126 32408 15136
rect 33610 14845 33670 14907
rect -2694 14605 -2598 14613
rect -2694 14528 -2684 14605
rect -2684 14528 -2605 14605
rect -2605 14528 -2598 14605
rect -2694 14516 -2598 14528
rect 8375 14198 8437 14256
rect 8437 14198 8439 14256
rect 8375 14194 8439 14198
rect 14924 14197 14986 14255
rect 14986 14197 14988 14255
rect 21578 14218 21640 14276
rect 21640 14218 21642 14276
rect 21578 14214 21642 14218
rect 14924 14193 14988 14197
rect -4065 13360 -3995 13372
rect -4065 13306 -4057 13360
rect -4057 13306 -4003 13360
rect -4003 13306 -3995 13360
rect -4065 13294 -3995 13306
rect 349 13982 465 14038
rect 34219 14217 34357 14229
rect 34219 14159 34232 14217
rect 34232 14159 34344 14217
rect 34344 14159 34357 14217
rect 34219 14147 34357 14159
rect 30231 14051 30293 14109
rect 30293 14051 30295 14109
rect 30231 14047 30295 14051
rect 1489 13500 1549 13562
rect -1835 13418 -1765 13424
rect -1835 13356 -1833 13418
rect -1833 13356 -1775 13418
rect -1775 13356 -1765 13418
rect -1835 13352 -1765 13356
rect -2692 12536 -2600 12543
rect -2692 12462 -2681 12536
rect -2681 12462 -2610 12536
rect -2610 12462 -2600 12536
rect -2692 12451 -2600 12462
rect -4063 11291 -3993 11303
rect -4063 11237 -4055 11291
rect -4055 11237 -4001 11291
rect -4001 11237 -3993 11291
rect -4063 11225 -3993 11237
rect -1833 11349 -1763 11355
rect -1833 11287 -1831 11349
rect -1831 11287 -1773 11349
rect -1773 11287 -1763 11349
rect -1833 11283 -1763 11287
rect -2686 10459 -2601 10471
rect -2686 10394 -2674 10459
rect -2674 10394 -2611 10459
rect -2611 10394 -2601 10459
rect -2686 10385 -2601 10394
rect -4065 9223 -3995 9235
rect -4065 9169 -4057 9223
rect -4057 9169 -4003 9223
rect -4003 9169 -3995 9223
rect -4065 9157 -3995 9169
rect -1835 9281 -1765 9287
rect -1835 9219 -1833 9281
rect -1833 9219 -1775 9281
rect -1775 9219 -1765 9281
rect -1835 9215 -1765 9219
rect -2691 8391 -2602 8401
rect -2691 8327 -2682 8391
rect -2682 8327 -2609 8391
rect -2609 8327 -2602 8391
rect -2691 8316 -2602 8327
rect -4065 7154 -3995 7166
rect -4065 7100 -4057 7154
rect -4057 7100 -4003 7154
rect -4003 7100 -3995 7154
rect -4065 7088 -3995 7100
rect -1835 7212 -1765 7218
rect -1835 7150 -1833 7212
rect -1833 7150 -1775 7212
rect -1775 7150 -1765 7212
rect -1835 7146 -1765 7150
rect -2688 6325 -2604 6332
rect -2688 6259 -2679 6325
rect -2679 6259 -2614 6325
rect -2614 6259 -2604 6325
rect -2688 6249 -2604 6259
rect -4067 5086 -3997 5098
rect -4067 5032 -4059 5086
rect -4059 5032 -4005 5086
rect -4005 5032 -3997 5086
rect -4067 5020 -3997 5032
rect -1837 5144 -1767 5150
rect -1837 5082 -1835 5144
rect -1835 5082 -1777 5144
rect -1777 5082 -1767 5144
rect -1837 5078 -1767 5082
rect -2689 4258 -2606 4265
rect -2689 4188 -2679 4258
rect -2679 4188 -2614 4258
rect -2614 4188 -2606 4258
rect -2689 4181 -2606 4188
rect 1711 12298 1773 12356
rect 1773 12298 1775 12356
rect 1711 12294 1775 12298
rect 1481 10915 1541 10977
rect 1703 9713 1765 9771
rect 1765 9713 1767 9771
rect 1703 9709 1767 9713
rect 356 4119 459 4127
rect 356 4056 369 4119
rect 369 4056 450 4119
rect 450 4056 459 4119
rect 356 4048 459 4056
rect -4065 3017 -3995 3029
rect -4065 2963 -4057 3017
rect -4057 2963 -4003 3017
rect -4003 2963 -3995 3017
rect -4065 2951 -3995 2963
rect -1835 3075 -1765 3081
rect -1835 3013 -1833 3075
rect -1833 3013 -1775 3075
rect -1775 3013 -1765 3075
rect -1835 3009 -1765 3013
rect -2691 2189 -2601 2196
rect -2691 2119 -2682 2189
rect -2682 2119 -2609 2189
rect -2609 2119 -2601 2189
rect -2691 2109 -2601 2119
rect -4067 949 -3997 961
rect -4067 895 -4059 949
rect -4059 895 -4005 949
rect -4005 895 -3997 949
rect -4067 883 -3997 895
rect -1837 1007 -1767 1013
rect -1837 945 -1835 1007
rect -1835 945 -1777 1007
rect -1777 945 -1767 1007
rect -1837 941 -1767 945
rect 1462 7637 1522 7699
rect 1684 6435 1746 6493
rect 1746 6435 1748 6493
rect 1684 6431 1748 6435
rect 1478 4877 1538 4939
rect 1700 3675 1762 3733
rect 1762 3675 1764 3733
rect 1700 3671 1764 3675
rect 33832 13643 33894 13701
rect 33894 13643 33896 13701
rect 33832 13639 33896 13643
rect 13499 13497 13652 13508
rect 11017 13443 11170 13454
rect 6950 13409 7103 13420
rect 4468 13355 4621 13366
rect 4468 13247 4479 13355
rect 4479 13247 4611 13355
rect 4611 13247 4621 13355
rect 6950 13301 6961 13409
rect 6961 13301 7093 13409
rect 7093 13301 7103 13409
rect 8097 13409 8250 13420
rect 6950 13291 7103 13301
rect 4468 13237 4621 13247
rect 8097 13301 8108 13409
rect 8108 13301 8240 13409
rect 8240 13301 8250 13409
rect 11017 13335 11028 13443
rect 11028 13335 11160 13443
rect 11160 13335 11170 13443
rect 13499 13389 13510 13497
rect 13510 13389 13642 13497
rect 13642 13389 13652 13497
rect 14646 13497 14799 13508
rect 13499 13379 13652 13389
rect 11017 13325 11170 13335
rect 14646 13389 14657 13497
rect 14657 13389 14789 13497
rect 14789 13389 14799 13497
rect 26778 13497 26931 13508
rect 20153 13429 20306 13440
rect 14646 13379 14799 13389
rect 17671 13375 17824 13386
rect 8097 13291 8250 13301
rect 4749 12316 4878 12327
rect 4749 12184 4759 12316
rect 4759 12184 4867 12316
rect 4867 12184 4878 12316
rect 4749 12174 4878 12184
rect 4482 11705 4635 11716
rect 4482 11597 4493 11705
rect 4493 11597 4625 11705
rect 4625 11597 4635 11705
rect 4482 11587 4635 11597
rect 4763 10666 4892 10677
rect 4763 10534 4773 10666
rect 4773 10534 4881 10666
rect 4881 10534 4892 10666
rect 4763 10524 4892 10534
rect 3515 10229 3630 10238
rect 3515 10150 3525 10229
rect 3525 10150 3618 10229
rect 3618 10150 3630 10229
rect 3515 10141 3630 10150
rect 4477 10101 4630 10112
rect 4477 9993 4488 10101
rect 4488 9993 4620 10101
rect 4620 9993 4630 10101
rect 4477 9983 4630 9993
rect 9187 12501 9332 12576
rect 11298 12404 11427 12415
rect 11298 12272 11308 12404
rect 11308 12272 11416 12404
rect 11416 12272 11427 12404
rect 11298 12262 11427 12272
rect 6297 12009 6450 12019
rect 6297 11901 6307 12009
rect 6307 11901 6439 12009
rect 6439 11901 6450 12009
rect 6297 11890 6450 11901
rect 7439 12007 7592 12017
rect 7439 11899 7449 12007
rect 7449 11899 7581 12007
rect 7581 11899 7592 12007
rect 7439 11888 7592 11899
rect 11031 11793 11184 11804
rect 11031 11685 11042 11793
rect 11042 11685 11174 11793
rect 11174 11685 11184 11793
rect 11031 11675 11184 11685
rect 6295 11362 6448 11373
rect 6295 11254 6306 11362
rect 6306 11254 6438 11362
rect 6438 11254 6448 11362
rect 6295 11244 6448 11254
rect 8193 11362 8346 11373
rect 8193 11254 8204 11362
rect 8204 11254 8336 11362
rect 8336 11254 8346 11362
rect 8193 11244 8346 11254
rect 11312 10754 11441 10765
rect 11312 10622 11322 10754
rect 11322 10622 11430 10754
rect 11430 10622 11441 10754
rect 11312 10612 11441 10622
rect 6936 10392 7014 10402
rect 6936 10326 6951 10392
rect 6951 10326 7014 10392
rect 6936 10316 7014 10326
rect 4758 9062 4887 9073
rect 4758 8930 4768 9062
rect 4768 8930 4876 9062
rect 4876 8930 4887 9062
rect 4758 8920 4887 8930
rect 6241 8966 6394 8976
rect 6241 8858 6251 8966
rect 6251 8858 6383 8966
rect 6383 8858 6394 8966
rect 6241 8847 6394 8858
rect 8139 8966 8292 8976
rect 8139 8858 8149 8966
rect 8149 8858 8281 8966
rect 8281 8858 8292 8966
rect 8139 8847 8292 8858
rect 10064 10317 10179 10326
rect 10064 10238 10074 10317
rect 10074 10238 10167 10317
rect 10167 10238 10179 10317
rect 10064 10229 10179 10238
rect 11026 10189 11179 10200
rect 11026 10081 11037 10189
rect 11037 10081 11169 10189
rect 11169 10081 11179 10189
rect 11026 10071 11179 10081
rect 17671 13267 17682 13375
rect 17682 13267 17814 13375
rect 17814 13267 17824 13375
rect 20153 13321 20164 13429
rect 20164 13321 20296 13429
rect 20296 13321 20306 13429
rect 21300 13429 21453 13440
rect 20153 13311 20306 13321
rect 17671 13257 17824 13267
rect 21300 13321 21311 13429
rect 21311 13321 21443 13429
rect 21443 13321 21453 13429
rect 21300 13311 21453 13321
rect 24296 13443 24449 13454
rect 24296 13335 24307 13443
rect 24307 13335 24439 13443
rect 24439 13335 24449 13443
rect 26778 13389 26789 13497
rect 26789 13389 26921 13497
rect 26921 13389 26931 13497
rect 27925 13497 28078 13508
rect 26778 13379 26931 13389
rect 24296 13325 24449 13335
rect 27925 13389 27936 13497
rect 27936 13389 28068 13497
rect 28068 13389 28078 13497
rect 27925 13379 28078 13389
rect 17952 12336 18081 12347
rect 17952 12204 17962 12336
rect 17962 12204 18070 12336
rect 18070 12204 18081 12336
rect 17952 12194 18081 12204
rect 12846 12097 12999 12107
rect 12846 11989 12856 12097
rect 12856 11989 12988 12097
rect 12988 11989 12999 12097
rect 12846 11978 12999 11989
rect 13988 12095 14141 12105
rect 13988 11987 13998 12095
rect 13998 11987 14130 12095
rect 14130 11987 14141 12095
rect 13988 11976 14141 11987
rect 17685 11725 17838 11736
rect 17685 11617 17696 11725
rect 17696 11617 17828 11725
rect 17828 11617 17838 11725
rect 12844 11450 12997 11461
rect 12844 11342 12855 11450
rect 12855 11342 12987 11450
rect 12987 11342 12997 11450
rect 12844 11332 12997 11342
rect 14742 11450 14895 11461
rect 14742 11342 14753 11450
rect 14753 11342 14885 11450
rect 14885 11342 14895 11450
rect 14742 11332 14895 11342
rect 13485 10480 13563 10490
rect 13485 10414 13500 10480
rect 13500 10414 13563 10480
rect 13485 10404 13563 10414
rect 17685 11607 17838 11617
rect 17966 10686 18095 10697
rect 17966 10554 17976 10686
rect 17976 10554 18084 10686
rect 18084 10554 18095 10686
rect 17966 10544 18095 10554
rect 16718 10249 16833 10258
rect 16718 10170 16728 10249
rect 16728 10170 16821 10249
rect 16821 10170 16833 10249
rect 16718 10161 16833 10170
rect 11307 9150 11436 9161
rect 11307 9018 11317 9150
rect 11317 9018 11425 9150
rect 11425 9018 11436 9150
rect 11307 9008 11436 9018
rect 12790 9054 12943 9064
rect 12790 8946 12800 9054
rect 12800 8946 12932 9054
rect 12932 8946 12943 9054
rect 12790 8935 12943 8946
rect 14688 9054 14841 9064
rect 14688 8946 14698 9054
rect 14698 8946 14830 9054
rect 14830 8946 14841 9054
rect 14688 8935 14841 8946
rect 17680 10121 17833 10132
rect 17680 10013 17691 10121
rect 17691 10013 17823 10121
rect 17823 10013 17833 10121
rect 17680 10003 17833 10013
rect 22321 12522 22418 12596
rect 24577 12404 24706 12415
rect 24577 12272 24587 12404
rect 24587 12272 24695 12404
rect 24695 12272 24706 12404
rect 24577 12262 24706 12272
rect 19500 12029 19653 12039
rect 19500 11921 19510 12029
rect 19510 11921 19642 12029
rect 19642 11921 19653 12029
rect 19500 11910 19653 11921
rect 20642 12027 20795 12037
rect 20642 11919 20652 12027
rect 20652 11919 20784 12027
rect 20784 11919 20795 12027
rect 20642 11908 20795 11919
rect 24310 11793 24463 11804
rect 24310 11685 24321 11793
rect 24321 11685 24453 11793
rect 24453 11685 24463 11793
rect 24310 11675 24463 11685
rect 19498 11382 19651 11393
rect 19498 11274 19509 11382
rect 19509 11274 19641 11382
rect 19641 11274 19651 11382
rect 19498 11264 19651 11274
rect 21396 11382 21549 11393
rect 21396 11274 21407 11382
rect 21407 11274 21539 11382
rect 21539 11274 21549 11382
rect 21396 11264 21549 11274
rect 24591 10754 24720 10765
rect 24591 10622 24601 10754
rect 24601 10622 24709 10754
rect 24709 10622 24720 10754
rect 24591 10612 24720 10622
rect 20139 10412 20217 10422
rect 20139 10346 20154 10412
rect 20154 10346 20217 10412
rect 20139 10336 20217 10346
rect 22874 9811 22970 9911
rect 17961 9082 18090 9093
rect 17961 8950 17971 9082
rect 17971 8950 18079 9082
rect 18079 8950 18090 9082
rect 17961 8940 18090 8950
rect 19444 8986 19597 8996
rect 19444 8878 19454 8986
rect 19454 8878 19586 8986
rect 19586 8878 19597 8986
rect 19444 8867 19597 8878
rect 21342 8986 21495 8996
rect 21342 8878 21352 8986
rect 21352 8878 21484 8986
rect 21484 8878 21495 8986
rect 21342 8867 21495 8878
rect 22394 8599 22536 8607
rect 22394 8485 22405 8599
rect 22405 8485 22528 8599
rect 22528 8485 22536 8599
rect 22394 8473 22536 8485
rect 23343 10317 23458 10326
rect 23343 10238 23353 10317
rect 23353 10238 23446 10317
rect 23446 10238 23458 10317
rect 23343 10229 23458 10238
rect 24305 10189 24458 10200
rect 24305 10081 24316 10189
rect 24316 10081 24448 10189
rect 24448 10081 24458 10189
rect 24305 10071 24458 10081
rect 26125 12097 26278 12107
rect 26125 11989 26135 12097
rect 26135 11989 26267 12097
rect 26267 11989 26278 12097
rect 26125 11978 26278 11989
rect 27267 12095 27420 12105
rect 27267 11987 27277 12095
rect 27277 11987 27409 12095
rect 27409 11987 27420 12095
rect 27267 11976 27420 11987
rect 32177 12909 32388 12925
rect 32177 12786 32196 12909
rect 32196 12786 32370 12909
rect 32370 12786 32388 12909
rect 32177 12768 32388 12786
rect 30004 12682 30064 12744
rect 30226 11480 30288 11538
rect 30288 11480 30290 11538
rect 30226 11476 30290 11480
rect 26123 11450 26276 11461
rect 26123 11342 26134 11450
rect 26134 11342 26266 11450
rect 26266 11342 26276 11450
rect 26123 11332 26276 11342
rect 28021 11450 28174 11461
rect 28021 11342 28032 11450
rect 28032 11342 28164 11450
rect 28164 11342 28174 11450
rect 28021 11332 28174 11342
rect 32257 11153 32410 11164
rect 32257 11045 32268 11153
rect 32268 11045 32400 11153
rect 32400 11045 32410 11153
rect 32257 11035 32410 11045
rect 33612 10754 33672 10816
rect 26764 10480 26842 10490
rect 26764 10414 26779 10480
rect 26779 10414 26842 10480
rect 26764 10404 26842 10414
rect 36483 23900 36575 23912
rect 36483 23820 36511 23900
rect 36511 23820 36571 23900
rect 36571 23820 36575 23900
rect 36483 23812 36575 23820
rect 38727 23886 38785 23892
rect 38727 23820 38729 23886
rect 38729 23820 38781 23886
rect 38781 23820 38785 23886
rect 38727 23816 38785 23820
rect 36483 20756 36575 20768
rect 36483 20676 36511 20756
rect 36511 20676 36571 20756
rect 36571 20676 36575 20756
rect 36483 20668 36575 20676
rect 38727 20742 38785 20748
rect 38727 20676 38729 20742
rect 38729 20676 38781 20742
rect 38781 20676 38785 20742
rect 38727 20672 38785 20676
rect 36479 17624 36571 17636
rect 36479 17544 36507 17624
rect 36507 17544 36567 17624
rect 36567 17544 36571 17624
rect 36479 17536 36571 17544
rect 38723 17610 38781 17616
rect 38723 17544 38725 17610
rect 38725 17544 38777 17610
rect 38777 17544 38781 17610
rect 38723 17540 38781 17544
rect 36479 14480 36571 14492
rect 36479 14400 36507 14480
rect 36507 14400 36567 14480
rect 36567 14400 36571 14480
rect 36479 14392 36571 14400
rect 37736 15778 37799 15875
rect 38723 14466 38781 14472
rect 38723 14400 38725 14466
rect 38725 14400 38777 14466
rect 38777 14400 38781 14466
rect 38723 14396 38781 14400
rect 30004 9649 30064 9711
rect 33834 9552 33896 9610
rect 33896 9552 33898 9610
rect 33834 9548 33898 9552
rect 36483 11278 36575 11290
rect 36483 11198 36511 11278
rect 36511 11198 36571 11278
rect 36571 11198 36575 11278
rect 36483 11190 36575 11198
rect 38727 11264 38785 11270
rect 38727 11198 38729 11264
rect 38729 11198 38781 11264
rect 38781 11198 38785 11264
rect 38727 11194 38785 11198
rect 24586 9150 24715 9161
rect 24586 9018 24596 9150
rect 24596 9018 24704 9150
rect 24704 9018 24715 9150
rect 24586 9008 24715 9018
rect 26069 9054 26222 9064
rect 26069 8946 26079 9054
rect 26079 8946 26211 9054
rect 26211 8946 26222 9054
rect 26069 8935 26222 8946
rect 27967 9054 28120 9064
rect 27967 8946 27977 9054
rect 27977 8946 28109 9054
rect 28109 8946 28120 9054
rect 27967 8935 28120 8946
rect 23503 8599 23645 8607
rect 23503 8485 23514 8599
rect 23514 8485 23637 8599
rect 23637 8485 23645 8599
rect 23503 8473 23645 8485
rect 6942 7629 7095 7640
rect 4460 7575 4613 7586
rect 4460 7467 4471 7575
rect 4471 7467 4603 7575
rect 4603 7467 4613 7575
rect 6942 7521 6953 7629
rect 6953 7521 7085 7629
rect 7085 7521 7095 7629
rect 8089 7629 8242 7640
rect 6942 7511 7095 7521
rect 4460 7457 4613 7467
rect 8089 7521 8100 7629
rect 8100 7521 8232 7629
rect 8232 7521 8242 7629
rect 13493 7627 13646 7638
rect 8089 7511 8242 7521
rect 11011 7573 11164 7584
rect 4741 6536 4870 6547
rect 4741 6404 4751 6536
rect 4751 6404 4859 6536
rect 4859 6404 4870 6536
rect 4741 6394 4870 6404
rect 4474 5925 4627 5936
rect 4474 5817 4485 5925
rect 4485 5817 4617 5925
rect 4617 5817 4627 5925
rect 4474 5807 4627 5817
rect 3127 4706 3361 4843
rect 4755 4886 4884 4897
rect 4755 4754 4765 4886
rect 4765 4754 4873 4886
rect 4873 4754 4884 4886
rect 4755 4744 4884 4754
rect 3507 4449 3622 4458
rect 3507 4370 3517 4449
rect 3517 4370 3610 4449
rect 3610 4370 3622 4449
rect 3507 4361 3622 4370
rect 4469 4321 4622 4332
rect 4469 4213 4480 4321
rect 4480 4213 4612 4321
rect 4612 4213 4622 4321
rect 4469 4203 4622 4213
rect 11011 7465 11022 7573
rect 11022 7465 11154 7573
rect 11154 7465 11164 7573
rect 13493 7519 13504 7627
rect 13504 7519 13636 7627
rect 13636 7519 13646 7627
rect 14640 7627 14793 7638
rect 13493 7509 13646 7519
rect 11011 7455 11164 7465
rect 14640 7519 14651 7627
rect 14651 7519 14783 7627
rect 14783 7519 14793 7627
rect 14640 7509 14793 7519
rect 11292 6534 11421 6545
rect 11292 6402 11302 6534
rect 11302 6402 11410 6534
rect 11410 6402 11421 6534
rect 11292 6392 11421 6402
rect 6289 6229 6442 6239
rect 6289 6121 6299 6229
rect 6299 6121 6431 6229
rect 6431 6121 6442 6229
rect 6289 6110 6442 6121
rect 7431 6227 7584 6237
rect 7431 6119 7441 6227
rect 7441 6119 7573 6227
rect 7573 6119 7584 6227
rect 7431 6108 7584 6119
rect 11025 5923 11178 5934
rect 11025 5815 11036 5923
rect 11036 5815 11168 5923
rect 11168 5815 11178 5923
rect 11025 5805 11178 5815
rect 6287 5582 6440 5593
rect 6287 5474 6298 5582
rect 6298 5474 6430 5582
rect 6430 5474 6440 5582
rect 6287 5464 6440 5474
rect 8185 5582 8338 5593
rect 8185 5474 8196 5582
rect 8196 5474 8328 5582
rect 8328 5474 8338 5582
rect 8185 5464 8338 5474
rect 9762 4700 9985 4836
rect 11306 4884 11435 4895
rect 11306 4752 11316 4884
rect 11316 4752 11424 4884
rect 11424 4752 11435 4884
rect 11306 4742 11435 4752
rect 6928 4612 7006 4622
rect 6928 4546 6943 4612
rect 6943 4546 7006 4612
rect 6928 4536 7006 4546
rect 10058 4447 10173 4456
rect 10058 4368 10068 4447
rect 10068 4368 10161 4447
rect 10161 4368 10173 4447
rect 10058 4359 10173 4368
rect 4750 3282 4879 3293
rect 4750 3150 4760 3282
rect 4760 3150 4868 3282
rect 4868 3150 4879 3282
rect 4750 3140 4879 3150
rect 6233 3186 6386 3196
rect 6233 3078 6243 3186
rect 6243 3078 6375 3186
rect 6375 3078 6386 3186
rect 6233 3067 6386 3078
rect 8131 3186 8284 3196
rect 8131 3078 8141 3186
rect 8141 3078 8273 3186
rect 8273 3078 8284 3186
rect 8131 3067 8284 3078
rect 11020 4319 11173 4330
rect 11020 4211 11031 4319
rect 11031 4211 11163 4319
rect 11163 4211 11173 4319
rect 11020 4201 11173 4211
rect 20148 7628 20301 7639
rect 17666 7574 17819 7585
rect 17666 7466 17677 7574
rect 17677 7466 17809 7574
rect 17809 7466 17819 7574
rect 20148 7520 20159 7628
rect 20159 7520 20291 7628
rect 20291 7520 20301 7628
rect 21295 7628 21448 7639
rect 20148 7510 20301 7520
rect 17666 7456 17819 7466
rect 21295 7520 21306 7628
rect 21306 7520 21438 7628
rect 21438 7520 21448 7628
rect 26770 7629 26923 7640
rect 21295 7510 21448 7520
rect 24288 7575 24441 7586
rect 17947 6535 18076 6546
rect 17947 6403 17957 6535
rect 17957 6403 18065 6535
rect 18065 6403 18076 6535
rect 17947 6393 18076 6403
rect 12840 6227 12993 6237
rect 12840 6119 12850 6227
rect 12850 6119 12982 6227
rect 12982 6119 12993 6227
rect 12840 6108 12993 6119
rect 13982 6225 14135 6235
rect 13982 6117 13992 6225
rect 13992 6117 14124 6225
rect 14124 6117 14135 6225
rect 13982 6106 14135 6117
rect 17680 5924 17833 5935
rect 17680 5816 17691 5924
rect 17691 5816 17823 5924
rect 17823 5816 17833 5924
rect 17680 5806 17833 5816
rect 12838 5580 12991 5591
rect 12838 5472 12849 5580
rect 12849 5472 12981 5580
rect 12981 5472 12991 5580
rect 12838 5462 12991 5472
rect 14736 5580 14889 5591
rect 14736 5472 14747 5580
rect 14747 5472 14879 5580
rect 14879 5472 14889 5580
rect 14736 5462 14889 5472
rect 16443 4709 16587 4821
rect 17961 4885 18090 4896
rect 17961 4753 17971 4885
rect 17971 4753 18079 4885
rect 18079 4753 18090 4885
rect 17961 4743 18090 4753
rect 13479 4610 13557 4620
rect 13479 4544 13494 4610
rect 13494 4544 13557 4610
rect 13479 4534 13557 4544
rect 16713 4448 16828 4457
rect 16713 4369 16723 4448
rect 16723 4369 16816 4448
rect 16816 4369 16828 4448
rect 16713 4360 16828 4369
rect 11301 3280 11430 3291
rect 11301 3148 11311 3280
rect 11311 3148 11419 3280
rect 11419 3148 11430 3280
rect 11301 3138 11430 3148
rect 12784 3184 12937 3194
rect 12784 3076 12794 3184
rect 12794 3076 12926 3184
rect 12926 3076 12937 3184
rect 12784 3065 12937 3076
rect 14682 3184 14835 3194
rect 14682 3076 14692 3184
rect 14692 3076 14824 3184
rect 14824 3076 14835 3184
rect 14682 3065 14835 3076
rect 17675 4320 17828 4331
rect 17675 4212 17686 4320
rect 17686 4212 17818 4320
rect 17818 4212 17828 4320
rect 17675 4202 17828 4212
rect 24288 7467 24299 7575
rect 24299 7467 24431 7575
rect 24431 7467 24441 7575
rect 26770 7521 26781 7629
rect 26781 7521 26913 7629
rect 26913 7521 26923 7629
rect 27917 7629 28070 7640
rect 26770 7511 26923 7521
rect 24288 7457 24441 7467
rect 27917 7521 27928 7629
rect 27928 7521 28060 7629
rect 28060 7521 28070 7629
rect 27917 7511 28070 7521
rect 24569 6536 24698 6547
rect 24569 6404 24579 6536
rect 24579 6404 24687 6536
rect 24687 6404 24698 6536
rect 24569 6394 24698 6404
rect 19495 6228 19648 6238
rect 19495 6120 19505 6228
rect 19505 6120 19637 6228
rect 19637 6120 19648 6228
rect 19495 6109 19648 6120
rect 20637 6226 20790 6236
rect 20637 6118 20647 6226
rect 20647 6118 20779 6226
rect 20779 6118 20790 6226
rect 20637 6107 20790 6118
rect 24302 5925 24455 5936
rect 24302 5817 24313 5925
rect 24313 5817 24445 5925
rect 24445 5817 24455 5925
rect 24302 5807 24455 5817
rect 19493 5581 19646 5592
rect 19493 5473 19504 5581
rect 19504 5473 19636 5581
rect 19636 5473 19646 5581
rect 19493 5463 19646 5473
rect 21391 5581 21544 5592
rect 21391 5473 21402 5581
rect 21402 5473 21534 5581
rect 21534 5473 21544 5581
rect 21391 5463 21544 5473
rect 24583 4886 24712 4897
rect 24583 4754 24593 4886
rect 24593 4754 24701 4886
rect 24701 4754 24712 4886
rect 24583 4744 24712 4754
rect 20134 4611 20212 4621
rect 20134 4545 20149 4611
rect 20149 4545 20212 4611
rect 20134 4535 20212 4545
rect 23335 4449 23450 4458
rect 23335 4370 23345 4449
rect 23345 4370 23438 4449
rect 23438 4370 23450 4449
rect 23335 4361 23450 4370
rect 17956 3281 18085 3292
rect 17956 3149 17966 3281
rect 17966 3149 18074 3281
rect 18074 3149 18085 3281
rect 17956 3139 18085 3149
rect 19439 3185 19592 3195
rect 19439 3077 19449 3185
rect 19449 3077 19581 3185
rect 19581 3077 19592 3185
rect 19439 3066 19592 3077
rect 21337 3185 21490 3195
rect 21337 3077 21347 3185
rect 21347 3077 21479 3185
rect 21479 3077 21490 3185
rect 21337 3066 21490 3077
rect 24297 4321 24450 4332
rect 24297 4213 24308 4321
rect 24308 4213 24440 4321
rect 24440 4213 24450 4321
rect 24297 4203 24450 4213
rect 26117 6229 26270 6239
rect 26117 6121 26127 6229
rect 26127 6121 26259 6229
rect 26259 6121 26270 6229
rect 26117 6110 26270 6121
rect 27259 6227 27412 6237
rect 27259 6119 27269 6227
rect 27269 6119 27401 6227
rect 27401 6119 27412 6227
rect 27259 6108 27412 6119
rect 26115 5582 26268 5593
rect 26115 5474 26126 5582
rect 26126 5474 26258 5582
rect 26258 5474 26268 5582
rect 26115 5464 26268 5474
rect 28013 5582 28166 5593
rect 28013 5474 28024 5582
rect 28024 5474 28156 5582
rect 28156 5474 28166 5582
rect 28013 5464 28166 5474
rect 26756 4612 26834 4622
rect 26756 4546 26771 4612
rect 26771 4546 26834 4612
rect 26756 4536 26834 4546
rect 29029 4104 29161 4110
rect 29029 4023 29037 4104
rect 29037 4023 29154 4104
rect 29154 4023 29161 4104
rect 29029 4014 29161 4023
rect 32179 8818 32390 8834
rect 32179 8695 32198 8818
rect 32198 8695 32372 8818
rect 32372 8695 32390 8818
rect 32179 8677 32390 8695
rect 30226 8447 30288 8505
rect 30288 8447 30290 8505
rect 30226 8443 30290 8447
rect 30075 7729 30135 7791
rect 32257 7658 32410 7669
rect 32257 7550 32268 7658
rect 32268 7550 32400 7658
rect 32400 7550 32410 7658
rect 32257 7540 32410 7550
rect 33612 7259 33672 7321
rect 29810 6678 29896 6779
rect 31458 6673 31551 6750
rect 29582 6545 29667 6605
rect 30297 6527 30359 6585
rect 30359 6527 30361 6585
rect 30297 6523 30361 6527
rect 37737 9455 37807 9528
rect 36483 8134 36575 8146
rect 36483 8054 36511 8134
rect 36511 8054 36571 8134
rect 36571 8054 36575 8134
rect 36483 8046 36575 8054
rect 38727 8120 38785 8126
rect 38727 8054 38729 8120
rect 38729 8054 38781 8120
rect 38781 8054 38785 8120
rect 38727 8050 38785 8054
rect 33834 6057 33896 6115
rect 33896 6057 33898 6115
rect 33834 6053 33898 6057
rect 32179 5323 32390 5339
rect 32179 5200 32198 5323
rect 32198 5200 32372 5323
rect 32372 5200 32390 5323
rect 32179 5182 32390 5200
rect 30072 4659 30132 4721
rect 29412 3695 29496 3785
rect 29846 3574 29912 3638
rect 30294 3457 30356 3515
rect 30356 3457 30358 3515
rect 30294 3453 30358 3457
rect 24578 3282 24707 3293
rect 24578 3150 24588 3282
rect 24588 3150 24696 3282
rect 24696 3150 24707 3282
rect 24578 3140 24707 3150
rect 26061 3186 26214 3196
rect 26061 3078 26071 3186
rect 26071 3078 26203 3186
rect 26203 3078 26214 3186
rect 26061 3067 26214 3078
rect 27959 3186 28112 3196
rect 27959 3078 27969 3186
rect 27969 3078 28101 3186
rect 28101 3078 28112 3186
rect 27959 3067 28112 3078
rect 32257 3310 32410 3321
rect 32257 3202 32268 3310
rect 32268 3202 32400 3310
rect 32400 3202 32410 3310
rect 32257 3192 32410 3202
rect 33612 2911 33672 2973
rect 8410 2370 8474 2374
rect 8410 2312 8472 2370
rect 8472 2312 8474 2370
rect 14964 2375 15028 2379
rect 14964 2317 15026 2375
rect 15026 2317 15028 2375
rect 21613 2363 21677 2367
rect 21613 2305 21675 2363
rect 21675 2305 21677 2363
rect 36479 5002 36571 5014
rect 36479 4922 36507 5002
rect 36507 4922 36567 5002
rect 36567 4922 36571 5002
rect 36479 4914 36571 4922
rect 38723 4988 38781 4994
rect 38723 4922 38725 4988
rect 38725 4922 38777 4988
rect 38777 4922 38781 4988
rect 38723 4918 38781 4922
rect 29826 2035 29910 2125
rect 34981 1961 35068 2034
rect 8188 1106 8248 1168
rect 14742 1111 14802 1173
rect 30079 1814 30139 1876
rect 36479 1858 36571 1870
rect 36479 1778 36507 1858
rect 36507 1778 36567 1858
rect 36567 1778 36571 1858
rect 36479 1770 36571 1778
rect 33834 1709 33896 1767
rect 33896 1709 33898 1767
rect 33834 1705 33898 1709
rect 38723 1844 38781 1850
rect 38723 1778 38725 1844
rect 38725 1778 38777 1844
rect 38777 1778 38781 1844
rect 38723 1774 38781 1778
rect 29243 1292 29325 1382
rect 21391 1099 21451 1161
rect 29410 976 29494 1066
rect 32179 975 32390 991
rect 32179 852 32198 975
rect 32198 852 32372 975
rect 32372 852 32390 975
rect 32179 834 32390 852
rect 29723 642 29784 717
rect 30301 612 30363 670
rect 30363 612 30365 670
rect 30301 608 30365 612
rect -2690 119 -2604 128
rect -2690 54 -2680 119
rect -2680 54 -2616 119
rect -2616 54 -2604 119
rect -2690 43 -2604 54
<< metal3 >>
rect 6240 27769 6250 27948
rect 6449 27769 6459 27948
rect 8722 27823 8732 28002
rect 8931 27823 8941 28002
rect 9869 27823 9879 28002
rect 10078 27823 10088 28002
rect 12753 27766 12763 27945
rect 12962 27766 12972 27945
rect 15235 27820 15245 27999
rect 15444 27820 15454 27999
rect 16382 27820 16392 27999
rect 16591 27820 16601 27999
rect 19287 27761 19297 27940
rect 19496 27761 19506 27940
rect 21769 27815 21779 27994
rect 21978 27815 21988 27994
rect 22916 27815 22926 27994
rect 23125 27815 23135 27994
rect 25845 27765 25855 27944
rect 26054 27765 26064 27944
rect 28327 27819 28337 27998
rect 28536 27819 28546 27998
rect 29474 27819 29484 27998
rect 29683 27819 29693 27998
rect 6534 26900 6713 26910
rect 6534 26692 6713 26701
rect 13047 26897 13226 26907
rect 13047 26689 13226 26698
rect 19581 26892 19760 26902
rect 19581 26684 19760 26693
rect 26139 26896 26318 26906
rect 26139 26688 26318 26697
rect 8068 26410 8077 26589
rect 8276 26410 8286 26589
rect 9210 26408 9219 26587
rect 9418 26408 9428 26587
rect 14581 26407 14590 26586
rect 14789 26407 14799 26586
rect 15723 26405 15732 26584
rect 15931 26405 15941 26584
rect 21115 26402 21124 26581
rect 21323 26402 21333 26581
rect 22257 26400 22266 26579
rect 22465 26400 22475 26579
rect 27673 26406 27682 26585
rect 27881 26406 27891 26585
rect 28815 26404 28824 26583
rect 29023 26404 29033 26583
rect 11393 26315 11776 26316
rect -1659 26268 5267 26291
rect -1659 26165 5091 26268
rect 5233 26165 5267 26268
rect -1659 26148 5267 26165
rect -1847 15530 -1749 15532
rect -4069 15450 -3991 15510
rect -1849 15502 -1739 15530
rect -4069 15440 -3988 15450
rect -4069 15364 -4065 15440
rect -4069 15362 -4063 15364
rect -3993 15362 -3988 15440
rect -1849 15408 -1843 15502
rect -1755 15408 -1739 15502
rect -1849 15378 -1739 15408
rect -4069 15352 -3988 15362
rect -4069 15296 -3991 15352
rect -1659 14620 -1567 26148
rect 6254 26119 6264 26298
rect 6463 26119 6473 26298
rect 11391 26294 11776 26315
rect 17897 26300 18332 26319
rect 11391 26170 11523 26294
rect 11752 26170 11776 26294
rect 11391 26145 11776 26170
rect 11391 26072 11558 26145
rect 12767 26116 12777 26295
rect 12976 26116 12986 26295
rect 17897 26161 18082 26300
rect 17899 26160 18082 26161
rect 18300 26160 18332 26300
rect 24476 26302 24884 26322
rect 17899 26137 18332 26160
rect 8067 25776 8077 25955
rect 8276 25776 8286 25955
rect 9965 25776 9975 25955
rect 10174 25776 10184 25955
rect 6548 25250 6727 25260
rect 637 25168 5193 25171
rect 637 25163 5199 25168
rect 637 25037 5051 25163
rect 5189 25037 5199 25163
rect 6548 25042 6727 25051
rect 637 25032 5199 25037
rect 637 25028 5193 25032
rect -855 23408 -651 23410
rect 637 23408 741 25028
rect 5330 24957 5422 24958
rect 8728 24957 8832 24959
rect 5330 24953 8832 24957
rect 5330 24867 8740 24953
rect 8818 24867 8832 24953
rect 5330 24854 8832 24867
rect 5330 24794 5422 24854
rect 5309 24789 5444 24794
rect 5309 24692 5319 24789
rect 5434 24692 5444 24789
rect 5309 24687 5444 24692
rect 6249 24515 6259 24694
rect 6458 24515 6468 24694
rect 6543 23646 6722 23656
rect 6543 23438 6722 23447
rect -855 23405 741 23408
rect -855 23244 -845 23405
rect -661 23244 741 23405
rect 8011 23367 8021 23546
rect 8220 23367 8230 23546
rect 9909 23367 9919 23546
rect 10118 23367 10128 23546
rect -855 23240 741 23244
rect -855 23239 -651 23240
rect 11391 23085 11557 26072
rect 14580 25773 14590 25952
rect 14789 25773 14799 25952
rect 16478 25773 16488 25952
rect 16687 25773 16697 25952
rect 13061 25247 13240 25257
rect 13061 25039 13240 25048
rect 11843 24954 11935 24955
rect 15241 24954 15345 24956
rect 11843 24950 15345 24954
rect 11843 24864 15253 24950
rect 15331 24864 15345 24950
rect 11843 24851 15345 24864
rect 11843 24791 11935 24851
rect 11822 24786 11957 24791
rect 11822 24689 11832 24786
rect 11947 24689 11957 24786
rect 11822 24684 11957 24689
rect 12762 24512 12772 24691
rect 12971 24512 12981 24691
rect 13056 23643 13235 23653
rect 13056 23435 13235 23444
rect 14524 23364 14534 23543
rect 14733 23364 14743 23543
rect 16422 23364 16432 23543
rect 16631 23364 16641 23543
rect -2704 14613 -1567 14620
rect -2704 14516 -2694 14613
rect -2598 14516 -1567 14613
rect -2704 14501 -1567 14516
rect -1659 14500 -1567 14501
rect -1495 22976 11557 23085
rect -1849 13462 -1751 13464
rect -4071 13382 -3993 13442
rect -1851 13434 -1741 13462
rect -4071 13372 -3990 13382
rect -4071 13296 -4067 13372
rect -4071 13294 -4065 13296
rect -3995 13294 -3990 13372
rect -1851 13340 -1845 13434
rect -1757 13340 -1741 13434
rect -1851 13310 -1741 13340
rect -4071 13284 -3990 13294
rect -4071 13228 -3993 13284
rect -1495 12548 -1415 22976
rect 17899 22906 18060 26137
rect 19301 26111 19311 26290
rect 19510 26111 19520 26290
rect 24476 26157 24606 26302
rect 24858 26157 24884 26302
rect 24476 26144 24884 26157
rect 21114 25768 21124 25947
rect 21323 25768 21333 25947
rect 23012 25768 23022 25947
rect 23221 25768 23231 25947
rect 19595 25242 19774 25252
rect 19595 25034 19774 25043
rect 18377 24949 18469 24950
rect 21775 24949 21879 24951
rect 18377 24945 21879 24949
rect 18377 24859 21787 24945
rect 21865 24859 21879 24945
rect 18377 24846 21879 24859
rect 18377 24786 18469 24846
rect 18356 24781 18491 24786
rect 18356 24684 18366 24781
rect 18481 24684 18491 24781
rect 18356 24679 18491 24684
rect 19296 24507 19306 24686
rect 19505 24507 19515 24686
rect 19590 23638 19769 23648
rect 19590 23430 19769 23439
rect 21058 23359 21068 23538
rect 21267 23359 21277 23538
rect 22956 23359 22966 23538
rect 23165 23359 23175 23538
rect -2702 12543 -1415 12548
rect -2702 12451 -2692 12543
rect -2600 12451 -1415 12543
rect -2702 12446 -1415 12451
rect -1351 22792 18060 22906
rect -1351 22791 -1272 22792
rect -1847 11393 -1749 11395
rect -4069 11313 -3991 11373
rect -1849 11365 -1739 11393
rect -4069 11303 -3988 11313
rect -4069 11227 -4065 11303
rect -4069 11225 -4063 11227
rect -3993 11225 -3988 11303
rect -1849 11271 -1843 11365
rect -1755 11271 -1739 11365
rect -1849 11241 -1739 11271
rect -4069 11215 -3988 11225
rect -4069 11159 -3991 11215
rect -1351 10479 -1275 22791
rect 24476 22732 24646 26144
rect 25859 26115 25869 26294
rect 26068 26115 26078 26294
rect 27672 25772 27682 25951
rect 27881 25772 27891 25951
rect 29570 25772 29580 25951
rect 29779 25772 29789 25951
rect 26153 25246 26332 25256
rect 26153 25038 26332 25047
rect 24935 24953 25027 24954
rect 28333 24953 28437 24955
rect 24935 24949 28437 24953
rect 24935 24863 28345 24949
rect 28423 24863 28437 24949
rect 24935 24850 28437 24863
rect 24935 24790 25027 24850
rect 24914 24785 25049 24790
rect 24914 24688 24924 24785
rect 25039 24688 25049 24785
rect 24914 24683 25049 24688
rect 25854 24511 25864 24690
rect 26063 24511 26073 24690
rect 36478 23912 36580 23922
rect 36478 23812 36483 23912
rect 36577 23812 36580 23912
rect 36478 23802 36580 23812
rect 38719 23898 38799 23932
rect 38719 23814 38727 23898
rect 38795 23814 38799 23898
rect 38719 23766 38799 23814
rect 26148 23642 26327 23652
rect 26148 23434 26327 23443
rect 27616 23363 27626 23542
rect 27825 23363 27835 23542
rect 29514 23363 29524 23542
rect 29723 23363 29733 23542
rect -2696 10471 -1275 10479
rect -2696 10385 -2686 10471
rect -2601 10385 -1275 10471
rect -2696 10367 -1275 10385
rect -1351 10364 -1275 10367
rect -1215 22622 24647 22732
rect -1849 9325 -1751 9327
rect -4071 9245 -3993 9305
rect -1851 9297 -1741 9325
rect -4071 9235 -3990 9245
rect -4071 9159 -4067 9235
rect -4071 9157 -4065 9159
rect -3995 9157 -3990 9235
rect -1851 9203 -1845 9297
rect -1757 9203 -1741 9297
rect -1851 9173 -1741 9203
rect -4071 9147 -3990 9157
rect -4071 9091 -3993 9147
rect -1215 8414 -1136 22622
rect 160 22621 372 22622
rect 5816 22215 5826 22394
rect 6025 22215 6035 22394
rect 6963 22215 6973 22394
rect 7172 22215 7182 22394
rect 9445 22161 9455 22340
rect 9654 22161 9664 22340
rect 12374 22211 12384 22390
rect 12583 22211 12593 22390
rect 13521 22211 13531 22390
rect 13730 22211 13740 22390
rect 16003 22157 16013 22336
rect 16212 22157 16222 22336
rect 18908 22216 18918 22395
rect 19117 22216 19127 22395
rect 20055 22216 20065 22395
rect 20264 22216 20274 22395
rect 22537 22162 22547 22341
rect 22746 22162 22756 22341
rect 25421 22219 25431 22398
rect 25630 22219 25640 22398
rect 26568 22219 26578 22398
rect 26777 22219 26787 22398
rect 29050 22165 29060 22344
rect 29259 22165 29269 22344
rect 9191 21292 9370 21302
rect 9191 21084 9370 21093
rect 15749 21288 15928 21298
rect 15749 21080 15928 21089
rect 22283 21293 22462 21303
rect 22283 21085 22462 21094
rect 28796 21296 28975 21306
rect 28796 21088 28975 21097
rect 6476 20800 6486 20979
rect 6685 20800 6694 20979
rect 7618 20802 7628 20981
rect 7827 20802 7836 20981
rect 13034 20796 13044 20975
rect 13243 20796 13252 20975
rect 14176 20798 14186 20977
rect 14385 20798 14394 20977
rect 19568 20801 19578 20980
rect 19777 20801 19786 20980
rect 20710 20803 20720 20982
rect 20919 20803 20928 20982
rect 26081 20804 26091 20983
rect 26290 20804 26299 20983
rect 27223 20806 27233 20985
rect 27432 20806 27441 20985
rect 36478 20768 36580 20778
rect 30247 20724 30649 20746
rect 9431 20511 9441 20690
rect 9640 20511 9650 20690
rect 15989 20507 15999 20686
rect 16198 20507 16208 20686
rect 22523 20512 22533 20691
rect 22732 20512 22742 20691
rect 29036 20515 29046 20694
rect 29245 20515 29255 20694
rect 30247 20568 30262 20724
rect 30480 20568 30649 20724
rect 36478 20668 36483 20768
rect 36577 20668 36580 20768
rect 36478 20658 36580 20668
rect 38719 20754 38799 20788
rect 38719 20670 38727 20754
rect 38795 20670 38799 20754
rect 38719 20622 38799 20670
rect 30247 20543 30649 20568
rect 5720 20168 5730 20347
rect 5929 20168 5939 20347
rect 7618 20168 7628 20347
rect 7827 20168 7837 20347
rect 12278 20164 12288 20343
rect 12487 20164 12497 20343
rect 14176 20164 14186 20343
rect 14385 20164 14395 20343
rect 18812 20169 18822 20348
rect 19021 20169 19031 20348
rect 20710 20169 20720 20348
rect 20919 20169 20929 20348
rect 25325 20172 25335 20351
rect 25534 20172 25544 20351
rect 27223 20172 27233 20351
rect 27432 20172 27442 20351
rect 9177 19642 9356 19652
rect 9177 19434 9356 19443
rect 15735 19638 15914 19648
rect 15735 19430 15914 19439
rect 22269 19643 22448 19653
rect 22269 19435 22448 19444
rect 28782 19646 28961 19656
rect 28782 19438 28961 19447
rect 26677 19353 26781 19355
rect 30087 19353 30179 19354
rect 7072 19349 7176 19351
rect 20164 19350 20268 19352
rect 23574 19350 23666 19351
rect 10482 19349 10574 19350
rect 7072 19345 10574 19349
rect 7072 19259 7086 19345
rect 7164 19259 10574 19345
rect 7072 19246 10574 19259
rect 10482 19186 10574 19246
rect 13630 19345 13734 19347
rect 20164 19346 23666 19350
rect 17040 19345 17132 19346
rect 13630 19341 17132 19345
rect 13630 19255 13644 19341
rect 13722 19255 17132 19341
rect 13630 19242 17132 19255
rect 20164 19260 20178 19346
rect 20256 19260 23666 19346
rect 20164 19247 23666 19260
rect 26677 19349 30179 19353
rect 26677 19263 26691 19349
rect 26769 19263 30179 19349
rect 26677 19250 30179 19263
rect 10460 19181 10595 19186
rect 17040 19182 17132 19242
rect 23574 19187 23666 19247
rect 30087 19190 30179 19250
rect 23552 19182 23687 19187
rect 9436 18907 9446 19086
rect 9645 18907 9655 19086
rect 10460 19084 10470 19181
rect 10585 19084 10595 19181
rect 10460 19079 10595 19084
rect 17018 19177 17153 19182
rect 15994 18903 16004 19082
rect 16203 18903 16213 19082
rect 17018 19080 17028 19177
rect 17143 19080 17153 19177
rect 17018 19075 17153 19080
rect 22528 18908 22538 19087
rect 22737 18908 22747 19087
rect 23552 19085 23562 19182
rect 23677 19085 23687 19182
rect 30065 19185 30200 19190
rect 23552 19080 23687 19085
rect 29041 18911 29051 19090
rect 29250 18911 29260 19090
rect 30065 19088 30075 19185
rect 30190 19088 30200 19185
rect 30065 19083 30200 19088
rect 9182 18038 9361 18048
rect 5776 17759 5786 17938
rect 5985 17759 5995 17938
rect 7674 17759 7684 17938
rect 7883 17759 7893 17938
rect 15740 18034 15919 18044
rect 9182 17830 9361 17839
rect 12334 17755 12344 17934
rect 12543 17755 12553 17934
rect 14232 17755 14242 17934
rect 14441 17755 14451 17934
rect 22274 18039 22453 18049
rect 15740 17826 15919 17835
rect 18868 17760 18878 17939
rect 19077 17760 19087 17939
rect 20766 17760 20776 17939
rect 20975 17760 20985 17939
rect 28787 18042 28966 18052
rect 22274 17831 22453 17840
rect 25381 17763 25391 17942
rect 25590 17763 25600 17942
rect 27279 17763 27289 17942
rect 27488 17763 27498 17942
rect 28787 17834 28966 17843
rect -1020 16602 -888 16603
rect 30468 16602 30649 20543
rect 36474 17636 36576 17646
rect 36474 17536 36479 17636
rect 36573 17536 36576 17636
rect 36474 17526 36576 17536
rect 38715 17622 38795 17656
rect 38715 17538 38723 17622
rect 38791 17538 38795 17622
rect 38715 17490 38795 17538
rect -2702 8401 -1136 8414
rect -2702 8316 -2691 8401
rect -2602 8316 -1136 8401
rect -2702 8305 -1136 8316
rect -1075 16485 30649 16602
rect -1849 7256 -1751 7258
rect -4071 7176 -3993 7236
rect -1851 7228 -1741 7256
rect -4071 7166 -3990 7176
rect -4071 7090 -4067 7166
rect -4071 7088 -4065 7090
rect -3995 7088 -3990 7166
rect -1851 7134 -1845 7228
rect -1757 7134 -1741 7228
rect -1851 7104 -1741 7134
rect -4071 7078 -3990 7088
rect -4071 7022 -3993 7078
rect -1075 6342 -996 16485
rect 23956 16423 24075 16425
rect -2702 6332 -996 6342
rect -2702 6249 -2688 6332
rect -2604 6249 -996 6332
rect -2702 6239 -996 6249
rect -931 16331 24075 16423
rect -1112 6238 -1034 6239
rect -1851 5188 -1753 5190
rect -4073 5108 -3995 5168
rect -1853 5160 -1743 5188
rect -4073 5098 -3992 5108
rect -4073 5022 -4069 5098
rect -4073 5020 -4067 5022
rect -3997 5020 -3992 5098
rect -1853 5066 -1847 5160
rect -1759 5066 -1743 5160
rect -1853 5036 -1743 5066
rect -4073 5010 -3992 5020
rect -4073 4954 -3995 5010
rect -931 4275 -858 16331
rect 17431 16268 17551 16269
rect -2699 4265 -858 4275
rect -2699 4181 -2689 4265
rect -2606 4181 -858 4265
rect -2699 4171 -858 4181
rect -798 16168 17552 16268
rect 23956 16267 24075 16331
rect -1849 3119 -1751 3121
rect -4071 3039 -3993 3099
rect -1851 3091 -1741 3119
rect -4071 3029 -3990 3039
rect -4071 2953 -4067 3029
rect -4071 2951 -4065 2953
rect -3995 2951 -3990 3029
rect -1851 2997 -1845 3091
rect -1757 2997 -1741 3091
rect -1851 2967 -1741 2997
rect -4071 2941 -3990 2951
rect -4071 2885 -3993 2941
rect -798 2205 -723 16168
rect 17431 16137 17551 16168
rect 23956 16165 23966 16267
rect 24065 16165 24075 16267
rect 23956 16156 24075 16165
rect -662 16005 10986 16106
rect 17431 16052 17441 16137
rect 17541 16052 17551 16137
rect 17431 16041 17551 16052
rect -662 15931 -586 16005
rect -2701 2196 -723 2205
rect -2701 2109 -2691 2196
rect -2601 2109 -723 2196
rect -2701 2098 -723 2109
rect -1851 1051 -1753 1053
rect -4073 971 -3995 1031
rect -1853 1023 -1743 1051
rect -4073 961 -3992 971
rect -4073 885 -4069 961
rect -4073 883 -4067 885
rect -3997 883 -3992 961
rect -1853 929 -1847 1023
rect -1759 929 -1743 1023
rect -1853 899 -1743 929
rect -4073 873 -3992 883
rect -4073 817 -3995 873
rect -661 144 -586 15931
rect 10854 15806 10986 16005
rect 34960 15982 37808 15985
rect 34959 15886 37808 15982
rect 10851 15801 10989 15806
rect 10851 15733 10861 15801
rect 10979 15733 10989 15801
rect 10851 15728 10989 15733
rect 10854 15723 10986 15728
rect 21340 15486 21438 15504
rect 8137 15466 8235 15484
rect 8137 15394 8147 15466
rect 8217 15394 8235 15466
rect 8137 15386 8235 15394
rect 14686 15465 14784 15483
rect 14686 15393 14696 15465
rect 14766 15393 14784 15465
rect 21340 15414 21350 15486
rect 21420 15414 21438 15486
rect 21340 15406 21438 15414
rect 14686 15385 14784 15393
rect 29993 15319 30091 15337
rect 29993 15247 30003 15319
rect 30073 15247 30091 15319
rect 29993 15239 30091 15247
rect 32223 15107 32233 15286
rect 32432 15107 32442 15286
rect 34959 15106 35086 15886
rect 37676 15885 37808 15886
rect 37725 15880 37808 15885
rect 37725 15875 37809 15880
rect 37725 15778 37736 15875
rect 37799 15778 37809 15875
rect 37725 15773 37809 15778
rect 37725 15769 37808 15773
rect 34959 15005 35087 15106
rect 33594 14911 33692 14929
rect 33594 14839 33604 14911
rect 33674 14839 33692 14911
rect 33594 14831 33692 14839
rect 21558 14282 21660 14298
rect 8355 14262 8457 14278
rect 8355 14194 8369 14262
rect 8443 14194 8457 14262
rect 8355 14180 8457 14194
rect 14904 14261 15006 14277
rect 14904 14193 14918 14261
rect 14992 14193 15006 14261
rect 21558 14214 21572 14282
rect 21646 14214 21660 14282
rect 21558 14200 21660 14214
rect 34209 14237 34568 14238
rect 34209 14229 34664 14237
rect 14904 14179 15006 14193
rect 34209 14147 34219 14229
rect 34357 14147 34664 14229
rect 34209 14138 34664 14147
rect 30211 14115 30313 14131
rect 30211 14047 30225 14115
rect 30299 14047 30313 14115
rect 339 14038 475 14043
rect 339 13982 349 14038
rect 465 13982 475 14038
rect 30211 14033 30313 14047
rect 339 13977 475 13982
rect 346 4127 469 13977
rect 34490 13808 34664 14138
rect 33689 13617 33699 13733
rect 34037 13617 34047 13733
rect 1473 13566 1571 13584
rect 1473 13494 1483 13566
rect 1553 13494 1571 13566
rect 1473 13486 1571 13494
rect 4436 13218 4446 13397
rect 4645 13218 4655 13397
rect 6918 13272 6928 13451
rect 7127 13272 7137 13451
rect 8065 13272 8075 13451
rect 8274 13272 8284 13451
rect 10985 13306 10995 13485
rect 11194 13306 11204 13485
rect 13467 13360 13477 13539
rect 13676 13360 13686 13539
rect 14614 13360 14624 13539
rect 14823 13360 14833 13539
rect 17639 13238 17649 13417
rect 17848 13238 17858 13417
rect 20121 13292 20131 13471
rect 20330 13292 20340 13471
rect 21268 13292 21278 13471
rect 21477 13292 21487 13471
rect 24264 13306 24274 13485
rect 24473 13306 24483 13485
rect 26746 13360 26756 13539
rect 26955 13360 26965 13539
rect 27893 13360 27903 13539
rect 28102 13360 28112 13539
rect 29988 12748 30086 12766
rect 29988 12676 29998 12748
rect 30068 12676 30086 12748
rect 32144 12746 32154 12941
rect 32420 12746 32430 12941
rect 29988 12668 30086 12676
rect 22519 12601 22776 12602
rect 22311 12596 22776 12601
rect 9177 12578 9342 12581
rect 9177 12576 9541 12578
rect 9177 12501 9187 12576
rect 9332 12501 9541 12576
rect 22311 12522 22321 12596
rect 22418 12522 22776 12596
rect 22311 12517 22776 12522
rect 9177 12496 9541 12501
rect 1691 12362 1793 12378
rect 1691 12294 1705 12362
rect 1779 12294 1793 12362
rect 1691 12280 1793 12294
rect 4730 12349 4909 12359
rect 4730 12141 4909 12150
rect 6264 11859 6273 12038
rect 6472 11859 6482 12038
rect 7406 11857 7415 12036
rect 7614 11857 7624 12036
rect 4450 11568 4460 11747
rect 4659 11568 4669 11747
rect 6263 11225 6273 11404
rect 6472 11225 6482 11404
rect 8161 11225 8171 11404
rect 8370 11225 8380 11404
rect 1465 10981 1563 10999
rect 1465 10909 1475 10981
rect 1545 10909 1563 10981
rect 1465 10901 1563 10909
rect 4744 10699 4923 10709
rect 4744 10491 4923 10500
rect 3526 10406 3618 10407
rect 6924 10406 7028 10408
rect 3526 10402 7028 10406
rect 3526 10316 6936 10402
rect 7014 10316 7028 10402
rect 3526 10303 7028 10316
rect 3526 10243 3618 10303
rect 3505 10238 3640 10243
rect 3505 10141 3515 10238
rect 3630 10141 3640 10238
rect 3505 10136 3640 10141
rect 4445 9964 4455 10143
rect 4654 9964 4664 10143
rect 1683 9777 1785 9793
rect 1683 9709 1697 9777
rect 1771 9709 1785 9777
rect 1683 9695 1785 9709
rect 4739 9095 4918 9105
rect 4739 8887 4918 8896
rect 6207 8816 6217 8995
rect 6416 8816 6426 8995
rect 8105 8816 8115 8995
rect 8314 8816 8324 8995
rect 2763 8093 2964 8094
rect 9397 8093 9541 12496
rect 11279 12437 11458 12447
rect 11279 12229 11458 12238
rect 17933 12369 18112 12379
rect 17933 12161 18112 12170
rect 12813 11947 12822 12126
rect 13021 11947 13031 12126
rect 13955 11945 13964 12124
rect 14163 11945 14173 12124
rect 19467 11879 19476 12058
rect 19675 11879 19685 12058
rect 20609 11877 20618 12056
rect 20817 11877 20827 12056
rect 10999 11656 11009 11835
rect 11208 11656 11218 11835
rect 17653 11588 17663 11767
rect 17862 11588 17872 11767
rect 12812 11313 12822 11492
rect 13021 11313 13031 11492
rect 14710 11313 14720 11492
rect 14919 11313 14929 11492
rect 19466 11245 19476 11424
rect 19675 11245 19685 11424
rect 21364 11245 21374 11424
rect 21573 11245 21583 11424
rect 11293 10787 11472 10797
rect 11293 10579 11472 10588
rect 17947 10719 18126 10729
rect 17947 10511 18126 10520
rect 10075 10494 10167 10495
rect 13473 10494 13577 10496
rect 10075 10490 13577 10494
rect 10075 10404 13485 10490
rect 13563 10404 13577 10490
rect 10075 10391 13577 10404
rect 16729 10426 16821 10427
rect 20127 10426 20231 10428
rect 16729 10422 20231 10426
rect 10075 10331 10167 10391
rect 16729 10336 20139 10422
rect 20217 10336 20231 10422
rect 10054 10326 10189 10331
rect 10054 10229 10064 10326
rect 10179 10229 10189 10326
rect 16729 10323 20231 10336
rect 16729 10263 16821 10323
rect 16708 10258 16843 10263
rect 10054 10224 10189 10229
rect 10994 10052 11004 10231
rect 11203 10052 11213 10231
rect 16708 10161 16718 10258
rect 16833 10161 16843 10258
rect 16708 10156 16843 10161
rect 17648 9984 17658 10163
rect 17857 9984 17867 10163
rect 11288 9183 11467 9193
rect 17942 9115 18121 9125
rect 11288 8975 11467 8984
rect 12756 8904 12766 9083
rect 12965 8904 12975 9083
rect 14654 8904 14664 9083
rect 14863 8904 14873 9083
rect 17942 8907 18121 8916
rect 19410 8836 19420 9015
rect 19619 8836 19629 9015
rect 21308 8836 21318 9015
rect 21517 8836 21527 9015
rect 22383 8607 22550 8617
rect 22383 8473 22394 8607
rect 22536 8473 22550 8607
rect 22383 8347 22550 8473
rect 10650 8346 22550 8347
rect 2763 7921 9541 8093
rect 9762 8175 22550 8346
rect 9762 8174 21661 8175
rect 1446 7703 1544 7721
rect 1446 7631 1456 7703
rect 1526 7631 1544 7703
rect 1446 7623 1544 7631
rect 1664 6499 1766 6515
rect 1664 6431 1678 6499
rect 1752 6431 1766 6499
rect 1664 6417 1766 6431
rect 1462 4943 1560 4961
rect 1462 4871 1472 4943
rect 1542 4871 1560 4943
rect 1462 4863 1560 4871
rect 2763 4848 2964 7921
rect 4428 7438 4438 7617
rect 4637 7438 4647 7617
rect 6910 7492 6920 7671
rect 7119 7492 7129 7671
rect 8057 7492 8067 7671
rect 8266 7492 8276 7671
rect 4722 6569 4901 6579
rect 4722 6361 4901 6370
rect 6256 6079 6265 6258
rect 6464 6079 6474 6258
rect 7398 6077 7407 6256
rect 7606 6077 7616 6256
rect 4442 5788 4452 5967
rect 4651 5788 4661 5967
rect 6255 5445 6265 5624
rect 6464 5445 6474 5624
rect 8153 5445 8163 5624
rect 8362 5445 8372 5624
rect 9762 5015 9948 8174
rect 22627 8093 22776 12517
rect 24558 12437 24737 12447
rect 24558 12229 24737 12238
rect 26092 11947 26101 12126
rect 26300 11947 26310 12126
rect 27234 11945 27243 12124
rect 27442 11945 27452 12124
rect 24278 11656 24288 11835
rect 24487 11656 24497 11835
rect 30206 11544 30308 11560
rect 26091 11313 26101 11492
rect 26300 11313 26310 11492
rect 27989 11313 27999 11492
rect 28198 11313 28208 11492
rect 30206 11476 30220 11544
rect 30294 11476 30308 11544
rect 30206 11462 30308 11476
rect 32225 11016 32235 11195
rect 32434 11016 32444 11195
rect 33596 10820 33694 10838
rect 24572 10787 24751 10797
rect 33596 10748 33606 10820
rect 33676 10748 33694 10820
rect 33596 10740 33694 10748
rect 24572 10579 24751 10588
rect 23354 10494 23446 10495
rect 26752 10494 26856 10496
rect 23354 10490 26856 10494
rect 23354 10404 26764 10490
rect 26842 10404 26856 10490
rect 23354 10391 26856 10404
rect 23354 10331 23446 10391
rect 23333 10326 23468 10331
rect 23333 10229 23343 10326
rect 23458 10229 23468 10326
rect 23333 10224 23468 10229
rect 24273 10052 24283 10231
rect 24482 10052 24492 10231
rect 22864 9911 23206 9916
rect 22864 9811 22874 9911
rect 22970 9811 23206 9911
rect 22864 9806 23206 9811
rect 22865 9803 23206 9806
rect 16167 7906 22776 8093
rect 23056 8097 23206 9803
rect 29988 9715 30086 9733
rect 29988 9643 29998 9715
rect 30068 9643 30086 9715
rect 29988 9635 30086 9643
rect 33691 9526 33701 9642
rect 34039 9526 34049 9642
rect 24567 9183 24746 9193
rect 24567 8975 24746 8984
rect 26035 8904 26045 9083
rect 26244 8904 26254 9083
rect 27933 8904 27943 9083
rect 28142 8904 28152 9083
rect 32146 8655 32156 8850
rect 32422 8655 32432 8850
rect 23492 8607 23659 8617
rect 23492 8473 23503 8607
rect 23645 8473 23659 8607
rect 23492 8345 23659 8473
rect 30206 8511 30308 8527
rect 30206 8443 30220 8511
rect 30294 8443 30308 8511
rect 30206 8429 30308 8443
rect 34490 8345 34663 13808
rect 23492 8259 34663 8345
rect 23493 8175 34663 8259
rect 34490 8172 34663 8175
rect 31205 8097 31324 8099
rect 10979 7436 10989 7615
rect 11188 7436 11198 7615
rect 13461 7490 13471 7669
rect 13670 7490 13680 7669
rect 14608 7490 14618 7669
rect 14817 7490 14827 7669
rect 11273 6567 11452 6577
rect 11273 6359 11452 6368
rect 12807 6077 12816 6256
rect 13015 6077 13025 6256
rect 13949 6075 13958 6254
rect 14157 6075 14167 6254
rect 10993 5786 11003 5965
rect 11202 5786 11212 5965
rect 12806 5443 12816 5622
rect 13015 5443 13025 5622
rect 14704 5443 14714 5622
rect 14913 5443 14923 5622
rect 4736 4919 4915 4929
rect 2762 4843 3374 4848
rect 2762 4706 3127 4843
rect 3361 4706 3374 4843
rect 9761 4890 9949 5015
rect 11287 4917 11466 4927
rect 9751 4836 9995 4890
rect 9751 4795 9762 4836
rect 4736 4711 4915 4720
rect 2762 4702 3374 4706
rect 3117 4701 3371 4702
rect 9752 4700 9762 4795
rect 9985 4700 9995 4836
rect 16167 4852 16368 7906
rect 23056 7902 31324 8097
rect 30059 7795 30157 7813
rect 30059 7723 30069 7795
rect 30139 7723 30157 7795
rect 30059 7715 30157 7723
rect 17634 7437 17644 7616
rect 17843 7437 17853 7616
rect 20116 7491 20126 7670
rect 20325 7491 20335 7670
rect 21263 7491 21273 7670
rect 21472 7491 21482 7670
rect 24256 7438 24266 7617
rect 24465 7438 24475 7617
rect 26738 7492 26748 7671
rect 26947 7492 26957 7671
rect 27885 7492 27895 7671
rect 28094 7492 28104 7671
rect 29238 6782 29906 6784
rect 29237 6779 29906 6782
rect 29237 6678 29810 6779
rect 29896 6678 29906 6779
rect 29237 6673 29906 6678
rect 31205 6755 31324 7902
rect 32225 7521 32235 7700
rect 32434 7521 32444 7700
rect 33596 7325 33694 7343
rect 33596 7253 33606 7325
rect 33676 7253 33694 7325
rect 33596 7245 33694 7253
rect 31205 6750 31561 6755
rect 31205 6673 31458 6750
rect 31551 6673 31561 6750
rect 17928 6568 18107 6578
rect 17928 6360 18107 6369
rect 24550 6569 24729 6579
rect 24550 6361 24729 6370
rect 19462 6078 19471 6257
rect 19670 6078 19680 6257
rect 20604 6076 20613 6255
rect 20812 6076 20822 6255
rect 26084 6079 26093 6258
rect 26292 6079 26302 6258
rect 27226 6077 27235 6256
rect 27434 6077 27444 6256
rect 17648 5787 17658 5966
rect 17857 5787 17867 5966
rect 24270 5788 24280 5967
rect 24479 5788 24489 5967
rect 19461 5444 19471 5623
rect 19670 5444 19680 5623
rect 21359 5444 21369 5623
rect 21568 5444 21578 5623
rect 26083 5445 26093 5624
rect 26292 5445 26302 5624
rect 27981 5445 27991 5624
rect 28190 5445 28200 5624
rect 17942 4918 18121 4928
rect 16167 4821 16615 4852
rect 16167 4799 16443 4821
rect 11287 4709 11466 4718
rect 16168 4709 16443 4799
rect 16587 4709 16615 4821
rect 17942 4710 18121 4719
rect 24564 4919 24743 4929
rect 24564 4711 24743 4720
rect 9752 4695 9995 4700
rect 16168 4691 16615 4709
rect 3518 4626 3610 4627
rect 6916 4626 7020 4628
rect 3518 4622 7020 4626
rect 3518 4536 6928 4622
rect 7006 4536 7020 4622
rect 3518 4523 7020 4536
rect 10069 4624 10161 4625
rect 13467 4624 13571 4626
rect 10069 4620 13571 4624
rect 10069 4534 13479 4620
rect 13557 4534 13571 4620
rect 3518 4463 3610 4523
rect 10069 4521 13571 4534
rect 16724 4625 16816 4626
rect 20122 4625 20226 4627
rect 16724 4621 20226 4625
rect 16724 4535 20134 4621
rect 20212 4535 20226 4621
rect 16724 4522 20226 4535
rect 23346 4626 23438 4627
rect 26744 4626 26848 4628
rect 23346 4622 26848 4626
rect 23346 4536 26756 4622
rect 26834 4536 26848 4622
rect 23346 4523 26848 4536
rect 3497 4458 3632 4463
rect 10069 4461 10161 4521
rect 16724 4462 16816 4522
rect 23346 4463 23438 4523
rect 3497 4361 3507 4458
rect 3622 4361 3632 4458
rect 10048 4456 10183 4461
rect 3497 4356 3632 4361
rect 4437 4184 4447 4363
rect 4646 4184 4656 4363
rect 10048 4359 10058 4456
rect 10173 4359 10183 4456
rect 16703 4457 16838 4462
rect 10048 4354 10183 4359
rect 10988 4182 10998 4361
rect 11197 4182 11207 4361
rect 16703 4360 16713 4457
rect 16828 4360 16838 4457
rect 23325 4458 23460 4463
rect 16703 4355 16838 4360
rect 17643 4183 17653 4362
rect 17852 4183 17862 4362
rect 23325 4361 23335 4458
rect 23450 4361 23460 4458
rect 23325 4356 23460 4361
rect 24265 4184 24275 4363
rect 24474 4184 24484 4363
rect 346 4048 356 4127
rect 459 4048 469 4127
rect 346 4043 469 4048
rect 29016 4110 29176 4116
rect 29016 4014 29029 4110
rect 29161 4014 29176 4110
rect 1680 3739 1782 3755
rect 1680 3671 1694 3739
rect 1768 3671 1782 3739
rect 1680 3657 1782 3671
rect 4731 3315 4910 3325
rect 11282 3313 11461 3323
rect 4731 3107 4910 3116
rect 6199 3036 6209 3215
rect 6408 3036 6418 3215
rect 8097 3036 8107 3215
rect 8306 3036 8316 3215
rect 17937 3314 18116 3324
rect 11282 3105 11461 3114
rect 12750 3034 12760 3213
rect 12959 3034 12969 3213
rect 14648 3034 14658 3213
rect 14857 3034 14867 3213
rect 24559 3315 24738 3325
rect 17937 3106 18116 3115
rect 19405 3035 19415 3214
rect 19614 3035 19624 3214
rect 21303 3035 21313 3214
rect 21512 3035 21522 3214
rect 24559 3107 24738 3116
rect 26027 3036 26037 3215
rect 26236 3036 26246 3215
rect 27925 3036 27935 3215
rect 28134 3036 28144 3215
rect 8390 2374 8492 2388
rect 8390 2306 8404 2374
rect 8478 2306 8492 2374
rect 8390 2290 8492 2306
rect 14944 2379 15046 2393
rect 14944 2311 14958 2379
rect 15032 2311 15046 2379
rect 14944 2295 15046 2311
rect 21593 2367 21695 2381
rect 21593 2299 21607 2367
rect 21681 2299 21695 2367
rect 21593 2283 21695 2299
rect 8172 1174 8270 1182
rect 8172 1102 8182 1174
rect 8252 1102 8270 1174
rect 8172 1084 8270 1102
rect 14726 1179 14824 1187
rect 14726 1107 14736 1179
rect 14806 1107 14824 1179
rect 14726 1089 14824 1107
rect 21375 1167 21473 1175
rect 21375 1095 21385 1167
rect 21455 1095 21473 1167
rect 21375 1077 21473 1095
rect 29016 508 29176 4014
rect 29237 4006 29337 6673
rect 31205 6668 31561 6673
rect 31205 6666 31524 6668
rect 29572 6605 29677 6610
rect 29572 6545 29582 6605
rect 29667 6545 29677 6605
rect 29572 6508 29677 6545
rect 30277 6591 30379 6607
rect 30277 6523 30291 6591
rect 30365 6523 30379 6591
rect 30277 6509 30379 6523
rect 29237 1382 29338 4006
rect 29406 3790 29508 3799
rect 29402 3785 29508 3790
rect 29402 3695 29412 3785
rect 29496 3695 29508 3785
rect 29402 3690 29508 3695
rect 29237 1292 29243 1382
rect 29325 1292 29338 1382
rect 29237 1282 29338 1292
rect 29406 3688 29508 3690
rect 29406 1071 29506 3688
rect 29400 1066 29506 1071
rect 29400 976 29410 1066
rect 29494 976 29506 1066
rect 29400 971 29506 976
rect 29406 969 29506 971
rect 29583 722 29660 6508
rect 33691 6031 33701 6147
rect 34039 6031 34049 6147
rect 32146 5160 32156 5355
rect 32422 5160 32432 5355
rect 30056 4725 30154 4743
rect 30056 4653 30066 4725
rect 30136 4653 30154 4725
rect 30056 4645 30154 4653
rect 29836 3638 29922 3643
rect 29836 3574 29846 3638
rect 29912 3574 29922 3638
rect 29836 2140 29922 3574
rect 30274 3521 30376 3537
rect 30274 3453 30288 3521
rect 30362 3453 30376 3521
rect 30274 3439 30376 3453
rect 32225 3173 32235 3352
rect 32434 3173 32444 3352
rect 33596 2977 33694 2995
rect 33596 2905 33606 2977
rect 33676 2905 33694 2977
rect 33596 2897 33694 2905
rect 29821 2125 29922 2140
rect 29821 2035 29826 2125
rect 29910 2035 29922 2125
rect 29821 2026 29922 2035
rect 34961 2034 35087 15005
rect 36474 14492 36576 14502
rect 36474 14392 36479 14492
rect 36573 14392 36576 14492
rect 36474 14382 36576 14392
rect 38715 14478 38795 14512
rect 38715 14394 38723 14478
rect 38791 14394 38795 14478
rect 38715 14346 38795 14394
rect 36478 11290 36580 11300
rect 36478 11190 36483 11290
rect 36577 11190 36580 11290
rect 36478 11180 36580 11190
rect 38719 11276 38799 11310
rect 38719 11192 38727 11276
rect 38795 11192 38799 11276
rect 38719 11144 38799 11192
rect 34961 1961 34981 2034
rect 35068 1961 35087 2034
rect 34961 1942 35087 1961
rect 35256 9545 37818 9662
rect 30063 1880 30161 1898
rect 30063 1808 30073 1880
rect 30143 1808 30161 1880
rect 30063 1800 30161 1808
rect 33691 1683 33701 1799
rect 34039 1683 34049 1799
rect 32146 812 32156 1007
rect 32422 812 32432 1007
rect 29583 717 29794 722
rect 29583 642 29723 717
rect 29784 642 29794 717
rect 29583 637 29794 642
rect 30281 676 30383 692
rect 30281 608 30295 676
rect 30369 608 30383 676
rect 30281 594 30383 608
rect 29015 377 29176 508
rect 35256 377 35360 9545
rect 37726 9528 37818 9545
rect 37726 9460 37737 9528
rect 37727 9455 37737 9460
rect 37807 9460 37818 9528
rect 37807 9455 37817 9460
rect 37727 9450 37817 9455
rect 36478 8146 36580 8156
rect 36478 8046 36483 8146
rect 36577 8046 36580 8146
rect 36478 8036 36580 8046
rect 38719 8132 38799 8166
rect 38719 8048 38727 8132
rect 38795 8048 38799 8132
rect 38719 8000 38799 8048
rect 36474 5014 36576 5024
rect 36474 4914 36479 5014
rect 36573 4914 36576 5014
rect 36474 4904 36576 4914
rect 38715 5000 38795 5034
rect 38715 4916 38723 5000
rect 38791 4916 38795 5000
rect 38715 4868 38795 4916
rect 36474 1870 36576 1880
rect 36474 1770 36479 1870
rect 36573 1770 36576 1870
rect 36474 1760 36576 1770
rect 38715 1856 38795 1890
rect 38715 1772 38723 1856
rect 38791 1772 38795 1856
rect 38715 1724 38795 1772
rect 29015 273 35360 377
rect -1320 142 -586 144
rect -2700 128 -586 142
rect -2700 43 -2690 128
rect -2604 43 -586 128
rect -2700 28 -586 43
rect -1464 27 -586 28
<< via3 >>
rect 6250 27917 6449 27948
rect 6250 27788 6272 27917
rect 6272 27788 6425 27917
rect 6425 27788 6449 27917
rect 6250 27769 6449 27788
rect 8732 27971 8931 28002
rect 8732 27842 8754 27971
rect 8754 27842 8907 27971
rect 8907 27842 8931 27971
rect 8732 27823 8931 27842
rect 9879 27971 10078 28002
rect 9879 27842 9901 27971
rect 9901 27842 10054 27971
rect 10054 27842 10078 27971
rect 9879 27823 10078 27842
rect 12763 27914 12962 27945
rect 12763 27785 12785 27914
rect 12785 27785 12938 27914
rect 12938 27785 12962 27914
rect 12763 27766 12962 27785
rect 15245 27968 15444 27999
rect 15245 27839 15267 27968
rect 15267 27839 15420 27968
rect 15420 27839 15444 27968
rect 15245 27820 15444 27839
rect 16392 27968 16591 27999
rect 16392 27839 16414 27968
rect 16414 27839 16567 27968
rect 16567 27839 16591 27968
rect 16392 27820 16591 27839
rect 19297 27909 19496 27940
rect 19297 27780 19319 27909
rect 19319 27780 19472 27909
rect 19472 27780 19496 27909
rect 19297 27761 19496 27780
rect 21779 27963 21978 27994
rect 21779 27834 21801 27963
rect 21801 27834 21954 27963
rect 21954 27834 21978 27963
rect 21779 27815 21978 27834
rect 22926 27963 23125 27994
rect 22926 27834 22948 27963
rect 22948 27834 23101 27963
rect 23101 27834 23125 27963
rect 22926 27815 23125 27834
rect 25855 27913 26054 27944
rect 25855 27784 25877 27913
rect 25877 27784 26030 27913
rect 26030 27784 26054 27913
rect 25855 27765 26054 27784
rect 28337 27967 28536 27998
rect 28337 27838 28359 27967
rect 28359 27838 28512 27967
rect 28512 27838 28536 27967
rect 28337 27819 28536 27838
rect 29484 27967 29683 27998
rect 29484 27838 29506 27967
rect 29506 27838 29659 27967
rect 29659 27838 29683 27967
rect 29484 27819 29683 27838
rect 6534 26878 6713 26900
rect 6534 26725 6553 26878
rect 6553 26725 6682 26878
rect 6682 26725 6713 26878
rect 6534 26701 6713 26725
rect 13047 26875 13226 26897
rect 13047 26722 13066 26875
rect 13066 26722 13195 26875
rect 13195 26722 13226 26875
rect 13047 26698 13226 26722
rect 19581 26870 19760 26892
rect 19581 26717 19600 26870
rect 19600 26717 19729 26870
rect 19729 26717 19760 26870
rect 19581 26693 19760 26717
rect 26139 26874 26318 26896
rect 26139 26721 26158 26874
rect 26158 26721 26287 26874
rect 26287 26721 26318 26874
rect 26139 26697 26318 26721
rect 8077 26570 8276 26589
rect 8077 26441 8101 26570
rect 8101 26441 8254 26570
rect 8254 26441 8276 26570
rect 8077 26410 8276 26441
rect 9219 26568 9418 26587
rect 9219 26439 9243 26568
rect 9243 26439 9396 26568
rect 9396 26439 9418 26568
rect 9219 26408 9418 26439
rect 14590 26567 14789 26586
rect 14590 26438 14614 26567
rect 14614 26438 14767 26567
rect 14767 26438 14789 26567
rect 14590 26407 14789 26438
rect 15732 26565 15931 26584
rect 15732 26436 15756 26565
rect 15756 26436 15909 26565
rect 15909 26436 15931 26565
rect 15732 26405 15931 26436
rect 21124 26562 21323 26581
rect 21124 26433 21148 26562
rect 21148 26433 21301 26562
rect 21301 26433 21323 26562
rect 21124 26402 21323 26433
rect 22266 26560 22465 26579
rect 22266 26431 22290 26560
rect 22290 26431 22443 26560
rect 22443 26431 22465 26560
rect 22266 26400 22465 26431
rect 27682 26566 27881 26585
rect 27682 26437 27706 26566
rect 27706 26437 27859 26566
rect 27859 26437 27881 26566
rect 27682 26406 27881 26437
rect 28824 26564 29023 26583
rect 28824 26435 28848 26564
rect 28848 26435 29001 26564
rect 29001 26435 29023 26564
rect 28824 26404 29023 26435
rect -4065 15364 -4063 15440
rect -4063 15364 -3999 15440
rect -1843 15492 -1755 15502
rect -1843 15420 -1833 15492
rect -1833 15420 -1763 15492
rect -1763 15420 -1755 15492
rect -1843 15408 -1755 15420
rect 6264 26267 6463 26298
rect 6264 26138 6286 26267
rect 6286 26138 6439 26267
rect 6439 26138 6463 26267
rect 6264 26119 6463 26138
rect 12777 26264 12976 26295
rect 12777 26135 12799 26264
rect 12799 26135 12952 26264
rect 12952 26135 12976 26264
rect 12777 26116 12976 26135
rect 8077 25924 8276 25955
rect 8077 25795 8099 25924
rect 8099 25795 8252 25924
rect 8252 25795 8276 25924
rect 8077 25776 8276 25795
rect 9975 25924 10174 25955
rect 9975 25795 9997 25924
rect 9997 25795 10150 25924
rect 10150 25795 10174 25924
rect 9975 25776 10174 25795
rect 6548 25228 6727 25250
rect 6548 25075 6567 25228
rect 6567 25075 6696 25228
rect 6696 25075 6727 25228
rect 6548 25051 6727 25075
rect 6259 24663 6458 24694
rect 6259 24534 6281 24663
rect 6281 24534 6434 24663
rect 6434 24534 6458 24663
rect 6259 24515 6458 24534
rect 6543 23624 6722 23646
rect 6543 23471 6562 23624
rect 6562 23471 6691 23624
rect 6691 23471 6722 23624
rect 6543 23447 6722 23471
rect 8021 23527 8220 23546
rect 8021 23398 8045 23527
rect 8045 23398 8198 23527
rect 8198 23398 8220 23527
rect 8021 23367 8220 23398
rect 9919 23527 10118 23546
rect 9919 23398 9943 23527
rect 9943 23398 10096 23527
rect 10096 23398 10118 23527
rect 9919 23367 10118 23398
rect 14590 25921 14789 25952
rect 14590 25792 14612 25921
rect 14612 25792 14765 25921
rect 14765 25792 14789 25921
rect 14590 25773 14789 25792
rect 16488 25921 16687 25952
rect 16488 25792 16510 25921
rect 16510 25792 16663 25921
rect 16663 25792 16687 25921
rect 16488 25773 16687 25792
rect 13061 25225 13240 25247
rect 13061 25072 13080 25225
rect 13080 25072 13209 25225
rect 13209 25072 13240 25225
rect 13061 25048 13240 25072
rect 12772 24660 12971 24691
rect 12772 24531 12794 24660
rect 12794 24531 12947 24660
rect 12947 24531 12971 24660
rect 12772 24512 12971 24531
rect 13056 23621 13235 23643
rect 13056 23468 13075 23621
rect 13075 23468 13204 23621
rect 13204 23468 13235 23621
rect 13056 23444 13235 23468
rect 14534 23524 14733 23543
rect 14534 23395 14558 23524
rect 14558 23395 14711 23524
rect 14711 23395 14733 23524
rect 14534 23364 14733 23395
rect 16432 23524 16631 23543
rect 16432 23395 16456 23524
rect 16456 23395 16609 23524
rect 16609 23395 16631 23524
rect 16432 23364 16631 23395
rect -4067 13296 -4065 13372
rect -4065 13296 -4001 13372
rect -1845 13424 -1757 13434
rect -1845 13352 -1835 13424
rect -1835 13352 -1765 13424
rect -1765 13352 -1757 13424
rect -1845 13340 -1757 13352
rect 19311 26259 19510 26290
rect 19311 26130 19333 26259
rect 19333 26130 19486 26259
rect 19486 26130 19510 26259
rect 19311 26111 19510 26130
rect 21124 25916 21323 25947
rect 21124 25787 21146 25916
rect 21146 25787 21299 25916
rect 21299 25787 21323 25916
rect 21124 25768 21323 25787
rect 23022 25916 23221 25947
rect 23022 25787 23044 25916
rect 23044 25787 23197 25916
rect 23197 25787 23221 25916
rect 23022 25768 23221 25787
rect 19595 25220 19774 25242
rect 19595 25067 19614 25220
rect 19614 25067 19743 25220
rect 19743 25067 19774 25220
rect 19595 25043 19774 25067
rect 19306 24655 19505 24686
rect 19306 24526 19328 24655
rect 19328 24526 19481 24655
rect 19481 24526 19505 24655
rect 19306 24507 19505 24526
rect 19590 23616 19769 23638
rect 19590 23463 19609 23616
rect 19609 23463 19738 23616
rect 19738 23463 19769 23616
rect 19590 23439 19769 23463
rect 21068 23519 21267 23538
rect 21068 23390 21092 23519
rect 21092 23390 21245 23519
rect 21245 23390 21267 23519
rect 21068 23359 21267 23390
rect 22966 23519 23165 23538
rect 22966 23390 22990 23519
rect 22990 23390 23143 23519
rect 23143 23390 23165 23519
rect 22966 23359 23165 23390
rect -4065 11227 -4063 11303
rect -4063 11227 -3999 11303
rect -1843 11355 -1755 11365
rect -1843 11283 -1833 11355
rect -1833 11283 -1763 11355
rect -1763 11283 -1755 11355
rect -1843 11271 -1755 11283
rect 25869 26263 26068 26294
rect 25869 26134 25891 26263
rect 25891 26134 26044 26263
rect 26044 26134 26068 26263
rect 25869 26115 26068 26134
rect 27682 25920 27881 25951
rect 27682 25791 27704 25920
rect 27704 25791 27857 25920
rect 27857 25791 27881 25920
rect 27682 25772 27881 25791
rect 29580 25920 29779 25951
rect 29580 25791 29602 25920
rect 29602 25791 29755 25920
rect 29755 25791 29779 25920
rect 29580 25772 29779 25791
rect 26153 25224 26332 25246
rect 26153 25071 26172 25224
rect 26172 25071 26301 25224
rect 26301 25071 26332 25224
rect 26153 25047 26332 25071
rect 25864 24659 26063 24690
rect 25864 24530 25886 24659
rect 25886 24530 26039 24659
rect 26039 24530 26063 24659
rect 25864 24511 26063 24530
rect 36485 23812 36575 23912
rect 36575 23812 36577 23912
rect 38727 23892 38795 23898
rect 38727 23816 38785 23892
rect 38785 23816 38795 23892
rect 38727 23814 38795 23816
rect 26148 23620 26327 23642
rect 26148 23467 26167 23620
rect 26167 23467 26296 23620
rect 26296 23467 26327 23620
rect 26148 23443 26327 23467
rect 27626 23523 27825 23542
rect 27626 23394 27650 23523
rect 27650 23394 27803 23523
rect 27803 23394 27825 23523
rect 27626 23363 27825 23394
rect 29524 23523 29723 23542
rect 29524 23394 29548 23523
rect 29548 23394 29701 23523
rect 29701 23394 29723 23523
rect 29524 23363 29723 23394
rect -4067 9159 -4065 9235
rect -4065 9159 -4001 9235
rect -1845 9287 -1757 9297
rect -1845 9215 -1835 9287
rect -1835 9215 -1765 9287
rect -1765 9215 -1757 9287
rect -1845 9203 -1757 9215
rect 5826 22363 6025 22394
rect 5826 22234 5850 22363
rect 5850 22234 6003 22363
rect 6003 22234 6025 22363
rect 5826 22215 6025 22234
rect 6973 22363 7172 22394
rect 6973 22234 6997 22363
rect 6997 22234 7150 22363
rect 7150 22234 7172 22363
rect 6973 22215 7172 22234
rect 9455 22309 9654 22340
rect 9455 22180 9479 22309
rect 9479 22180 9632 22309
rect 9632 22180 9654 22309
rect 9455 22161 9654 22180
rect 12384 22359 12583 22390
rect 12384 22230 12408 22359
rect 12408 22230 12561 22359
rect 12561 22230 12583 22359
rect 12384 22211 12583 22230
rect 13531 22359 13730 22390
rect 13531 22230 13555 22359
rect 13555 22230 13708 22359
rect 13708 22230 13730 22359
rect 13531 22211 13730 22230
rect 16013 22305 16212 22336
rect 16013 22176 16037 22305
rect 16037 22176 16190 22305
rect 16190 22176 16212 22305
rect 16013 22157 16212 22176
rect 18918 22364 19117 22395
rect 18918 22235 18942 22364
rect 18942 22235 19095 22364
rect 19095 22235 19117 22364
rect 18918 22216 19117 22235
rect 20065 22364 20264 22395
rect 20065 22235 20089 22364
rect 20089 22235 20242 22364
rect 20242 22235 20264 22364
rect 20065 22216 20264 22235
rect 22547 22310 22746 22341
rect 22547 22181 22571 22310
rect 22571 22181 22724 22310
rect 22724 22181 22746 22310
rect 22547 22162 22746 22181
rect 25431 22367 25630 22398
rect 25431 22238 25455 22367
rect 25455 22238 25608 22367
rect 25608 22238 25630 22367
rect 25431 22219 25630 22238
rect 26578 22367 26777 22398
rect 26578 22238 26602 22367
rect 26602 22238 26755 22367
rect 26755 22238 26777 22367
rect 26578 22219 26777 22238
rect 29060 22313 29259 22344
rect 29060 22184 29084 22313
rect 29084 22184 29237 22313
rect 29237 22184 29259 22313
rect 29060 22165 29259 22184
rect 9191 21270 9370 21292
rect 9191 21117 9222 21270
rect 9222 21117 9351 21270
rect 9351 21117 9370 21270
rect 9191 21093 9370 21117
rect 15749 21266 15928 21288
rect 15749 21113 15780 21266
rect 15780 21113 15909 21266
rect 15909 21113 15928 21266
rect 15749 21089 15928 21113
rect 22283 21271 22462 21293
rect 22283 21118 22314 21271
rect 22314 21118 22443 21271
rect 22443 21118 22462 21271
rect 22283 21094 22462 21118
rect 28796 21274 28975 21296
rect 28796 21121 28827 21274
rect 28827 21121 28956 21274
rect 28956 21121 28975 21274
rect 28796 21097 28975 21121
rect 6486 20960 6685 20979
rect 6486 20831 6508 20960
rect 6508 20831 6661 20960
rect 6661 20831 6685 20960
rect 6486 20800 6685 20831
rect 7628 20962 7827 20981
rect 7628 20833 7650 20962
rect 7650 20833 7803 20962
rect 7803 20833 7827 20962
rect 7628 20802 7827 20833
rect 13044 20956 13243 20975
rect 13044 20827 13066 20956
rect 13066 20827 13219 20956
rect 13219 20827 13243 20956
rect 13044 20796 13243 20827
rect 14186 20958 14385 20977
rect 14186 20829 14208 20958
rect 14208 20829 14361 20958
rect 14361 20829 14385 20958
rect 14186 20798 14385 20829
rect 19578 20961 19777 20980
rect 19578 20832 19600 20961
rect 19600 20832 19753 20961
rect 19753 20832 19777 20961
rect 19578 20801 19777 20832
rect 20720 20963 20919 20982
rect 20720 20834 20742 20963
rect 20742 20834 20895 20963
rect 20895 20834 20919 20963
rect 20720 20803 20919 20834
rect 26091 20964 26290 20983
rect 26091 20835 26113 20964
rect 26113 20835 26266 20964
rect 26266 20835 26290 20964
rect 26091 20804 26290 20835
rect 27233 20966 27432 20985
rect 27233 20837 27255 20966
rect 27255 20837 27408 20966
rect 27408 20837 27432 20966
rect 27233 20806 27432 20837
rect 9441 20659 9640 20690
rect 9441 20530 9465 20659
rect 9465 20530 9618 20659
rect 9618 20530 9640 20659
rect 9441 20511 9640 20530
rect 15999 20655 16198 20686
rect 15999 20526 16023 20655
rect 16023 20526 16176 20655
rect 16176 20526 16198 20655
rect 15999 20507 16198 20526
rect 22533 20660 22732 20691
rect 22533 20531 22557 20660
rect 22557 20531 22710 20660
rect 22710 20531 22732 20660
rect 22533 20512 22732 20531
rect 29046 20663 29245 20694
rect 29046 20534 29070 20663
rect 29070 20534 29223 20663
rect 29223 20534 29245 20663
rect 29046 20515 29245 20534
rect 36485 20668 36575 20768
rect 36575 20668 36577 20768
rect 38727 20748 38795 20754
rect 38727 20672 38785 20748
rect 38785 20672 38795 20748
rect 38727 20670 38795 20672
rect 5730 20316 5929 20347
rect 5730 20187 5754 20316
rect 5754 20187 5907 20316
rect 5907 20187 5929 20316
rect 5730 20168 5929 20187
rect 7628 20316 7827 20347
rect 7628 20187 7652 20316
rect 7652 20187 7805 20316
rect 7805 20187 7827 20316
rect 7628 20168 7827 20187
rect 12288 20312 12487 20343
rect 12288 20183 12312 20312
rect 12312 20183 12465 20312
rect 12465 20183 12487 20312
rect 12288 20164 12487 20183
rect 14186 20312 14385 20343
rect 14186 20183 14210 20312
rect 14210 20183 14363 20312
rect 14363 20183 14385 20312
rect 14186 20164 14385 20183
rect 18822 20317 19021 20348
rect 18822 20188 18846 20317
rect 18846 20188 18999 20317
rect 18999 20188 19021 20317
rect 18822 20169 19021 20188
rect 20720 20317 20919 20348
rect 20720 20188 20744 20317
rect 20744 20188 20897 20317
rect 20897 20188 20919 20317
rect 20720 20169 20919 20188
rect 25335 20320 25534 20351
rect 25335 20191 25359 20320
rect 25359 20191 25512 20320
rect 25512 20191 25534 20320
rect 25335 20172 25534 20191
rect 27233 20320 27432 20351
rect 27233 20191 27257 20320
rect 27257 20191 27410 20320
rect 27410 20191 27432 20320
rect 27233 20172 27432 20191
rect 9177 19620 9356 19642
rect 9177 19467 9208 19620
rect 9208 19467 9337 19620
rect 9337 19467 9356 19620
rect 9177 19443 9356 19467
rect 15735 19616 15914 19638
rect 15735 19463 15766 19616
rect 15766 19463 15895 19616
rect 15895 19463 15914 19616
rect 15735 19439 15914 19463
rect 22269 19621 22448 19643
rect 22269 19468 22300 19621
rect 22300 19468 22429 19621
rect 22429 19468 22448 19621
rect 22269 19444 22448 19468
rect 28782 19624 28961 19646
rect 28782 19471 28813 19624
rect 28813 19471 28942 19624
rect 28942 19471 28961 19624
rect 28782 19447 28961 19471
rect 9446 19055 9645 19086
rect 9446 18926 9470 19055
rect 9470 18926 9623 19055
rect 9623 18926 9645 19055
rect 9446 18907 9645 18926
rect 16004 19051 16203 19082
rect 16004 18922 16028 19051
rect 16028 18922 16181 19051
rect 16181 18922 16203 19051
rect 16004 18903 16203 18922
rect 22538 19056 22737 19087
rect 22538 18927 22562 19056
rect 22562 18927 22715 19056
rect 22715 18927 22737 19056
rect 22538 18908 22737 18927
rect 29051 19059 29250 19090
rect 29051 18930 29075 19059
rect 29075 18930 29228 19059
rect 29228 18930 29250 19059
rect 29051 18911 29250 18930
rect 9182 18016 9361 18038
rect 5786 17919 5985 17938
rect 5786 17790 5808 17919
rect 5808 17790 5961 17919
rect 5961 17790 5985 17919
rect 5786 17759 5985 17790
rect 7684 17919 7883 17938
rect 7684 17790 7706 17919
rect 7706 17790 7859 17919
rect 7859 17790 7883 17919
rect 7684 17759 7883 17790
rect 9182 17863 9213 18016
rect 9213 17863 9342 18016
rect 9342 17863 9361 18016
rect 15740 18012 15919 18034
rect 9182 17839 9361 17863
rect 12344 17915 12543 17934
rect 12344 17786 12366 17915
rect 12366 17786 12519 17915
rect 12519 17786 12543 17915
rect 12344 17755 12543 17786
rect 14242 17915 14441 17934
rect 14242 17786 14264 17915
rect 14264 17786 14417 17915
rect 14417 17786 14441 17915
rect 14242 17755 14441 17786
rect 15740 17859 15771 18012
rect 15771 17859 15900 18012
rect 15900 17859 15919 18012
rect 22274 18017 22453 18039
rect 15740 17835 15919 17859
rect 18878 17920 19077 17939
rect 18878 17791 18900 17920
rect 18900 17791 19053 17920
rect 19053 17791 19077 17920
rect 18878 17760 19077 17791
rect 20776 17920 20975 17939
rect 20776 17791 20798 17920
rect 20798 17791 20951 17920
rect 20951 17791 20975 17920
rect 20776 17760 20975 17791
rect 22274 17864 22305 18017
rect 22305 17864 22434 18017
rect 22434 17864 22453 18017
rect 28787 18020 28966 18042
rect 22274 17840 22453 17864
rect 25391 17923 25590 17942
rect 25391 17794 25413 17923
rect 25413 17794 25566 17923
rect 25566 17794 25590 17923
rect 25391 17763 25590 17794
rect 27289 17923 27488 17942
rect 27289 17794 27311 17923
rect 27311 17794 27464 17923
rect 27464 17794 27488 17923
rect 27289 17763 27488 17794
rect 28787 17867 28818 18020
rect 28818 17867 28947 18020
rect 28947 17867 28966 18020
rect 28787 17843 28966 17867
rect 36481 17536 36571 17636
rect 36571 17536 36573 17636
rect 38723 17616 38791 17622
rect 38723 17540 38781 17616
rect 38781 17540 38791 17616
rect 38723 17538 38791 17540
rect -4067 7090 -4065 7166
rect -4065 7090 -4001 7166
rect -1845 7218 -1757 7228
rect -1845 7146 -1835 7218
rect -1835 7146 -1765 7218
rect -1765 7146 -1757 7218
rect -1845 7134 -1757 7146
rect -4069 5022 -4067 5098
rect -4067 5022 -4003 5098
rect -1847 5150 -1759 5160
rect -1847 5078 -1837 5150
rect -1837 5078 -1767 5150
rect -1767 5078 -1759 5150
rect -1847 5066 -1759 5078
rect -4067 2953 -4065 3029
rect -4065 2953 -4001 3029
rect -1845 3081 -1757 3091
rect -1845 3009 -1835 3081
rect -1835 3009 -1765 3081
rect -1765 3009 -1757 3081
rect -1845 2997 -1757 3009
rect -4069 885 -4067 961
rect -4067 885 -4003 961
rect -1847 1013 -1759 1023
rect -1847 941 -1837 1013
rect -1837 941 -1767 1013
rect -1767 941 -1759 1013
rect -1847 929 -1759 941
rect 8147 15462 8217 15466
rect 8147 15400 8153 15462
rect 8153 15400 8213 15462
rect 8213 15400 8217 15462
rect 8147 15394 8217 15400
rect 14696 15461 14766 15465
rect 14696 15399 14702 15461
rect 14702 15399 14762 15461
rect 14762 15399 14766 15461
rect 14696 15393 14766 15399
rect 21350 15482 21420 15486
rect 21350 15420 21356 15482
rect 21356 15420 21416 15482
rect 21416 15420 21420 15482
rect 21350 15414 21420 15420
rect 30003 15315 30073 15319
rect 30003 15253 30009 15315
rect 30009 15253 30069 15315
rect 30069 15253 30073 15315
rect 30003 15247 30073 15253
rect 32233 15255 32432 15286
rect 32233 15126 32255 15255
rect 32255 15126 32408 15255
rect 32408 15126 32432 15255
rect 32233 15107 32432 15126
rect 33604 14907 33674 14911
rect 33604 14845 33610 14907
rect 33610 14845 33670 14907
rect 33670 14845 33674 14907
rect 33604 14839 33674 14845
rect 8369 14256 8443 14262
rect 8369 14194 8375 14256
rect 8375 14194 8439 14256
rect 8439 14194 8443 14256
rect 14918 14255 14992 14261
rect 14918 14193 14924 14255
rect 14924 14193 14988 14255
rect 14988 14193 14992 14255
rect 21572 14276 21646 14282
rect 21572 14214 21578 14276
rect 21578 14214 21642 14276
rect 21642 14214 21646 14276
rect 30225 14109 30299 14115
rect 30225 14047 30231 14109
rect 30231 14047 30295 14109
rect 30295 14047 30299 14109
rect 33699 13701 34037 13733
rect 33699 13639 33832 13701
rect 33832 13639 33896 13701
rect 33896 13639 34037 13701
rect 33699 13617 34037 13639
rect 1483 13562 1553 13566
rect 1483 13500 1489 13562
rect 1489 13500 1549 13562
rect 1549 13500 1553 13562
rect 1483 13494 1553 13500
rect 4446 13366 4645 13397
rect 4446 13237 4468 13366
rect 4468 13237 4621 13366
rect 4621 13237 4645 13366
rect 4446 13218 4645 13237
rect 6928 13420 7127 13451
rect 6928 13291 6950 13420
rect 6950 13291 7103 13420
rect 7103 13291 7127 13420
rect 6928 13272 7127 13291
rect 8075 13420 8274 13451
rect 8075 13291 8097 13420
rect 8097 13291 8250 13420
rect 8250 13291 8274 13420
rect 8075 13272 8274 13291
rect 10995 13454 11194 13485
rect 10995 13325 11017 13454
rect 11017 13325 11170 13454
rect 11170 13325 11194 13454
rect 10995 13306 11194 13325
rect 13477 13508 13676 13539
rect 13477 13379 13499 13508
rect 13499 13379 13652 13508
rect 13652 13379 13676 13508
rect 13477 13360 13676 13379
rect 14624 13508 14823 13539
rect 14624 13379 14646 13508
rect 14646 13379 14799 13508
rect 14799 13379 14823 13508
rect 14624 13360 14823 13379
rect 17649 13386 17848 13417
rect 17649 13257 17671 13386
rect 17671 13257 17824 13386
rect 17824 13257 17848 13386
rect 17649 13238 17848 13257
rect 20131 13440 20330 13471
rect 20131 13311 20153 13440
rect 20153 13311 20306 13440
rect 20306 13311 20330 13440
rect 20131 13292 20330 13311
rect 21278 13440 21477 13471
rect 21278 13311 21300 13440
rect 21300 13311 21453 13440
rect 21453 13311 21477 13440
rect 21278 13292 21477 13311
rect 24274 13454 24473 13485
rect 24274 13325 24296 13454
rect 24296 13325 24449 13454
rect 24449 13325 24473 13454
rect 24274 13306 24473 13325
rect 26756 13508 26955 13539
rect 26756 13379 26778 13508
rect 26778 13379 26931 13508
rect 26931 13379 26955 13508
rect 26756 13360 26955 13379
rect 27903 13508 28102 13539
rect 27903 13379 27925 13508
rect 27925 13379 28078 13508
rect 28078 13379 28102 13508
rect 27903 13360 28102 13379
rect 29998 12744 30068 12748
rect 29998 12682 30004 12744
rect 30004 12682 30064 12744
rect 30064 12682 30068 12744
rect 29998 12676 30068 12682
rect 32154 12925 32420 12941
rect 32154 12768 32177 12925
rect 32177 12768 32388 12925
rect 32388 12768 32420 12925
rect 32154 12746 32420 12768
rect 1705 12356 1779 12362
rect 1705 12294 1711 12356
rect 1711 12294 1775 12356
rect 1775 12294 1779 12356
rect 4730 12327 4909 12349
rect 4730 12174 4749 12327
rect 4749 12174 4878 12327
rect 4878 12174 4909 12327
rect 4730 12150 4909 12174
rect 6273 12019 6472 12038
rect 6273 11890 6297 12019
rect 6297 11890 6450 12019
rect 6450 11890 6472 12019
rect 6273 11859 6472 11890
rect 7415 12017 7614 12036
rect 7415 11888 7439 12017
rect 7439 11888 7592 12017
rect 7592 11888 7614 12017
rect 7415 11857 7614 11888
rect 4460 11716 4659 11747
rect 4460 11587 4482 11716
rect 4482 11587 4635 11716
rect 4635 11587 4659 11716
rect 4460 11568 4659 11587
rect 6273 11373 6472 11404
rect 6273 11244 6295 11373
rect 6295 11244 6448 11373
rect 6448 11244 6472 11373
rect 6273 11225 6472 11244
rect 8171 11373 8370 11404
rect 8171 11244 8193 11373
rect 8193 11244 8346 11373
rect 8346 11244 8370 11373
rect 8171 11225 8370 11244
rect 1475 10977 1545 10981
rect 1475 10915 1481 10977
rect 1481 10915 1541 10977
rect 1541 10915 1545 10977
rect 1475 10909 1545 10915
rect 4744 10677 4923 10699
rect 4744 10524 4763 10677
rect 4763 10524 4892 10677
rect 4892 10524 4923 10677
rect 4744 10500 4923 10524
rect 4455 10112 4654 10143
rect 4455 9983 4477 10112
rect 4477 9983 4630 10112
rect 4630 9983 4654 10112
rect 4455 9964 4654 9983
rect 1697 9771 1771 9777
rect 1697 9709 1703 9771
rect 1703 9709 1767 9771
rect 1767 9709 1771 9771
rect 4739 9073 4918 9095
rect 4739 8920 4758 9073
rect 4758 8920 4887 9073
rect 4887 8920 4918 9073
rect 4739 8896 4918 8920
rect 6217 8976 6416 8995
rect 6217 8847 6241 8976
rect 6241 8847 6394 8976
rect 6394 8847 6416 8976
rect 6217 8816 6416 8847
rect 8115 8976 8314 8995
rect 8115 8847 8139 8976
rect 8139 8847 8292 8976
rect 8292 8847 8314 8976
rect 8115 8816 8314 8847
rect 11279 12415 11458 12437
rect 11279 12262 11298 12415
rect 11298 12262 11427 12415
rect 11427 12262 11458 12415
rect 11279 12238 11458 12262
rect 17933 12347 18112 12369
rect 17933 12194 17952 12347
rect 17952 12194 18081 12347
rect 18081 12194 18112 12347
rect 17933 12170 18112 12194
rect 12822 12107 13021 12126
rect 12822 11978 12846 12107
rect 12846 11978 12999 12107
rect 12999 11978 13021 12107
rect 12822 11947 13021 11978
rect 13964 12105 14163 12124
rect 13964 11976 13988 12105
rect 13988 11976 14141 12105
rect 14141 11976 14163 12105
rect 13964 11945 14163 11976
rect 19476 12039 19675 12058
rect 19476 11910 19500 12039
rect 19500 11910 19653 12039
rect 19653 11910 19675 12039
rect 19476 11879 19675 11910
rect 20618 12037 20817 12056
rect 20618 11908 20642 12037
rect 20642 11908 20795 12037
rect 20795 11908 20817 12037
rect 20618 11877 20817 11908
rect 11009 11804 11208 11835
rect 11009 11675 11031 11804
rect 11031 11675 11184 11804
rect 11184 11675 11208 11804
rect 11009 11656 11208 11675
rect 17663 11736 17862 11767
rect 17663 11607 17685 11736
rect 17685 11607 17838 11736
rect 17838 11607 17862 11736
rect 17663 11588 17862 11607
rect 12822 11461 13021 11492
rect 12822 11332 12844 11461
rect 12844 11332 12997 11461
rect 12997 11332 13021 11461
rect 12822 11313 13021 11332
rect 14720 11461 14919 11492
rect 14720 11332 14742 11461
rect 14742 11332 14895 11461
rect 14895 11332 14919 11461
rect 14720 11313 14919 11332
rect 19476 11393 19675 11424
rect 19476 11264 19498 11393
rect 19498 11264 19651 11393
rect 19651 11264 19675 11393
rect 19476 11245 19675 11264
rect 21374 11393 21573 11424
rect 21374 11264 21396 11393
rect 21396 11264 21549 11393
rect 21549 11264 21573 11393
rect 21374 11245 21573 11264
rect 11293 10765 11472 10787
rect 11293 10612 11312 10765
rect 11312 10612 11441 10765
rect 11441 10612 11472 10765
rect 11293 10588 11472 10612
rect 17947 10697 18126 10719
rect 17947 10544 17966 10697
rect 17966 10544 18095 10697
rect 18095 10544 18126 10697
rect 17947 10520 18126 10544
rect 11004 10200 11203 10231
rect 11004 10071 11026 10200
rect 11026 10071 11179 10200
rect 11179 10071 11203 10200
rect 11004 10052 11203 10071
rect 17658 10132 17857 10163
rect 17658 10003 17680 10132
rect 17680 10003 17833 10132
rect 17833 10003 17857 10132
rect 17658 9984 17857 10003
rect 11288 9161 11467 9183
rect 11288 9008 11307 9161
rect 11307 9008 11436 9161
rect 11436 9008 11467 9161
rect 17942 9093 18121 9115
rect 11288 8984 11467 9008
rect 12766 9064 12965 9083
rect 12766 8935 12790 9064
rect 12790 8935 12943 9064
rect 12943 8935 12965 9064
rect 12766 8904 12965 8935
rect 14664 9064 14863 9083
rect 14664 8935 14688 9064
rect 14688 8935 14841 9064
rect 14841 8935 14863 9064
rect 14664 8904 14863 8935
rect 17942 8940 17961 9093
rect 17961 8940 18090 9093
rect 18090 8940 18121 9093
rect 17942 8916 18121 8940
rect 19420 8996 19619 9015
rect 19420 8867 19444 8996
rect 19444 8867 19597 8996
rect 19597 8867 19619 8996
rect 19420 8836 19619 8867
rect 21318 8996 21517 9015
rect 21318 8867 21342 8996
rect 21342 8867 21495 8996
rect 21495 8867 21517 8996
rect 21318 8836 21517 8867
rect 1456 7699 1526 7703
rect 1456 7637 1462 7699
rect 1462 7637 1522 7699
rect 1522 7637 1526 7699
rect 1456 7631 1526 7637
rect 1678 6493 1752 6499
rect 1678 6431 1684 6493
rect 1684 6431 1748 6493
rect 1748 6431 1752 6493
rect 1472 4939 1542 4943
rect 1472 4877 1478 4939
rect 1478 4877 1538 4939
rect 1538 4877 1542 4939
rect 1472 4871 1542 4877
rect 4438 7586 4637 7617
rect 4438 7457 4460 7586
rect 4460 7457 4613 7586
rect 4613 7457 4637 7586
rect 4438 7438 4637 7457
rect 6920 7640 7119 7671
rect 6920 7511 6942 7640
rect 6942 7511 7095 7640
rect 7095 7511 7119 7640
rect 6920 7492 7119 7511
rect 8067 7640 8266 7671
rect 8067 7511 8089 7640
rect 8089 7511 8242 7640
rect 8242 7511 8266 7640
rect 8067 7492 8266 7511
rect 4722 6547 4901 6569
rect 4722 6394 4741 6547
rect 4741 6394 4870 6547
rect 4870 6394 4901 6547
rect 4722 6370 4901 6394
rect 6265 6239 6464 6258
rect 6265 6110 6289 6239
rect 6289 6110 6442 6239
rect 6442 6110 6464 6239
rect 6265 6079 6464 6110
rect 7407 6237 7606 6256
rect 7407 6108 7431 6237
rect 7431 6108 7584 6237
rect 7584 6108 7606 6237
rect 7407 6077 7606 6108
rect 4452 5936 4651 5967
rect 4452 5807 4474 5936
rect 4474 5807 4627 5936
rect 4627 5807 4651 5936
rect 4452 5788 4651 5807
rect 6265 5593 6464 5624
rect 6265 5464 6287 5593
rect 6287 5464 6440 5593
rect 6440 5464 6464 5593
rect 6265 5445 6464 5464
rect 8163 5593 8362 5624
rect 8163 5464 8185 5593
rect 8185 5464 8338 5593
rect 8338 5464 8362 5593
rect 8163 5445 8362 5464
rect 24558 12415 24737 12437
rect 24558 12262 24577 12415
rect 24577 12262 24706 12415
rect 24706 12262 24737 12415
rect 24558 12238 24737 12262
rect 26101 12107 26300 12126
rect 26101 11978 26125 12107
rect 26125 11978 26278 12107
rect 26278 11978 26300 12107
rect 26101 11947 26300 11978
rect 27243 12105 27442 12124
rect 27243 11976 27267 12105
rect 27267 11976 27420 12105
rect 27420 11976 27442 12105
rect 27243 11945 27442 11976
rect 24288 11804 24487 11835
rect 24288 11675 24310 11804
rect 24310 11675 24463 11804
rect 24463 11675 24487 11804
rect 24288 11656 24487 11675
rect 26101 11461 26300 11492
rect 26101 11332 26123 11461
rect 26123 11332 26276 11461
rect 26276 11332 26300 11461
rect 26101 11313 26300 11332
rect 27999 11461 28198 11492
rect 27999 11332 28021 11461
rect 28021 11332 28174 11461
rect 28174 11332 28198 11461
rect 27999 11313 28198 11332
rect 30220 11538 30294 11544
rect 30220 11476 30226 11538
rect 30226 11476 30290 11538
rect 30290 11476 30294 11538
rect 32235 11164 32434 11195
rect 32235 11035 32257 11164
rect 32257 11035 32410 11164
rect 32410 11035 32434 11164
rect 32235 11016 32434 11035
rect 24572 10765 24751 10787
rect 24572 10612 24591 10765
rect 24591 10612 24720 10765
rect 24720 10612 24751 10765
rect 33606 10816 33676 10820
rect 33606 10754 33612 10816
rect 33612 10754 33672 10816
rect 33672 10754 33676 10816
rect 33606 10748 33676 10754
rect 24572 10588 24751 10612
rect 24283 10200 24482 10231
rect 24283 10071 24305 10200
rect 24305 10071 24458 10200
rect 24458 10071 24482 10200
rect 24283 10052 24482 10071
rect 29998 9711 30068 9715
rect 29998 9649 30004 9711
rect 30004 9649 30064 9711
rect 30064 9649 30068 9711
rect 29998 9643 30068 9649
rect 33701 9610 34039 9642
rect 33701 9548 33834 9610
rect 33834 9548 33898 9610
rect 33898 9548 34039 9610
rect 33701 9526 34039 9548
rect 24567 9161 24746 9183
rect 24567 9008 24586 9161
rect 24586 9008 24715 9161
rect 24715 9008 24746 9161
rect 24567 8984 24746 9008
rect 26045 9064 26244 9083
rect 26045 8935 26069 9064
rect 26069 8935 26222 9064
rect 26222 8935 26244 9064
rect 26045 8904 26244 8935
rect 27943 9064 28142 9083
rect 27943 8935 27967 9064
rect 27967 8935 28120 9064
rect 28120 8935 28142 9064
rect 27943 8904 28142 8935
rect 32156 8834 32422 8850
rect 32156 8677 32179 8834
rect 32179 8677 32390 8834
rect 32390 8677 32422 8834
rect 32156 8655 32422 8677
rect 30220 8505 30294 8511
rect 30220 8443 30226 8505
rect 30226 8443 30290 8505
rect 30290 8443 30294 8505
rect 10989 7584 11188 7615
rect 10989 7455 11011 7584
rect 11011 7455 11164 7584
rect 11164 7455 11188 7584
rect 10989 7436 11188 7455
rect 13471 7638 13670 7669
rect 13471 7509 13493 7638
rect 13493 7509 13646 7638
rect 13646 7509 13670 7638
rect 13471 7490 13670 7509
rect 14618 7638 14817 7669
rect 14618 7509 14640 7638
rect 14640 7509 14793 7638
rect 14793 7509 14817 7638
rect 14618 7490 14817 7509
rect 11273 6545 11452 6567
rect 11273 6392 11292 6545
rect 11292 6392 11421 6545
rect 11421 6392 11452 6545
rect 11273 6368 11452 6392
rect 12816 6237 13015 6256
rect 12816 6108 12840 6237
rect 12840 6108 12993 6237
rect 12993 6108 13015 6237
rect 12816 6077 13015 6108
rect 13958 6235 14157 6254
rect 13958 6106 13982 6235
rect 13982 6106 14135 6235
rect 14135 6106 14157 6235
rect 13958 6075 14157 6106
rect 11003 5934 11202 5965
rect 11003 5805 11025 5934
rect 11025 5805 11178 5934
rect 11178 5805 11202 5934
rect 11003 5786 11202 5805
rect 12816 5591 13015 5622
rect 12816 5462 12838 5591
rect 12838 5462 12991 5591
rect 12991 5462 13015 5591
rect 12816 5443 13015 5462
rect 14714 5591 14913 5622
rect 14714 5462 14736 5591
rect 14736 5462 14889 5591
rect 14889 5462 14913 5591
rect 14714 5443 14913 5462
rect 4736 4897 4915 4919
rect 4736 4744 4755 4897
rect 4755 4744 4884 4897
rect 4884 4744 4915 4897
rect 11287 4895 11466 4917
rect 4736 4720 4915 4744
rect 11287 4742 11306 4895
rect 11306 4742 11435 4895
rect 11435 4742 11466 4895
rect 30069 7791 30139 7795
rect 30069 7729 30075 7791
rect 30075 7729 30135 7791
rect 30135 7729 30139 7791
rect 30069 7723 30139 7729
rect 17644 7585 17843 7616
rect 17644 7456 17666 7585
rect 17666 7456 17819 7585
rect 17819 7456 17843 7585
rect 17644 7437 17843 7456
rect 20126 7639 20325 7670
rect 20126 7510 20148 7639
rect 20148 7510 20301 7639
rect 20301 7510 20325 7639
rect 20126 7491 20325 7510
rect 21273 7639 21472 7670
rect 21273 7510 21295 7639
rect 21295 7510 21448 7639
rect 21448 7510 21472 7639
rect 21273 7491 21472 7510
rect 24266 7586 24465 7617
rect 24266 7457 24288 7586
rect 24288 7457 24441 7586
rect 24441 7457 24465 7586
rect 24266 7438 24465 7457
rect 26748 7640 26947 7671
rect 26748 7511 26770 7640
rect 26770 7511 26923 7640
rect 26923 7511 26947 7640
rect 26748 7492 26947 7511
rect 27895 7640 28094 7671
rect 27895 7511 27917 7640
rect 27917 7511 28070 7640
rect 28070 7511 28094 7640
rect 27895 7492 28094 7511
rect 32235 7669 32434 7700
rect 32235 7540 32257 7669
rect 32257 7540 32410 7669
rect 32410 7540 32434 7669
rect 32235 7521 32434 7540
rect 33606 7321 33676 7325
rect 33606 7259 33612 7321
rect 33612 7259 33672 7321
rect 33672 7259 33676 7321
rect 33606 7253 33676 7259
rect 17928 6546 18107 6568
rect 17928 6393 17947 6546
rect 17947 6393 18076 6546
rect 18076 6393 18107 6546
rect 17928 6369 18107 6393
rect 24550 6547 24729 6569
rect 24550 6394 24569 6547
rect 24569 6394 24698 6547
rect 24698 6394 24729 6547
rect 24550 6370 24729 6394
rect 19471 6238 19670 6257
rect 19471 6109 19495 6238
rect 19495 6109 19648 6238
rect 19648 6109 19670 6238
rect 19471 6078 19670 6109
rect 20613 6236 20812 6255
rect 20613 6107 20637 6236
rect 20637 6107 20790 6236
rect 20790 6107 20812 6236
rect 20613 6076 20812 6107
rect 26093 6239 26292 6258
rect 26093 6110 26117 6239
rect 26117 6110 26270 6239
rect 26270 6110 26292 6239
rect 26093 6079 26292 6110
rect 27235 6237 27434 6256
rect 27235 6108 27259 6237
rect 27259 6108 27412 6237
rect 27412 6108 27434 6237
rect 27235 6077 27434 6108
rect 17658 5935 17857 5966
rect 17658 5806 17680 5935
rect 17680 5806 17833 5935
rect 17833 5806 17857 5935
rect 17658 5787 17857 5806
rect 24280 5936 24479 5967
rect 24280 5807 24302 5936
rect 24302 5807 24455 5936
rect 24455 5807 24479 5936
rect 24280 5788 24479 5807
rect 19471 5592 19670 5623
rect 19471 5463 19493 5592
rect 19493 5463 19646 5592
rect 19646 5463 19670 5592
rect 19471 5444 19670 5463
rect 21369 5592 21568 5623
rect 21369 5463 21391 5592
rect 21391 5463 21544 5592
rect 21544 5463 21568 5592
rect 21369 5444 21568 5463
rect 26093 5593 26292 5624
rect 26093 5464 26115 5593
rect 26115 5464 26268 5593
rect 26268 5464 26292 5593
rect 26093 5445 26292 5464
rect 27991 5593 28190 5624
rect 27991 5464 28013 5593
rect 28013 5464 28166 5593
rect 28166 5464 28190 5593
rect 27991 5445 28190 5464
rect 17942 4896 18121 4918
rect 11287 4718 11466 4742
rect 17942 4743 17961 4896
rect 17961 4743 18090 4896
rect 18090 4743 18121 4896
rect 17942 4719 18121 4743
rect 24564 4897 24743 4919
rect 24564 4744 24583 4897
rect 24583 4744 24712 4897
rect 24712 4744 24743 4897
rect 24564 4720 24743 4744
rect 4447 4332 4646 4363
rect 4447 4203 4469 4332
rect 4469 4203 4622 4332
rect 4622 4203 4646 4332
rect 4447 4184 4646 4203
rect 10998 4330 11197 4361
rect 10998 4201 11020 4330
rect 11020 4201 11173 4330
rect 11173 4201 11197 4330
rect 10998 4182 11197 4201
rect 17653 4331 17852 4362
rect 17653 4202 17675 4331
rect 17675 4202 17828 4331
rect 17828 4202 17852 4331
rect 17653 4183 17852 4202
rect 24275 4332 24474 4363
rect 24275 4203 24297 4332
rect 24297 4203 24450 4332
rect 24450 4203 24474 4332
rect 24275 4184 24474 4203
rect 1694 3733 1768 3739
rect 1694 3671 1700 3733
rect 1700 3671 1764 3733
rect 1764 3671 1768 3733
rect 4731 3293 4910 3315
rect 4731 3140 4750 3293
rect 4750 3140 4879 3293
rect 4879 3140 4910 3293
rect 11282 3291 11461 3313
rect 4731 3116 4910 3140
rect 6209 3196 6408 3215
rect 6209 3067 6233 3196
rect 6233 3067 6386 3196
rect 6386 3067 6408 3196
rect 6209 3036 6408 3067
rect 8107 3196 8306 3215
rect 8107 3067 8131 3196
rect 8131 3067 8284 3196
rect 8284 3067 8306 3196
rect 8107 3036 8306 3067
rect 11282 3138 11301 3291
rect 11301 3138 11430 3291
rect 11430 3138 11461 3291
rect 17937 3292 18116 3314
rect 11282 3114 11461 3138
rect 12760 3194 12959 3213
rect 12760 3065 12784 3194
rect 12784 3065 12937 3194
rect 12937 3065 12959 3194
rect 12760 3034 12959 3065
rect 14658 3194 14857 3213
rect 14658 3065 14682 3194
rect 14682 3065 14835 3194
rect 14835 3065 14857 3194
rect 14658 3034 14857 3065
rect 17937 3139 17956 3292
rect 17956 3139 18085 3292
rect 18085 3139 18116 3292
rect 24559 3293 24738 3315
rect 17937 3115 18116 3139
rect 19415 3195 19614 3214
rect 19415 3066 19439 3195
rect 19439 3066 19592 3195
rect 19592 3066 19614 3195
rect 19415 3035 19614 3066
rect 21313 3195 21512 3214
rect 21313 3066 21337 3195
rect 21337 3066 21490 3195
rect 21490 3066 21512 3195
rect 21313 3035 21512 3066
rect 24559 3140 24578 3293
rect 24578 3140 24707 3293
rect 24707 3140 24738 3293
rect 24559 3116 24738 3140
rect 26037 3196 26236 3215
rect 26037 3067 26061 3196
rect 26061 3067 26214 3196
rect 26214 3067 26236 3196
rect 26037 3036 26236 3067
rect 27935 3196 28134 3215
rect 27935 3067 27959 3196
rect 27959 3067 28112 3196
rect 28112 3067 28134 3196
rect 27935 3036 28134 3067
rect 8404 2312 8410 2374
rect 8410 2312 8474 2374
rect 8474 2312 8478 2374
rect 8404 2306 8478 2312
rect 14958 2317 14964 2379
rect 14964 2317 15028 2379
rect 15028 2317 15032 2379
rect 14958 2311 15032 2317
rect 21607 2305 21613 2367
rect 21613 2305 21677 2367
rect 21677 2305 21681 2367
rect 21607 2299 21681 2305
rect 8182 1168 8252 1174
rect 8182 1106 8188 1168
rect 8188 1106 8248 1168
rect 8248 1106 8252 1168
rect 8182 1102 8252 1106
rect 14736 1173 14806 1179
rect 14736 1111 14742 1173
rect 14742 1111 14802 1173
rect 14802 1111 14806 1173
rect 14736 1107 14806 1111
rect 21385 1161 21455 1167
rect 21385 1099 21391 1161
rect 21391 1099 21451 1161
rect 21451 1099 21455 1161
rect 21385 1095 21455 1099
rect 30291 6585 30365 6591
rect 30291 6523 30297 6585
rect 30297 6523 30361 6585
rect 30361 6523 30365 6585
rect 33701 6115 34039 6147
rect 33701 6053 33834 6115
rect 33834 6053 33898 6115
rect 33898 6053 34039 6115
rect 33701 6031 34039 6053
rect 32156 5339 32422 5355
rect 32156 5182 32179 5339
rect 32179 5182 32390 5339
rect 32390 5182 32422 5339
rect 32156 5160 32422 5182
rect 30066 4721 30136 4725
rect 30066 4659 30072 4721
rect 30072 4659 30132 4721
rect 30132 4659 30136 4721
rect 30066 4653 30136 4659
rect 30288 3515 30362 3521
rect 30288 3453 30294 3515
rect 30294 3453 30358 3515
rect 30358 3453 30362 3515
rect 32235 3321 32434 3352
rect 32235 3192 32257 3321
rect 32257 3192 32410 3321
rect 32410 3192 32434 3321
rect 32235 3173 32434 3192
rect 33606 2973 33676 2977
rect 33606 2911 33612 2973
rect 33612 2911 33672 2973
rect 33672 2911 33676 2973
rect 33606 2905 33676 2911
rect 36481 14392 36571 14492
rect 36571 14392 36573 14492
rect 38723 14472 38791 14478
rect 38723 14396 38781 14472
rect 38781 14396 38791 14472
rect 38723 14394 38791 14396
rect 36485 11190 36575 11290
rect 36575 11190 36577 11290
rect 38727 11270 38795 11276
rect 38727 11194 38785 11270
rect 38785 11194 38795 11270
rect 38727 11192 38795 11194
rect 30073 1876 30143 1880
rect 30073 1814 30079 1876
rect 30079 1814 30139 1876
rect 30139 1814 30143 1876
rect 30073 1808 30143 1814
rect 33701 1767 34039 1799
rect 33701 1705 33834 1767
rect 33834 1705 33898 1767
rect 33898 1705 34039 1767
rect 33701 1683 34039 1705
rect 32156 991 32422 1007
rect 32156 834 32179 991
rect 32179 834 32390 991
rect 32390 834 32422 991
rect 32156 812 32422 834
rect 30295 670 30369 676
rect 30295 608 30301 670
rect 30301 608 30365 670
rect 30365 608 30369 670
rect 36485 8046 36575 8146
rect 36575 8046 36577 8146
rect 38727 8126 38795 8132
rect 38727 8050 38785 8126
rect 38785 8050 38795 8126
rect 38727 8048 38795 8050
rect 36481 4914 36571 5014
rect 36571 4914 36573 5014
rect 38723 4994 38791 5000
rect 38723 4918 38781 4994
rect 38781 4918 38791 4994
rect 38723 4916 38791 4918
rect 36481 1770 36571 1870
rect 36571 1770 36573 1870
rect 38723 1850 38791 1856
rect 38723 1774 38781 1850
rect 38781 1774 38791 1850
rect 38723 1772 38791 1774
<< metal4 >>
rect 2374 28310 5801 28315
rect 2374 28299 6236 28310
rect 16860 28299 19771 29436
rect 2374 28269 27084 28299
rect 30076 28269 36611 28277
rect 2374 28002 36611 28269
rect 2374 27959 8732 28002
rect 2370 27948 8732 27959
rect 2370 27769 6250 27948
rect 6449 27823 8732 27948
rect 8931 27823 9879 28002
rect 10078 27999 36611 28002
rect 10078 27945 15245 27999
rect 10078 27823 12763 27945
rect 6449 27769 12763 27823
rect 2370 27766 12763 27769
rect 12962 27820 15245 27945
rect 15444 27820 16392 27999
rect 16591 27998 36611 27999
rect 16591 27994 28337 27998
rect 16591 27940 21779 27994
rect 16591 27820 19297 27940
rect 12962 27766 19297 27820
rect 2370 27761 19297 27766
rect 19496 27815 21779 27940
rect 21978 27815 22926 27994
rect 23125 27944 28337 27994
rect 23125 27815 25855 27944
rect 19496 27765 25855 27815
rect 26054 27819 28337 27944
rect 28536 27819 29484 27998
rect 29683 27819 36611 27998
rect 26054 27765 36611 27819
rect 19496 27761 36611 27765
rect 2370 27564 36611 27761
rect 2370 22660 3884 27564
rect 4052 27563 4788 27564
rect 5384 27559 36611 27564
rect 5384 26512 6236 27559
rect 5384 26298 6604 26512
rect 5384 26119 6264 26298
rect 6463 26130 6604 26298
rect 6463 26125 6949 26130
rect 8827 26125 9174 26128
rect 10041 26125 10657 27559
rect 6463 26119 10657 26125
rect 5384 25955 10657 26119
rect 5384 25776 8077 25955
rect 8276 25776 9975 25955
rect 10174 25776 10657 25955
rect 5384 25620 10657 25776
rect 5384 24890 6236 25620
rect 10041 25615 10657 25620
rect 12222 26295 13117 26509
rect 12222 26116 12777 26295
rect 12976 26127 13117 26295
rect 12976 26122 13462 26127
rect 15340 26122 15687 26125
rect 16554 26122 17170 27559
rect 19276 27555 23704 27559
rect 12976 26116 17170 26122
rect 12222 25952 17170 26116
rect 12222 25773 14590 25952
rect 14789 25773 16488 25952
rect 16687 25773 17170 25952
rect 12222 25617 17170 25773
rect 5384 24694 6977 24890
rect 5384 24515 6259 24694
rect 6458 24515 6977 24694
rect 5384 24246 6977 24515
rect 12222 24887 12392 25617
rect 16554 25612 17170 25617
rect 18756 26290 19651 26504
rect 18756 26111 19311 26290
rect 19510 26122 19651 26290
rect 19510 26117 19996 26122
rect 21874 26117 22221 26120
rect 23088 26117 23704 27555
rect 19510 26111 23704 26117
rect 18756 25947 23704 26111
rect 18756 25768 21124 25947
rect 21323 25768 23022 25947
rect 23221 25768 23704 25947
rect 18756 25612 23704 25768
rect 12222 24691 13490 24887
rect 12222 24512 12772 24691
rect 12971 24512 13490 24691
rect 5384 22959 6236 24246
rect 12222 24243 13490 24512
rect 18756 24882 18926 25612
rect 23088 25607 23704 25612
rect 25314 26294 26209 26508
rect 25314 26115 25869 26294
rect 26068 26126 26209 26294
rect 26068 26121 26554 26126
rect 28432 26121 28779 26124
rect 29646 26121 36611 27559
rect 26068 26115 36611 26121
rect 25314 26035 36611 26115
rect 25314 25951 30262 26035
rect 25314 25772 27682 25951
rect 27881 25772 29580 25951
rect 29779 25772 30262 25951
rect 25314 25616 30262 25772
rect 25314 24886 25484 25616
rect 29646 25611 30262 25616
rect 18756 24686 20024 24882
rect 18756 24507 19306 24686
rect 19505 24507 20024 24686
rect 18756 24238 20024 24507
rect 25314 24690 26582 24886
rect 34620 24768 36611 26035
rect 25314 24511 25864 24690
rect 26063 24511 26582 24690
rect 25314 24242 26582 24511
rect 34612 24607 36611 24768
rect 34612 23912 36609 24607
rect 34612 23812 36485 23912
rect 36577 23812 36609 23912
rect 7997 23546 8242 23549
rect 7997 23528 8021 23546
rect 8220 23528 8242 23546
rect 9895 23546 10140 23549
rect 9895 23528 9919 23546
rect 10118 23528 10140 23546
rect 7893 23224 7917 23461
rect 8427 23224 9763 23410
rect 14510 23543 14755 23546
rect 14510 23525 14534 23543
rect 14733 23525 14755 23543
rect 16408 23543 16653 23546
rect 16408 23525 16432 23543
rect 16631 23525 16653 23543
rect 7893 23219 10260 23224
rect 14406 23221 14430 23458
rect 14940 23221 16276 23407
rect 21044 23538 21289 23541
rect 21044 23520 21068 23538
rect 21267 23520 21289 23538
rect 22942 23538 23187 23541
rect 22942 23520 22966 23538
rect 23165 23520 23187 23538
rect 8281 23217 9952 23219
rect 14406 23216 16773 23221
rect 20940 23216 20964 23453
rect 21474 23216 22810 23402
rect 27602 23542 27847 23545
rect 27602 23524 27626 23542
rect 27825 23524 27847 23542
rect 29500 23542 29745 23545
rect 29500 23524 29524 23542
rect 29723 23524 29745 23542
rect 27498 23220 27522 23457
rect 28032 23220 29368 23406
rect 14794 23214 16465 23216
rect 20940 23211 23307 23216
rect 27498 23215 29865 23220
rect 27886 23213 29557 23215
rect 21328 23209 22999 23211
rect 5380 22665 6237 22959
rect 29273 22690 30125 22695
rect 34612 22690 36609 23812
rect 38715 23639 38895 23672
rect 29273 22683 36609 22690
rect 8437 22665 36609 22683
rect 5376 22660 36609 22665
rect 2370 22398 36609 22660
rect 2370 22395 25431 22398
rect 2370 22394 18918 22395
rect 2370 22215 5826 22394
rect 6025 22215 6973 22394
rect 7172 22390 18918 22394
rect 7172 22340 12384 22390
rect 7172 22215 9455 22340
rect 2370 22161 9455 22215
rect 9654 22211 12384 22340
rect 12583 22211 13531 22390
rect 13730 22336 18918 22390
rect 13730 22211 16013 22336
rect 9654 22161 16013 22211
rect 2370 22157 16013 22161
rect 16212 22216 18918 22336
rect 19117 22216 20065 22395
rect 20264 22341 25431 22395
rect 20264 22216 22547 22341
rect 16212 22162 22547 22216
rect 22746 22219 25431 22341
rect 25630 22219 26578 22398
rect 26777 22344 36609 22398
rect 26777 22219 29060 22344
rect 22746 22165 29060 22219
rect 29259 22165 36609 22344
rect 22746 22162 36609 22165
rect 16212 22157 36609 22162
rect 2370 21955 36609 22157
rect 2370 21945 5863 21955
rect 2370 19450 3884 21945
rect 5376 20517 5863 21945
rect 8437 21943 36609 21955
rect 8919 21363 9429 21370
rect 9300 20690 10195 20904
rect 9300 20522 9441 20690
rect 6730 20517 7077 20520
rect 8955 20517 9441 20522
rect 5376 20511 9441 20517
rect 9640 20511 10195 20690
rect 5376 20347 10195 20511
rect 5376 20168 5730 20347
rect 5929 20168 7628 20347
rect 7827 20168 10195 20347
rect 5376 20012 10195 20168
rect 5376 20007 5863 20012
rect -4169 19448 3884 19450
rect -4203 16975 3884 19448
rect 10025 19282 10195 20012
rect 11805 20513 12421 21943
rect 15858 20686 16753 20900
rect 15858 20518 15999 20686
rect 13288 20513 13635 20516
rect 15513 20513 15999 20518
rect 11805 20507 15999 20513
rect 16198 20507 16753 20686
rect 11805 20343 16753 20507
rect 11805 20164 12288 20343
rect 12487 20164 14186 20343
rect 14385 20164 16753 20343
rect 11805 20008 16753 20164
rect 18339 20518 18955 21943
rect 22392 20691 23287 20905
rect 22392 20523 22533 20691
rect 19822 20518 20169 20521
rect 22047 20518 22533 20523
rect 18339 20512 22533 20518
rect 22732 20512 23287 20691
rect 18339 20348 23287 20512
rect 18339 20169 18822 20348
rect 19021 20169 20720 20348
rect 20919 20169 23287 20348
rect 18339 20013 23287 20169
rect 18339 20008 18955 20013
rect 11805 20003 12421 20008
rect 8927 19086 10195 19282
rect 16583 19278 16753 20008
rect 23117 19283 23287 20013
rect 24852 20521 25468 21943
rect 29273 21910 36609 21943
rect 30048 21908 36609 21910
rect 28905 20694 29800 20908
rect 28905 20526 29046 20694
rect 26335 20521 26682 20524
rect 28560 20521 29046 20526
rect 24852 20515 29046 20521
rect 29245 20515 29800 20694
rect 24852 20351 29800 20515
rect 24852 20172 25335 20351
rect 25534 20172 27233 20351
rect 27432 20172 29800 20351
rect 24852 20016 29800 20172
rect 24852 20011 25468 20016
rect 29630 19286 29800 20016
rect 8927 18907 9446 19086
rect 9645 18907 10195 19086
rect 8927 18638 10195 18907
rect 15485 19082 16753 19278
rect 15485 18903 16004 19082
rect 16203 18903 16753 19082
rect 15485 18634 16753 18903
rect 22019 19087 23287 19283
rect 22019 18908 22538 19087
rect 22737 18908 23287 19087
rect 22019 18639 23287 18908
rect 28532 19090 29800 19286
rect 28532 18911 29051 19090
rect 29250 18911 29800 19090
rect 28532 18642 29800 18911
rect 34612 20768 36609 21908
rect 38715 20845 38895 20908
rect 34612 20668 36485 20768
rect 36577 20668 36609 20768
rect 5764 17938 6009 17941
rect 5764 17920 5786 17938
rect 5985 17920 6009 17938
rect 7662 17938 7907 17941
rect 7662 17920 7684 17938
rect 7883 17920 7907 17938
rect 6141 17616 7477 17802
rect 7987 17616 8011 17853
rect 12322 17934 12567 17937
rect 12322 17916 12344 17934
rect 12543 17916 12567 17934
rect 14220 17934 14465 17937
rect 14220 17916 14242 17934
rect 14441 17916 14465 17934
rect 5644 17611 8011 17616
rect 12699 17612 14035 17798
rect 14545 17612 14569 17849
rect 18856 17939 19101 17942
rect 18856 17921 18878 17939
rect 19077 17921 19101 17939
rect 20754 17939 20999 17942
rect 20754 17921 20776 17939
rect 20975 17921 20999 17939
rect 19233 17617 20569 17803
rect 21079 17617 21103 17854
rect 25369 17942 25614 17945
rect 25369 17924 25391 17942
rect 25590 17924 25614 17942
rect 27267 17942 27512 17945
rect 27267 17924 27289 17942
rect 27488 17924 27512 17942
rect 25746 17620 27082 17806
rect 27592 17620 27616 17857
rect 18736 17612 21103 17617
rect 25249 17615 27616 17620
rect 34612 17636 36609 20668
rect 38715 20459 38895 20514
rect 38715 17712 38895 17775
rect 25557 17613 27228 17615
rect 5952 17609 7623 17611
rect 12202 17607 14569 17612
rect 19044 17610 20715 17612
rect 12510 17605 14181 17607
rect -4203 16123 -3727 16975
rect -4201 15440 -3957 16123
rect -4201 15364 -4065 15440
rect -3999 15364 -3957 15440
rect -4201 13372 -3957 15364
rect 2370 15647 3884 16975
rect 34612 17536 36481 17636
rect 36573 17536 36609 17636
rect 34612 15655 36609 17536
rect 38715 17371 38895 17381
rect 32684 15654 36609 15655
rect 29281 15653 36609 15654
rect 2363 15646 8015 15647
rect 14414 15646 36609 15653
rect 2363 15486 36609 15646
rect 2363 15466 21350 15486
rect 2363 15394 8147 15466
rect 8217 15465 21350 15466
rect 8217 15394 14696 15465
rect 2363 15393 14696 15394
rect 14766 15414 21350 15465
rect 21420 15414 36609 15486
rect 14766 15393 36609 15414
rect 2363 15355 36609 15393
rect 2363 15348 22915 15355
rect 2363 15347 8015 15348
rect -1849 15245 -1659 15281
rect 2363 13726 2769 15347
rect 29068 15319 36609 15355
rect 29068 15247 30003 15319
rect 30073 15286 36609 15319
rect 30073 15247 32233 15286
rect 29068 15195 32233 15247
rect 8681 14161 8682 14369
rect 14713 14345 15223 14346
rect 14713 14164 14714 14345
rect 21380 14153 21381 14329
rect 8676 13727 12233 13759
rect 14989 13732 18546 13759
rect 21824 13732 25381 13759
rect 29068 13739 29535 15195
rect 32091 15192 32233 15195
rect 32211 15107 32233 15192
rect 32432 15193 36609 15286
rect 32432 15192 32560 15193
rect 32432 15107 32456 15192
rect 32211 15104 32456 15107
rect 33444 14911 33830 15193
rect 33444 14870 33604 14911
rect 33446 14839 33604 14870
rect 33674 14870 33830 14911
rect 33674 14839 33828 14870
rect 33446 14817 33828 14839
rect 34173 14492 36609 15193
rect 34173 14392 36481 14492
rect 36573 14392 36609 14492
rect 30442 13985 30443 14156
rect 28443 13732 29535 13739
rect 33698 13734 33754 13735
rect 14989 13727 29535 13732
rect 1247 13722 5404 13726
rect 8676 13722 29535 13727
rect -1851 13589 -1659 13595
rect -4201 13296 -4067 13372
rect -4001 13296 -3957 13372
rect -4201 11303 -3957 13296
rect 1247 13566 29535 13722
rect 1247 13494 1483 13566
rect 1553 13539 29535 13566
rect 1553 13494 13477 13539
rect 1247 13485 13477 13494
rect 1247 13472 10995 13485
rect 2368 13451 10995 13472
rect 2368 13397 6928 13451
rect 2368 13218 4446 13397
rect 4645 13272 6928 13397
rect 7127 13272 8075 13451
rect 8274 13306 10995 13451
rect 11194 13360 13477 13485
rect 13676 13360 14624 13539
rect 14823 13485 26756 13539
rect 14823 13471 24274 13485
rect 14823 13417 20131 13471
rect 14823 13360 17649 13417
rect 11194 13306 17649 13360
rect 8274 13272 17649 13306
rect 4645 13238 17649 13272
rect 17848 13292 20131 13417
rect 20330 13292 21278 13471
rect 21477 13306 24274 13471
rect 24473 13360 26756 13485
rect 26955 13360 27903 13539
rect 28102 13360 29535 13539
rect 33694 13733 33754 13734
rect 33991 13734 34030 13735
rect 33991 13733 34045 13734
rect 33694 13617 33699 13733
rect 34037 13617 34045 13733
rect 33694 13476 33754 13617
rect 24473 13306 29535 13360
rect 33991 13476 34045 13617
rect 21477 13292 29535 13306
rect 17848 13238 29535 13292
rect 4645 13218 29535 13238
rect -1851 13105 -1659 13187
rect 2368 13100 29535 13218
rect 2368 13099 12233 13100
rect 14786 13099 25381 13100
rect 2368 13012 8853 13099
rect 2368 12997 6262 13012
rect -1849 11521 -1659 11553
rect -4201 11227 -4065 11303
rect -3999 11227 -3957 11303
rect -4201 9235 -3957 11227
rect 2368 11128 3046 12997
rect -1849 11088 -1659 11119
rect 1234 10981 3046 11128
rect 1234 10909 1475 10981
rect 1545 10909 3046 10981
rect 1234 10887 3046 10909
rect -1851 9458 -1659 9572
rect -4201 9159 -4067 9235
rect -4001 9159 -3957 9235
rect -4201 7166 -3957 9159
rect -1851 9010 -1659 9056
rect 2368 7873 3046 10887
rect 3905 11747 4800 11961
rect 3905 11568 4460 11747
rect 4659 11579 4800 11747
rect 4659 11574 5145 11579
rect 7023 11574 7370 11577
rect 8237 11574 8853 13012
rect 4659 11568 8853 11574
rect 3905 11404 8853 11568
rect 3905 11225 6273 11404
rect 6472 11225 8171 11404
rect 8370 11225 8853 11404
rect 3905 11069 8853 11225
rect 3905 10339 4075 11069
rect 8237 11064 8853 11069
rect 10454 11835 11349 12049
rect 10454 11656 11009 11835
rect 11208 11667 11349 11835
rect 11208 11662 11694 11667
rect 13572 11662 13919 11665
rect 14786 11662 15402 13099
rect 17628 13032 22056 13099
rect 11208 11656 15402 11662
rect 10454 11492 15402 11656
rect 10454 11313 12822 11492
rect 13021 11313 14720 11492
rect 14919 11313 15402 11492
rect 10454 11157 15402 11313
rect 10454 10427 10624 11157
rect 14786 11152 15402 11157
rect 17108 11767 18003 11981
rect 17108 11588 17663 11767
rect 17862 11599 18003 11767
rect 17862 11594 18348 11599
rect 20226 11594 20573 11597
rect 21440 11594 22056 13032
rect 28065 13077 29535 13100
rect 17862 11588 22056 11594
rect 17108 11424 22056 11588
rect 17108 11245 19476 11424
rect 19675 11245 21374 11424
rect 21573 11245 22056 11424
rect 17108 11089 22056 11245
rect 3905 10143 5173 10339
rect 3905 9964 4455 10143
rect 4654 9964 5173 10143
rect 3905 9695 5173 9964
rect 10454 10231 11722 10427
rect 10454 10052 11004 10231
rect 11203 10052 11722 10231
rect 10454 9783 11722 10052
rect 17108 10359 17278 11089
rect 21440 11084 22056 11089
rect 23733 11835 24628 12049
rect 23733 11656 24288 11835
rect 24487 11667 24628 11835
rect 24487 11662 24973 11667
rect 26851 11662 27198 11665
rect 28065 11662 28681 13077
rect 24487 11656 28681 11662
rect 23733 11492 28681 11656
rect 23733 11313 26101 11492
rect 26300 11313 27999 11492
rect 28198 11313 28681 11492
rect 23733 11157 28681 11313
rect 23733 10427 23903 11157
rect 28065 11152 28681 11157
rect 29068 12846 29535 13077
rect 29068 12748 30550 12846
rect 29068 12676 29998 12748
rect 30068 12676 30550 12748
rect 29068 12608 30550 12676
rect 17108 10163 18376 10359
rect 17108 9984 17658 10163
rect 17857 9984 18376 10163
rect 17108 9715 18376 9984
rect 23733 10231 25001 10427
rect 23733 10052 24283 10231
rect 24482 10052 25001 10231
rect 23733 9783 25001 10052
rect 29068 9830 29535 12608
rect 30088 11593 30447 11595
rect 31976 11360 33329 11371
rect 34173 11360 36609 14392
rect 38715 14243 38895 14263
rect 38715 11403 38895 11436
rect 31976 11290 36609 11360
rect 31976 11195 36485 11290
rect 31976 11101 32235 11195
rect 32213 11016 32235 11101
rect 32434 11190 36485 11195
rect 36577 11190 36609 11290
rect 32434 11101 36609 11190
rect 32434 11016 32458 11101
rect 33131 11099 36609 11101
rect 32213 11013 32458 11016
rect 33446 10820 33832 11099
rect 33446 10779 33606 10820
rect 33448 10748 33606 10779
rect 33676 10779 33832 10820
rect 33676 10748 33830 10779
rect 33448 10726 33830 10748
rect 29068 9715 30553 9830
rect 29068 9643 29998 9715
rect 30068 9643 30553 9715
rect 33700 9643 33756 9644
rect 29068 9592 30553 9643
rect 33696 9642 33756 9643
rect 33993 9643 34032 9644
rect 33993 9642 34047 9643
rect 6193 8995 6438 8998
rect 6193 8977 6217 8995
rect 6416 8977 6438 8995
rect 8091 8995 8336 8998
rect 8091 8977 8115 8995
rect 8314 8977 8336 8995
rect 12742 9083 12987 9086
rect 12742 9065 12766 9083
rect 12965 9065 12987 9083
rect 14640 9083 14885 9086
rect 14640 9065 14664 9083
rect 14863 9065 14885 9083
rect 6089 8673 6113 8910
rect 6623 8673 7959 8859
rect 12638 8761 12662 8998
rect 13172 8761 14508 8947
rect 19396 9015 19641 9018
rect 19396 8997 19420 9015
rect 19619 8997 19641 9015
rect 21294 9015 21539 9018
rect 21294 8997 21318 9015
rect 21517 8997 21539 9015
rect 12638 8756 15005 8761
rect 13026 8754 14697 8756
rect 19292 8693 19316 8930
rect 19826 8693 21162 8879
rect 26021 9083 26266 9086
rect 26021 9065 26045 9083
rect 26244 9065 26266 9083
rect 27919 9083 28164 9086
rect 27919 9065 27943 9083
rect 28142 9065 28164 9083
rect 25917 8761 25941 8998
rect 26451 8761 27787 8947
rect 25917 8756 28284 8761
rect 26305 8754 27976 8756
rect 19292 8688 21659 8693
rect 19680 8686 21351 8688
rect 6089 8668 8456 8673
rect 6477 8666 8148 8668
rect 29068 8135 29535 9592
rect 33696 9526 33701 9642
rect 34039 9526 34047 9642
rect 33696 9385 33756 9526
rect 33993 9385 34047 9526
rect 30089 8555 30450 8557
rect 30088 8400 30089 8555
rect 30449 8397 30450 8555
rect 34173 8146 36609 11099
rect 38715 11067 38895 11072
rect 38715 8237 38895 8255
rect 34173 8138 36485 8146
rect 33354 8135 36485 8138
rect 29068 8046 36485 8135
rect 36577 8046 36609 8146
rect 10967 7873 15400 7879
rect 17622 7873 22055 7887
rect 24244 7873 28677 7889
rect 29068 7873 36609 8046
rect 2368 7832 36609 7873
rect 1227 7795 36609 7832
rect 1227 7723 30069 7795
rect 30139 7723 36609 7795
rect 1227 7703 36609 7723
rect 1227 7631 1456 7703
rect 1526 7700 36609 7703
rect 1526 7671 32235 7700
rect 1526 7631 6920 7671
rect 1227 7617 6920 7631
rect 1227 7591 4438 7617
rect 2368 7438 4438 7591
rect 4637 7492 6920 7617
rect 7119 7492 8067 7671
rect 8266 7670 26748 7671
rect 8266 7669 20126 7670
rect 8266 7615 13471 7669
rect 8266 7492 10989 7615
rect 4637 7438 10989 7492
rect 2368 7436 10989 7438
rect 11188 7490 13471 7615
rect 13670 7490 14618 7669
rect 14817 7616 20126 7669
rect 14817 7490 17644 7616
rect 11188 7437 17644 7490
rect 17843 7491 20126 7616
rect 20325 7491 21273 7670
rect 21472 7617 26748 7670
rect 21472 7491 24266 7617
rect 17843 7438 24266 7491
rect 24465 7492 26748 7617
rect 26947 7492 27895 7671
rect 28094 7598 32235 7671
rect 28094 7492 29535 7598
rect 32213 7521 32235 7598
rect 32434 7598 36609 7700
rect 32434 7521 32458 7598
rect 33354 7593 36609 7598
rect 32213 7518 32458 7521
rect 24465 7438 29535 7492
rect 17843 7437 29535 7438
rect 11188 7436 29535 7437
rect -1851 7359 -1659 7411
rect -4201 7090 -4067 7166
rect -4001 7090 -3957 7166
rect -4201 5098 -3957 7090
rect 2368 7210 29535 7436
rect 33446 7325 33832 7593
rect 33446 7284 33606 7325
rect 33448 7253 33606 7284
rect 33676 7284 33832 7325
rect 33676 7253 33830 7284
rect 33448 7231 33830 7253
rect -1851 6906 -1659 6957
rect -1853 5296 -1659 5384
rect -4201 5022 -4069 5098
rect -4003 5022 -3957 5098
rect -4201 3029 -3957 5022
rect 2368 5075 3046 7210
rect 1221 4943 3046 5075
rect -1853 4770 -1659 4894
rect 1221 4871 1472 4943
rect 1542 4871 3046 4943
rect 1221 4834 3046 4871
rect -1851 3254 -1659 3285
rect -4201 2953 -4067 3029
rect -4001 2953 -3957 3029
rect -4201 961 -3957 2953
rect -1851 2718 -1659 2852
rect 2368 1219 3046 4834
rect 3897 5967 4792 6181
rect 3897 5788 4452 5967
rect 4651 5799 4792 5967
rect 4651 5794 5137 5799
rect 7015 5794 7362 5797
rect 8229 5794 8845 7210
rect 4651 5788 8845 5794
rect 3897 5624 8845 5788
rect 3897 5445 6265 5624
rect 6464 5445 8163 5624
rect 8362 5445 8845 5624
rect 3897 5289 8845 5445
rect 3897 4559 4067 5289
rect 8229 5284 8845 5289
rect 10448 5965 11343 6179
rect 10448 5786 11003 5965
rect 11202 5797 11343 5965
rect 11202 5792 11688 5797
rect 13566 5792 13913 5795
rect 14780 5792 15396 7210
rect 11202 5786 15396 5792
rect 10448 5622 15396 5786
rect 10448 5443 12816 5622
rect 13015 5443 14714 5622
rect 14913 5443 15396 5622
rect 10448 5287 15396 5443
rect 3897 4363 5165 4559
rect 3897 4184 4447 4363
rect 4646 4184 5165 4363
rect 3897 3915 5165 4184
rect 10448 4557 10618 5287
rect 14780 5282 15396 5287
rect 17103 5966 17998 6180
rect 17103 5787 17658 5966
rect 17857 5798 17998 5966
rect 17857 5793 18343 5798
rect 20221 5793 20568 5796
rect 21435 5793 22051 7210
rect 17857 5787 22051 5793
rect 17103 5623 22051 5787
rect 17103 5444 19471 5623
rect 19670 5444 21369 5623
rect 21568 5444 22051 5623
rect 17103 5288 22051 5444
rect 17103 4558 17273 5288
rect 21435 5283 22051 5288
rect 23725 5967 24620 6181
rect 23725 5788 24280 5967
rect 24479 5799 24620 5967
rect 24479 5794 24965 5799
rect 26843 5794 27190 5797
rect 28057 5794 28673 7210
rect 24479 5788 28673 5794
rect 23725 5624 28673 5788
rect 23725 5445 26093 5624
rect 26292 5445 27991 5624
rect 28190 5445 28673 5624
rect 23725 5289 28673 5445
rect 23725 4559 23895 5289
rect 28057 5284 28673 5289
rect 29068 4818 29535 7210
rect 30149 6634 30512 6635
rect 30509 6474 30512 6634
rect 33700 6148 33756 6149
rect 33696 6147 33756 6148
rect 33993 6148 34032 6149
rect 33993 6147 34047 6148
rect 33696 6031 33701 6147
rect 34039 6031 34047 6147
rect 33696 5890 33756 6031
rect 33993 5890 34047 6031
rect 32093 5018 32466 5088
rect 34173 5014 36609 7593
rect 38715 5094 38895 5137
rect 34173 4914 36481 5014
rect 36573 4914 36609 5014
rect 29068 4725 30553 4818
rect 29068 4653 30066 4725
rect 30136 4653 30553 4725
rect 29068 4580 30553 4653
rect 10448 4361 11716 4557
rect 10448 4182 10998 4361
rect 11197 4182 11716 4361
rect 10448 3913 11716 4182
rect 17103 4362 18371 4558
rect 17103 4183 17653 4362
rect 17852 4183 18371 4362
rect 17103 3914 18371 4183
rect 23725 4363 24993 4559
rect 23725 4184 24275 4363
rect 24474 4184 24993 4363
rect 23725 3915 24993 4184
rect 6185 3215 6430 3218
rect 6185 3197 6209 3215
rect 6408 3197 6430 3215
rect 8083 3215 8328 3218
rect 8083 3197 8107 3215
rect 8306 3197 8328 3215
rect 6081 2893 6105 3130
rect 6615 2893 7951 3079
rect 12736 3213 12981 3216
rect 12736 3195 12760 3213
rect 12959 3195 12981 3213
rect 14634 3213 14879 3216
rect 14634 3195 14658 3213
rect 14857 3195 14879 3213
rect 6081 2888 8448 2893
rect 12632 2891 12656 3128
rect 13166 2891 14502 3077
rect 19391 3214 19636 3217
rect 19391 3196 19415 3214
rect 19614 3196 19636 3214
rect 21289 3214 21534 3217
rect 21289 3196 21313 3214
rect 21512 3196 21534 3214
rect 19287 2892 19311 3129
rect 19821 2892 21157 3078
rect 26013 3215 26258 3218
rect 26013 3197 26037 3215
rect 26236 3197 26258 3215
rect 27911 3215 28156 3218
rect 27911 3197 27935 3215
rect 28134 3197 28156 3215
rect 25909 2893 25933 3130
rect 26443 2893 27779 3079
rect 6469 2886 8140 2888
rect 12632 2886 14999 2891
rect 19287 2887 21654 2892
rect 25909 2888 28276 2893
rect 13020 2884 14691 2886
rect 19675 2885 21346 2887
rect 26297 2886 27968 2888
rect 29068 2006 29535 4580
rect 30144 3566 30506 3567
rect 30144 3392 30145 3566
rect 30505 3392 30506 3566
rect 32502 3501 33640 3503
rect 34173 3501 36609 4914
rect 38715 4756 38895 4763
rect 32502 3500 36609 3501
rect 32028 3352 36609 3500
rect 32028 3254 32235 3352
rect 32213 3173 32235 3254
rect 32434 3259 36609 3352
rect 32434 3254 32885 3259
rect 33446 3257 36609 3259
rect 32434 3173 32458 3254
rect 32213 3170 32458 3173
rect 33446 2977 33832 3257
rect 34612 3248 36609 3257
rect 33446 2936 33606 2977
rect 33448 2905 33606 2936
rect 33676 2936 33832 2977
rect 33676 2905 33830 2936
rect 33448 2883 33830 2905
rect 29068 1880 30547 2006
rect 29068 1808 30073 1880
rect 30143 1808 30547 1880
rect 36375 1870 36609 3248
rect 38715 1976 38895 2004
rect 29068 1768 30547 1808
rect 33700 1800 33756 1801
rect 33696 1799 33756 1800
rect 33993 1800 34032 1801
rect 33993 1799 34047 1800
rect 29068 1219 29535 1768
rect 33696 1683 33701 1799
rect 34039 1683 34047 1799
rect 33696 1542 33756 1683
rect 33993 1542 34047 1683
rect 36375 1770 36481 1870
rect 36573 1770 36609 1870
rect -1853 1165 -1659 1201
rect 2363 1179 29537 1219
rect 2363 1174 14736 1179
rect -4201 885 -4069 961
rect -4003 885 -3957 961
rect -4201 46 -3957 885
rect 2363 1102 8182 1174
rect 8252 1107 14736 1174
rect 14806 1167 29537 1179
rect 14806 1107 21385 1167
rect 8252 1102 21385 1107
rect 2363 1095 21385 1102
rect 21455 1095 29537 1167
rect 2363 965 29537 1095
rect 36375 838 36609 1770
rect 30154 555 30155 713
rect 30515 555 30516 713
<< via4 >>
rect 6475 26900 6985 26978
rect 6475 26701 6534 26900
rect 6534 26701 6713 26900
rect 6713 26701 6985 26900
rect 6475 26674 6985 26701
rect 8043 26589 8347 26740
rect 8043 26410 8077 26589
rect 8077 26410 8276 26589
rect 8276 26410 8347 26589
rect 8043 26230 8347 26410
rect 9177 26587 9481 26750
rect 9177 26408 9219 26587
rect 9219 26408 9418 26587
rect 9418 26408 9481 26587
rect 9177 26240 9481 26408
rect 12988 26897 13498 26975
rect 12988 26698 13047 26897
rect 13047 26698 13226 26897
rect 13226 26698 13498 26897
rect 12988 26671 13498 26698
rect 14556 26586 14860 26737
rect 14556 26407 14590 26586
rect 14590 26407 14789 26586
rect 14789 26407 14860 26586
rect 14556 26227 14860 26407
rect 15690 26584 15994 26747
rect 15690 26405 15732 26584
rect 15732 26405 15931 26584
rect 15931 26405 15994 26584
rect 15690 26237 15994 26405
rect 19522 26892 20032 26970
rect 19522 26693 19581 26892
rect 19581 26693 19760 26892
rect 19760 26693 20032 26892
rect 19522 26666 20032 26693
rect 21090 26581 21394 26732
rect 6469 25250 6979 25318
rect 6469 25051 6548 25250
rect 6548 25051 6727 25250
rect 6727 25051 6979 25250
rect 6469 25014 6979 25051
rect 21090 26402 21124 26581
rect 21124 26402 21323 26581
rect 21323 26402 21394 26581
rect 21090 26222 21394 26402
rect 22224 26579 22528 26742
rect 22224 26400 22266 26579
rect 22266 26400 22465 26579
rect 22465 26400 22528 26579
rect 22224 26232 22528 26400
rect 26080 26896 26590 26974
rect 26080 26697 26139 26896
rect 26139 26697 26318 26896
rect 26318 26697 26590 26896
rect 26080 26670 26590 26697
rect 27648 26585 27952 26736
rect 12982 25247 13492 25315
rect 12982 25048 13061 25247
rect 13061 25048 13240 25247
rect 13240 25048 13492 25247
rect 12982 25011 13492 25048
rect 27648 26406 27682 26585
rect 27682 26406 27881 26585
rect 27881 26406 27952 26585
rect 27648 26226 27952 26406
rect 28782 26583 29086 26746
rect 28782 26404 28824 26583
rect 28824 26404 29023 26583
rect 29023 26404 29086 26583
rect 28782 26236 29086 26404
rect 19516 25242 20026 25310
rect 19516 25043 19595 25242
rect 19595 25043 19774 25242
rect 19774 25043 20026 25242
rect 19516 25006 20026 25043
rect 26074 25246 26584 25314
rect 26074 25047 26153 25246
rect 26153 25047 26332 25246
rect 26332 25047 26584 25246
rect 26074 25010 26584 25047
rect 6468 23646 6978 23713
rect 6468 23447 6543 23646
rect 6543 23447 6722 23646
rect 6722 23447 6978 23646
rect 12981 23643 13491 23710
rect 6468 23409 6978 23447
rect 7917 23367 8021 23528
rect 8021 23367 8220 23528
rect 8220 23367 8427 23528
rect 7917 23224 8427 23367
rect 9763 23367 9919 23528
rect 9919 23367 10118 23528
rect 10118 23367 10273 23528
rect 12981 23444 13056 23643
rect 13056 23444 13235 23643
rect 13235 23444 13491 23643
rect 19515 23638 20025 23705
rect 12981 23406 13491 23444
rect 9763 23224 10273 23367
rect 14430 23364 14534 23525
rect 14534 23364 14733 23525
rect 14733 23364 14940 23525
rect 14430 23221 14940 23364
rect 16276 23364 16432 23525
rect 16432 23364 16631 23525
rect 16631 23364 16786 23525
rect 19515 23439 19590 23638
rect 19590 23439 19769 23638
rect 19769 23439 20025 23638
rect 26073 23642 26583 23709
rect 19515 23401 20025 23439
rect 16276 23221 16786 23364
rect 20964 23359 21068 23520
rect 21068 23359 21267 23520
rect 21267 23359 21474 23520
rect 20964 23216 21474 23359
rect 22810 23359 22966 23520
rect 22966 23359 23165 23520
rect 23165 23359 23320 23520
rect 26073 23443 26148 23642
rect 26148 23443 26327 23642
rect 26327 23443 26583 23642
rect 26073 23405 26583 23443
rect 22810 23216 23320 23359
rect 27522 23363 27626 23524
rect 27626 23363 27825 23524
rect 27825 23363 28032 23524
rect 27522 23220 28032 23363
rect 29368 23363 29524 23524
rect 29524 23363 29723 23524
rect 29723 23363 29878 23524
rect 29368 23220 29878 23363
rect 38705 23898 38949 24003
rect 38705 23814 38727 23898
rect 38727 23814 38795 23898
rect 38795 23814 38949 23898
rect 38705 23672 38949 23814
rect 8919 21292 9429 21363
rect 6423 20979 6727 21142
rect 6423 20800 6486 20979
rect 6486 20800 6685 20979
rect 6685 20800 6727 20979
rect 6423 20632 6727 20800
rect 7557 20981 7861 21132
rect 8919 21093 9191 21292
rect 9191 21093 9370 21292
rect 9370 21093 9429 21292
rect 8919 21066 9429 21093
rect 7557 20802 7628 20981
rect 7628 20802 7827 20981
rect 7827 20802 7861 20981
rect 7557 20622 7861 20802
rect 8925 19642 9435 19710
rect 8925 19443 9177 19642
rect 9177 19443 9356 19642
rect 9356 19443 9435 19642
rect 8925 19406 9435 19443
rect 15477 21288 15987 21366
rect 12981 20975 13285 21138
rect 12981 20796 13044 20975
rect 13044 20796 13243 20975
rect 13243 20796 13285 20975
rect 12981 20628 13285 20796
rect 14115 20977 14419 21128
rect 15477 21089 15749 21288
rect 15749 21089 15928 21288
rect 15928 21089 15987 21288
rect 15477 21062 15987 21089
rect 14115 20798 14186 20977
rect 14186 20798 14385 20977
rect 14385 20798 14419 20977
rect 14115 20618 14419 20798
rect 22011 21293 22521 21371
rect 19515 20980 19819 21143
rect 19515 20801 19578 20980
rect 19578 20801 19777 20980
rect 19777 20801 19819 20980
rect 19515 20633 19819 20801
rect 20649 20982 20953 21133
rect 22011 21094 22283 21293
rect 22283 21094 22462 21293
rect 22462 21094 22521 21293
rect 22011 21067 22521 21094
rect 20649 20803 20720 20982
rect 20720 20803 20919 20982
rect 20919 20803 20953 20982
rect 20649 20623 20953 20803
rect 15483 19638 15993 19706
rect 15483 19439 15735 19638
rect 15735 19439 15914 19638
rect 15914 19439 15993 19638
rect 15483 19402 15993 19439
rect 22017 19643 22527 19711
rect 22017 19444 22269 19643
rect 22269 19444 22448 19643
rect 22448 19444 22527 19643
rect 22017 19407 22527 19444
rect 28524 21296 29034 21374
rect 26028 20983 26332 21146
rect 26028 20804 26091 20983
rect 26091 20804 26290 20983
rect 26290 20804 26332 20983
rect 26028 20636 26332 20804
rect 27162 20985 27466 21136
rect 28524 21097 28796 21296
rect 28796 21097 28975 21296
rect 28975 21097 29034 21296
rect 28524 21070 29034 21097
rect 27162 20806 27233 20985
rect 27233 20806 27432 20985
rect 27432 20806 27466 20985
rect 27162 20626 27466 20806
rect 28530 19646 29040 19714
rect 28530 19447 28782 19646
rect 28782 19447 28961 19646
rect 28961 19447 29040 19646
rect 28530 19410 29040 19447
rect 8926 18038 9436 18105
rect 5631 17759 5786 17920
rect 5786 17759 5985 17920
rect 5985 17759 6141 17920
rect 5631 17616 6141 17759
rect 7477 17759 7684 17920
rect 7684 17759 7883 17920
rect 7883 17759 7987 17920
rect 7477 17616 7987 17759
rect 8926 17839 9182 18038
rect 9182 17839 9361 18038
rect 9361 17839 9436 18038
rect 15484 18034 15994 18101
rect 8926 17801 9436 17839
rect 12189 17755 12344 17916
rect 12344 17755 12543 17916
rect 12543 17755 12699 17916
rect 12189 17612 12699 17755
rect 14035 17755 14242 17916
rect 14242 17755 14441 17916
rect 14441 17755 14545 17916
rect 14035 17612 14545 17755
rect 15484 17835 15740 18034
rect 15740 17835 15919 18034
rect 15919 17835 15994 18034
rect 22018 18039 22528 18106
rect 15484 17797 15994 17835
rect 18723 17760 18878 17921
rect 18878 17760 19077 17921
rect 19077 17760 19233 17921
rect 18723 17617 19233 17760
rect 20569 17760 20776 17921
rect 20776 17760 20975 17921
rect 20975 17760 21079 17921
rect 20569 17617 21079 17760
rect 22018 17840 22274 18039
rect 22274 17840 22453 18039
rect 22453 17840 22528 18039
rect 28531 18042 29041 18109
rect 22018 17802 22528 17840
rect 25236 17763 25391 17924
rect 25391 17763 25590 17924
rect 25590 17763 25746 17924
rect 25236 17620 25746 17763
rect 27082 17763 27289 17924
rect 27289 17763 27488 17924
rect 27488 17763 27592 17924
rect 27082 17620 27592 17763
rect 28531 17843 28787 18042
rect 28787 17843 28966 18042
rect 28966 17843 29041 18042
rect 28531 17805 29041 17843
rect 38707 20754 38951 20845
rect 38707 20670 38727 20754
rect 38727 20670 38795 20754
rect 38795 20670 38951 20754
rect 38707 20514 38951 20670
rect -1878 15502 -1455 15683
rect 38705 17622 38949 17712
rect 38705 17538 38723 17622
rect 38723 17538 38791 17622
rect 38791 17538 38949 17622
rect 38705 17381 38949 17538
rect -1878 15408 -1843 15502
rect -1843 15408 -1755 15502
rect -1755 15408 -1455 15502
rect -1878 15281 -1455 15408
rect 8172 14262 8681 14370
rect 8172 14194 8369 14262
rect 8369 14194 8443 14262
rect 8443 14194 8681 14262
rect 8172 14062 8681 14194
rect 14714 14261 15223 14345
rect 14714 14193 14918 14261
rect 14918 14193 14992 14261
rect 14992 14193 15223 14261
rect 14714 14037 15223 14193
rect 21381 14282 21890 14330
rect 21381 14214 21572 14282
rect 21572 14214 21646 14282
rect 21646 14214 21890 14282
rect 21381 14023 21890 14214
rect 30082 14115 30442 14156
rect 30082 14047 30225 14115
rect 30225 14047 30299 14115
rect 30299 14047 30442 14115
rect 30082 13883 30442 14047
rect -1883 13434 -1460 13589
rect -1883 13340 -1845 13434
rect -1845 13340 -1757 13434
rect -1757 13340 -1460 13434
rect -1883 13187 -1460 13340
rect 33754 13733 33991 13792
rect 33754 13617 33991 13733
rect 33754 13335 33991 13617
rect 1509 12362 2017 12432
rect 1509 12294 1705 12362
rect 1705 12294 1779 12362
rect 1779 12294 2017 12362
rect 1509 12124 2017 12294
rect -1893 11365 -1470 11521
rect -1893 11271 -1843 11365
rect -1843 11271 -1755 11365
rect -1755 11271 -1470 11365
rect -1893 11119 -1470 11271
rect 4671 12349 5181 12427
rect 4671 12150 4730 12349
rect 4730 12150 4909 12349
rect 4909 12150 5181 12349
rect 4671 12123 5181 12150
rect 6239 12038 6543 12189
rect 1484 9777 1992 9850
rect 1484 9709 1697 9777
rect 1697 9709 1771 9777
rect 1771 9709 1992 9777
rect 1484 9542 1992 9709
rect -1867 9297 -1444 9458
rect -1867 9203 -1845 9297
rect -1845 9203 -1757 9297
rect -1757 9203 -1444 9297
rect -1867 9056 -1444 9203
rect 6239 11859 6273 12038
rect 6273 11859 6472 12038
rect 6472 11859 6543 12038
rect 6239 11679 6543 11859
rect 7373 12036 7677 12199
rect 7373 11857 7415 12036
rect 7415 11857 7614 12036
rect 7614 11857 7677 12036
rect 7373 11689 7677 11857
rect 11220 12437 11730 12515
rect 11220 12238 11279 12437
rect 11279 12238 11458 12437
rect 11458 12238 11730 12437
rect 11220 12211 11730 12238
rect 12788 12126 13092 12277
rect 12788 11947 12822 12126
rect 12822 11947 13021 12126
rect 13021 11947 13092 12126
rect 12788 11767 13092 11947
rect 13922 12124 14226 12287
rect 13922 11945 13964 12124
rect 13964 11945 14163 12124
rect 14163 11945 14226 12124
rect 13922 11777 14226 11945
rect 17874 12369 18384 12447
rect 17874 12170 17933 12369
rect 17933 12170 18112 12369
rect 18112 12170 18384 12369
rect 17874 12143 18384 12170
rect 19442 12058 19746 12209
rect 4665 10699 5175 10767
rect 4665 10500 4744 10699
rect 4744 10500 4923 10699
rect 4923 10500 5175 10699
rect 4665 10463 5175 10500
rect 19442 11879 19476 12058
rect 19476 11879 19675 12058
rect 19675 11879 19746 12058
rect 19442 11699 19746 11879
rect 20576 12056 20880 12219
rect 20576 11877 20618 12056
rect 20618 11877 20817 12056
rect 20817 11877 20880 12056
rect 20576 11709 20880 11877
rect 24499 12437 25009 12515
rect 24499 12238 24558 12437
rect 24558 12238 24737 12437
rect 24737 12238 25009 12437
rect 24499 12211 25009 12238
rect 26067 12126 26371 12277
rect 11214 10787 11724 10855
rect 11214 10588 11293 10787
rect 11293 10588 11472 10787
rect 11472 10588 11724 10787
rect 11214 10551 11724 10588
rect 26067 11947 26101 12126
rect 26101 11947 26300 12126
rect 26300 11947 26371 12126
rect 26067 11767 26371 11947
rect 27201 12124 27505 12287
rect 27201 11945 27243 12124
rect 27243 11945 27442 12124
rect 27442 11945 27505 12124
rect 27201 11777 27505 11945
rect 17868 10719 18378 10787
rect 17868 10520 17947 10719
rect 17947 10520 18126 10719
rect 18126 10520 18378 10719
rect 17868 10483 18378 10520
rect 32091 12941 32464 12943
rect 32091 12746 32154 12941
rect 32154 12746 32420 12941
rect 32420 12746 32464 12941
rect 24493 10787 25003 10855
rect 24493 10588 24572 10787
rect 24572 10588 24751 10787
rect 24751 10588 25003 10787
rect 24493 10551 25003 10588
rect 32091 12604 32464 12746
rect 30088 11544 30448 11593
rect 30088 11476 30220 11544
rect 30220 11476 30294 11544
rect 30294 11476 30448 11544
rect 30088 11320 30448 11476
rect 38707 14478 38951 14594
rect 38707 14394 38723 14478
rect 38723 14394 38791 14478
rect 38791 14394 38951 14478
rect 38707 14263 38951 14394
rect 33756 9642 33993 9701
rect 11213 9183 11723 9250
rect 4664 9095 5174 9162
rect 4664 8896 4739 9095
rect 4739 8896 4918 9095
rect 4918 8896 5174 9095
rect 11213 8984 11288 9183
rect 11288 8984 11467 9183
rect 11467 8984 11723 9183
rect 24492 9183 25002 9250
rect 17867 9115 18377 9182
rect 4664 8858 5174 8896
rect 6113 8816 6217 8977
rect 6217 8816 6416 8977
rect 6416 8816 6623 8977
rect 6113 8673 6623 8816
rect 7959 8816 8115 8977
rect 8115 8816 8314 8977
rect 8314 8816 8469 8977
rect 11213 8946 11723 8984
rect 7959 8673 8469 8816
rect 12662 8904 12766 9065
rect 12766 8904 12965 9065
rect 12965 8904 13172 9065
rect 12662 8761 13172 8904
rect 14508 8904 14664 9065
rect 14664 8904 14863 9065
rect 14863 8904 15018 9065
rect 14508 8761 15018 8904
rect 17867 8916 17942 9115
rect 17942 8916 18121 9115
rect 18121 8916 18377 9115
rect 17867 8878 18377 8916
rect 19316 8836 19420 8997
rect 19420 8836 19619 8997
rect 19619 8836 19826 8997
rect 19316 8693 19826 8836
rect 21162 8836 21318 8997
rect 21318 8836 21517 8997
rect 21517 8836 21672 8997
rect 24492 8984 24567 9183
rect 24567 8984 24746 9183
rect 24746 8984 25002 9183
rect 24492 8946 25002 8984
rect 21162 8693 21672 8836
rect 25941 8904 26045 9065
rect 26045 8904 26244 9065
rect 26244 8904 26451 9065
rect 25941 8761 26451 8904
rect 27787 8904 27943 9065
rect 27943 8904 28142 9065
rect 28142 8904 28297 9065
rect 27787 8761 28297 8904
rect 33756 9526 33993 9642
rect 33756 9244 33993 9526
rect 32093 8850 32466 8852
rect 32093 8655 32156 8850
rect 32156 8655 32422 8850
rect 32422 8655 32466 8850
rect 30089 8511 30449 8555
rect 30089 8443 30220 8511
rect 30220 8443 30294 8511
rect 30294 8443 30449 8511
rect 30089 8282 30449 8443
rect 32093 8513 32466 8655
rect 38707 11276 38951 11403
rect 38707 11192 38727 11276
rect 38727 11192 38795 11276
rect 38795 11192 38951 11276
rect 38707 11072 38951 11192
rect 38707 8132 38951 8237
rect 38707 8048 38727 8132
rect 38727 8048 38795 8132
rect 38795 8048 38951 8132
rect 38707 7906 38951 8048
rect -1883 7228 -1460 7359
rect -1883 7134 -1845 7228
rect -1845 7134 -1757 7228
rect -1757 7134 -1460 7228
rect -1883 6957 -1460 7134
rect 1460 6499 1968 6545
rect 1460 6431 1678 6499
rect 1678 6431 1752 6499
rect 1752 6431 1968 6499
rect 1460 6237 1968 6431
rect -1878 5160 -1455 5296
rect -1878 5066 -1847 5160
rect -1847 5066 -1759 5160
rect -1759 5066 -1455 5160
rect 4663 6569 5173 6647
rect 4663 6370 4722 6569
rect 4722 6370 4901 6569
rect 4901 6370 5173 6569
rect 4663 6343 5173 6370
rect 6231 6258 6535 6409
rect -1878 4894 -1455 5066
rect 1435 3739 1943 3781
rect 1435 3671 1694 3739
rect 1694 3671 1768 3739
rect 1768 3671 1943 3739
rect 1435 3473 1943 3671
rect -1873 3091 -1450 3254
rect -1873 2997 -1845 3091
rect -1845 2997 -1757 3091
rect -1757 2997 -1450 3091
rect -1873 2852 -1450 2997
rect 6231 6079 6265 6258
rect 6265 6079 6464 6258
rect 6464 6079 6535 6258
rect 6231 5899 6535 6079
rect 7365 6256 7669 6419
rect 7365 6077 7407 6256
rect 7407 6077 7606 6256
rect 7606 6077 7669 6256
rect 7365 5909 7669 6077
rect 11214 6567 11724 6645
rect 11214 6368 11273 6567
rect 11273 6368 11452 6567
rect 11452 6368 11724 6567
rect 11214 6341 11724 6368
rect 12782 6256 13086 6407
rect 12782 6077 12816 6256
rect 12816 6077 13015 6256
rect 13015 6077 13086 6256
rect 12782 5897 13086 6077
rect 13916 6254 14220 6417
rect 13916 6075 13958 6254
rect 13958 6075 14157 6254
rect 14157 6075 14220 6254
rect 13916 5907 14220 6075
rect 17869 6568 18379 6646
rect 17869 6369 17928 6568
rect 17928 6369 18107 6568
rect 18107 6369 18379 6568
rect 17869 6342 18379 6369
rect 19437 6257 19741 6408
rect 4657 4919 5167 4987
rect 4657 4720 4736 4919
rect 4736 4720 4915 4919
rect 4915 4720 5167 4919
rect 4657 4683 5167 4720
rect 19437 6078 19471 6257
rect 19471 6078 19670 6257
rect 19670 6078 19741 6257
rect 19437 5898 19741 6078
rect 20571 6255 20875 6418
rect 20571 6076 20613 6255
rect 20613 6076 20812 6255
rect 20812 6076 20875 6255
rect 20571 5908 20875 6076
rect 24491 6569 25001 6647
rect 24491 6370 24550 6569
rect 24550 6370 24729 6569
rect 24729 6370 25001 6569
rect 24491 6343 25001 6370
rect 26059 6258 26363 6409
rect 11208 4917 11718 4985
rect 11208 4718 11287 4917
rect 11287 4718 11466 4917
rect 11466 4718 11718 4917
rect 11208 4681 11718 4718
rect 26059 6079 26093 6258
rect 26093 6079 26292 6258
rect 26292 6079 26363 6258
rect 26059 5899 26363 6079
rect 27193 6256 27497 6419
rect 27193 6077 27235 6256
rect 27235 6077 27434 6256
rect 27434 6077 27497 6256
rect 27193 5909 27497 6077
rect 17863 4918 18373 4986
rect 17863 4719 17942 4918
rect 17942 4719 18121 4918
rect 18121 4719 18373 4918
rect 17863 4682 18373 4719
rect 24485 4919 24995 4987
rect 24485 4720 24564 4919
rect 24564 4720 24743 4919
rect 24743 4720 24995 4919
rect 24485 4683 24995 4720
rect 30149 6591 30509 6634
rect 30149 6523 30291 6591
rect 30291 6523 30365 6591
rect 30365 6523 30509 6591
rect 30149 6361 30509 6523
rect 33756 6147 33993 6206
rect 33756 6031 33993 6147
rect 33756 5749 33993 6031
rect 32093 5355 32466 5357
rect 32093 5160 32156 5355
rect 32156 5160 32422 5355
rect 32422 5160 32466 5355
rect 32093 5088 32466 5160
rect 4656 3315 5166 3382
rect 4656 3116 4731 3315
rect 4731 3116 4910 3315
rect 4910 3116 5166 3315
rect 11207 3313 11717 3380
rect 4656 3078 5166 3116
rect 6105 3036 6209 3197
rect 6209 3036 6408 3197
rect 6408 3036 6615 3197
rect 6105 2893 6615 3036
rect 7951 3036 8107 3197
rect 8107 3036 8306 3197
rect 8306 3036 8461 3197
rect 11207 3114 11282 3313
rect 11282 3114 11461 3313
rect 11461 3114 11717 3313
rect 17862 3314 18372 3381
rect 11207 3076 11717 3114
rect 7951 2893 8461 3036
rect 12656 3034 12760 3195
rect 12760 3034 12959 3195
rect 12959 3034 13166 3195
rect 12656 2891 13166 3034
rect 14502 3034 14658 3195
rect 14658 3034 14857 3195
rect 14857 3034 15012 3195
rect 17862 3115 17937 3314
rect 17937 3115 18116 3314
rect 18116 3115 18372 3314
rect 24484 3315 24994 3382
rect 17862 3077 18372 3115
rect 14502 2891 15012 3034
rect 19311 3035 19415 3196
rect 19415 3035 19614 3196
rect 19614 3035 19821 3196
rect 19311 2892 19821 3035
rect 21157 3035 21313 3196
rect 21313 3035 21512 3196
rect 21512 3035 21667 3196
rect 24484 3116 24559 3315
rect 24559 3116 24738 3315
rect 24738 3116 24994 3315
rect 24484 3078 24994 3116
rect 21157 2892 21667 3035
rect 25933 3036 26037 3197
rect 26037 3036 26236 3197
rect 26236 3036 26443 3197
rect 25933 2893 26443 3036
rect 27779 3036 27935 3197
rect 27935 3036 28134 3197
rect 28134 3036 28289 3197
rect 27779 2893 28289 3036
rect 8134 2374 8642 2564
rect 8134 2306 8404 2374
rect 8404 2306 8478 2374
rect 8478 2306 8642 2374
rect 8134 2256 8642 2306
rect 14673 2379 15181 2545
rect 14673 2311 14958 2379
rect 14958 2311 15032 2379
rect 15032 2311 15181 2379
rect 14673 2237 15181 2311
rect 21379 2367 21887 2520
rect 21379 2299 21607 2367
rect 21607 2299 21681 2367
rect 21681 2299 21887 2367
rect 21379 2212 21887 2299
rect 30145 3521 30505 3566
rect 30145 3453 30288 3521
rect 30288 3453 30362 3521
rect 30362 3453 30505 3521
rect 30145 3293 30505 3453
rect 38705 5000 38949 5094
rect 38705 4916 38723 5000
rect 38723 4916 38791 5000
rect 38791 4916 38949 5000
rect 38705 4763 38949 4916
rect 33756 1799 33993 1858
rect 33756 1683 33993 1799
rect 33756 1401 33993 1683
rect -1873 1023 -1450 1165
rect -1873 929 -1847 1023
rect -1847 929 -1759 1023
rect -1759 929 -1450 1023
rect 32093 1007 32466 1009
rect -1873 763 -1450 929
rect 32093 812 32156 1007
rect 32156 812 32422 1007
rect 32422 812 32466 1007
rect 38707 1856 38951 1976
rect 38707 1772 38723 1856
rect 38723 1772 38791 1856
rect 38791 1772 38951 1856
rect 38707 1645 38951 1772
rect 30155 676 30515 713
rect 30155 608 30295 676
rect 30295 608 30369 676
rect 30369 608 30515 676
rect 30155 440 30515 608
rect 32093 670 32466 812
<< metal5 >>
rect 2853 27341 4987 27344
rect -2561 26978 39070 27341
rect -2561 26674 6475 26978
rect 6985 26975 39070 26978
rect 6985 26750 12988 26975
rect 6985 26740 9177 26750
rect 6985 26674 8043 26740
rect -2561 26230 8043 26674
rect 8347 26240 9177 26740
rect 9481 26671 12988 26750
rect 13498 26974 39070 26975
rect 13498 26970 26080 26974
rect 13498 26747 19522 26970
rect 13498 26737 15690 26747
rect 13498 26671 14556 26737
rect 9481 26240 14556 26671
rect 8347 26230 14556 26240
rect -2561 26227 14556 26230
rect 14860 26237 15690 26737
rect 15994 26666 19522 26747
rect 20032 26742 26080 26970
rect 20032 26732 22224 26742
rect 20032 26666 21090 26732
rect 15994 26237 21090 26666
rect 14860 26227 21090 26237
rect -2561 26222 21090 26227
rect 21394 26232 22224 26732
rect 22528 26670 26080 26742
rect 26590 26746 39070 26974
rect 26590 26736 28782 26746
rect 26590 26670 27648 26736
rect 22528 26232 27648 26670
rect 21394 26226 27648 26232
rect 27952 26236 28782 26736
rect 29086 26236 39070 26746
rect 27952 26226 39070 26236
rect 21394 26222 39070 26226
rect -2561 25318 39070 26222
rect -2561 25014 6469 25318
rect 6979 25315 39070 25318
rect 6979 25014 12982 25315
rect -2561 25011 12982 25014
rect 13492 25314 39070 25315
rect 13492 25310 26074 25314
rect 13492 25011 19516 25310
rect -2561 25006 19516 25011
rect 20026 25010 26074 25310
rect 26584 25010 39070 25314
rect 20026 25006 39070 25010
rect -2561 24985 39070 25006
rect -2592 24003 39070 24985
rect -2592 23713 38705 24003
rect -2592 23409 6468 23713
rect 6978 23710 38705 23713
rect 6978 23528 12981 23710
rect 6978 23409 7917 23528
rect -2592 23224 7917 23409
rect 8427 23224 9763 23528
rect 10273 23406 12981 23528
rect 13491 23709 38705 23710
rect 13491 23705 26073 23709
rect 13491 23525 19515 23705
rect 13491 23406 14430 23525
rect 10273 23224 14430 23406
rect -2592 23221 14430 23224
rect 14940 23221 16276 23525
rect 16786 23401 19515 23525
rect 20025 23520 26073 23705
rect 20025 23401 20964 23520
rect 16786 23221 20964 23401
rect -2592 23216 20964 23221
rect 21474 23216 22810 23520
rect 23320 23405 26073 23520
rect 26583 23672 38705 23709
rect 38949 23672 39070 24003
rect 26583 23524 39070 23672
rect 26583 23405 27522 23524
rect 23320 23220 27522 23405
rect 28032 23220 29368 23524
rect 29878 23220 39070 23524
rect 23320 23216 39070 23220
rect -2592 21877 39070 23216
rect -2561 21374 39070 21877
rect -2561 21371 28524 21374
rect -2561 21366 22011 21371
rect -2561 21363 15477 21366
rect -2561 21142 8919 21363
rect -2561 20632 6423 21142
rect 6727 21132 8919 21142
rect 6727 20632 7557 21132
rect -2561 20622 7557 20632
rect 7861 21066 8919 21132
rect 9429 21138 15477 21363
rect 9429 21066 12981 21138
rect 7861 20628 12981 21066
rect 13285 21128 15477 21138
rect 13285 20628 14115 21128
rect 7861 20622 14115 20628
rect -2561 20618 14115 20622
rect 14419 21062 15477 21128
rect 15987 21143 22011 21366
rect 15987 21062 19515 21143
rect 14419 20633 19515 21062
rect 19819 21133 22011 21143
rect 19819 20633 20649 21133
rect 14419 20623 20649 20633
rect 20953 21067 22011 21133
rect 22521 21146 28524 21371
rect 22521 21067 26028 21146
rect 20953 20636 26028 21067
rect 26332 21136 28524 21146
rect 26332 20636 27162 21136
rect 20953 20626 27162 20636
rect 27466 21070 28524 21136
rect 29034 21070 39070 21374
rect 27466 20845 39070 21070
rect 27466 20626 38707 20845
rect 20953 20623 38707 20626
rect 14419 20618 38707 20623
rect -2561 20514 38707 20618
rect 38951 20514 39070 20845
rect -2561 19714 39070 20514
rect -2561 19711 28530 19714
rect -2561 19710 22017 19711
rect -2561 19406 8925 19710
rect 9435 19706 22017 19710
rect 9435 19406 15483 19706
rect -2561 19402 15483 19406
rect 15993 19407 22017 19706
rect 22527 19410 28530 19711
rect 29040 19410 39070 19714
rect 22527 19407 39070 19410
rect 15993 19402 39070 19407
rect -2561 18109 39070 19402
rect -2561 18106 28531 18109
rect -2561 18105 22018 18106
rect -2561 17920 8926 18105
rect -2561 17616 5631 17920
rect 6141 17616 7477 17920
rect 7987 17801 8926 17920
rect 9436 18101 22018 18105
rect 9436 17916 15484 18101
rect 9436 17801 12189 17916
rect 7987 17616 12189 17801
rect -2561 17612 12189 17616
rect 12699 17612 14035 17916
rect 14545 17797 15484 17916
rect 15994 17921 22018 18101
rect 15994 17797 18723 17921
rect 14545 17617 18723 17797
rect 19233 17617 20569 17921
rect 21079 17802 22018 17921
rect 22528 17924 28531 18106
rect 22528 17802 25236 17924
rect 21079 17620 25236 17802
rect 25746 17620 27082 17924
rect 27592 17805 28531 17924
rect 29041 17805 39070 18109
rect 27592 17712 39070 17805
rect 27592 17620 38705 17712
rect 21079 17617 38705 17620
rect 14545 17612 38705 17617
rect -2561 17381 38705 17612
rect 38949 17381 39070 17712
rect -2561 15683 39070 17381
rect -2561 15281 -1878 15683
rect -1455 15281 39070 15683
rect -2561 14594 39070 15281
rect -2561 14370 38707 14594
rect -2561 14062 8172 14370
rect 8681 14345 38707 14370
rect 8681 14062 14714 14345
rect -2561 14037 14714 14062
rect 15223 14330 38707 14345
rect 15223 14037 21381 14330
rect -2561 14023 21381 14037
rect 21890 14263 38707 14330
rect 38951 14263 39070 14594
rect 21890 14156 39070 14263
rect 21890 14023 30082 14156
rect -2561 13883 30082 14023
rect 30442 13883 39070 14156
rect -2561 13792 39070 13883
rect -2561 13589 33754 13792
rect -2561 13187 -1883 13589
rect -1460 13335 33754 13589
rect 33991 13335 39070 13792
rect -1460 13187 39070 13335
rect -2561 12943 39070 13187
rect -2561 12604 32091 12943
rect 32464 12604 39070 12943
rect -2561 12515 39070 12604
rect -2561 12432 11220 12515
rect -2561 12124 1509 12432
rect 2017 12427 11220 12432
rect 2017 12124 4671 12427
rect -2561 12123 4671 12124
rect 5181 12211 11220 12427
rect 11730 12447 24499 12515
rect 11730 12287 17874 12447
rect 11730 12277 13922 12287
rect 11730 12211 12788 12277
rect 5181 12199 12788 12211
rect 5181 12189 7373 12199
rect 5181 12123 6239 12189
rect -2561 11679 6239 12123
rect 6543 11689 7373 12189
rect 7677 11767 12788 12199
rect 13092 11777 13922 12277
rect 14226 12143 17874 12287
rect 18384 12219 24499 12447
rect 18384 12209 20576 12219
rect 18384 12143 19442 12209
rect 14226 11777 19442 12143
rect 13092 11767 19442 11777
rect 7677 11699 19442 11767
rect 19746 11709 20576 12209
rect 20880 12211 24499 12219
rect 25009 12287 39070 12515
rect 25009 12277 27201 12287
rect 25009 12211 26067 12277
rect 20880 11767 26067 12211
rect 26371 11777 27201 12277
rect 27505 11777 39070 12287
rect 26371 11767 39070 11777
rect 20880 11709 39070 11767
rect 19746 11699 39070 11709
rect 7677 11689 39070 11699
rect 6543 11679 39070 11689
rect -2561 11593 39070 11679
rect -2561 11521 30088 11593
rect -2561 11119 -1893 11521
rect -1470 11320 30088 11521
rect 30448 11403 39070 11593
rect 30448 11320 38707 11403
rect -1470 11119 38707 11320
rect -2561 11072 38707 11119
rect 38951 11072 39070 11403
rect -2561 10855 39070 11072
rect -2561 10767 11214 10855
rect -2561 10463 4665 10767
rect 5175 10551 11214 10767
rect 11724 10787 24493 10855
rect 11724 10551 17868 10787
rect 5175 10483 17868 10551
rect 18378 10551 24493 10787
rect 25003 10551 39070 10855
rect 18378 10483 39070 10551
rect 5175 10463 39070 10483
rect -2561 9850 39070 10463
rect -2561 9542 1484 9850
rect 1992 9701 39070 9850
rect 1992 9542 33756 9701
rect -2561 9458 33756 9542
rect -2561 9056 -1867 9458
rect -1444 9250 33756 9458
rect -1444 9162 11213 9250
rect -1444 9056 4664 9162
rect -2561 8858 4664 9056
rect 5174 8977 11213 9162
rect 5174 8858 6113 8977
rect -2561 8673 6113 8858
rect 6623 8673 7959 8977
rect 8469 8946 11213 8977
rect 11723 9182 24492 9250
rect 11723 9065 17867 9182
rect 11723 8946 12662 9065
rect 8469 8761 12662 8946
rect 13172 8761 14508 9065
rect 15018 8878 17867 9065
rect 18377 8997 24492 9182
rect 18377 8878 19316 8997
rect 15018 8761 19316 8878
rect 8469 8693 19316 8761
rect 19826 8693 21162 8997
rect 21672 8946 24492 8997
rect 25002 9244 33756 9250
rect 33993 9244 39070 9701
rect 25002 9065 39070 9244
rect 25002 8946 25941 9065
rect 21672 8761 25941 8946
rect 26451 8761 27787 9065
rect 28297 8852 39070 9065
rect 28297 8761 32093 8852
rect 21672 8693 32093 8761
rect 8469 8673 32093 8693
rect -2561 8555 32093 8673
rect -2561 8282 30089 8555
rect 30449 8513 32093 8555
rect 32466 8513 39070 8852
rect 30449 8282 39070 8513
rect -2561 8237 39070 8282
rect -2561 7906 38707 8237
rect 38951 7906 39070 8237
rect -2561 7359 39070 7906
rect -2561 6957 -1883 7359
rect -1460 6957 39070 7359
rect -2561 6647 39070 6957
rect -2561 6545 4663 6647
rect -2561 6237 1460 6545
rect 1968 6343 4663 6545
rect 5173 6646 24491 6647
rect 5173 6645 17869 6646
rect 5173 6419 11214 6645
rect 5173 6409 7365 6419
rect 5173 6343 6231 6409
rect 1968 6237 6231 6343
rect -2561 5899 6231 6237
rect 6535 5909 7365 6409
rect 7669 6341 11214 6419
rect 11724 6417 17869 6645
rect 11724 6407 13916 6417
rect 11724 6341 12782 6407
rect 7669 5909 12782 6341
rect 6535 5899 12782 5909
rect -2561 5897 12782 5899
rect 13086 5907 13916 6407
rect 14220 6342 17869 6417
rect 18379 6418 24491 6646
rect 18379 6408 20571 6418
rect 18379 6342 19437 6408
rect 14220 5907 19437 6342
rect 13086 5898 19437 5907
rect 19741 5908 20571 6408
rect 20875 6343 24491 6418
rect 25001 6634 39070 6647
rect 25001 6419 30149 6634
rect 25001 6409 27193 6419
rect 25001 6343 26059 6409
rect 20875 5908 26059 6343
rect 19741 5899 26059 5908
rect 26363 5909 27193 6409
rect 27497 6361 30149 6419
rect 30509 6361 39070 6634
rect 27497 6206 39070 6361
rect 27497 5909 33756 6206
rect 26363 5899 33756 5909
rect 19741 5898 33756 5899
rect 13086 5897 33756 5898
rect -2561 5749 33756 5897
rect 33993 5749 39070 6206
rect -2561 5357 39070 5749
rect -2561 5296 32093 5357
rect -2561 4894 -1878 5296
rect -1455 5088 32093 5296
rect 32466 5094 39070 5357
rect 32466 5088 38705 5094
rect -1455 4987 38705 5088
rect -1455 4894 4657 4987
rect -2561 4683 4657 4894
rect 5167 4986 24485 4987
rect 5167 4985 17863 4986
rect 5167 4683 11208 4985
rect -2561 4681 11208 4683
rect 11718 4682 17863 4985
rect 18373 4683 24485 4986
rect 24995 4763 38705 4987
rect 38949 4763 39070 5094
rect 24995 4683 39070 4763
rect 18373 4682 39070 4683
rect 11718 4681 39070 4682
rect -2561 3781 39070 4681
rect -2561 3473 1435 3781
rect 1943 3566 39070 3781
rect 1943 3473 30145 3566
rect -2561 3382 30145 3473
rect -2561 3254 4656 3382
rect -2561 2852 -1873 3254
rect -1450 3078 4656 3254
rect 5166 3381 24484 3382
rect 5166 3380 17862 3381
rect 5166 3197 11207 3380
rect 5166 3078 6105 3197
rect -1450 2893 6105 3078
rect 6615 2893 7951 3197
rect 8461 3076 11207 3197
rect 11717 3195 17862 3380
rect 11717 3076 12656 3195
rect 8461 2893 12656 3076
rect -1450 2891 12656 2893
rect 13166 2891 14502 3195
rect 15012 3077 17862 3195
rect 18372 3196 24484 3381
rect 18372 3077 19311 3196
rect 15012 2892 19311 3077
rect 19821 2892 21157 3196
rect 21667 3078 24484 3196
rect 24994 3293 30145 3382
rect 30505 3293 39070 3566
rect 24994 3197 39070 3293
rect 24994 3078 25933 3197
rect 21667 2893 25933 3078
rect 26443 2893 27779 3197
rect 28289 2893 39070 3197
rect 21667 2892 39070 2893
rect 15012 2891 39070 2892
rect -1450 2852 39070 2891
rect -2561 2564 39070 2852
rect -2561 2256 8134 2564
rect 8642 2545 39070 2564
rect 8642 2256 14673 2545
rect -2561 2237 14673 2256
rect 15181 2520 39070 2545
rect 15181 2237 21379 2520
rect -2561 2212 21379 2237
rect 21887 2212 39070 2520
rect -2561 1976 39070 2212
rect -2561 1858 38707 1976
rect -2561 1401 33756 1858
rect 33993 1645 38707 1858
rect 38951 1645 39070 1976
rect 33993 1401 39070 1645
rect -2561 1165 39070 1401
rect -2561 763 -1873 1165
rect -1450 1009 39070 1165
rect -1450 763 32093 1009
rect -2561 713 32093 763
rect -2561 440 30155 713
rect 30515 670 32093 713
rect 32466 670 39070 1009
rect 30515 440 39070 670
rect -2561 164 39070 440
rect -2561 149 -862 164
rect -453 149 39070 164
rect 16859 -805 19778 149
<< labels >>
flabel metal1 -4163 19834 -3932 19972 1 FreeSans 800 0 0 0 B[0]
port 1 n
flabel metal1 -4161 20248 -3930 20386 1 FreeSans 800 0 0 0 B[1]
port 2 n
flabel metal1 -4161 20685 -3930 20823 1 FreeSans 800 0 0 0 B[2]
port 3 n
flabel metal1 -4163 21110 -3932 21248 1 FreeSans 800 0 0 0 B[3]
port 4 n
flabel metal1 -4163 21527 -3932 21665 1 FreeSans 800 0 0 0 B[4]
port 5 n
flabel metal1 -4163 21966 -3932 22104 1 FreeSans 800 0 0 0 B[5]
port 6 n
flabel metal1 -4163 22399 -3932 22537 1 FreeSans 800 0 0 0 B[6]
port 7 n
flabel metal1 -4161 22830 -3930 22968 1 FreeSans 800 0 0 0 B[7]
port 8 n
flabel metal1 -4161 23255 -3655 23392 1 FreeSans 800 0 0 0 opcode[0]
port 9 n
flabel metal1 -4161 23668 -3655 23805 1 FreeSans 800 0 0 0 opcode[1]
port 10 n
flabel metal1 -4160 24095 -3929 24233 1 FreeSans 800 0 0 0 A[7]
port 11 n
flabel metal1 -4160 24527 -3929 24665 1 FreeSans 800 0 0 0 A[6]
port 12 n
flabel metal1 -4160 24974 -3929 25112 1 FreeSans 800 0 0 0 A[5]
port 13 n
flabel metal1 -4156 25396 -3925 25534 1 FreeSans 800 0 0 0 A[4]
port 14 n
flabel metal1 -4156 25829 -3925 25967 1 FreeSans 800 0 0 0 A[3]
port 15 n
flabel metal1 -4156 26251 -3925 26389 1 FreeSans 800 0 0 0 A[2]
port 16 n
flabel metal1 -4156 26669 -3925 26807 1 FreeSans 800 0 0 0 A[1]
port 17 n
flabel metal1 -4156 27099 -3925 27237 1 FreeSans 800 0 0 0 A[0]
port 18 n
flabel metal1 4387 28457 4526 28562 1 FreeSans 800 0 0 0 Cout
port 19 n
flabel metal4 17228 28311 19525 29269 1 FreeSans 4000 0 0 0 VDD
port 20 n
flabel metal5 17064 -707 19575 278 1 FreeSans 4000 0 0 0 VSS
port 21 n
flabel metal1 39227 297 39561 609 1 FreeSans 1600 0 0 0 Y[7]
port 22 n
flabel metal1 39227 3437 39561 3749 1 FreeSans 1600 0 0 0 Y[6]
port 23 n
flabel metal1 39231 22332 39565 22644 1 FreeSans 1600 0 0 0 Y[0]
port 24 n
flabel metal1 39232 19190 39566 19502 1 FreeSans 1600 0 0 0 Y[1]
port 25 n
flabel metal1 39229 16057 39563 16369 1 FreeSans 1600 0 0 0 Y[2]
port 26 n
flabel metal1 39228 12913 39562 13225 1 FreeSans 1600 0 0 0 Y[3]
port 27 n
flabel metal1 39231 9712 39565 10024 1 FreeSans 1600 0 0 0 Y[4]
port 28 n
flabel metal1 39231 6567 39565 6879 1 FreeSans 1600 0 0 0 Y[5]
port 29 n
<< end >>
