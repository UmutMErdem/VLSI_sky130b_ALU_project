magic
tech sky130B
timestamp 1735468497
<< nwell >>
rect -298 -81 298 81
<< pmos >>
rect -251 -50 -221 50
rect -192 -50 -162 50
rect -133 -50 -103 50
rect -74 -50 -44 50
rect -15 -50 15 50
rect 44 -50 74 50
rect 103 -50 133 50
rect 162 -50 192 50
rect 221 -50 251 50
<< pdiff >>
rect -280 44 -251 50
rect -280 -44 -274 44
rect -257 -44 -251 44
rect -280 -50 -251 -44
rect -221 44 -192 50
rect -221 -44 -215 44
rect -198 -44 -192 44
rect -221 -50 -192 -44
rect -162 44 -133 50
rect -162 -44 -156 44
rect -139 -44 -133 44
rect -162 -50 -133 -44
rect -103 44 -74 50
rect -103 -44 -97 44
rect -80 -44 -74 44
rect -103 -50 -74 -44
rect -44 44 -15 50
rect -44 -44 -38 44
rect -21 -44 -15 44
rect -44 -50 -15 -44
rect 15 44 44 50
rect 15 -44 21 44
rect 38 -44 44 44
rect 15 -50 44 -44
rect 74 44 103 50
rect 74 -44 80 44
rect 97 -44 103 44
rect 74 -50 103 -44
rect 133 44 162 50
rect 133 -44 139 44
rect 156 -44 162 44
rect 133 -50 162 -44
rect 192 44 221 50
rect 192 -44 198 44
rect 215 -44 221 44
rect 192 -50 221 -44
rect 251 44 280 50
rect 251 -44 257 44
rect 274 -44 280 44
rect 251 -50 280 -44
<< pdiffc >>
rect -274 -44 -257 44
rect -215 -44 -198 44
rect -156 -44 -139 44
rect -97 -44 -80 44
rect -38 -44 -21 44
rect 21 -44 38 44
rect 80 -44 97 44
rect 139 -44 156 44
rect 198 -44 215 44
rect 257 -44 274 44
<< poly >>
rect -251 50 -221 63
rect -192 50 -162 63
rect -133 50 -103 63
rect -74 50 -44 63
rect -15 50 15 63
rect 44 50 74 63
rect 103 50 133 63
rect 162 50 192 63
rect 221 50 251 63
rect -251 -63 -221 -50
rect -192 -63 -162 -50
rect -133 -63 -103 -50
rect -74 -63 -44 -50
rect -15 -63 15 -50
rect 44 -63 74 -50
rect 103 -63 133 -50
rect 162 -63 192 -50
rect 221 -63 251 -50
<< locali >>
rect -274 44 -257 52
rect -274 -52 -257 -44
rect -215 44 -198 52
rect -215 -52 -198 -44
rect -156 44 -139 52
rect -156 -52 -139 -44
rect -97 44 -80 52
rect -97 -52 -80 -44
rect -38 44 -21 52
rect -38 -52 -21 -44
rect 21 44 38 52
rect 21 -52 38 -44
rect 80 44 97 52
rect 80 -52 97 -44
rect 139 44 156 52
rect 139 -52 156 -44
rect 198 44 215 52
rect 198 -52 215 -44
rect 257 44 274 52
rect 257 -52 274 -44
<< viali >>
rect -274 -44 -257 44
rect -215 -44 -198 44
rect -156 -44 -139 44
rect -97 -44 -80 44
rect -38 -44 -21 44
rect 21 -44 38 44
rect 80 -44 97 44
rect 139 -44 156 44
rect 198 -44 215 44
rect 257 -44 274 44
<< metal1 >>
rect -277 44 -254 50
rect -277 -44 -274 44
rect -257 -44 -254 44
rect -277 -50 -254 -44
rect -218 44 -195 50
rect -218 -44 -215 44
rect -198 -44 -195 44
rect -218 -50 -195 -44
rect -159 44 -136 50
rect -159 -44 -156 44
rect -139 -44 -136 44
rect -159 -50 -136 -44
rect -100 44 -77 50
rect -100 -44 -97 44
rect -80 -44 -77 44
rect -100 -50 -77 -44
rect -41 44 -18 50
rect -41 -44 -38 44
rect -21 -44 -18 44
rect -41 -50 -18 -44
rect 18 44 41 50
rect 18 -44 21 44
rect 38 -44 41 44
rect 18 -50 41 -44
rect 77 44 100 50
rect 77 -44 80 44
rect 97 -44 100 44
rect 77 -50 100 -44
rect 136 44 159 50
rect 136 -44 139 44
rect 156 -44 159 44
rect 136 -50 159 -44
rect 195 44 218 50
rect 195 -44 198 44
rect 215 -44 218 44
rect 195 -50 218 -44
rect 254 44 277 50
rect 254 -44 257 44
rect 274 -44 277 44
rect 254 -50 277 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
