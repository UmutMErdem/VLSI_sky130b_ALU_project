magic
tech sky130B
magscale 1 2
timestamp 1736541398
use and2  and2_0
timestamp 1736444617
transform 1 0 -30 0 1 3475
box 0 -794 1193 576
use and2  and2_1
timestamp 1736444617
transform 1 0 -38 0 1 890
box 0 -794 1193 576
use and2  and2_2
timestamp 1736444617
transform 1 0 -38 0 1 -3412
box 0 -794 1193 576
use and2  and2_3
timestamp 1736444617
transform 1 0 -49 0 1 -6457
box 0 -794 1193 576
use and2  and2_4
timestamp 1736444617
transform 1 0 9465 0 1 5317
box 0 -794 1193 576
use and2  and2_5
timestamp 1736444617
transform 1 0 9437 0 1 -8070
box 0 -794 1193 576
use and2  and2_6
timestamp 1736444617
transform 1 0 2486 0 1 -8127
box 0 -794 1193 576
use and2  and2_7
timestamp 1736444617
transform 1 0 2514 0 1 5260
box 0 -794 1193 576
use and2  and2_8
timestamp 1736444617
transform 1 0 32745 0 1 -6645
box 0 -794 1193 576
use and2  and2_9
timestamp 1736444617
transform 1 0 32745 0 1 2533
box 0 -794 1193 576
use and2  and2_10
timestamp 1736444617
transform 1 0 16731 0 1 5317
box 0 -794 1193 576
use and2  and2_11
timestamp 1736444617
transform 1 0 16703 0 1 -8070
box 0 -794 1193 576
use and2  and2_12
timestamp 1736444617
transform 1 0 32747 0 1 5663
box 0 -794 1193 576
use and2  and2_13
timestamp 1736444617
transform 1 0 32748 0 1 -9720
box 0 -794 1193 576
use and2  and2_14
timestamp 1736444617
transform 1 0 32748 0 1 -3575
box 0 -794 1193 576
use and2  and2_15
timestamp 1736444617
transform 1 0 32745 0 1 -500
box 0 -794 1193 576
use fulladder  fulladder_0
timestamp 1735941024
transform 1 0 11806 0 1 -961
box -2361 -464 3896 5054
use fulladder  fulladder_1
timestamp 1735941024
transform 1 0 11798 0 1 -6741
box -2361 -464 3896 5054
use fulladder  fulladder_2
timestamp 1735941024
transform 1 0 4847 0 1 -6798
box -2361 -464 3896 5054
use fulladder  fulladder_3
timestamp 1735941024
transform 1 0 4855 0 1 -1018
box -2361 -464 3896 5054
use fulladder  fulladder_6
timestamp 1735941024
transform 1 0 19072 0 1 -961
box -2361 -464 3896 5054
use fulladder  fulladder_7
timestamp 1735941024
transform 1 0 19064 0 1 -6741
box -2361 -464 3896 5054
use fulladder  fulladder_8
timestamp 1735941024
transform 1 0 26309 0 1 -961
box -2361 -464 3896 5054
use fulladder  fulladder_9
timestamp 1735941024
transform 1 0 26301 0 1 -6741
box -2361 -464 3896 5054
use half_adder  half_adder_0
timestamp 1736520155
transform 1 0 38348 0 1 -9392
box -1792 -1094 1193 1827
use half_adder  half_adder_1
timestamp 1736520155
transform 1 0 38348 0 1 3595
box -1792 -1094 1193 1827
use half_adder  half_adder_2
timestamp 1736520155
transform 1 0 38291 0 1 -496
box -1792 -1094 1193 1827
use half_adder  half_adder_3
timestamp 1736520155
transform 1 0 38320 0 1 -5044
box -1792 -1094 1193 1827
<< end >>
