magic
tech sky130B
magscale 1 2
timestamp 1736810822
<< nwell >>
rect 859 22054 2636 22344
rect 4003 22054 5780 22344
rect 7135 22058 8912 22348
rect 10279 22058 12056 22348
rect 859 21854 2637 22054
rect 4003 21854 5781 22054
rect 7135 21858 8913 22058
rect 10279 21858 12057 22058
rect 13481 22054 15258 22344
rect 16625 22054 18402 22344
rect 19757 22058 21534 22348
rect 22901 22058 24678 22348
rect 418 21530 3110 21854
rect 3562 21530 6254 21854
rect 6694 21534 9386 21858
rect 9838 21534 12530 21858
rect 13481 21854 15259 22054
rect 16625 21854 18403 22054
rect 19757 21858 21535 22058
rect 22901 21858 24679 22058
rect 13040 21530 15732 21854
rect 16184 21530 18876 21854
rect 19316 21534 22008 21858
rect 22460 21534 25152 21858
rect 2860 16673 4052 16919
rect 4308 16673 5500 16919
rect 5806 16675 6998 16921
rect 7254 16675 8446 16921
rect 2860 16661 4053 16673
rect 4308 16661 5501 16673
rect 5806 16663 6999 16675
rect 7254 16663 8447 16675
rect 2861 16349 4053 16661
rect 4309 16349 5501 16661
rect 5807 16351 6999 16663
rect 7255 16351 8447 16663
rect 8774 16673 9966 16919
rect 10222 16673 11414 16919
rect 11720 16675 12912 16921
rect 13168 16675 14360 16921
rect 8774 16661 9967 16673
rect 10222 16661 11415 16673
rect 11720 16663 12913 16675
rect 13168 16663 14361 16675
rect 8775 16349 9967 16661
rect 10223 16349 11415 16661
rect 11721 16351 12913 16663
rect 13169 16351 14361 16663
rect 14624 16346 15538 17124
rect 15792 16346 16706 17124
rect 15054 15756 15538 16346
rect 16222 16086 16706 16346
rect 16960 16344 17874 17124
rect 18128 16346 19042 17124
rect 19302 16348 20216 17126
rect 17390 16086 17874 16344
rect 16221 16038 16706 16086
rect 17389 16038 17874 16086
rect 16221 15762 16705 16038
rect 17389 15762 17873 16038
rect 18558 15762 19042 16346
rect 19732 16082 20216 16348
rect 20470 16346 21384 17126
rect 21638 16348 22552 17126
rect 19730 16040 20216 16082
rect 20900 16081 21384 16346
rect 22068 16081 22552 16348
rect 22806 16346 23720 17126
rect 23236 16082 23720 16346
rect 20899 16040 21384 16081
rect 22067 16040 22552 16081
rect 23235 16040 23720 16082
rect 19730 15758 20214 16040
rect 20899 15757 21383 16040
rect 22067 15757 22551 16040
rect 23235 15758 23719 16040
rect 3361 14916 5138 15206
rect 6505 14916 8282 15206
rect 9637 14920 11414 15210
rect 12781 14920 14558 15210
rect 3361 14716 5139 14916
rect 6505 14716 8283 14916
rect 9637 14720 11415 14920
rect 12781 14720 14559 14920
rect 15983 14916 17760 15206
rect 19127 14916 20904 15206
rect 22259 14920 24036 15210
rect 25403 14920 27180 15210
rect 2920 14392 5612 14716
rect 6064 14392 8756 14716
rect 9196 14396 11888 14720
rect 12340 14396 15032 14720
rect 15983 14716 17761 14916
rect 19127 14716 20905 14916
rect 22259 14720 24037 14920
rect 25403 14720 27181 14920
rect 15542 14392 18234 14716
rect 18686 14392 21378 14716
rect 21818 14396 24510 14720
rect 24962 14396 27654 14720
rect 3361 12182 5138 12472
rect 6505 12182 8282 12472
rect 9637 12186 11414 12476
rect 12781 12186 14558 12476
rect 3361 11982 5139 12182
rect 6505 11982 8283 12182
rect 9637 11986 11415 12186
rect 12781 11986 14559 12186
rect 15983 12182 17760 12472
rect 19127 12182 20904 12472
rect 22259 12186 24036 12476
rect 25403 12186 27180 12476
rect 2920 11658 5612 11982
rect 6064 11658 8756 11982
rect 9196 11662 11888 11986
rect 12340 11662 15032 11986
rect 15983 11982 17761 12182
rect 19127 11982 20905 12182
rect 22259 11986 24037 12186
rect 25403 11986 27181 12186
rect 15542 11658 18234 11982
rect 18686 11658 21378 11982
rect 21818 11662 24510 11986
rect 24962 11662 27654 11986
rect 3351 9450 5128 9740
rect 6495 9450 8272 9740
rect 9627 9454 11404 9744
rect 12771 9454 14548 9744
rect 3351 9250 5129 9450
rect 6495 9250 8273 9450
rect 9627 9254 11405 9454
rect 12771 9254 14549 9454
rect 15973 9450 17750 9740
rect 19117 9450 20894 9740
rect 22249 9454 24026 9744
rect 25393 9454 27170 9744
rect 2910 8926 5602 9250
rect 6054 8926 8746 9250
rect 9186 8930 11878 9254
rect 12330 8930 15022 9254
rect 15973 9250 17751 9450
rect 19117 9250 20895 9450
rect 22249 9254 24027 9454
rect 25393 9254 27171 9454
rect 15532 8926 18224 9250
rect 18676 8926 21368 9250
rect 21808 8930 24500 9254
rect 24952 8930 27644 9254
rect 3318 6600 3794 6792
rect 5386 6602 5862 6792
rect 3128 6305 3972 6600
rect 5196 6307 6040 6602
rect 7455 6600 7931 6792
rect 9523 6602 9999 6792
rect 11592 6602 12068 6794
rect 13660 6604 14136 6794
rect 2647 5981 4452 6305
rect 4715 5983 6520 6307
rect 7265 6305 8109 6600
rect 9333 6307 10177 6602
rect 11402 6307 12246 6602
rect 13470 6309 14314 6604
rect 15729 6602 16205 6794
rect 17797 6604 18273 6794
rect 3074 5288 3912 5981
rect 5142 5290 5980 5983
rect 6784 5981 8589 6305
rect 8852 5983 10657 6307
rect 10921 5983 12726 6307
rect 12989 5985 14794 6309
rect 15539 6307 16383 6602
rect 17607 6309 18451 6604
rect 7211 5288 8049 5981
rect 9279 5290 10117 5983
rect 11348 5290 12186 5983
rect 13416 5292 14254 5985
rect 15058 5983 16863 6307
rect 17126 5985 18931 6309
rect 19379 6297 19863 6849
rect 20117 6301 20601 6847
rect 20855 6297 21339 6847
rect 21597 6295 22081 6847
rect 22337 6295 22821 6847
rect 23075 6295 23559 6847
rect 23813 6295 24297 6847
rect 24551 6295 25035 6847
rect 15485 5290 16323 5983
rect 17553 5292 18391 5985
rect 653 2202 2430 2492
rect 3797 2202 5574 2492
rect 6929 2206 8706 2496
rect 10073 2206 11850 2496
rect 653 2002 2431 2202
rect 3797 2002 5575 2202
rect 6929 2006 8707 2206
rect 10073 2006 11851 2206
rect 13275 2202 15052 2492
rect 16419 2202 18196 2492
rect 19551 2206 21328 2496
rect 22695 2206 24472 2496
rect 212 1678 2904 2002
rect 3356 1678 6048 2002
rect 6488 1682 9180 2006
rect 9632 1682 12324 2006
rect 13275 2002 15053 2202
rect 16419 2002 18197 2202
rect 19551 2006 21329 2206
rect 22695 2006 24473 2206
rect 12834 1678 15526 2002
rect 15978 1678 18670 2002
rect 19110 1682 21802 2006
rect 22254 1682 24946 2006
rect 685 -1690 2462 -1400
rect 3829 -1690 5606 -1400
rect 6961 -1686 8738 -1396
rect 10105 -1686 11882 -1396
rect 685 -1890 2463 -1690
rect 3829 -1890 5607 -1690
rect 6961 -1886 8739 -1686
rect 10105 -1886 11883 -1686
rect 13307 -1690 15084 -1400
rect 16451 -1690 18228 -1400
rect 19583 -1686 21360 -1396
rect 22727 -1686 24504 -1396
rect 244 -2214 2936 -1890
rect 3388 -2214 6080 -1890
rect 6520 -2210 9212 -1886
rect 9664 -2210 12356 -1886
rect 13307 -1890 15085 -1690
rect 16451 -1890 18229 -1690
rect 19583 -1886 21361 -1686
rect 22727 -1886 24505 -1686
rect 12866 -2214 15558 -1890
rect 16010 -2214 18702 -1890
rect 19142 -2210 21834 -1886
rect 22286 -2210 24978 -1886
<< nmos >>
rect 1346 20459 1406 20659
rect 1538 20259 1598 20659
rect 1656 20259 1716 20659
rect 1774 20259 1834 20659
rect 1892 20259 1952 20659
rect 2088 20459 2148 20659
rect 4490 20459 4550 20659
rect 4682 20259 4742 20659
rect 4800 20259 4860 20659
rect 4918 20259 4978 20659
rect 5036 20259 5096 20659
rect 5232 20459 5292 20659
rect 7622 20463 7682 20663
rect 7814 20263 7874 20663
rect 7932 20263 7992 20663
rect 8050 20263 8110 20663
rect 8168 20263 8228 20663
rect 8364 20463 8424 20663
rect 10766 20463 10826 20663
rect 10958 20263 11018 20663
rect 11076 20263 11136 20663
rect 11194 20263 11254 20663
rect 11312 20263 11372 20663
rect 11508 20463 11568 20663
rect 13968 20459 14028 20659
rect 14160 20259 14220 20659
rect 14278 20259 14338 20659
rect 14396 20259 14456 20659
rect 14514 20259 14574 20659
rect 14710 20459 14770 20659
rect 17112 20459 17172 20659
rect 17304 20259 17364 20659
rect 17422 20259 17482 20659
rect 17540 20259 17600 20659
rect 17658 20259 17718 20659
rect 17854 20459 17914 20659
rect 20244 20463 20304 20663
rect 20436 20263 20496 20663
rect 20554 20263 20614 20663
rect 20672 20263 20732 20663
rect 20790 20263 20850 20663
rect 20986 20463 21046 20663
rect 23388 20463 23448 20663
rect 23580 20263 23640 20663
rect 23698 20263 23758 20663
rect 23816 20263 23876 20663
rect 23934 20263 23994 20663
rect 24130 20463 24190 20663
rect 3192 15774 3252 16174
rect 3310 15774 3370 16174
rect 3545 15974 3605 16174
rect 4640 15774 4700 16174
rect 4758 15774 4818 16174
rect 4993 15974 5053 16174
rect 6138 15776 6198 16176
rect 6256 15776 6316 16176
rect 6491 15976 6551 16176
rect 7586 15776 7646 16176
rect 7704 15776 7764 16176
rect 7939 15976 7999 16176
rect 9106 15774 9166 16174
rect 9224 15774 9284 16174
rect 9459 15974 9519 16174
rect 10554 15774 10614 16174
rect 10672 15774 10732 16174
rect 10907 15974 10967 16174
rect 12052 15776 12112 16176
rect 12170 15776 12230 16176
rect 12405 15976 12465 16176
rect 13500 15776 13560 16176
rect 13618 15776 13678 16176
rect 13853 15976 13913 16176
rect 14628 15822 14688 16022
rect 14746 15822 14806 16022
rect 14864 15822 14924 16022
rect 15796 15824 15856 16024
rect 15914 15824 15974 16024
rect 16032 15824 16092 16024
rect 16964 15824 17024 16024
rect 17082 15824 17142 16024
rect 17200 15824 17260 16024
rect 18132 15824 18192 16024
rect 18250 15824 18310 16024
rect 18368 15824 18428 16024
rect 19306 15824 19366 16024
rect 19424 15824 19484 16024
rect 19542 15824 19602 16024
rect 20474 15824 20534 16024
rect 20592 15824 20652 16024
rect 20710 15824 20770 16024
rect 21642 15826 21702 16026
rect 21760 15826 21820 16026
rect 21878 15826 21938 16026
rect 22810 15826 22870 16026
rect 22928 15826 22988 16026
rect 23046 15826 23106 16026
rect 3848 13321 3908 13521
rect 4040 13121 4100 13521
rect 4158 13121 4218 13521
rect 4276 13121 4336 13521
rect 4394 13121 4454 13521
rect 4590 13321 4650 13521
rect 6992 13321 7052 13521
rect 7184 13121 7244 13521
rect 7302 13121 7362 13521
rect 7420 13121 7480 13521
rect 7538 13121 7598 13521
rect 7734 13321 7794 13521
rect 10124 13325 10184 13525
rect 10316 13125 10376 13525
rect 10434 13125 10494 13525
rect 10552 13125 10612 13525
rect 10670 13125 10730 13525
rect 10866 13325 10926 13525
rect 13268 13325 13328 13525
rect 13460 13125 13520 13525
rect 13578 13125 13638 13525
rect 13696 13125 13756 13525
rect 13814 13125 13874 13525
rect 14010 13325 14070 13525
rect 16470 13321 16530 13521
rect 16662 13121 16722 13521
rect 16780 13121 16840 13521
rect 16898 13121 16958 13521
rect 17016 13121 17076 13521
rect 17212 13321 17272 13521
rect 19614 13321 19674 13521
rect 19806 13121 19866 13521
rect 19924 13121 19984 13521
rect 20042 13121 20102 13521
rect 20160 13121 20220 13521
rect 20356 13321 20416 13521
rect 22746 13325 22806 13525
rect 22938 13125 22998 13525
rect 23056 13125 23116 13525
rect 23174 13125 23234 13525
rect 23292 13125 23352 13525
rect 23488 13325 23548 13525
rect 25890 13325 25950 13525
rect 26082 13125 26142 13525
rect 26200 13125 26260 13525
rect 26318 13125 26378 13525
rect 26436 13125 26496 13525
rect 26632 13325 26692 13525
rect 3848 10587 3908 10787
rect 4040 10387 4100 10787
rect 4158 10387 4218 10787
rect 4276 10387 4336 10787
rect 4394 10387 4454 10787
rect 4590 10587 4650 10787
rect 6992 10587 7052 10787
rect 7184 10387 7244 10787
rect 7302 10387 7362 10787
rect 7420 10387 7480 10787
rect 7538 10387 7598 10787
rect 7734 10587 7794 10787
rect 10124 10591 10184 10791
rect 10316 10391 10376 10791
rect 10434 10391 10494 10791
rect 10552 10391 10612 10791
rect 10670 10391 10730 10791
rect 10866 10591 10926 10791
rect 13268 10591 13328 10791
rect 13460 10391 13520 10791
rect 13578 10391 13638 10791
rect 13696 10391 13756 10791
rect 13814 10391 13874 10791
rect 14010 10591 14070 10791
rect 16470 10587 16530 10787
rect 16662 10387 16722 10787
rect 16780 10387 16840 10787
rect 16898 10387 16958 10787
rect 17016 10387 17076 10787
rect 17212 10587 17272 10787
rect 19614 10587 19674 10787
rect 19806 10387 19866 10787
rect 19924 10387 19984 10787
rect 20042 10387 20102 10787
rect 20160 10387 20220 10787
rect 20356 10587 20416 10787
rect 22746 10591 22806 10791
rect 22938 10391 22998 10791
rect 23056 10391 23116 10791
rect 23174 10391 23234 10791
rect 23292 10391 23352 10791
rect 23488 10591 23548 10791
rect 25890 10591 25950 10791
rect 26082 10391 26142 10791
rect 26200 10391 26260 10791
rect 26318 10391 26378 10791
rect 26436 10391 26496 10791
rect 26632 10591 26692 10791
rect 3838 7855 3898 8055
rect 4030 7655 4090 8055
rect 4148 7655 4208 8055
rect 4266 7655 4326 8055
rect 4384 7655 4444 8055
rect 4580 7855 4640 8055
rect 6982 7855 7042 8055
rect 7174 7655 7234 8055
rect 7292 7655 7352 8055
rect 7410 7655 7470 8055
rect 7528 7655 7588 8055
rect 7724 7855 7784 8055
rect 10114 7859 10174 8059
rect 10306 7659 10366 8059
rect 10424 7659 10484 8059
rect 10542 7659 10602 8059
rect 10660 7659 10720 8059
rect 10856 7859 10916 8059
rect 13258 7859 13318 8059
rect 13450 7659 13510 8059
rect 13568 7659 13628 8059
rect 13686 7659 13746 8059
rect 13804 7659 13864 8059
rect 14000 7859 14060 8059
rect 16460 7855 16520 8055
rect 16652 7655 16712 8055
rect 16770 7655 16830 8055
rect 16888 7655 16948 8055
rect 17006 7655 17066 8055
rect 17202 7855 17262 8055
rect 19604 7855 19664 8055
rect 19796 7655 19856 8055
rect 19914 7655 19974 8055
rect 20032 7655 20092 8055
rect 20150 7655 20210 8055
rect 20346 7855 20406 8055
rect 22736 7859 22796 8059
rect 22928 7659 22988 8059
rect 23046 7659 23106 8059
rect 23164 7659 23224 8059
rect 23282 7659 23342 8059
rect 23478 7859 23538 8059
rect 25880 7859 25940 8059
rect 26072 7659 26132 8059
rect 26190 7659 26250 8059
rect 26308 7659 26368 8059
rect 26426 7659 26486 8059
rect 26622 7859 26682 8059
rect 2866 4818 2926 5018
rect 3286 4618 3346 5018
rect 3404 4618 3464 5018
rect 3522 4618 3582 5018
rect 3640 4618 3700 5018
rect 4164 4818 4224 5018
rect 4934 4820 4994 5020
rect 5354 4620 5414 5020
rect 5472 4620 5532 5020
rect 5590 4620 5650 5020
rect 5708 4620 5768 5020
rect 6232 4820 6292 5020
rect 7003 4818 7063 5018
rect 7423 4618 7483 5018
rect 7541 4618 7601 5018
rect 7659 4618 7719 5018
rect 7777 4618 7837 5018
rect 8301 4818 8361 5018
rect 9071 4820 9131 5020
rect 9491 4620 9551 5020
rect 9609 4620 9669 5020
rect 9727 4620 9787 5020
rect 9845 4620 9905 5020
rect 10369 4820 10429 5020
rect 11140 4820 11200 5020
rect 11560 4620 11620 5020
rect 11678 4620 11738 5020
rect 11796 4620 11856 5020
rect 11914 4620 11974 5020
rect 12438 4820 12498 5020
rect 13208 4822 13268 5022
rect 13628 4622 13688 5022
rect 13746 4622 13806 5022
rect 13864 4622 13924 5022
rect 13982 4622 14042 5022
rect 14506 4822 14566 5022
rect 19591 5973 19651 6173
rect 20329 5975 20389 6175
rect 21067 5971 21127 6171
rect 21809 5971 21869 6171
rect 22549 5971 22609 6171
rect 23287 5971 23347 6171
rect 24025 5975 24085 6175
rect 24763 5975 24823 6175
rect 15277 4820 15337 5020
rect 15697 4620 15757 5020
rect 15815 4620 15875 5020
rect 15933 4620 15993 5020
rect 16051 4620 16111 5020
rect 16575 4820 16635 5020
rect 17345 4822 17405 5022
rect 17765 4622 17825 5022
rect 17883 4622 17943 5022
rect 18001 4622 18061 5022
rect 18119 4622 18179 5022
rect 18643 4822 18703 5022
rect 1140 607 1200 807
rect 1332 407 1392 807
rect 1450 407 1510 807
rect 1568 407 1628 807
rect 1686 407 1746 807
rect 1882 607 1942 807
rect 4284 607 4344 807
rect 4476 407 4536 807
rect 4594 407 4654 807
rect 4712 407 4772 807
rect 4830 407 4890 807
rect 5026 607 5086 807
rect 7416 611 7476 811
rect 7608 411 7668 811
rect 7726 411 7786 811
rect 7844 411 7904 811
rect 7962 411 8022 811
rect 8158 611 8218 811
rect 10560 611 10620 811
rect 10752 411 10812 811
rect 10870 411 10930 811
rect 10988 411 11048 811
rect 11106 411 11166 811
rect 11302 611 11362 811
rect 13762 607 13822 807
rect 13954 407 14014 807
rect 14072 407 14132 807
rect 14190 407 14250 807
rect 14308 407 14368 807
rect 14504 607 14564 807
rect 16906 607 16966 807
rect 17098 407 17158 807
rect 17216 407 17276 807
rect 17334 407 17394 807
rect 17452 407 17512 807
rect 17648 607 17708 807
rect 20038 611 20098 811
rect 20230 411 20290 811
rect 20348 411 20408 811
rect 20466 411 20526 811
rect 20584 411 20644 811
rect 20780 611 20840 811
rect 23182 611 23242 811
rect 23374 411 23434 811
rect 23492 411 23552 811
rect 23610 411 23670 811
rect 23728 411 23788 811
rect 23924 611 23984 811
rect 1172 -3285 1232 -3085
rect 1364 -3485 1424 -3085
rect 1482 -3485 1542 -3085
rect 1600 -3485 1660 -3085
rect 1718 -3485 1778 -3085
rect 1914 -3285 1974 -3085
rect 4316 -3285 4376 -3085
rect 4508 -3485 4568 -3085
rect 4626 -3485 4686 -3085
rect 4744 -3485 4804 -3085
rect 4862 -3485 4922 -3085
rect 5058 -3285 5118 -3085
rect 7448 -3281 7508 -3081
rect 7640 -3481 7700 -3081
rect 7758 -3481 7818 -3081
rect 7876 -3481 7936 -3081
rect 7994 -3481 8054 -3081
rect 8190 -3281 8250 -3081
rect 10592 -3281 10652 -3081
rect 10784 -3481 10844 -3081
rect 10902 -3481 10962 -3081
rect 11020 -3481 11080 -3081
rect 11138 -3481 11198 -3081
rect 11334 -3281 11394 -3081
rect 13794 -3285 13854 -3085
rect 13986 -3485 14046 -3085
rect 14104 -3485 14164 -3085
rect 14222 -3485 14282 -3085
rect 14340 -3485 14400 -3085
rect 14536 -3285 14596 -3085
rect 16938 -3285 16998 -3085
rect 17130 -3485 17190 -3085
rect 17248 -3485 17308 -3085
rect 17366 -3485 17426 -3085
rect 17484 -3485 17544 -3085
rect 17680 -3285 17740 -3085
rect 20070 -3281 20130 -3081
rect 20262 -3481 20322 -3081
rect 20380 -3481 20440 -3081
rect 20498 -3481 20558 -3081
rect 20616 -3481 20676 -3081
rect 20812 -3281 20872 -3081
rect 23214 -3281 23274 -3081
rect 23406 -3481 23466 -3081
rect 23524 -3481 23584 -3081
rect 23642 -3481 23702 -3081
rect 23760 -3481 23820 -3081
rect 23956 -3281 24016 -3081
<< pmos >>
rect 512 21592 572 21792
rect 630 21592 690 21792
rect 748 21592 808 21792
rect 953 21592 1013 21992
rect 1071 21592 1131 21992
rect 1189 21592 1249 21992
rect 1420 21592 1480 21992
rect 1538 21592 1598 21992
rect 1656 21592 1716 21992
rect 1774 21592 1834 21992
rect 1892 21592 1952 21992
rect 2010 21592 2070 21992
rect 2247 21592 2307 21992
rect 2365 21592 2425 21992
rect 2483 21592 2543 21992
rect 2720 21592 2780 21792
rect 2838 21592 2898 21792
rect 2956 21592 3016 21792
rect 3656 21592 3716 21792
rect 3774 21592 3834 21792
rect 3892 21592 3952 21792
rect 4097 21592 4157 21992
rect 4215 21592 4275 21992
rect 4333 21592 4393 21992
rect 4564 21592 4624 21992
rect 4682 21592 4742 21992
rect 4800 21592 4860 21992
rect 4918 21592 4978 21992
rect 5036 21592 5096 21992
rect 5154 21592 5214 21992
rect 5391 21592 5451 21992
rect 5509 21592 5569 21992
rect 5627 21592 5687 21992
rect 5864 21592 5924 21792
rect 5982 21592 6042 21792
rect 6100 21592 6160 21792
rect 6788 21596 6848 21796
rect 6906 21596 6966 21796
rect 7024 21596 7084 21796
rect 7229 21596 7289 21996
rect 7347 21596 7407 21996
rect 7465 21596 7525 21996
rect 7696 21596 7756 21996
rect 7814 21596 7874 21996
rect 7932 21596 7992 21996
rect 8050 21596 8110 21996
rect 8168 21596 8228 21996
rect 8286 21596 8346 21996
rect 8523 21596 8583 21996
rect 8641 21596 8701 21996
rect 8759 21596 8819 21996
rect 8996 21596 9056 21796
rect 9114 21596 9174 21796
rect 9232 21596 9292 21796
rect 9932 21596 9992 21796
rect 10050 21596 10110 21796
rect 10168 21596 10228 21796
rect 10373 21596 10433 21996
rect 10491 21596 10551 21996
rect 10609 21596 10669 21996
rect 10840 21596 10900 21996
rect 10958 21596 11018 21996
rect 11076 21596 11136 21996
rect 11194 21596 11254 21996
rect 11312 21596 11372 21996
rect 11430 21596 11490 21996
rect 11667 21596 11727 21996
rect 11785 21596 11845 21996
rect 11903 21596 11963 21996
rect 12140 21596 12200 21796
rect 12258 21596 12318 21796
rect 12376 21596 12436 21796
rect 13134 21592 13194 21792
rect 13252 21592 13312 21792
rect 13370 21592 13430 21792
rect 13575 21592 13635 21992
rect 13693 21592 13753 21992
rect 13811 21592 13871 21992
rect 14042 21592 14102 21992
rect 14160 21592 14220 21992
rect 14278 21592 14338 21992
rect 14396 21592 14456 21992
rect 14514 21592 14574 21992
rect 14632 21592 14692 21992
rect 14869 21592 14929 21992
rect 14987 21592 15047 21992
rect 15105 21592 15165 21992
rect 15342 21592 15402 21792
rect 15460 21592 15520 21792
rect 15578 21592 15638 21792
rect 16278 21592 16338 21792
rect 16396 21592 16456 21792
rect 16514 21592 16574 21792
rect 16719 21592 16779 21992
rect 16837 21592 16897 21992
rect 16955 21592 17015 21992
rect 17186 21592 17246 21992
rect 17304 21592 17364 21992
rect 17422 21592 17482 21992
rect 17540 21592 17600 21992
rect 17658 21592 17718 21992
rect 17776 21592 17836 21992
rect 18013 21592 18073 21992
rect 18131 21592 18191 21992
rect 18249 21592 18309 21992
rect 18486 21592 18546 21792
rect 18604 21592 18664 21792
rect 18722 21592 18782 21792
rect 19410 21596 19470 21796
rect 19528 21596 19588 21796
rect 19646 21596 19706 21796
rect 19851 21596 19911 21996
rect 19969 21596 20029 21996
rect 20087 21596 20147 21996
rect 20318 21596 20378 21996
rect 20436 21596 20496 21996
rect 20554 21596 20614 21996
rect 20672 21596 20732 21996
rect 20790 21596 20850 21996
rect 20908 21596 20968 21996
rect 21145 21596 21205 21996
rect 21263 21596 21323 21996
rect 21381 21596 21441 21996
rect 21618 21596 21678 21796
rect 21736 21596 21796 21796
rect 21854 21596 21914 21796
rect 22554 21596 22614 21796
rect 22672 21596 22732 21796
rect 22790 21596 22850 21796
rect 22995 21596 23055 21996
rect 23113 21596 23173 21996
rect 23231 21596 23291 21996
rect 23462 21596 23522 21996
rect 23580 21596 23640 21996
rect 23698 21596 23758 21996
rect 23816 21596 23876 21996
rect 23934 21596 23994 21996
rect 24052 21596 24112 21996
rect 24289 21596 24349 21996
rect 24407 21596 24467 21996
rect 24525 21596 24585 21996
rect 24762 21596 24822 21796
rect 24880 21596 24940 21796
rect 24998 21596 25058 21796
rect 2955 16411 3015 16611
rect 3073 16411 3133 16611
rect 3191 16411 3251 16611
rect 3309 16411 3369 16611
rect 3427 16411 3487 16611
rect 3545 16411 3605 16611
rect 3663 16411 3723 16611
rect 3781 16411 3841 16611
rect 3899 16411 3959 16611
rect 4403 16411 4463 16611
rect 4521 16411 4581 16611
rect 4639 16411 4699 16611
rect 4757 16411 4817 16611
rect 4875 16411 4935 16611
rect 4993 16411 5053 16611
rect 5111 16411 5171 16611
rect 5229 16411 5289 16611
rect 5347 16411 5407 16611
rect 5901 16413 5961 16613
rect 6019 16413 6079 16613
rect 6137 16413 6197 16613
rect 6255 16413 6315 16613
rect 6373 16413 6433 16613
rect 6491 16413 6551 16613
rect 6609 16413 6669 16613
rect 6727 16413 6787 16613
rect 6845 16413 6905 16613
rect 7349 16413 7409 16613
rect 7467 16413 7527 16613
rect 7585 16413 7645 16613
rect 7703 16413 7763 16613
rect 7821 16413 7881 16613
rect 7939 16413 7999 16613
rect 8057 16413 8117 16613
rect 8175 16413 8235 16613
rect 8293 16413 8353 16613
rect 8869 16411 8929 16611
rect 8987 16411 9047 16611
rect 9105 16411 9165 16611
rect 9223 16411 9283 16611
rect 9341 16411 9401 16611
rect 9459 16411 9519 16611
rect 9577 16411 9637 16611
rect 9695 16411 9755 16611
rect 9813 16411 9873 16611
rect 10317 16411 10377 16611
rect 10435 16411 10495 16611
rect 10553 16411 10613 16611
rect 10671 16411 10731 16611
rect 10789 16411 10849 16611
rect 10907 16411 10967 16611
rect 11025 16411 11085 16611
rect 11143 16411 11203 16611
rect 11261 16411 11321 16611
rect 11815 16413 11875 16613
rect 11933 16413 11993 16613
rect 12051 16413 12111 16613
rect 12169 16413 12229 16613
rect 12287 16413 12347 16613
rect 12405 16413 12465 16613
rect 12523 16413 12583 16613
rect 12641 16413 12701 16613
rect 12759 16413 12819 16613
rect 13263 16413 13323 16613
rect 13381 16413 13441 16613
rect 13499 16413 13559 16613
rect 13617 16413 13677 16613
rect 13735 16413 13795 16613
rect 13853 16413 13913 16613
rect 13971 16413 14031 16613
rect 14089 16413 14149 16613
rect 14207 16413 14267 16613
rect 14718 16408 14778 16808
rect 14836 16408 14896 16808
rect 14954 16408 15014 16808
rect 15072 16408 15132 16808
rect 15190 16408 15250 16808
rect 15308 16408 15368 16808
rect 15886 16408 15946 16808
rect 16004 16408 16064 16808
rect 16122 16408 16182 16808
rect 16240 16408 16300 16808
rect 16358 16408 16418 16808
rect 16476 16408 16536 16808
rect 17054 16406 17114 16806
rect 17172 16406 17232 16806
rect 17290 16406 17350 16806
rect 17408 16406 17468 16806
rect 17526 16406 17586 16806
rect 17644 16406 17704 16806
rect 18222 16408 18282 16808
rect 18340 16408 18400 16808
rect 18458 16408 18518 16808
rect 18576 16408 18636 16808
rect 18694 16408 18754 16808
rect 18812 16408 18872 16808
rect 19396 16410 19456 16810
rect 19514 16410 19574 16810
rect 19632 16410 19692 16810
rect 19750 16410 19810 16810
rect 19868 16410 19928 16810
rect 19986 16410 20046 16810
rect 20564 16408 20624 16808
rect 20682 16408 20742 16808
rect 20800 16408 20860 16808
rect 20918 16408 20978 16808
rect 21036 16408 21096 16808
rect 21154 16408 21214 16808
rect 21732 16410 21792 16810
rect 21850 16410 21910 16810
rect 21968 16410 22028 16810
rect 22086 16410 22146 16810
rect 22204 16410 22264 16810
rect 22322 16410 22382 16810
rect 15148 15818 15208 16018
rect 15266 15818 15326 16018
rect 15384 15818 15444 16018
rect 16315 15824 16375 16024
rect 16433 15824 16493 16024
rect 16551 15824 16611 16024
rect 17483 15824 17543 16024
rect 17601 15824 17661 16024
rect 17719 15824 17779 16024
rect 18652 15824 18712 16024
rect 18770 15824 18830 16024
rect 18888 15824 18948 16024
rect 19824 15820 19884 16020
rect 19942 15820 20002 16020
rect 20060 15820 20120 16020
rect 22900 16408 22960 16808
rect 23018 16408 23078 16808
rect 23136 16408 23196 16808
rect 23254 16408 23314 16808
rect 23372 16408 23432 16808
rect 23490 16408 23550 16808
rect 20993 15819 21053 16019
rect 21111 15819 21171 16019
rect 21229 15819 21289 16019
rect 22161 15819 22221 16019
rect 22279 15819 22339 16019
rect 22397 15819 22457 16019
rect 23329 15820 23389 16020
rect 23447 15820 23507 16020
rect 23565 15820 23625 16020
rect 3014 14454 3074 14654
rect 3132 14454 3192 14654
rect 3250 14454 3310 14654
rect 3455 14454 3515 14854
rect 3573 14454 3633 14854
rect 3691 14454 3751 14854
rect 3922 14454 3982 14854
rect 4040 14454 4100 14854
rect 4158 14454 4218 14854
rect 4276 14454 4336 14854
rect 4394 14454 4454 14854
rect 4512 14454 4572 14854
rect 4749 14454 4809 14854
rect 4867 14454 4927 14854
rect 4985 14454 5045 14854
rect 5222 14454 5282 14654
rect 5340 14454 5400 14654
rect 5458 14454 5518 14654
rect 6158 14454 6218 14654
rect 6276 14454 6336 14654
rect 6394 14454 6454 14654
rect 6599 14454 6659 14854
rect 6717 14454 6777 14854
rect 6835 14454 6895 14854
rect 7066 14454 7126 14854
rect 7184 14454 7244 14854
rect 7302 14454 7362 14854
rect 7420 14454 7480 14854
rect 7538 14454 7598 14854
rect 7656 14454 7716 14854
rect 7893 14454 7953 14854
rect 8011 14454 8071 14854
rect 8129 14454 8189 14854
rect 8366 14454 8426 14654
rect 8484 14454 8544 14654
rect 8602 14454 8662 14654
rect 9290 14458 9350 14658
rect 9408 14458 9468 14658
rect 9526 14458 9586 14658
rect 9731 14458 9791 14858
rect 9849 14458 9909 14858
rect 9967 14458 10027 14858
rect 10198 14458 10258 14858
rect 10316 14458 10376 14858
rect 10434 14458 10494 14858
rect 10552 14458 10612 14858
rect 10670 14458 10730 14858
rect 10788 14458 10848 14858
rect 11025 14458 11085 14858
rect 11143 14458 11203 14858
rect 11261 14458 11321 14858
rect 11498 14458 11558 14658
rect 11616 14458 11676 14658
rect 11734 14458 11794 14658
rect 12434 14458 12494 14658
rect 12552 14458 12612 14658
rect 12670 14458 12730 14658
rect 12875 14458 12935 14858
rect 12993 14458 13053 14858
rect 13111 14458 13171 14858
rect 13342 14458 13402 14858
rect 13460 14458 13520 14858
rect 13578 14458 13638 14858
rect 13696 14458 13756 14858
rect 13814 14458 13874 14858
rect 13932 14458 13992 14858
rect 14169 14458 14229 14858
rect 14287 14458 14347 14858
rect 14405 14458 14465 14858
rect 14642 14458 14702 14658
rect 14760 14458 14820 14658
rect 14878 14458 14938 14658
rect 15636 14454 15696 14654
rect 15754 14454 15814 14654
rect 15872 14454 15932 14654
rect 16077 14454 16137 14854
rect 16195 14454 16255 14854
rect 16313 14454 16373 14854
rect 16544 14454 16604 14854
rect 16662 14454 16722 14854
rect 16780 14454 16840 14854
rect 16898 14454 16958 14854
rect 17016 14454 17076 14854
rect 17134 14454 17194 14854
rect 17371 14454 17431 14854
rect 17489 14454 17549 14854
rect 17607 14454 17667 14854
rect 17844 14454 17904 14654
rect 17962 14454 18022 14654
rect 18080 14454 18140 14654
rect 18780 14454 18840 14654
rect 18898 14454 18958 14654
rect 19016 14454 19076 14654
rect 19221 14454 19281 14854
rect 19339 14454 19399 14854
rect 19457 14454 19517 14854
rect 19688 14454 19748 14854
rect 19806 14454 19866 14854
rect 19924 14454 19984 14854
rect 20042 14454 20102 14854
rect 20160 14454 20220 14854
rect 20278 14454 20338 14854
rect 20515 14454 20575 14854
rect 20633 14454 20693 14854
rect 20751 14454 20811 14854
rect 20988 14454 21048 14654
rect 21106 14454 21166 14654
rect 21224 14454 21284 14654
rect 21912 14458 21972 14658
rect 22030 14458 22090 14658
rect 22148 14458 22208 14658
rect 22353 14458 22413 14858
rect 22471 14458 22531 14858
rect 22589 14458 22649 14858
rect 22820 14458 22880 14858
rect 22938 14458 22998 14858
rect 23056 14458 23116 14858
rect 23174 14458 23234 14858
rect 23292 14458 23352 14858
rect 23410 14458 23470 14858
rect 23647 14458 23707 14858
rect 23765 14458 23825 14858
rect 23883 14458 23943 14858
rect 24120 14458 24180 14658
rect 24238 14458 24298 14658
rect 24356 14458 24416 14658
rect 25056 14458 25116 14658
rect 25174 14458 25234 14658
rect 25292 14458 25352 14658
rect 25497 14458 25557 14858
rect 25615 14458 25675 14858
rect 25733 14458 25793 14858
rect 25964 14458 26024 14858
rect 26082 14458 26142 14858
rect 26200 14458 26260 14858
rect 26318 14458 26378 14858
rect 26436 14458 26496 14858
rect 26554 14458 26614 14858
rect 26791 14458 26851 14858
rect 26909 14458 26969 14858
rect 27027 14458 27087 14858
rect 27264 14458 27324 14658
rect 27382 14458 27442 14658
rect 27500 14458 27560 14658
rect 3014 11720 3074 11920
rect 3132 11720 3192 11920
rect 3250 11720 3310 11920
rect 3455 11720 3515 12120
rect 3573 11720 3633 12120
rect 3691 11720 3751 12120
rect 3922 11720 3982 12120
rect 4040 11720 4100 12120
rect 4158 11720 4218 12120
rect 4276 11720 4336 12120
rect 4394 11720 4454 12120
rect 4512 11720 4572 12120
rect 4749 11720 4809 12120
rect 4867 11720 4927 12120
rect 4985 11720 5045 12120
rect 5222 11720 5282 11920
rect 5340 11720 5400 11920
rect 5458 11720 5518 11920
rect 6158 11720 6218 11920
rect 6276 11720 6336 11920
rect 6394 11720 6454 11920
rect 6599 11720 6659 12120
rect 6717 11720 6777 12120
rect 6835 11720 6895 12120
rect 7066 11720 7126 12120
rect 7184 11720 7244 12120
rect 7302 11720 7362 12120
rect 7420 11720 7480 12120
rect 7538 11720 7598 12120
rect 7656 11720 7716 12120
rect 7893 11720 7953 12120
rect 8011 11720 8071 12120
rect 8129 11720 8189 12120
rect 8366 11720 8426 11920
rect 8484 11720 8544 11920
rect 8602 11720 8662 11920
rect 9290 11724 9350 11924
rect 9408 11724 9468 11924
rect 9526 11724 9586 11924
rect 9731 11724 9791 12124
rect 9849 11724 9909 12124
rect 9967 11724 10027 12124
rect 10198 11724 10258 12124
rect 10316 11724 10376 12124
rect 10434 11724 10494 12124
rect 10552 11724 10612 12124
rect 10670 11724 10730 12124
rect 10788 11724 10848 12124
rect 11025 11724 11085 12124
rect 11143 11724 11203 12124
rect 11261 11724 11321 12124
rect 11498 11724 11558 11924
rect 11616 11724 11676 11924
rect 11734 11724 11794 11924
rect 12434 11724 12494 11924
rect 12552 11724 12612 11924
rect 12670 11724 12730 11924
rect 12875 11724 12935 12124
rect 12993 11724 13053 12124
rect 13111 11724 13171 12124
rect 13342 11724 13402 12124
rect 13460 11724 13520 12124
rect 13578 11724 13638 12124
rect 13696 11724 13756 12124
rect 13814 11724 13874 12124
rect 13932 11724 13992 12124
rect 14169 11724 14229 12124
rect 14287 11724 14347 12124
rect 14405 11724 14465 12124
rect 14642 11724 14702 11924
rect 14760 11724 14820 11924
rect 14878 11724 14938 11924
rect 15636 11720 15696 11920
rect 15754 11720 15814 11920
rect 15872 11720 15932 11920
rect 16077 11720 16137 12120
rect 16195 11720 16255 12120
rect 16313 11720 16373 12120
rect 16544 11720 16604 12120
rect 16662 11720 16722 12120
rect 16780 11720 16840 12120
rect 16898 11720 16958 12120
rect 17016 11720 17076 12120
rect 17134 11720 17194 12120
rect 17371 11720 17431 12120
rect 17489 11720 17549 12120
rect 17607 11720 17667 12120
rect 17844 11720 17904 11920
rect 17962 11720 18022 11920
rect 18080 11720 18140 11920
rect 18780 11720 18840 11920
rect 18898 11720 18958 11920
rect 19016 11720 19076 11920
rect 19221 11720 19281 12120
rect 19339 11720 19399 12120
rect 19457 11720 19517 12120
rect 19688 11720 19748 12120
rect 19806 11720 19866 12120
rect 19924 11720 19984 12120
rect 20042 11720 20102 12120
rect 20160 11720 20220 12120
rect 20278 11720 20338 12120
rect 20515 11720 20575 12120
rect 20633 11720 20693 12120
rect 20751 11720 20811 12120
rect 20988 11720 21048 11920
rect 21106 11720 21166 11920
rect 21224 11720 21284 11920
rect 21912 11724 21972 11924
rect 22030 11724 22090 11924
rect 22148 11724 22208 11924
rect 22353 11724 22413 12124
rect 22471 11724 22531 12124
rect 22589 11724 22649 12124
rect 22820 11724 22880 12124
rect 22938 11724 22998 12124
rect 23056 11724 23116 12124
rect 23174 11724 23234 12124
rect 23292 11724 23352 12124
rect 23410 11724 23470 12124
rect 23647 11724 23707 12124
rect 23765 11724 23825 12124
rect 23883 11724 23943 12124
rect 24120 11724 24180 11924
rect 24238 11724 24298 11924
rect 24356 11724 24416 11924
rect 25056 11724 25116 11924
rect 25174 11724 25234 11924
rect 25292 11724 25352 11924
rect 25497 11724 25557 12124
rect 25615 11724 25675 12124
rect 25733 11724 25793 12124
rect 25964 11724 26024 12124
rect 26082 11724 26142 12124
rect 26200 11724 26260 12124
rect 26318 11724 26378 12124
rect 26436 11724 26496 12124
rect 26554 11724 26614 12124
rect 26791 11724 26851 12124
rect 26909 11724 26969 12124
rect 27027 11724 27087 12124
rect 27264 11724 27324 11924
rect 27382 11724 27442 11924
rect 27500 11724 27560 11924
rect 3004 8988 3064 9188
rect 3122 8988 3182 9188
rect 3240 8988 3300 9188
rect 3445 8988 3505 9388
rect 3563 8988 3623 9388
rect 3681 8988 3741 9388
rect 3912 8988 3972 9388
rect 4030 8988 4090 9388
rect 4148 8988 4208 9388
rect 4266 8988 4326 9388
rect 4384 8988 4444 9388
rect 4502 8988 4562 9388
rect 4739 8988 4799 9388
rect 4857 8988 4917 9388
rect 4975 8988 5035 9388
rect 5212 8988 5272 9188
rect 5330 8988 5390 9188
rect 5448 8988 5508 9188
rect 6148 8988 6208 9188
rect 6266 8988 6326 9188
rect 6384 8988 6444 9188
rect 6589 8988 6649 9388
rect 6707 8988 6767 9388
rect 6825 8988 6885 9388
rect 7056 8988 7116 9388
rect 7174 8988 7234 9388
rect 7292 8988 7352 9388
rect 7410 8988 7470 9388
rect 7528 8988 7588 9388
rect 7646 8988 7706 9388
rect 7883 8988 7943 9388
rect 8001 8988 8061 9388
rect 8119 8988 8179 9388
rect 8356 8988 8416 9188
rect 8474 8988 8534 9188
rect 8592 8988 8652 9188
rect 9280 8992 9340 9192
rect 9398 8992 9458 9192
rect 9516 8992 9576 9192
rect 9721 8992 9781 9392
rect 9839 8992 9899 9392
rect 9957 8992 10017 9392
rect 10188 8992 10248 9392
rect 10306 8992 10366 9392
rect 10424 8992 10484 9392
rect 10542 8992 10602 9392
rect 10660 8992 10720 9392
rect 10778 8992 10838 9392
rect 11015 8992 11075 9392
rect 11133 8992 11193 9392
rect 11251 8992 11311 9392
rect 11488 8992 11548 9192
rect 11606 8992 11666 9192
rect 11724 8992 11784 9192
rect 12424 8992 12484 9192
rect 12542 8992 12602 9192
rect 12660 8992 12720 9192
rect 12865 8992 12925 9392
rect 12983 8992 13043 9392
rect 13101 8992 13161 9392
rect 13332 8992 13392 9392
rect 13450 8992 13510 9392
rect 13568 8992 13628 9392
rect 13686 8992 13746 9392
rect 13804 8992 13864 9392
rect 13922 8992 13982 9392
rect 14159 8992 14219 9392
rect 14277 8992 14337 9392
rect 14395 8992 14455 9392
rect 14632 8992 14692 9192
rect 14750 8992 14810 9192
rect 14868 8992 14928 9192
rect 15626 8988 15686 9188
rect 15744 8988 15804 9188
rect 15862 8988 15922 9188
rect 16067 8988 16127 9388
rect 16185 8988 16245 9388
rect 16303 8988 16363 9388
rect 16534 8988 16594 9388
rect 16652 8988 16712 9388
rect 16770 8988 16830 9388
rect 16888 8988 16948 9388
rect 17006 8988 17066 9388
rect 17124 8988 17184 9388
rect 17361 8988 17421 9388
rect 17479 8988 17539 9388
rect 17597 8988 17657 9388
rect 17834 8988 17894 9188
rect 17952 8988 18012 9188
rect 18070 8988 18130 9188
rect 18770 8988 18830 9188
rect 18888 8988 18948 9188
rect 19006 8988 19066 9188
rect 19211 8988 19271 9388
rect 19329 8988 19389 9388
rect 19447 8988 19507 9388
rect 19678 8988 19738 9388
rect 19796 8988 19856 9388
rect 19914 8988 19974 9388
rect 20032 8988 20092 9388
rect 20150 8988 20210 9388
rect 20268 8988 20328 9388
rect 20505 8988 20565 9388
rect 20623 8988 20683 9388
rect 20741 8988 20801 9388
rect 20978 8988 21038 9188
rect 21096 8988 21156 9188
rect 21214 8988 21274 9188
rect 21902 8992 21962 9192
rect 22020 8992 22080 9192
rect 22138 8992 22198 9192
rect 22343 8992 22403 9392
rect 22461 8992 22521 9392
rect 22579 8992 22639 9392
rect 22810 8992 22870 9392
rect 22928 8992 22988 9392
rect 23046 8992 23106 9392
rect 23164 8992 23224 9392
rect 23282 8992 23342 9392
rect 23400 8992 23460 9392
rect 23637 8992 23697 9392
rect 23755 8992 23815 9392
rect 23873 8992 23933 9392
rect 24110 8992 24170 9192
rect 24228 8992 24288 9192
rect 24346 8992 24406 9192
rect 25046 8992 25106 9192
rect 25164 8992 25224 9192
rect 25282 8992 25342 9192
rect 25487 8992 25547 9392
rect 25605 8992 25665 9392
rect 25723 8992 25783 9392
rect 25954 8992 26014 9392
rect 26072 8992 26132 9392
rect 26190 8992 26250 9392
rect 26308 8992 26368 9392
rect 26426 8992 26486 9392
rect 26544 8992 26604 9392
rect 26781 8992 26841 9392
rect 26899 8992 26959 9392
rect 27017 8992 27077 9392
rect 27254 8992 27314 9192
rect 27372 8992 27432 9192
rect 27490 8992 27550 9192
rect 2741 6043 2801 6243
rect 2859 6043 2919 6243
rect 2977 6043 3037 6243
rect 3225 6043 3285 6443
rect 3343 6043 3403 6443
rect 3461 6043 3521 6443
rect 3579 6043 3639 6443
rect 3697 6043 3757 6443
rect 3815 6043 3875 6443
rect 4062 6043 4122 6243
rect 4180 6043 4240 6243
rect 4298 6043 4358 6243
rect 4809 6045 4869 6245
rect 4927 6045 4987 6245
rect 5045 6045 5105 6245
rect 5293 6045 5353 6445
rect 5411 6045 5471 6445
rect 5529 6045 5589 6445
rect 5647 6045 5707 6445
rect 5765 6045 5825 6445
rect 5883 6045 5943 6445
rect 6130 6045 6190 6245
rect 6248 6045 6308 6245
rect 6366 6045 6426 6245
rect 3168 5350 3228 5750
rect 3286 5350 3346 5750
rect 3404 5350 3464 5750
rect 3522 5350 3582 5750
rect 3640 5350 3700 5750
rect 3758 5350 3818 5750
rect 6878 6043 6938 6243
rect 6996 6043 7056 6243
rect 7114 6043 7174 6243
rect 7362 6043 7422 6443
rect 7480 6043 7540 6443
rect 7598 6043 7658 6443
rect 7716 6043 7776 6443
rect 7834 6043 7894 6443
rect 7952 6043 8012 6443
rect 8199 6043 8259 6243
rect 8317 6043 8377 6243
rect 8435 6043 8495 6243
rect 8946 6045 9006 6245
rect 9064 6045 9124 6245
rect 9182 6045 9242 6245
rect 9430 6045 9490 6445
rect 9548 6045 9608 6445
rect 9666 6045 9726 6445
rect 9784 6045 9844 6445
rect 9902 6045 9962 6445
rect 10020 6045 10080 6445
rect 10267 6045 10327 6245
rect 10385 6045 10445 6245
rect 10503 6045 10563 6245
rect 11015 6045 11075 6245
rect 11133 6045 11193 6245
rect 11251 6045 11311 6245
rect 11499 6045 11559 6445
rect 11617 6045 11677 6445
rect 11735 6045 11795 6445
rect 11853 6045 11913 6445
rect 11971 6045 12031 6445
rect 12089 6045 12149 6445
rect 12336 6045 12396 6245
rect 12454 6045 12514 6245
rect 12572 6045 12632 6245
rect 13083 6047 13143 6247
rect 13201 6047 13261 6247
rect 13319 6047 13379 6247
rect 13567 6047 13627 6447
rect 13685 6047 13745 6447
rect 13803 6047 13863 6447
rect 13921 6047 13981 6447
rect 14039 6047 14099 6447
rect 14157 6047 14217 6447
rect 14404 6047 14464 6247
rect 14522 6047 14582 6247
rect 14640 6047 14700 6247
rect 5236 5352 5296 5752
rect 5354 5352 5414 5752
rect 5472 5352 5532 5752
rect 5590 5352 5650 5752
rect 5708 5352 5768 5752
rect 5826 5352 5886 5752
rect 7305 5350 7365 5750
rect 7423 5350 7483 5750
rect 7541 5350 7601 5750
rect 7659 5350 7719 5750
rect 7777 5350 7837 5750
rect 7895 5350 7955 5750
rect 9373 5352 9433 5752
rect 9491 5352 9551 5752
rect 9609 5352 9669 5752
rect 9727 5352 9787 5752
rect 9845 5352 9905 5752
rect 9963 5352 10023 5752
rect 11442 5352 11502 5752
rect 11560 5352 11620 5752
rect 11678 5352 11738 5752
rect 11796 5352 11856 5752
rect 11914 5352 11974 5752
rect 12032 5352 12092 5752
rect 15152 6045 15212 6245
rect 15270 6045 15330 6245
rect 15388 6045 15448 6245
rect 15636 6045 15696 6445
rect 15754 6045 15814 6445
rect 15872 6045 15932 6445
rect 15990 6045 16050 6445
rect 16108 6045 16168 6445
rect 16226 6045 16286 6445
rect 16473 6045 16533 6245
rect 16591 6045 16651 6245
rect 16709 6045 16769 6245
rect 17220 6047 17280 6247
rect 17338 6047 17398 6247
rect 17456 6047 17516 6247
rect 17704 6047 17764 6447
rect 17822 6047 17882 6447
rect 17940 6047 18000 6447
rect 18058 6047 18118 6447
rect 18176 6047 18236 6447
rect 18294 6047 18354 6447
rect 19473 6359 19533 6559
rect 19591 6359 19651 6559
rect 19709 6359 19769 6559
rect 20211 6363 20271 6563
rect 20329 6363 20389 6563
rect 20447 6363 20507 6563
rect 20949 6359 21009 6559
rect 21067 6359 21127 6559
rect 21185 6359 21245 6559
rect 21691 6357 21751 6557
rect 21809 6357 21869 6557
rect 21927 6357 21987 6557
rect 22431 6357 22491 6557
rect 22549 6357 22609 6557
rect 22667 6357 22727 6557
rect 23169 6357 23229 6557
rect 23287 6357 23347 6557
rect 23405 6357 23465 6557
rect 23907 6357 23967 6557
rect 24025 6357 24085 6557
rect 24143 6357 24203 6557
rect 24645 6357 24705 6557
rect 24763 6357 24823 6557
rect 24881 6357 24941 6557
rect 18541 6047 18601 6247
rect 18659 6047 18719 6247
rect 18777 6047 18837 6247
rect 13510 5354 13570 5754
rect 13628 5354 13688 5754
rect 13746 5354 13806 5754
rect 13864 5354 13924 5754
rect 13982 5354 14042 5754
rect 14100 5354 14160 5754
rect 15579 5352 15639 5752
rect 15697 5352 15757 5752
rect 15815 5352 15875 5752
rect 15933 5352 15993 5752
rect 16051 5352 16111 5752
rect 16169 5352 16229 5752
rect 17647 5354 17707 5754
rect 17765 5354 17825 5754
rect 17883 5354 17943 5754
rect 18001 5354 18061 5754
rect 18119 5354 18179 5754
rect 18237 5354 18297 5754
rect 306 1740 366 1940
rect 424 1740 484 1940
rect 542 1740 602 1940
rect 747 1740 807 2140
rect 865 1740 925 2140
rect 983 1740 1043 2140
rect 1214 1740 1274 2140
rect 1332 1740 1392 2140
rect 1450 1740 1510 2140
rect 1568 1740 1628 2140
rect 1686 1740 1746 2140
rect 1804 1740 1864 2140
rect 2041 1740 2101 2140
rect 2159 1740 2219 2140
rect 2277 1740 2337 2140
rect 2514 1740 2574 1940
rect 2632 1740 2692 1940
rect 2750 1740 2810 1940
rect 3450 1740 3510 1940
rect 3568 1740 3628 1940
rect 3686 1740 3746 1940
rect 3891 1740 3951 2140
rect 4009 1740 4069 2140
rect 4127 1740 4187 2140
rect 4358 1740 4418 2140
rect 4476 1740 4536 2140
rect 4594 1740 4654 2140
rect 4712 1740 4772 2140
rect 4830 1740 4890 2140
rect 4948 1740 5008 2140
rect 5185 1740 5245 2140
rect 5303 1740 5363 2140
rect 5421 1740 5481 2140
rect 5658 1740 5718 1940
rect 5776 1740 5836 1940
rect 5894 1740 5954 1940
rect 6582 1744 6642 1944
rect 6700 1744 6760 1944
rect 6818 1744 6878 1944
rect 7023 1744 7083 2144
rect 7141 1744 7201 2144
rect 7259 1744 7319 2144
rect 7490 1744 7550 2144
rect 7608 1744 7668 2144
rect 7726 1744 7786 2144
rect 7844 1744 7904 2144
rect 7962 1744 8022 2144
rect 8080 1744 8140 2144
rect 8317 1744 8377 2144
rect 8435 1744 8495 2144
rect 8553 1744 8613 2144
rect 8790 1744 8850 1944
rect 8908 1744 8968 1944
rect 9026 1744 9086 1944
rect 9726 1744 9786 1944
rect 9844 1744 9904 1944
rect 9962 1744 10022 1944
rect 10167 1744 10227 2144
rect 10285 1744 10345 2144
rect 10403 1744 10463 2144
rect 10634 1744 10694 2144
rect 10752 1744 10812 2144
rect 10870 1744 10930 2144
rect 10988 1744 11048 2144
rect 11106 1744 11166 2144
rect 11224 1744 11284 2144
rect 11461 1744 11521 2144
rect 11579 1744 11639 2144
rect 11697 1744 11757 2144
rect 11934 1744 11994 1944
rect 12052 1744 12112 1944
rect 12170 1744 12230 1944
rect 12928 1740 12988 1940
rect 13046 1740 13106 1940
rect 13164 1740 13224 1940
rect 13369 1740 13429 2140
rect 13487 1740 13547 2140
rect 13605 1740 13665 2140
rect 13836 1740 13896 2140
rect 13954 1740 14014 2140
rect 14072 1740 14132 2140
rect 14190 1740 14250 2140
rect 14308 1740 14368 2140
rect 14426 1740 14486 2140
rect 14663 1740 14723 2140
rect 14781 1740 14841 2140
rect 14899 1740 14959 2140
rect 15136 1740 15196 1940
rect 15254 1740 15314 1940
rect 15372 1740 15432 1940
rect 16072 1740 16132 1940
rect 16190 1740 16250 1940
rect 16308 1740 16368 1940
rect 16513 1740 16573 2140
rect 16631 1740 16691 2140
rect 16749 1740 16809 2140
rect 16980 1740 17040 2140
rect 17098 1740 17158 2140
rect 17216 1740 17276 2140
rect 17334 1740 17394 2140
rect 17452 1740 17512 2140
rect 17570 1740 17630 2140
rect 17807 1740 17867 2140
rect 17925 1740 17985 2140
rect 18043 1740 18103 2140
rect 18280 1740 18340 1940
rect 18398 1740 18458 1940
rect 18516 1740 18576 1940
rect 19204 1744 19264 1944
rect 19322 1744 19382 1944
rect 19440 1744 19500 1944
rect 19645 1744 19705 2144
rect 19763 1744 19823 2144
rect 19881 1744 19941 2144
rect 20112 1744 20172 2144
rect 20230 1744 20290 2144
rect 20348 1744 20408 2144
rect 20466 1744 20526 2144
rect 20584 1744 20644 2144
rect 20702 1744 20762 2144
rect 20939 1744 20999 2144
rect 21057 1744 21117 2144
rect 21175 1744 21235 2144
rect 21412 1744 21472 1944
rect 21530 1744 21590 1944
rect 21648 1744 21708 1944
rect 22348 1744 22408 1944
rect 22466 1744 22526 1944
rect 22584 1744 22644 1944
rect 22789 1744 22849 2144
rect 22907 1744 22967 2144
rect 23025 1744 23085 2144
rect 23256 1744 23316 2144
rect 23374 1744 23434 2144
rect 23492 1744 23552 2144
rect 23610 1744 23670 2144
rect 23728 1744 23788 2144
rect 23846 1744 23906 2144
rect 24083 1744 24143 2144
rect 24201 1744 24261 2144
rect 24319 1744 24379 2144
rect 24556 1744 24616 1944
rect 24674 1744 24734 1944
rect 24792 1744 24852 1944
rect 338 -2152 398 -1952
rect 456 -2152 516 -1952
rect 574 -2152 634 -1952
rect 779 -2152 839 -1752
rect 897 -2152 957 -1752
rect 1015 -2152 1075 -1752
rect 1246 -2152 1306 -1752
rect 1364 -2152 1424 -1752
rect 1482 -2152 1542 -1752
rect 1600 -2152 1660 -1752
rect 1718 -2152 1778 -1752
rect 1836 -2152 1896 -1752
rect 2073 -2152 2133 -1752
rect 2191 -2152 2251 -1752
rect 2309 -2152 2369 -1752
rect 2546 -2152 2606 -1952
rect 2664 -2152 2724 -1952
rect 2782 -2152 2842 -1952
rect 3482 -2152 3542 -1952
rect 3600 -2152 3660 -1952
rect 3718 -2152 3778 -1952
rect 3923 -2152 3983 -1752
rect 4041 -2152 4101 -1752
rect 4159 -2152 4219 -1752
rect 4390 -2152 4450 -1752
rect 4508 -2152 4568 -1752
rect 4626 -2152 4686 -1752
rect 4744 -2152 4804 -1752
rect 4862 -2152 4922 -1752
rect 4980 -2152 5040 -1752
rect 5217 -2152 5277 -1752
rect 5335 -2152 5395 -1752
rect 5453 -2152 5513 -1752
rect 5690 -2152 5750 -1952
rect 5808 -2152 5868 -1952
rect 5926 -2152 5986 -1952
rect 6614 -2148 6674 -1948
rect 6732 -2148 6792 -1948
rect 6850 -2148 6910 -1948
rect 7055 -2148 7115 -1748
rect 7173 -2148 7233 -1748
rect 7291 -2148 7351 -1748
rect 7522 -2148 7582 -1748
rect 7640 -2148 7700 -1748
rect 7758 -2148 7818 -1748
rect 7876 -2148 7936 -1748
rect 7994 -2148 8054 -1748
rect 8112 -2148 8172 -1748
rect 8349 -2148 8409 -1748
rect 8467 -2148 8527 -1748
rect 8585 -2148 8645 -1748
rect 8822 -2148 8882 -1948
rect 8940 -2148 9000 -1948
rect 9058 -2148 9118 -1948
rect 9758 -2148 9818 -1948
rect 9876 -2148 9936 -1948
rect 9994 -2148 10054 -1948
rect 10199 -2148 10259 -1748
rect 10317 -2148 10377 -1748
rect 10435 -2148 10495 -1748
rect 10666 -2148 10726 -1748
rect 10784 -2148 10844 -1748
rect 10902 -2148 10962 -1748
rect 11020 -2148 11080 -1748
rect 11138 -2148 11198 -1748
rect 11256 -2148 11316 -1748
rect 11493 -2148 11553 -1748
rect 11611 -2148 11671 -1748
rect 11729 -2148 11789 -1748
rect 11966 -2148 12026 -1948
rect 12084 -2148 12144 -1948
rect 12202 -2148 12262 -1948
rect 12960 -2152 13020 -1952
rect 13078 -2152 13138 -1952
rect 13196 -2152 13256 -1952
rect 13401 -2152 13461 -1752
rect 13519 -2152 13579 -1752
rect 13637 -2152 13697 -1752
rect 13868 -2152 13928 -1752
rect 13986 -2152 14046 -1752
rect 14104 -2152 14164 -1752
rect 14222 -2152 14282 -1752
rect 14340 -2152 14400 -1752
rect 14458 -2152 14518 -1752
rect 14695 -2152 14755 -1752
rect 14813 -2152 14873 -1752
rect 14931 -2152 14991 -1752
rect 15168 -2152 15228 -1952
rect 15286 -2152 15346 -1952
rect 15404 -2152 15464 -1952
rect 16104 -2152 16164 -1952
rect 16222 -2152 16282 -1952
rect 16340 -2152 16400 -1952
rect 16545 -2152 16605 -1752
rect 16663 -2152 16723 -1752
rect 16781 -2152 16841 -1752
rect 17012 -2152 17072 -1752
rect 17130 -2152 17190 -1752
rect 17248 -2152 17308 -1752
rect 17366 -2152 17426 -1752
rect 17484 -2152 17544 -1752
rect 17602 -2152 17662 -1752
rect 17839 -2152 17899 -1752
rect 17957 -2152 18017 -1752
rect 18075 -2152 18135 -1752
rect 18312 -2152 18372 -1952
rect 18430 -2152 18490 -1952
rect 18548 -2152 18608 -1952
rect 19236 -2148 19296 -1948
rect 19354 -2148 19414 -1948
rect 19472 -2148 19532 -1948
rect 19677 -2148 19737 -1748
rect 19795 -2148 19855 -1748
rect 19913 -2148 19973 -1748
rect 20144 -2148 20204 -1748
rect 20262 -2148 20322 -1748
rect 20380 -2148 20440 -1748
rect 20498 -2148 20558 -1748
rect 20616 -2148 20676 -1748
rect 20734 -2148 20794 -1748
rect 20971 -2148 21031 -1748
rect 21089 -2148 21149 -1748
rect 21207 -2148 21267 -1748
rect 21444 -2148 21504 -1948
rect 21562 -2148 21622 -1948
rect 21680 -2148 21740 -1948
rect 22380 -2148 22440 -1948
rect 22498 -2148 22558 -1948
rect 22616 -2148 22676 -1948
rect 22821 -2148 22881 -1748
rect 22939 -2148 22999 -1748
rect 23057 -2148 23117 -1748
rect 23288 -2148 23348 -1748
rect 23406 -2148 23466 -1748
rect 23524 -2148 23584 -1748
rect 23642 -2148 23702 -1748
rect 23760 -2148 23820 -1748
rect 23878 -2148 23938 -1748
rect 24115 -2148 24175 -1748
rect 24233 -2148 24293 -1748
rect 24351 -2148 24411 -1748
rect 24588 -2148 24648 -1948
rect 24706 -2148 24766 -1948
rect 24824 -2148 24884 -1948
<< ndiff >>
rect 1288 20647 1346 20659
rect 1288 20471 1300 20647
rect 1334 20471 1346 20647
rect 1288 20459 1346 20471
rect 1406 20647 1538 20659
rect 1406 20471 1418 20647
rect 1452 20471 1492 20647
rect 1406 20459 1492 20471
rect 1480 20271 1492 20459
rect 1526 20271 1538 20647
rect 1480 20259 1538 20271
rect 1598 20647 1656 20659
rect 1598 20271 1610 20647
rect 1644 20271 1656 20647
rect 1598 20259 1656 20271
rect 1716 20647 1774 20659
rect 1716 20271 1728 20647
rect 1762 20271 1774 20647
rect 1716 20259 1774 20271
rect 1834 20647 1892 20659
rect 1834 20271 1846 20647
rect 1880 20271 1892 20647
rect 1834 20259 1892 20271
rect 1952 20647 2088 20659
rect 1952 20271 1964 20647
rect 1998 20471 2042 20647
rect 2076 20471 2088 20647
rect 1998 20459 2088 20471
rect 2148 20647 2206 20659
rect 2148 20471 2160 20647
rect 2194 20471 2206 20647
rect 2148 20459 2206 20471
rect 4432 20647 4490 20659
rect 4432 20471 4444 20647
rect 4478 20471 4490 20647
rect 4432 20459 4490 20471
rect 4550 20647 4682 20659
rect 4550 20471 4562 20647
rect 4596 20471 4636 20647
rect 4550 20459 4636 20471
rect 1998 20271 2010 20459
rect 1952 20259 2010 20271
rect 4624 20271 4636 20459
rect 4670 20271 4682 20647
rect 4624 20259 4682 20271
rect 4742 20647 4800 20659
rect 4742 20271 4754 20647
rect 4788 20271 4800 20647
rect 4742 20259 4800 20271
rect 4860 20647 4918 20659
rect 4860 20271 4872 20647
rect 4906 20271 4918 20647
rect 4860 20259 4918 20271
rect 4978 20647 5036 20659
rect 4978 20271 4990 20647
rect 5024 20271 5036 20647
rect 4978 20259 5036 20271
rect 5096 20647 5232 20659
rect 5096 20271 5108 20647
rect 5142 20471 5186 20647
rect 5220 20471 5232 20647
rect 5142 20459 5232 20471
rect 5292 20647 5350 20659
rect 5292 20471 5304 20647
rect 5338 20471 5350 20647
rect 5292 20459 5350 20471
rect 7564 20651 7622 20663
rect 7564 20475 7576 20651
rect 7610 20475 7622 20651
rect 7564 20463 7622 20475
rect 7682 20651 7814 20663
rect 7682 20475 7694 20651
rect 7728 20475 7768 20651
rect 7682 20463 7768 20475
rect 5142 20271 5154 20459
rect 5096 20259 5154 20271
rect 7756 20275 7768 20463
rect 7802 20275 7814 20651
rect 7756 20263 7814 20275
rect 7874 20651 7932 20663
rect 7874 20275 7886 20651
rect 7920 20275 7932 20651
rect 7874 20263 7932 20275
rect 7992 20651 8050 20663
rect 7992 20275 8004 20651
rect 8038 20275 8050 20651
rect 7992 20263 8050 20275
rect 8110 20651 8168 20663
rect 8110 20275 8122 20651
rect 8156 20275 8168 20651
rect 8110 20263 8168 20275
rect 8228 20651 8364 20663
rect 8228 20275 8240 20651
rect 8274 20475 8318 20651
rect 8352 20475 8364 20651
rect 8274 20463 8364 20475
rect 8424 20651 8482 20663
rect 8424 20475 8436 20651
rect 8470 20475 8482 20651
rect 8424 20463 8482 20475
rect 10708 20651 10766 20663
rect 10708 20475 10720 20651
rect 10754 20475 10766 20651
rect 10708 20463 10766 20475
rect 10826 20651 10958 20663
rect 10826 20475 10838 20651
rect 10872 20475 10912 20651
rect 10826 20463 10912 20475
rect 8274 20275 8286 20463
rect 8228 20263 8286 20275
rect 10900 20275 10912 20463
rect 10946 20275 10958 20651
rect 10900 20263 10958 20275
rect 11018 20651 11076 20663
rect 11018 20275 11030 20651
rect 11064 20275 11076 20651
rect 11018 20263 11076 20275
rect 11136 20651 11194 20663
rect 11136 20275 11148 20651
rect 11182 20275 11194 20651
rect 11136 20263 11194 20275
rect 11254 20651 11312 20663
rect 11254 20275 11266 20651
rect 11300 20275 11312 20651
rect 11254 20263 11312 20275
rect 11372 20651 11508 20663
rect 11372 20275 11384 20651
rect 11418 20475 11462 20651
rect 11496 20475 11508 20651
rect 11418 20463 11508 20475
rect 11568 20651 11626 20663
rect 11568 20475 11580 20651
rect 11614 20475 11626 20651
rect 11568 20463 11626 20475
rect 13910 20647 13968 20659
rect 13910 20471 13922 20647
rect 13956 20471 13968 20647
rect 11418 20275 11430 20463
rect 11372 20263 11430 20275
rect 13910 20459 13968 20471
rect 14028 20647 14160 20659
rect 14028 20471 14040 20647
rect 14074 20471 14114 20647
rect 14028 20459 14114 20471
rect 14102 20271 14114 20459
rect 14148 20271 14160 20647
rect 14102 20259 14160 20271
rect 14220 20647 14278 20659
rect 14220 20271 14232 20647
rect 14266 20271 14278 20647
rect 14220 20259 14278 20271
rect 14338 20647 14396 20659
rect 14338 20271 14350 20647
rect 14384 20271 14396 20647
rect 14338 20259 14396 20271
rect 14456 20647 14514 20659
rect 14456 20271 14468 20647
rect 14502 20271 14514 20647
rect 14456 20259 14514 20271
rect 14574 20647 14710 20659
rect 14574 20271 14586 20647
rect 14620 20471 14664 20647
rect 14698 20471 14710 20647
rect 14620 20459 14710 20471
rect 14770 20647 14828 20659
rect 14770 20471 14782 20647
rect 14816 20471 14828 20647
rect 14770 20459 14828 20471
rect 17054 20647 17112 20659
rect 17054 20471 17066 20647
rect 17100 20471 17112 20647
rect 17054 20459 17112 20471
rect 17172 20647 17304 20659
rect 17172 20471 17184 20647
rect 17218 20471 17258 20647
rect 17172 20459 17258 20471
rect 14620 20271 14632 20459
rect 14574 20259 14632 20271
rect 17246 20271 17258 20459
rect 17292 20271 17304 20647
rect 17246 20259 17304 20271
rect 17364 20647 17422 20659
rect 17364 20271 17376 20647
rect 17410 20271 17422 20647
rect 17364 20259 17422 20271
rect 17482 20647 17540 20659
rect 17482 20271 17494 20647
rect 17528 20271 17540 20647
rect 17482 20259 17540 20271
rect 17600 20647 17658 20659
rect 17600 20271 17612 20647
rect 17646 20271 17658 20647
rect 17600 20259 17658 20271
rect 17718 20647 17854 20659
rect 17718 20271 17730 20647
rect 17764 20471 17808 20647
rect 17842 20471 17854 20647
rect 17764 20459 17854 20471
rect 17914 20647 17972 20659
rect 17914 20471 17926 20647
rect 17960 20471 17972 20647
rect 17914 20459 17972 20471
rect 20186 20651 20244 20663
rect 20186 20475 20198 20651
rect 20232 20475 20244 20651
rect 20186 20463 20244 20475
rect 20304 20651 20436 20663
rect 20304 20475 20316 20651
rect 20350 20475 20390 20651
rect 20304 20463 20390 20475
rect 17764 20271 17776 20459
rect 17718 20259 17776 20271
rect 20378 20275 20390 20463
rect 20424 20275 20436 20651
rect 20378 20263 20436 20275
rect 20496 20651 20554 20663
rect 20496 20275 20508 20651
rect 20542 20275 20554 20651
rect 20496 20263 20554 20275
rect 20614 20651 20672 20663
rect 20614 20275 20626 20651
rect 20660 20275 20672 20651
rect 20614 20263 20672 20275
rect 20732 20651 20790 20663
rect 20732 20275 20744 20651
rect 20778 20275 20790 20651
rect 20732 20263 20790 20275
rect 20850 20651 20986 20663
rect 20850 20275 20862 20651
rect 20896 20475 20940 20651
rect 20974 20475 20986 20651
rect 20896 20463 20986 20475
rect 21046 20651 21104 20663
rect 21046 20475 21058 20651
rect 21092 20475 21104 20651
rect 21046 20463 21104 20475
rect 23330 20651 23388 20663
rect 23330 20475 23342 20651
rect 23376 20475 23388 20651
rect 23330 20463 23388 20475
rect 23448 20651 23580 20663
rect 23448 20475 23460 20651
rect 23494 20475 23534 20651
rect 23448 20463 23534 20475
rect 20896 20275 20908 20463
rect 20850 20263 20908 20275
rect 23522 20275 23534 20463
rect 23568 20275 23580 20651
rect 23522 20263 23580 20275
rect 23640 20651 23698 20663
rect 23640 20275 23652 20651
rect 23686 20275 23698 20651
rect 23640 20263 23698 20275
rect 23758 20651 23816 20663
rect 23758 20275 23770 20651
rect 23804 20275 23816 20651
rect 23758 20263 23816 20275
rect 23876 20651 23934 20663
rect 23876 20275 23888 20651
rect 23922 20275 23934 20651
rect 23876 20263 23934 20275
rect 23994 20651 24130 20663
rect 23994 20275 24006 20651
rect 24040 20475 24084 20651
rect 24118 20475 24130 20651
rect 24040 20463 24130 20475
rect 24190 20651 24248 20663
rect 24190 20475 24202 20651
rect 24236 20475 24248 20651
rect 24190 20463 24248 20475
rect 24040 20275 24052 20463
rect 23994 20263 24052 20275
rect 3134 16162 3192 16174
rect 3134 15786 3146 16162
rect 3180 15786 3192 16162
rect 3134 15774 3192 15786
rect 3252 16162 3310 16174
rect 3252 15786 3264 16162
rect 3298 15786 3310 16162
rect 3252 15774 3310 15786
rect 3370 16162 3428 16174
rect 3370 15786 3382 16162
rect 3416 15786 3428 16162
rect 3487 16162 3545 16174
rect 3487 15986 3499 16162
rect 3533 15986 3545 16162
rect 3487 15974 3545 15986
rect 3605 16162 3663 16174
rect 3605 15986 3617 16162
rect 3651 15986 3663 16162
rect 3605 15974 3663 15986
rect 4582 16162 4640 16174
rect 3370 15774 3428 15786
rect 4582 15786 4594 16162
rect 4628 15786 4640 16162
rect 4582 15774 4640 15786
rect 4700 16162 4758 16174
rect 4700 15786 4712 16162
rect 4746 15786 4758 16162
rect 4700 15774 4758 15786
rect 4818 16162 4876 16174
rect 4818 15786 4830 16162
rect 4864 15786 4876 16162
rect 4935 16162 4993 16174
rect 4935 15986 4947 16162
rect 4981 15986 4993 16162
rect 4935 15974 4993 15986
rect 5053 16162 5111 16174
rect 5053 15986 5065 16162
rect 5099 15986 5111 16162
rect 5053 15974 5111 15986
rect 6080 16164 6138 16176
rect 4818 15774 4876 15786
rect 6080 15788 6092 16164
rect 6126 15788 6138 16164
rect 6080 15776 6138 15788
rect 6198 16164 6256 16176
rect 6198 15788 6210 16164
rect 6244 15788 6256 16164
rect 6198 15776 6256 15788
rect 6316 16164 6374 16176
rect 6316 15788 6328 16164
rect 6362 15788 6374 16164
rect 6433 16164 6491 16176
rect 6433 15988 6445 16164
rect 6479 15988 6491 16164
rect 6433 15976 6491 15988
rect 6551 16164 6609 16176
rect 6551 15988 6563 16164
rect 6597 15988 6609 16164
rect 6551 15976 6609 15988
rect 7528 16164 7586 16176
rect 6316 15776 6374 15788
rect 7528 15788 7540 16164
rect 7574 15788 7586 16164
rect 7528 15776 7586 15788
rect 7646 16164 7704 16176
rect 7646 15788 7658 16164
rect 7692 15788 7704 16164
rect 7646 15776 7704 15788
rect 7764 16164 7822 16176
rect 7764 15788 7776 16164
rect 7810 15788 7822 16164
rect 7881 16164 7939 16176
rect 7881 15988 7893 16164
rect 7927 15988 7939 16164
rect 7881 15976 7939 15988
rect 7999 16164 8057 16176
rect 7999 15988 8011 16164
rect 8045 15988 8057 16164
rect 7999 15976 8057 15988
rect 9048 16162 9106 16174
rect 7764 15776 7822 15788
rect 9048 15786 9060 16162
rect 9094 15786 9106 16162
rect 9048 15774 9106 15786
rect 9166 16162 9224 16174
rect 9166 15786 9178 16162
rect 9212 15786 9224 16162
rect 9166 15774 9224 15786
rect 9284 16162 9342 16174
rect 9284 15786 9296 16162
rect 9330 15786 9342 16162
rect 9401 16162 9459 16174
rect 9401 15986 9413 16162
rect 9447 15986 9459 16162
rect 9401 15974 9459 15986
rect 9519 16162 9577 16174
rect 9519 15986 9531 16162
rect 9565 15986 9577 16162
rect 9519 15974 9577 15986
rect 10496 16162 10554 16174
rect 9284 15774 9342 15786
rect 10496 15786 10508 16162
rect 10542 15786 10554 16162
rect 10496 15774 10554 15786
rect 10614 16162 10672 16174
rect 10614 15786 10626 16162
rect 10660 15786 10672 16162
rect 10614 15774 10672 15786
rect 10732 16162 10790 16174
rect 10732 15786 10744 16162
rect 10778 15786 10790 16162
rect 10849 16162 10907 16174
rect 10849 15986 10861 16162
rect 10895 15986 10907 16162
rect 10849 15974 10907 15986
rect 10967 16162 11025 16174
rect 10967 15986 10979 16162
rect 11013 15986 11025 16162
rect 10967 15974 11025 15986
rect 11994 16164 12052 16176
rect 10732 15774 10790 15786
rect 11994 15788 12006 16164
rect 12040 15788 12052 16164
rect 11994 15776 12052 15788
rect 12112 16164 12170 16176
rect 12112 15788 12124 16164
rect 12158 15788 12170 16164
rect 12112 15776 12170 15788
rect 12230 16164 12288 16176
rect 12230 15788 12242 16164
rect 12276 15788 12288 16164
rect 12347 16164 12405 16176
rect 12347 15988 12359 16164
rect 12393 15988 12405 16164
rect 12347 15976 12405 15988
rect 12465 16164 12523 16176
rect 12465 15988 12477 16164
rect 12511 15988 12523 16164
rect 12465 15976 12523 15988
rect 13442 16164 13500 16176
rect 12230 15776 12288 15788
rect 13442 15788 13454 16164
rect 13488 15788 13500 16164
rect 13442 15776 13500 15788
rect 13560 16164 13618 16176
rect 13560 15788 13572 16164
rect 13606 15788 13618 16164
rect 13560 15776 13618 15788
rect 13678 16164 13736 16176
rect 13678 15788 13690 16164
rect 13724 15788 13736 16164
rect 13795 16164 13853 16176
rect 13795 15988 13807 16164
rect 13841 15988 13853 16164
rect 13795 15976 13853 15988
rect 13913 16164 13971 16176
rect 13913 15988 13925 16164
rect 13959 15988 13971 16164
rect 13913 15976 13971 15988
rect 14570 16010 14628 16022
rect 14570 15834 14582 16010
rect 14616 15834 14628 16010
rect 14570 15822 14628 15834
rect 14688 16010 14746 16022
rect 14688 15834 14700 16010
rect 14734 15834 14746 16010
rect 14688 15822 14746 15834
rect 14806 16010 14864 16022
rect 14806 15834 14818 16010
rect 14852 15834 14864 16010
rect 14806 15822 14864 15834
rect 14924 16010 14982 16022
rect 14924 15834 14936 16010
rect 14970 15834 14982 16010
rect 14924 15822 14982 15834
rect 13678 15776 13736 15788
rect 15738 16012 15796 16024
rect 15738 15836 15750 16012
rect 15784 15836 15796 16012
rect 15738 15824 15796 15836
rect 15856 16012 15914 16024
rect 15856 15836 15868 16012
rect 15902 15836 15914 16012
rect 15856 15824 15914 15836
rect 15974 16012 16032 16024
rect 15974 15836 15986 16012
rect 16020 15836 16032 16012
rect 15974 15824 16032 15836
rect 16092 16012 16150 16024
rect 16092 15836 16104 16012
rect 16138 15836 16150 16012
rect 16092 15824 16150 15836
rect 16906 16012 16964 16024
rect 16906 15836 16918 16012
rect 16952 15836 16964 16012
rect 16906 15824 16964 15836
rect 17024 16012 17082 16024
rect 17024 15836 17036 16012
rect 17070 15836 17082 16012
rect 17024 15824 17082 15836
rect 17142 16012 17200 16024
rect 17142 15836 17154 16012
rect 17188 15836 17200 16012
rect 17142 15824 17200 15836
rect 17260 16012 17318 16024
rect 17260 15836 17272 16012
rect 17306 15836 17318 16012
rect 17260 15824 17318 15836
rect 18074 16012 18132 16024
rect 18074 15836 18086 16012
rect 18120 15836 18132 16012
rect 18074 15824 18132 15836
rect 18192 16012 18250 16024
rect 18192 15836 18204 16012
rect 18238 15836 18250 16012
rect 18192 15824 18250 15836
rect 18310 16012 18368 16024
rect 18310 15836 18322 16012
rect 18356 15836 18368 16012
rect 18310 15824 18368 15836
rect 18428 16012 18486 16024
rect 18428 15836 18440 16012
rect 18474 15836 18486 16012
rect 18428 15824 18486 15836
rect 19248 16012 19306 16024
rect 19248 15836 19260 16012
rect 19294 15836 19306 16012
rect 19248 15824 19306 15836
rect 19366 16012 19424 16024
rect 19366 15836 19378 16012
rect 19412 15836 19424 16012
rect 19366 15824 19424 15836
rect 19484 16012 19542 16024
rect 19484 15836 19496 16012
rect 19530 15836 19542 16012
rect 19484 15824 19542 15836
rect 19602 16012 19660 16024
rect 19602 15836 19614 16012
rect 19648 15836 19660 16012
rect 19602 15824 19660 15836
rect 20416 16012 20474 16024
rect 20416 15836 20428 16012
rect 20462 15836 20474 16012
rect 20416 15824 20474 15836
rect 20534 16012 20592 16024
rect 20534 15836 20546 16012
rect 20580 15836 20592 16012
rect 20534 15824 20592 15836
rect 20652 16012 20710 16024
rect 20652 15836 20664 16012
rect 20698 15836 20710 16012
rect 20652 15824 20710 15836
rect 20770 16012 20828 16024
rect 20770 15836 20782 16012
rect 20816 15836 20828 16012
rect 20770 15824 20828 15836
rect 21584 16014 21642 16026
rect 21584 15838 21596 16014
rect 21630 15838 21642 16014
rect 21584 15826 21642 15838
rect 21702 16014 21760 16026
rect 21702 15838 21714 16014
rect 21748 15838 21760 16014
rect 21702 15826 21760 15838
rect 21820 16014 21878 16026
rect 21820 15838 21832 16014
rect 21866 15838 21878 16014
rect 21820 15826 21878 15838
rect 21938 16014 21996 16026
rect 21938 15838 21950 16014
rect 21984 15838 21996 16014
rect 21938 15826 21996 15838
rect 22752 16014 22810 16026
rect 22752 15838 22764 16014
rect 22798 15838 22810 16014
rect 22752 15826 22810 15838
rect 22870 16014 22928 16026
rect 22870 15838 22882 16014
rect 22916 15838 22928 16014
rect 22870 15826 22928 15838
rect 22988 16014 23046 16026
rect 22988 15838 23000 16014
rect 23034 15838 23046 16014
rect 22988 15826 23046 15838
rect 23106 16014 23164 16026
rect 23106 15838 23118 16014
rect 23152 15838 23164 16014
rect 23106 15826 23164 15838
rect 3790 13509 3848 13521
rect 3790 13333 3802 13509
rect 3836 13333 3848 13509
rect 3790 13321 3848 13333
rect 3908 13509 4040 13521
rect 3908 13333 3920 13509
rect 3954 13333 3994 13509
rect 3908 13321 3994 13333
rect 3982 13133 3994 13321
rect 4028 13133 4040 13509
rect 3982 13121 4040 13133
rect 4100 13509 4158 13521
rect 4100 13133 4112 13509
rect 4146 13133 4158 13509
rect 4100 13121 4158 13133
rect 4218 13509 4276 13521
rect 4218 13133 4230 13509
rect 4264 13133 4276 13509
rect 4218 13121 4276 13133
rect 4336 13509 4394 13521
rect 4336 13133 4348 13509
rect 4382 13133 4394 13509
rect 4336 13121 4394 13133
rect 4454 13509 4590 13521
rect 4454 13133 4466 13509
rect 4500 13333 4544 13509
rect 4578 13333 4590 13509
rect 4500 13321 4590 13333
rect 4650 13509 4708 13521
rect 4650 13333 4662 13509
rect 4696 13333 4708 13509
rect 4650 13321 4708 13333
rect 6934 13509 6992 13521
rect 6934 13333 6946 13509
rect 6980 13333 6992 13509
rect 6934 13321 6992 13333
rect 7052 13509 7184 13521
rect 7052 13333 7064 13509
rect 7098 13333 7138 13509
rect 7052 13321 7138 13333
rect 4500 13133 4512 13321
rect 4454 13121 4512 13133
rect 7126 13133 7138 13321
rect 7172 13133 7184 13509
rect 7126 13121 7184 13133
rect 7244 13509 7302 13521
rect 7244 13133 7256 13509
rect 7290 13133 7302 13509
rect 7244 13121 7302 13133
rect 7362 13509 7420 13521
rect 7362 13133 7374 13509
rect 7408 13133 7420 13509
rect 7362 13121 7420 13133
rect 7480 13509 7538 13521
rect 7480 13133 7492 13509
rect 7526 13133 7538 13509
rect 7480 13121 7538 13133
rect 7598 13509 7734 13521
rect 7598 13133 7610 13509
rect 7644 13333 7688 13509
rect 7722 13333 7734 13509
rect 7644 13321 7734 13333
rect 7794 13509 7852 13521
rect 7794 13333 7806 13509
rect 7840 13333 7852 13509
rect 7794 13321 7852 13333
rect 10066 13513 10124 13525
rect 10066 13337 10078 13513
rect 10112 13337 10124 13513
rect 10066 13325 10124 13337
rect 10184 13513 10316 13525
rect 10184 13337 10196 13513
rect 10230 13337 10270 13513
rect 10184 13325 10270 13337
rect 7644 13133 7656 13321
rect 7598 13121 7656 13133
rect 10258 13137 10270 13325
rect 10304 13137 10316 13513
rect 10258 13125 10316 13137
rect 10376 13513 10434 13525
rect 10376 13137 10388 13513
rect 10422 13137 10434 13513
rect 10376 13125 10434 13137
rect 10494 13513 10552 13525
rect 10494 13137 10506 13513
rect 10540 13137 10552 13513
rect 10494 13125 10552 13137
rect 10612 13513 10670 13525
rect 10612 13137 10624 13513
rect 10658 13137 10670 13513
rect 10612 13125 10670 13137
rect 10730 13513 10866 13525
rect 10730 13137 10742 13513
rect 10776 13337 10820 13513
rect 10854 13337 10866 13513
rect 10776 13325 10866 13337
rect 10926 13513 10984 13525
rect 10926 13337 10938 13513
rect 10972 13337 10984 13513
rect 10926 13325 10984 13337
rect 13210 13513 13268 13525
rect 13210 13337 13222 13513
rect 13256 13337 13268 13513
rect 13210 13325 13268 13337
rect 13328 13513 13460 13525
rect 13328 13337 13340 13513
rect 13374 13337 13414 13513
rect 13328 13325 13414 13337
rect 10776 13137 10788 13325
rect 10730 13125 10788 13137
rect 13402 13137 13414 13325
rect 13448 13137 13460 13513
rect 13402 13125 13460 13137
rect 13520 13513 13578 13525
rect 13520 13137 13532 13513
rect 13566 13137 13578 13513
rect 13520 13125 13578 13137
rect 13638 13513 13696 13525
rect 13638 13137 13650 13513
rect 13684 13137 13696 13513
rect 13638 13125 13696 13137
rect 13756 13513 13814 13525
rect 13756 13137 13768 13513
rect 13802 13137 13814 13513
rect 13756 13125 13814 13137
rect 13874 13513 14010 13525
rect 13874 13137 13886 13513
rect 13920 13337 13964 13513
rect 13998 13337 14010 13513
rect 13920 13325 14010 13337
rect 14070 13513 14128 13525
rect 14070 13337 14082 13513
rect 14116 13337 14128 13513
rect 14070 13325 14128 13337
rect 16412 13509 16470 13521
rect 16412 13333 16424 13509
rect 16458 13333 16470 13509
rect 13920 13137 13932 13325
rect 13874 13125 13932 13137
rect 16412 13321 16470 13333
rect 16530 13509 16662 13521
rect 16530 13333 16542 13509
rect 16576 13333 16616 13509
rect 16530 13321 16616 13333
rect 16604 13133 16616 13321
rect 16650 13133 16662 13509
rect 16604 13121 16662 13133
rect 16722 13509 16780 13521
rect 16722 13133 16734 13509
rect 16768 13133 16780 13509
rect 16722 13121 16780 13133
rect 16840 13509 16898 13521
rect 16840 13133 16852 13509
rect 16886 13133 16898 13509
rect 16840 13121 16898 13133
rect 16958 13509 17016 13521
rect 16958 13133 16970 13509
rect 17004 13133 17016 13509
rect 16958 13121 17016 13133
rect 17076 13509 17212 13521
rect 17076 13133 17088 13509
rect 17122 13333 17166 13509
rect 17200 13333 17212 13509
rect 17122 13321 17212 13333
rect 17272 13509 17330 13521
rect 17272 13333 17284 13509
rect 17318 13333 17330 13509
rect 17272 13321 17330 13333
rect 19556 13509 19614 13521
rect 19556 13333 19568 13509
rect 19602 13333 19614 13509
rect 19556 13321 19614 13333
rect 19674 13509 19806 13521
rect 19674 13333 19686 13509
rect 19720 13333 19760 13509
rect 19674 13321 19760 13333
rect 17122 13133 17134 13321
rect 17076 13121 17134 13133
rect 19748 13133 19760 13321
rect 19794 13133 19806 13509
rect 19748 13121 19806 13133
rect 19866 13509 19924 13521
rect 19866 13133 19878 13509
rect 19912 13133 19924 13509
rect 19866 13121 19924 13133
rect 19984 13509 20042 13521
rect 19984 13133 19996 13509
rect 20030 13133 20042 13509
rect 19984 13121 20042 13133
rect 20102 13509 20160 13521
rect 20102 13133 20114 13509
rect 20148 13133 20160 13509
rect 20102 13121 20160 13133
rect 20220 13509 20356 13521
rect 20220 13133 20232 13509
rect 20266 13333 20310 13509
rect 20344 13333 20356 13509
rect 20266 13321 20356 13333
rect 20416 13509 20474 13521
rect 20416 13333 20428 13509
rect 20462 13333 20474 13509
rect 20416 13321 20474 13333
rect 22688 13513 22746 13525
rect 22688 13337 22700 13513
rect 22734 13337 22746 13513
rect 22688 13325 22746 13337
rect 22806 13513 22938 13525
rect 22806 13337 22818 13513
rect 22852 13337 22892 13513
rect 22806 13325 22892 13337
rect 20266 13133 20278 13321
rect 20220 13121 20278 13133
rect 22880 13137 22892 13325
rect 22926 13137 22938 13513
rect 22880 13125 22938 13137
rect 22998 13513 23056 13525
rect 22998 13137 23010 13513
rect 23044 13137 23056 13513
rect 22998 13125 23056 13137
rect 23116 13513 23174 13525
rect 23116 13137 23128 13513
rect 23162 13137 23174 13513
rect 23116 13125 23174 13137
rect 23234 13513 23292 13525
rect 23234 13137 23246 13513
rect 23280 13137 23292 13513
rect 23234 13125 23292 13137
rect 23352 13513 23488 13525
rect 23352 13137 23364 13513
rect 23398 13337 23442 13513
rect 23476 13337 23488 13513
rect 23398 13325 23488 13337
rect 23548 13513 23606 13525
rect 23548 13337 23560 13513
rect 23594 13337 23606 13513
rect 23548 13325 23606 13337
rect 25832 13513 25890 13525
rect 25832 13337 25844 13513
rect 25878 13337 25890 13513
rect 25832 13325 25890 13337
rect 25950 13513 26082 13525
rect 25950 13337 25962 13513
rect 25996 13337 26036 13513
rect 25950 13325 26036 13337
rect 23398 13137 23410 13325
rect 23352 13125 23410 13137
rect 26024 13137 26036 13325
rect 26070 13137 26082 13513
rect 26024 13125 26082 13137
rect 26142 13513 26200 13525
rect 26142 13137 26154 13513
rect 26188 13137 26200 13513
rect 26142 13125 26200 13137
rect 26260 13513 26318 13525
rect 26260 13137 26272 13513
rect 26306 13137 26318 13513
rect 26260 13125 26318 13137
rect 26378 13513 26436 13525
rect 26378 13137 26390 13513
rect 26424 13137 26436 13513
rect 26378 13125 26436 13137
rect 26496 13513 26632 13525
rect 26496 13137 26508 13513
rect 26542 13337 26586 13513
rect 26620 13337 26632 13513
rect 26542 13325 26632 13337
rect 26692 13513 26750 13525
rect 26692 13337 26704 13513
rect 26738 13337 26750 13513
rect 26692 13325 26750 13337
rect 26542 13137 26554 13325
rect 26496 13125 26554 13137
rect 3790 10775 3848 10787
rect 3790 10599 3802 10775
rect 3836 10599 3848 10775
rect 3790 10587 3848 10599
rect 3908 10775 4040 10787
rect 3908 10599 3920 10775
rect 3954 10599 3994 10775
rect 3908 10587 3994 10599
rect 3982 10399 3994 10587
rect 4028 10399 4040 10775
rect 3982 10387 4040 10399
rect 4100 10775 4158 10787
rect 4100 10399 4112 10775
rect 4146 10399 4158 10775
rect 4100 10387 4158 10399
rect 4218 10775 4276 10787
rect 4218 10399 4230 10775
rect 4264 10399 4276 10775
rect 4218 10387 4276 10399
rect 4336 10775 4394 10787
rect 4336 10399 4348 10775
rect 4382 10399 4394 10775
rect 4336 10387 4394 10399
rect 4454 10775 4590 10787
rect 4454 10399 4466 10775
rect 4500 10599 4544 10775
rect 4578 10599 4590 10775
rect 4500 10587 4590 10599
rect 4650 10775 4708 10787
rect 4650 10599 4662 10775
rect 4696 10599 4708 10775
rect 4650 10587 4708 10599
rect 6934 10775 6992 10787
rect 6934 10599 6946 10775
rect 6980 10599 6992 10775
rect 6934 10587 6992 10599
rect 7052 10775 7184 10787
rect 7052 10599 7064 10775
rect 7098 10599 7138 10775
rect 7052 10587 7138 10599
rect 4500 10399 4512 10587
rect 4454 10387 4512 10399
rect 7126 10399 7138 10587
rect 7172 10399 7184 10775
rect 7126 10387 7184 10399
rect 7244 10775 7302 10787
rect 7244 10399 7256 10775
rect 7290 10399 7302 10775
rect 7244 10387 7302 10399
rect 7362 10775 7420 10787
rect 7362 10399 7374 10775
rect 7408 10399 7420 10775
rect 7362 10387 7420 10399
rect 7480 10775 7538 10787
rect 7480 10399 7492 10775
rect 7526 10399 7538 10775
rect 7480 10387 7538 10399
rect 7598 10775 7734 10787
rect 7598 10399 7610 10775
rect 7644 10599 7688 10775
rect 7722 10599 7734 10775
rect 7644 10587 7734 10599
rect 7794 10775 7852 10787
rect 7794 10599 7806 10775
rect 7840 10599 7852 10775
rect 7794 10587 7852 10599
rect 10066 10779 10124 10791
rect 10066 10603 10078 10779
rect 10112 10603 10124 10779
rect 10066 10591 10124 10603
rect 10184 10779 10316 10791
rect 10184 10603 10196 10779
rect 10230 10603 10270 10779
rect 10184 10591 10270 10603
rect 7644 10399 7656 10587
rect 7598 10387 7656 10399
rect 10258 10403 10270 10591
rect 10304 10403 10316 10779
rect 10258 10391 10316 10403
rect 10376 10779 10434 10791
rect 10376 10403 10388 10779
rect 10422 10403 10434 10779
rect 10376 10391 10434 10403
rect 10494 10779 10552 10791
rect 10494 10403 10506 10779
rect 10540 10403 10552 10779
rect 10494 10391 10552 10403
rect 10612 10779 10670 10791
rect 10612 10403 10624 10779
rect 10658 10403 10670 10779
rect 10612 10391 10670 10403
rect 10730 10779 10866 10791
rect 10730 10403 10742 10779
rect 10776 10603 10820 10779
rect 10854 10603 10866 10779
rect 10776 10591 10866 10603
rect 10926 10779 10984 10791
rect 10926 10603 10938 10779
rect 10972 10603 10984 10779
rect 10926 10591 10984 10603
rect 13210 10779 13268 10791
rect 13210 10603 13222 10779
rect 13256 10603 13268 10779
rect 13210 10591 13268 10603
rect 13328 10779 13460 10791
rect 13328 10603 13340 10779
rect 13374 10603 13414 10779
rect 13328 10591 13414 10603
rect 10776 10403 10788 10591
rect 10730 10391 10788 10403
rect 13402 10403 13414 10591
rect 13448 10403 13460 10779
rect 13402 10391 13460 10403
rect 13520 10779 13578 10791
rect 13520 10403 13532 10779
rect 13566 10403 13578 10779
rect 13520 10391 13578 10403
rect 13638 10779 13696 10791
rect 13638 10403 13650 10779
rect 13684 10403 13696 10779
rect 13638 10391 13696 10403
rect 13756 10779 13814 10791
rect 13756 10403 13768 10779
rect 13802 10403 13814 10779
rect 13756 10391 13814 10403
rect 13874 10779 14010 10791
rect 13874 10403 13886 10779
rect 13920 10603 13964 10779
rect 13998 10603 14010 10779
rect 13920 10591 14010 10603
rect 14070 10779 14128 10791
rect 14070 10603 14082 10779
rect 14116 10603 14128 10779
rect 14070 10591 14128 10603
rect 16412 10775 16470 10787
rect 16412 10599 16424 10775
rect 16458 10599 16470 10775
rect 13920 10403 13932 10591
rect 13874 10391 13932 10403
rect 16412 10587 16470 10599
rect 16530 10775 16662 10787
rect 16530 10599 16542 10775
rect 16576 10599 16616 10775
rect 16530 10587 16616 10599
rect 16604 10399 16616 10587
rect 16650 10399 16662 10775
rect 16604 10387 16662 10399
rect 16722 10775 16780 10787
rect 16722 10399 16734 10775
rect 16768 10399 16780 10775
rect 16722 10387 16780 10399
rect 16840 10775 16898 10787
rect 16840 10399 16852 10775
rect 16886 10399 16898 10775
rect 16840 10387 16898 10399
rect 16958 10775 17016 10787
rect 16958 10399 16970 10775
rect 17004 10399 17016 10775
rect 16958 10387 17016 10399
rect 17076 10775 17212 10787
rect 17076 10399 17088 10775
rect 17122 10599 17166 10775
rect 17200 10599 17212 10775
rect 17122 10587 17212 10599
rect 17272 10775 17330 10787
rect 17272 10599 17284 10775
rect 17318 10599 17330 10775
rect 17272 10587 17330 10599
rect 19556 10775 19614 10787
rect 19556 10599 19568 10775
rect 19602 10599 19614 10775
rect 19556 10587 19614 10599
rect 19674 10775 19806 10787
rect 19674 10599 19686 10775
rect 19720 10599 19760 10775
rect 19674 10587 19760 10599
rect 17122 10399 17134 10587
rect 17076 10387 17134 10399
rect 19748 10399 19760 10587
rect 19794 10399 19806 10775
rect 19748 10387 19806 10399
rect 19866 10775 19924 10787
rect 19866 10399 19878 10775
rect 19912 10399 19924 10775
rect 19866 10387 19924 10399
rect 19984 10775 20042 10787
rect 19984 10399 19996 10775
rect 20030 10399 20042 10775
rect 19984 10387 20042 10399
rect 20102 10775 20160 10787
rect 20102 10399 20114 10775
rect 20148 10399 20160 10775
rect 20102 10387 20160 10399
rect 20220 10775 20356 10787
rect 20220 10399 20232 10775
rect 20266 10599 20310 10775
rect 20344 10599 20356 10775
rect 20266 10587 20356 10599
rect 20416 10775 20474 10787
rect 20416 10599 20428 10775
rect 20462 10599 20474 10775
rect 20416 10587 20474 10599
rect 22688 10779 22746 10791
rect 22688 10603 22700 10779
rect 22734 10603 22746 10779
rect 22688 10591 22746 10603
rect 22806 10779 22938 10791
rect 22806 10603 22818 10779
rect 22852 10603 22892 10779
rect 22806 10591 22892 10603
rect 20266 10399 20278 10587
rect 20220 10387 20278 10399
rect 22880 10403 22892 10591
rect 22926 10403 22938 10779
rect 22880 10391 22938 10403
rect 22998 10779 23056 10791
rect 22998 10403 23010 10779
rect 23044 10403 23056 10779
rect 22998 10391 23056 10403
rect 23116 10779 23174 10791
rect 23116 10403 23128 10779
rect 23162 10403 23174 10779
rect 23116 10391 23174 10403
rect 23234 10779 23292 10791
rect 23234 10403 23246 10779
rect 23280 10403 23292 10779
rect 23234 10391 23292 10403
rect 23352 10779 23488 10791
rect 23352 10403 23364 10779
rect 23398 10603 23442 10779
rect 23476 10603 23488 10779
rect 23398 10591 23488 10603
rect 23548 10779 23606 10791
rect 23548 10603 23560 10779
rect 23594 10603 23606 10779
rect 23548 10591 23606 10603
rect 25832 10779 25890 10791
rect 25832 10603 25844 10779
rect 25878 10603 25890 10779
rect 25832 10591 25890 10603
rect 25950 10779 26082 10791
rect 25950 10603 25962 10779
rect 25996 10603 26036 10779
rect 25950 10591 26036 10603
rect 23398 10403 23410 10591
rect 23352 10391 23410 10403
rect 26024 10403 26036 10591
rect 26070 10403 26082 10779
rect 26024 10391 26082 10403
rect 26142 10779 26200 10791
rect 26142 10403 26154 10779
rect 26188 10403 26200 10779
rect 26142 10391 26200 10403
rect 26260 10779 26318 10791
rect 26260 10403 26272 10779
rect 26306 10403 26318 10779
rect 26260 10391 26318 10403
rect 26378 10779 26436 10791
rect 26378 10403 26390 10779
rect 26424 10403 26436 10779
rect 26378 10391 26436 10403
rect 26496 10779 26632 10791
rect 26496 10403 26508 10779
rect 26542 10603 26586 10779
rect 26620 10603 26632 10779
rect 26542 10591 26632 10603
rect 26692 10779 26750 10791
rect 26692 10603 26704 10779
rect 26738 10603 26750 10779
rect 26692 10591 26750 10603
rect 26542 10403 26554 10591
rect 26496 10391 26554 10403
rect 3780 8043 3838 8055
rect 3780 7867 3792 8043
rect 3826 7867 3838 8043
rect 3780 7855 3838 7867
rect 3898 8043 4030 8055
rect 3898 7867 3910 8043
rect 3944 7867 3984 8043
rect 3898 7855 3984 7867
rect 3972 7667 3984 7855
rect 4018 7667 4030 8043
rect 3972 7655 4030 7667
rect 4090 8043 4148 8055
rect 4090 7667 4102 8043
rect 4136 7667 4148 8043
rect 4090 7655 4148 7667
rect 4208 8043 4266 8055
rect 4208 7667 4220 8043
rect 4254 7667 4266 8043
rect 4208 7655 4266 7667
rect 4326 8043 4384 8055
rect 4326 7667 4338 8043
rect 4372 7667 4384 8043
rect 4326 7655 4384 7667
rect 4444 8043 4580 8055
rect 4444 7667 4456 8043
rect 4490 7867 4534 8043
rect 4568 7867 4580 8043
rect 4490 7855 4580 7867
rect 4640 8043 4698 8055
rect 4640 7867 4652 8043
rect 4686 7867 4698 8043
rect 4640 7855 4698 7867
rect 6924 8043 6982 8055
rect 6924 7867 6936 8043
rect 6970 7867 6982 8043
rect 6924 7855 6982 7867
rect 7042 8043 7174 8055
rect 7042 7867 7054 8043
rect 7088 7867 7128 8043
rect 7042 7855 7128 7867
rect 4490 7667 4502 7855
rect 4444 7655 4502 7667
rect 7116 7667 7128 7855
rect 7162 7667 7174 8043
rect 7116 7655 7174 7667
rect 7234 8043 7292 8055
rect 7234 7667 7246 8043
rect 7280 7667 7292 8043
rect 7234 7655 7292 7667
rect 7352 8043 7410 8055
rect 7352 7667 7364 8043
rect 7398 7667 7410 8043
rect 7352 7655 7410 7667
rect 7470 8043 7528 8055
rect 7470 7667 7482 8043
rect 7516 7667 7528 8043
rect 7470 7655 7528 7667
rect 7588 8043 7724 8055
rect 7588 7667 7600 8043
rect 7634 7867 7678 8043
rect 7712 7867 7724 8043
rect 7634 7855 7724 7867
rect 7784 8043 7842 8055
rect 7784 7867 7796 8043
rect 7830 7867 7842 8043
rect 7784 7855 7842 7867
rect 10056 8047 10114 8059
rect 10056 7871 10068 8047
rect 10102 7871 10114 8047
rect 10056 7859 10114 7871
rect 10174 8047 10306 8059
rect 10174 7871 10186 8047
rect 10220 7871 10260 8047
rect 10174 7859 10260 7871
rect 7634 7667 7646 7855
rect 7588 7655 7646 7667
rect 10248 7671 10260 7859
rect 10294 7671 10306 8047
rect 10248 7659 10306 7671
rect 10366 8047 10424 8059
rect 10366 7671 10378 8047
rect 10412 7671 10424 8047
rect 10366 7659 10424 7671
rect 10484 8047 10542 8059
rect 10484 7671 10496 8047
rect 10530 7671 10542 8047
rect 10484 7659 10542 7671
rect 10602 8047 10660 8059
rect 10602 7671 10614 8047
rect 10648 7671 10660 8047
rect 10602 7659 10660 7671
rect 10720 8047 10856 8059
rect 10720 7671 10732 8047
rect 10766 7871 10810 8047
rect 10844 7871 10856 8047
rect 10766 7859 10856 7871
rect 10916 8047 10974 8059
rect 10916 7871 10928 8047
rect 10962 7871 10974 8047
rect 10916 7859 10974 7871
rect 13200 8047 13258 8059
rect 13200 7871 13212 8047
rect 13246 7871 13258 8047
rect 13200 7859 13258 7871
rect 13318 8047 13450 8059
rect 13318 7871 13330 8047
rect 13364 7871 13404 8047
rect 13318 7859 13404 7871
rect 10766 7671 10778 7859
rect 10720 7659 10778 7671
rect 13392 7671 13404 7859
rect 13438 7671 13450 8047
rect 13392 7659 13450 7671
rect 13510 8047 13568 8059
rect 13510 7671 13522 8047
rect 13556 7671 13568 8047
rect 13510 7659 13568 7671
rect 13628 8047 13686 8059
rect 13628 7671 13640 8047
rect 13674 7671 13686 8047
rect 13628 7659 13686 7671
rect 13746 8047 13804 8059
rect 13746 7671 13758 8047
rect 13792 7671 13804 8047
rect 13746 7659 13804 7671
rect 13864 8047 14000 8059
rect 13864 7671 13876 8047
rect 13910 7871 13954 8047
rect 13988 7871 14000 8047
rect 13910 7859 14000 7871
rect 14060 8047 14118 8059
rect 14060 7871 14072 8047
rect 14106 7871 14118 8047
rect 14060 7859 14118 7871
rect 16402 8043 16460 8055
rect 16402 7867 16414 8043
rect 16448 7867 16460 8043
rect 13910 7671 13922 7859
rect 13864 7659 13922 7671
rect 16402 7855 16460 7867
rect 16520 8043 16652 8055
rect 16520 7867 16532 8043
rect 16566 7867 16606 8043
rect 16520 7855 16606 7867
rect 16594 7667 16606 7855
rect 16640 7667 16652 8043
rect 16594 7655 16652 7667
rect 16712 8043 16770 8055
rect 16712 7667 16724 8043
rect 16758 7667 16770 8043
rect 16712 7655 16770 7667
rect 16830 8043 16888 8055
rect 16830 7667 16842 8043
rect 16876 7667 16888 8043
rect 16830 7655 16888 7667
rect 16948 8043 17006 8055
rect 16948 7667 16960 8043
rect 16994 7667 17006 8043
rect 16948 7655 17006 7667
rect 17066 8043 17202 8055
rect 17066 7667 17078 8043
rect 17112 7867 17156 8043
rect 17190 7867 17202 8043
rect 17112 7855 17202 7867
rect 17262 8043 17320 8055
rect 17262 7867 17274 8043
rect 17308 7867 17320 8043
rect 17262 7855 17320 7867
rect 19546 8043 19604 8055
rect 19546 7867 19558 8043
rect 19592 7867 19604 8043
rect 19546 7855 19604 7867
rect 19664 8043 19796 8055
rect 19664 7867 19676 8043
rect 19710 7867 19750 8043
rect 19664 7855 19750 7867
rect 17112 7667 17124 7855
rect 17066 7655 17124 7667
rect 19738 7667 19750 7855
rect 19784 7667 19796 8043
rect 19738 7655 19796 7667
rect 19856 8043 19914 8055
rect 19856 7667 19868 8043
rect 19902 7667 19914 8043
rect 19856 7655 19914 7667
rect 19974 8043 20032 8055
rect 19974 7667 19986 8043
rect 20020 7667 20032 8043
rect 19974 7655 20032 7667
rect 20092 8043 20150 8055
rect 20092 7667 20104 8043
rect 20138 7667 20150 8043
rect 20092 7655 20150 7667
rect 20210 8043 20346 8055
rect 20210 7667 20222 8043
rect 20256 7867 20300 8043
rect 20334 7867 20346 8043
rect 20256 7855 20346 7867
rect 20406 8043 20464 8055
rect 20406 7867 20418 8043
rect 20452 7867 20464 8043
rect 20406 7855 20464 7867
rect 22678 8047 22736 8059
rect 22678 7871 22690 8047
rect 22724 7871 22736 8047
rect 22678 7859 22736 7871
rect 22796 8047 22928 8059
rect 22796 7871 22808 8047
rect 22842 7871 22882 8047
rect 22796 7859 22882 7871
rect 20256 7667 20268 7855
rect 20210 7655 20268 7667
rect 22870 7671 22882 7859
rect 22916 7671 22928 8047
rect 22870 7659 22928 7671
rect 22988 8047 23046 8059
rect 22988 7671 23000 8047
rect 23034 7671 23046 8047
rect 22988 7659 23046 7671
rect 23106 8047 23164 8059
rect 23106 7671 23118 8047
rect 23152 7671 23164 8047
rect 23106 7659 23164 7671
rect 23224 8047 23282 8059
rect 23224 7671 23236 8047
rect 23270 7671 23282 8047
rect 23224 7659 23282 7671
rect 23342 8047 23478 8059
rect 23342 7671 23354 8047
rect 23388 7871 23432 8047
rect 23466 7871 23478 8047
rect 23388 7859 23478 7871
rect 23538 8047 23596 8059
rect 23538 7871 23550 8047
rect 23584 7871 23596 8047
rect 23538 7859 23596 7871
rect 25822 8047 25880 8059
rect 25822 7871 25834 8047
rect 25868 7871 25880 8047
rect 25822 7859 25880 7871
rect 25940 8047 26072 8059
rect 25940 7871 25952 8047
rect 25986 7871 26026 8047
rect 25940 7859 26026 7871
rect 23388 7671 23400 7859
rect 23342 7659 23400 7671
rect 26014 7671 26026 7859
rect 26060 7671 26072 8047
rect 26014 7659 26072 7671
rect 26132 8047 26190 8059
rect 26132 7671 26144 8047
rect 26178 7671 26190 8047
rect 26132 7659 26190 7671
rect 26250 8047 26308 8059
rect 26250 7671 26262 8047
rect 26296 7671 26308 8047
rect 26250 7659 26308 7671
rect 26368 8047 26426 8059
rect 26368 7671 26380 8047
rect 26414 7671 26426 8047
rect 26368 7659 26426 7671
rect 26486 8047 26622 8059
rect 26486 7671 26498 8047
rect 26532 7871 26576 8047
rect 26610 7871 26622 8047
rect 26532 7859 26622 7871
rect 26682 8047 26740 8059
rect 26682 7871 26694 8047
rect 26728 7871 26740 8047
rect 26682 7859 26740 7871
rect 26532 7671 26544 7859
rect 26486 7659 26544 7671
rect 2808 5006 2866 5018
rect 2808 4830 2820 5006
rect 2854 4830 2866 5006
rect 2808 4818 2866 4830
rect 2926 5006 2984 5018
rect 2926 4830 2938 5006
rect 2972 4830 2984 5006
rect 2926 4818 2984 4830
rect 3228 5006 3286 5018
rect 3228 4630 3240 5006
rect 3274 4630 3286 5006
rect 3228 4618 3286 4630
rect 3346 5006 3404 5018
rect 3346 4630 3358 5006
rect 3392 4630 3404 5006
rect 3346 4618 3404 4630
rect 3464 5006 3522 5018
rect 3464 4630 3476 5006
rect 3510 4630 3522 5006
rect 3464 4618 3522 4630
rect 3582 5006 3640 5018
rect 3582 4630 3594 5006
rect 3628 4630 3640 5006
rect 3582 4618 3640 4630
rect 3700 5006 3758 5018
rect 3700 4630 3712 5006
rect 3746 4630 3758 5006
rect 4106 5006 4164 5018
rect 4106 4830 4118 5006
rect 4152 4830 4164 5006
rect 4106 4818 4164 4830
rect 4224 5006 4282 5018
rect 4224 4830 4236 5006
rect 4270 4830 4282 5006
rect 4224 4818 4282 4830
rect 4876 5008 4934 5020
rect 4876 4832 4888 5008
rect 4922 4832 4934 5008
rect 4876 4820 4934 4832
rect 4994 5008 5052 5020
rect 4994 4832 5006 5008
rect 5040 4832 5052 5008
rect 4994 4820 5052 4832
rect 5296 5008 5354 5020
rect 3700 4618 3758 4630
rect 5296 4632 5308 5008
rect 5342 4632 5354 5008
rect 5296 4620 5354 4632
rect 5414 5008 5472 5020
rect 5414 4632 5426 5008
rect 5460 4632 5472 5008
rect 5414 4620 5472 4632
rect 5532 5008 5590 5020
rect 5532 4632 5544 5008
rect 5578 4632 5590 5008
rect 5532 4620 5590 4632
rect 5650 5008 5708 5020
rect 5650 4632 5662 5008
rect 5696 4632 5708 5008
rect 5650 4620 5708 4632
rect 5768 5008 5826 5020
rect 5768 4632 5780 5008
rect 5814 4632 5826 5008
rect 6174 5008 6232 5020
rect 6174 4832 6186 5008
rect 6220 4832 6232 5008
rect 6174 4820 6232 4832
rect 6292 5008 6350 5020
rect 19533 6161 19591 6173
rect 6292 4832 6304 5008
rect 6338 4832 6350 5008
rect 6292 4820 6350 4832
rect 6945 5006 7003 5018
rect 6945 4830 6957 5006
rect 6991 4830 7003 5006
rect 6945 4818 7003 4830
rect 7063 5006 7121 5018
rect 7063 4830 7075 5006
rect 7109 4830 7121 5006
rect 7063 4818 7121 4830
rect 7365 5006 7423 5018
rect 5768 4620 5826 4632
rect 7365 4630 7377 5006
rect 7411 4630 7423 5006
rect 7365 4618 7423 4630
rect 7483 5006 7541 5018
rect 7483 4630 7495 5006
rect 7529 4630 7541 5006
rect 7483 4618 7541 4630
rect 7601 5006 7659 5018
rect 7601 4630 7613 5006
rect 7647 4630 7659 5006
rect 7601 4618 7659 4630
rect 7719 5006 7777 5018
rect 7719 4630 7731 5006
rect 7765 4630 7777 5006
rect 7719 4618 7777 4630
rect 7837 5006 7895 5018
rect 7837 4630 7849 5006
rect 7883 4630 7895 5006
rect 8243 5006 8301 5018
rect 8243 4830 8255 5006
rect 8289 4830 8301 5006
rect 8243 4818 8301 4830
rect 8361 5006 8419 5018
rect 8361 4830 8373 5006
rect 8407 4830 8419 5006
rect 8361 4818 8419 4830
rect 9013 5008 9071 5020
rect 9013 4832 9025 5008
rect 9059 4832 9071 5008
rect 9013 4820 9071 4832
rect 9131 5008 9189 5020
rect 9131 4832 9143 5008
rect 9177 4832 9189 5008
rect 9131 4820 9189 4832
rect 9433 5008 9491 5020
rect 7837 4618 7895 4630
rect 9433 4632 9445 5008
rect 9479 4632 9491 5008
rect 9433 4620 9491 4632
rect 9551 5008 9609 5020
rect 9551 4632 9563 5008
rect 9597 4632 9609 5008
rect 9551 4620 9609 4632
rect 9669 5008 9727 5020
rect 9669 4632 9681 5008
rect 9715 4632 9727 5008
rect 9669 4620 9727 4632
rect 9787 5008 9845 5020
rect 9787 4632 9799 5008
rect 9833 4632 9845 5008
rect 9787 4620 9845 4632
rect 9905 5008 9963 5020
rect 9905 4632 9917 5008
rect 9951 4632 9963 5008
rect 10311 5008 10369 5020
rect 10311 4832 10323 5008
rect 10357 4832 10369 5008
rect 10311 4820 10369 4832
rect 10429 5008 10487 5020
rect 10429 4832 10441 5008
rect 10475 4832 10487 5008
rect 10429 4820 10487 4832
rect 11082 5008 11140 5020
rect 11082 4832 11094 5008
rect 11128 4832 11140 5008
rect 11082 4820 11140 4832
rect 11200 5008 11258 5020
rect 11200 4832 11212 5008
rect 11246 4832 11258 5008
rect 11200 4820 11258 4832
rect 11502 5008 11560 5020
rect 9905 4620 9963 4632
rect 11502 4632 11514 5008
rect 11548 4632 11560 5008
rect 11502 4620 11560 4632
rect 11620 5008 11678 5020
rect 11620 4632 11632 5008
rect 11666 4632 11678 5008
rect 11620 4620 11678 4632
rect 11738 5008 11796 5020
rect 11738 4632 11750 5008
rect 11784 4632 11796 5008
rect 11738 4620 11796 4632
rect 11856 5008 11914 5020
rect 11856 4632 11868 5008
rect 11902 4632 11914 5008
rect 11856 4620 11914 4632
rect 11974 5008 12032 5020
rect 11974 4632 11986 5008
rect 12020 4632 12032 5008
rect 12380 5008 12438 5020
rect 12380 4832 12392 5008
rect 12426 4832 12438 5008
rect 12380 4820 12438 4832
rect 12498 5008 12556 5020
rect 12498 4832 12510 5008
rect 12544 4832 12556 5008
rect 12498 4820 12556 4832
rect 13150 5010 13208 5022
rect 13150 4834 13162 5010
rect 13196 4834 13208 5010
rect 13150 4822 13208 4834
rect 13268 5010 13326 5022
rect 13268 4834 13280 5010
rect 13314 4834 13326 5010
rect 13268 4822 13326 4834
rect 13570 5010 13628 5022
rect 11974 4620 12032 4632
rect 13570 4634 13582 5010
rect 13616 4634 13628 5010
rect 13570 4622 13628 4634
rect 13688 5010 13746 5022
rect 13688 4634 13700 5010
rect 13734 4634 13746 5010
rect 13688 4622 13746 4634
rect 13806 5010 13864 5022
rect 13806 4634 13818 5010
rect 13852 4634 13864 5010
rect 13806 4622 13864 4634
rect 13924 5010 13982 5022
rect 13924 4634 13936 5010
rect 13970 4634 13982 5010
rect 13924 4622 13982 4634
rect 14042 5010 14100 5022
rect 14042 4634 14054 5010
rect 14088 4634 14100 5010
rect 14448 5010 14506 5022
rect 14448 4834 14460 5010
rect 14494 4834 14506 5010
rect 14448 4822 14506 4834
rect 14566 5010 14624 5022
rect 19533 5985 19545 6161
rect 19579 5985 19591 6161
rect 19533 5973 19591 5985
rect 19651 6161 19709 6173
rect 19651 5985 19663 6161
rect 19697 5985 19709 6161
rect 19651 5973 19709 5985
rect 20271 6163 20329 6175
rect 20271 5987 20283 6163
rect 20317 5987 20329 6163
rect 20271 5975 20329 5987
rect 20389 6163 20447 6175
rect 20389 5987 20401 6163
rect 20435 5987 20447 6163
rect 20389 5975 20447 5987
rect 21009 6159 21067 6171
rect 21009 5983 21021 6159
rect 21055 5983 21067 6159
rect 21009 5971 21067 5983
rect 21127 6159 21185 6171
rect 21127 5983 21139 6159
rect 21173 5983 21185 6159
rect 21127 5971 21185 5983
rect 21751 6159 21809 6171
rect 21751 5983 21763 6159
rect 21797 5983 21809 6159
rect 21751 5971 21809 5983
rect 21869 6159 21927 6171
rect 21869 5983 21881 6159
rect 21915 5983 21927 6159
rect 21869 5971 21927 5983
rect 22491 6159 22549 6171
rect 22491 5983 22503 6159
rect 22537 5983 22549 6159
rect 22491 5971 22549 5983
rect 22609 6159 22667 6171
rect 22609 5983 22621 6159
rect 22655 5983 22667 6159
rect 22609 5971 22667 5983
rect 23229 6159 23287 6171
rect 23229 5983 23241 6159
rect 23275 5983 23287 6159
rect 23229 5971 23287 5983
rect 23347 6159 23405 6171
rect 23347 5983 23359 6159
rect 23393 5983 23405 6159
rect 23347 5971 23405 5983
rect 23967 6163 24025 6175
rect 23967 5987 23979 6163
rect 24013 5987 24025 6163
rect 23967 5975 24025 5987
rect 24085 6163 24143 6175
rect 24085 5987 24097 6163
rect 24131 5987 24143 6163
rect 24085 5975 24143 5987
rect 24705 6163 24763 6175
rect 24705 5987 24717 6163
rect 24751 5987 24763 6163
rect 24705 5975 24763 5987
rect 24823 6163 24881 6175
rect 24823 5987 24835 6163
rect 24869 5987 24881 6163
rect 24823 5975 24881 5987
rect 14566 4834 14578 5010
rect 14612 4834 14624 5010
rect 14566 4822 14624 4834
rect 15219 5008 15277 5020
rect 15219 4832 15231 5008
rect 15265 4832 15277 5008
rect 15219 4820 15277 4832
rect 15337 5008 15395 5020
rect 15337 4832 15349 5008
rect 15383 4832 15395 5008
rect 15337 4820 15395 4832
rect 15639 5008 15697 5020
rect 14042 4622 14100 4634
rect 15639 4632 15651 5008
rect 15685 4632 15697 5008
rect 15639 4620 15697 4632
rect 15757 5008 15815 5020
rect 15757 4632 15769 5008
rect 15803 4632 15815 5008
rect 15757 4620 15815 4632
rect 15875 5008 15933 5020
rect 15875 4632 15887 5008
rect 15921 4632 15933 5008
rect 15875 4620 15933 4632
rect 15993 5008 16051 5020
rect 15993 4632 16005 5008
rect 16039 4632 16051 5008
rect 15993 4620 16051 4632
rect 16111 5008 16169 5020
rect 16111 4632 16123 5008
rect 16157 4632 16169 5008
rect 16517 5008 16575 5020
rect 16517 4832 16529 5008
rect 16563 4832 16575 5008
rect 16517 4820 16575 4832
rect 16635 5008 16693 5020
rect 16635 4832 16647 5008
rect 16681 4832 16693 5008
rect 16635 4820 16693 4832
rect 17287 5010 17345 5022
rect 17287 4834 17299 5010
rect 17333 4834 17345 5010
rect 17287 4822 17345 4834
rect 17405 5010 17463 5022
rect 17405 4834 17417 5010
rect 17451 4834 17463 5010
rect 17405 4822 17463 4834
rect 17707 5010 17765 5022
rect 16111 4620 16169 4632
rect 17707 4634 17719 5010
rect 17753 4634 17765 5010
rect 17707 4622 17765 4634
rect 17825 5010 17883 5022
rect 17825 4634 17837 5010
rect 17871 4634 17883 5010
rect 17825 4622 17883 4634
rect 17943 5010 18001 5022
rect 17943 4634 17955 5010
rect 17989 4634 18001 5010
rect 17943 4622 18001 4634
rect 18061 5010 18119 5022
rect 18061 4634 18073 5010
rect 18107 4634 18119 5010
rect 18061 4622 18119 4634
rect 18179 5010 18237 5022
rect 18179 4634 18191 5010
rect 18225 4634 18237 5010
rect 18585 5010 18643 5022
rect 18585 4834 18597 5010
rect 18631 4834 18643 5010
rect 18585 4822 18643 4834
rect 18703 5010 18761 5022
rect 18703 4834 18715 5010
rect 18749 4834 18761 5010
rect 18703 4822 18761 4834
rect 18179 4622 18237 4634
rect 1082 795 1140 807
rect 1082 619 1094 795
rect 1128 619 1140 795
rect 1082 607 1140 619
rect 1200 795 1332 807
rect 1200 619 1212 795
rect 1246 619 1286 795
rect 1200 607 1286 619
rect 1274 419 1286 607
rect 1320 419 1332 795
rect 1274 407 1332 419
rect 1392 795 1450 807
rect 1392 419 1404 795
rect 1438 419 1450 795
rect 1392 407 1450 419
rect 1510 795 1568 807
rect 1510 419 1522 795
rect 1556 419 1568 795
rect 1510 407 1568 419
rect 1628 795 1686 807
rect 1628 419 1640 795
rect 1674 419 1686 795
rect 1628 407 1686 419
rect 1746 795 1882 807
rect 1746 419 1758 795
rect 1792 619 1836 795
rect 1870 619 1882 795
rect 1792 607 1882 619
rect 1942 795 2000 807
rect 1942 619 1954 795
rect 1988 619 2000 795
rect 1942 607 2000 619
rect 4226 795 4284 807
rect 4226 619 4238 795
rect 4272 619 4284 795
rect 4226 607 4284 619
rect 4344 795 4476 807
rect 4344 619 4356 795
rect 4390 619 4430 795
rect 4344 607 4430 619
rect 1792 419 1804 607
rect 1746 407 1804 419
rect 4418 419 4430 607
rect 4464 419 4476 795
rect 4418 407 4476 419
rect 4536 795 4594 807
rect 4536 419 4548 795
rect 4582 419 4594 795
rect 4536 407 4594 419
rect 4654 795 4712 807
rect 4654 419 4666 795
rect 4700 419 4712 795
rect 4654 407 4712 419
rect 4772 795 4830 807
rect 4772 419 4784 795
rect 4818 419 4830 795
rect 4772 407 4830 419
rect 4890 795 5026 807
rect 4890 419 4902 795
rect 4936 619 4980 795
rect 5014 619 5026 795
rect 4936 607 5026 619
rect 5086 795 5144 807
rect 5086 619 5098 795
rect 5132 619 5144 795
rect 5086 607 5144 619
rect 7358 799 7416 811
rect 7358 623 7370 799
rect 7404 623 7416 799
rect 7358 611 7416 623
rect 7476 799 7608 811
rect 7476 623 7488 799
rect 7522 623 7562 799
rect 7476 611 7562 623
rect 4936 419 4948 607
rect 4890 407 4948 419
rect 7550 423 7562 611
rect 7596 423 7608 799
rect 7550 411 7608 423
rect 7668 799 7726 811
rect 7668 423 7680 799
rect 7714 423 7726 799
rect 7668 411 7726 423
rect 7786 799 7844 811
rect 7786 423 7798 799
rect 7832 423 7844 799
rect 7786 411 7844 423
rect 7904 799 7962 811
rect 7904 423 7916 799
rect 7950 423 7962 799
rect 7904 411 7962 423
rect 8022 799 8158 811
rect 8022 423 8034 799
rect 8068 623 8112 799
rect 8146 623 8158 799
rect 8068 611 8158 623
rect 8218 799 8276 811
rect 8218 623 8230 799
rect 8264 623 8276 799
rect 8218 611 8276 623
rect 10502 799 10560 811
rect 10502 623 10514 799
rect 10548 623 10560 799
rect 10502 611 10560 623
rect 10620 799 10752 811
rect 10620 623 10632 799
rect 10666 623 10706 799
rect 10620 611 10706 623
rect 8068 423 8080 611
rect 8022 411 8080 423
rect 10694 423 10706 611
rect 10740 423 10752 799
rect 10694 411 10752 423
rect 10812 799 10870 811
rect 10812 423 10824 799
rect 10858 423 10870 799
rect 10812 411 10870 423
rect 10930 799 10988 811
rect 10930 423 10942 799
rect 10976 423 10988 799
rect 10930 411 10988 423
rect 11048 799 11106 811
rect 11048 423 11060 799
rect 11094 423 11106 799
rect 11048 411 11106 423
rect 11166 799 11302 811
rect 11166 423 11178 799
rect 11212 623 11256 799
rect 11290 623 11302 799
rect 11212 611 11302 623
rect 11362 799 11420 811
rect 11362 623 11374 799
rect 11408 623 11420 799
rect 11362 611 11420 623
rect 13704 795 13762 807
rect 13704 619 13716 795
rect 13750 619 13762 795
rect 11212 423 11224 611
rect 11166 411 11224 423
rect 13704 607 13762 619
rect 13822 795 13954 807
rect 13822 619 13834 795
rect 13868 619 13908 795
rect 13822 607 13908 619
rect 13896 419 13908 607
rect 13942 419 13954 795
rect 13896 407 13954 419
rect 14014 795 14072 807
rect 14014 419 14026 795
rect 14060 419 14072 795
rect 14014 407 14072 419
rect 14132 795 14190 807
rect 14132 419 14144 795
rect 14178 419 14190 795
rect 14132 407 14190 419
rect 14250 795 14308 807
rect 14250 419 14262 795
rect 14296 419 14308 795
rect 14250 407 14308 419
rect 14368 795 14504 807
rect 14368 419 14380 795
rect 14414 619 14458 795
rect 14492 619 14504 795
rect 14414 607 14504 619
rect 14564 795 14622 807
rect 14564 619 14576 795
rect 14610 619 14622 795
rect 14564 607 14622 619
rect 16848 795 16906 807
rect 16848 619 16860 795
rect 16894 619 16906 795
rect 16848 607 16906 619
rect 16966 795 17098 807
rect 16966 619 16978 795
rect 17012 619 17052 795
rect 16966 607 17052 619
rect 14414 419 14426 607
rect 14368 407 14426 419
rect 17040 419 17052 607
rect 17086 419 17098 795
rect 17040 407 17098 419
rect 17158 795 17216 807
rect 17158 419 17170 795
rect 17204 419 17216 795
rect 17158 407 17216 419
rect 17276 795 17334 807
rect 17276 419 17288 795
rect 17322 419 17334 795
rect 17276 407 17334 419
rect 17394 795 17452 807
rect 17394 419 17406 795
rect 17440 419 17452 795
rect 17394 407 17452 419
rect 17512 795 17648 807
rect 17512 419 17524 795
rect 17558 619 17602 795
rect 17636 619 17648 795
rect 17558 607 17648 619
rect 17708 795 17766 807
rect 17708 619 17720 795
rect 17754 619 17766 795
rect 17708 607 17766 619
rect 19980 799 20038 811
rect 19980 623 19992 799
rect 20026 623 20038 799
rect 19980 611 20038 623
rect 20098 799 20230 811
rect 20098 623 20110 799
rect 20144 623 20184 799
rect 20098 611 20184 623
rect 17558 419 17570 607
rect 17512 407 17570 419
rect 20172 423 20184 611
rect 20218 423 20230 799
rect 20172 411 20230 423
rect 20290 799 20348 811
rect 20290 423 20302 799
rect 20336 423 20348 799
rect 20290 411 20348 423
rect 20408 799 20466 811
rect 20408 423 20420 799
rect 20454 423 20466 799
rect 20408 411 20466 423
rect 20526 799 20584 811
rect 20526 423 20538 799
rect 20572 423 20584 799
rect 20526 411 20584 423
rect 20644 799 20780 811
rect 20644 423 20656 799
rect 20690 623 20734 799
rect 20768 623 20780 799
rect 20690 611 20780 623
rect 20840 799 20898 811
rect 20840 623 20852 799
rect 20886 623 20898 799
rect 20840 611 20898 623
rect 23124 799 23182 811
rect 23124 623 23136 799
rect 23170 623 23182 799
rect 23124 611 23182 623
rect 23242 799 23374 811
rect 23242 623 23254 799
rect 23288 623 23328 799
rect 23242 611 23328 623
rect 20690 423 20702 611
rect 20644 411 20702 423
rect 23316 423 23328 611
rect 23362 423 23374 799
rect 23316 411 23374 423
rect 23434 799 23492 811
rect 23434 423 23446 799
rect 23480 423 23492 799
rect 23434 411 23492 423
rect 23552 799 23610 811
rect 23552 423 23564 799
rect 23598 423 23610 799
rect 23552 411 23610 423
rect 23670 799 23728 811
rect 23670 423 23682 799
rect 23716 423 23728 799
rect 23670 411 23728 423
rect 23788 799 23924 811
rect 23788 423 23800 799
rect 23834 623 23878 799
rect 23912 623 23924 799
rect 23834 611 23924 623
rect 23984 799 24042 811
rect 23984 623 23996 799
rect 24030 623 24042 799
rect 23984 611 24042 623
rect 23834 423 23846 611
rect 23788 411 23846 423
rect 1114 -3097 1172 -3085
rect 1114 -3273 1126 -3097
rect 1160 -3273 1172 -3097
rect 1114 -3285 1172 -3273
rect 1232 -3097 1364 -3085
rect 1232 -3273 1244 -3097
rect 1278 -3273 1318 -3097
rect 1232 -3285 1318 -3273
rect 1306 -3473 1318 -3285
rect 1352 -3473 1364 -3097
rect 1306 -3485 1364 -3473
rect 1424 -3097 1482 -3085
rect 1424 -3473 1436 -3097
rect 1470 -3473 1482 -3097
rect 1424 -3485 1482 -3473
rect 1542 -3097 1600 -3085
rect 1542 -3473 1554 -3097
rect 1588 -3473 1600 -3097
rect 1542 -3485 1600 -3473
rect 1660 -3097 1718 -3085
rect 1660 -3473 1672 -3097
rect 1706 -3473 1718 -3097
rect 1660 -3485 1718 -3473
rect 1778 -3097 1914 -3085
rect 1778 -3473 1790 -3097
rect 1824 -3273 1868 -3097
rect 1902 -3273 1914 -3097
rect 1824 -3285 1914 -3273
rect 1974 -3097 2032 -3085
rect 1974 -3273 1986 -3097
rect 2020 -3273 2032 -3097
rect 1974 -3285 2032 -3273
rect 4258 -3097 4316 -3085
rect 4258 -3273 4270 -3097
rect 4304 -3273 4316 -3097
rect 4258 -3285 4316 -3273
rect 4376 -3097 4508 -3085
rect 4376 -3273 4388 -3097
rect 4422 -3273 4462 -3097
rect 4376 -3285 4462 -3273
rect 1824 -3473 1836 -3285
rect 1778 -3485 1836 -3473
rect 4450 -3473 4462 -3285
rect 4496 -3473 4508 -3097
rect 4450 -3485 4508 -3473
rect 4568 -3097 4626 -3085
rect 4568 -3473 4580 -3097
rect 4614 -3473 4626 -3097
rect 4568 -3485 4626 -3473
rect 4686 -3097 4744 -3085
rect 4686 -3473 4698 -3097
rect 4732 -3473 4744 -3097
rect 4686 -3485 4744 -3473
rect 4804 -3097 4862 -3085
rect 4804 -3473 4816 -3097
rect 4850 -3473 4862 -3097
rect 4804 -3485 4862 -3473
rect 4922 -3097 5058 -3085
rect 4922 -3473 4934 -3097
rect 4968 -3273 5012 -3097
rect 5046 -3273 5058 -3097
rect 4968 -3285 5058 -3273
rect 5118 -3097 5176 -3085
rect 5118 -3273 5130 -3097
rect 5164 -3273 5176 -3097
rect 5118 -3285 5176 -3273
rect 7390 -3093 7448 -3081
rect 7390 -3269 7402 -3093
rect 7436 -3269 7448 -3093
rect 7390 -3281 7448 -3269
rect 7508 -3093 7640 -3081
rect 7508 -3269 7520 -3093
rect 7554 -3269 7594 -3093
rect 7508 -3281 7594 -3269
rect 4968 -3473 4980 -3285
rect 4922 -3485 4980 -3473
rect 7582 -3469 7594 -3281
rect 7628 -3469 7640 -3093
rect 7582 -3481 7640 -3469
rect 7700 -3093 7758 -3081
rect 7700 -3469 7712 -3093
rect 7746 -3469 7758 -3093
rect 7700 -3481 7758 -3469
rect 7818 -3093 7876 -3081
rect 7818 -3469 7830 -3093
rect 7864 -3469 7876 -3093
rect 7818 -3481 7876 -3469
rect 7936 -3093 7994 -3081
rect 7936 -3469 7948 -3093
rect 7982 -3469 7994 -3093
rect 7936 -3481 7994 -3469
rect 8054 -3093 8190 -3081
rect 8054 -3469 8066 -3093
rect 8100 -3269 8144 -3093
rect 8178 -3269 8190 -3093
rect 8100 -3281 8190 -3269
rect 8250 -3093 8308 -3081
rect 8250 -3269 8262 -3093
rect 8296 -3269 8308 -3093
rect 8250 -3281 8308 -3269
rect 10534 -3093 10592 -3081
rect 10534 -3269 10546 -3093
rect 10580 -3269 10592 -3093
rect 10534 -3281 10592 -3269
rect 10652 -3093 10784 -3081
rect 10652 -3269 10664 -3093
rect 10698 -3269 10738 -3093
rect 10652 -3281 10738 -3269
rect 8100 -3469 8112 -3281
rect 8054 -3481 8112 -3469
rect 10726 -3469 10738 -3281
rect 10772 -3469 10784 -3093
rect 10726 -3481 10784 -3469
rect 10844 -3093 10902 -3081
rect 10844 -3469 10856 -3093
rect 10890 -3469 10902 -3093
rect 10844 -3481 10902 -3469
rect 10962 -3093 11020 -3081
rect 10962 -3469 10974 -3093
rect 11008 -3469 11020 -3093
rect 10962 -3481 11020 -3469
rect 11080 -3093 11138 -3081
rect 11080 -3469 11092 -3093
rect 11126 -3469 11138 -3093
rect 11080 -3481 11138 -3469
rect 11198 -3093 11334 -3081
rect 11198 -3469 11210 -3093
rect 11244 -3269 11288 -3093
rect 11322 -3269 11334 -3093
rect 11244 -3281 11334 -3269
rect 11394 -3093 11452 -3081
rect 11394 -3269 11406 -3093
rect 11440 -3269 11452 -3093
rect 11394 -3281 11452 -3269
rect 13736 -3097 13794 -3085
rect 13736 -3273 13748 -3097
rect 13782 -3273 13794 -3097
rect 11244 -3469 11256 -3281
rect 11198 -3481 11256 -3469
rect 13736 -3285 13794 -3273
rect 13854 -3097 13986 -3085
rect 13854 -3273 13866 -3097
rect 13900 -3273 13940 -3097
rect 13854 -3285 13940 -3273
rect 13928 -3473 13940 -3285
rect 13974 -3473 13986 -3097
rect 13928 -3485 13986 -3473
rect 14046 -3097 14104 -3085
rect 14046 -3473 14058 -3097
rect 14092 -3473 14104 -3097
rect 14046 -3485 14104 -3473
rect 14164 -3097 14222 -3085
rect 14164 -3473 14176 -3097
rect 14210 -3473 14222 -3097
rect 14164 -3485 14222 -3473
rect 14282 -3097 14340 -3085
rect 14282 -3473 14294 -3097
rect 14328 -3473 14340 -3097
rect 14282 -3485 14340 -3473
rect 14400 -3097 14536 -3085
rect 14400 -3473 14412 -3097
rect 14446 -3273 14490 -3097
rect 14524 -3273 14536 -3097
rect 14446 -3285 14536 -3273
rect 14596 -3097 14654 -3085
rect 14596 -3273 14608 -3097
rect 14642 -3273 14654 -3097
rect 14596 -3285 14654 -3273
rect 16880 -3097 16938 -3085
rect 16880 -3273 16892 -3097
rect 16926 -3273 16938 -3097
rect 16880 -3285 16938 -3273
rect 16998 -3097 17130 -3085
rect 16998 -3273 17010 -3097
rect 17044 -3273 17084 -3097
rect 16998 -3285 17084 -3273
rect 14446 -3473 14458 -3285
rect 14400 -3485 14458 -3473
rect 17072 -3473 17084 -3285
rect 17118 -3473 17130 -3097
rect 17072 -3485 17130 -3473
rect 17190 -3097 17248 -3085
rect 17190 -3473 17202 -3097
rect 17236 -3473 17248 -3097
rect 17190 -3485 17248 -3473
rect 17308 -3097 17366 -3085
rect 17308 -3473 17320 -3097
rect 17354 -3473 17366 -3097
rect 17308 -3485 17366 -3473
rect 17426 -3097 17484 -3085
rect 17426 -3473 17438 -3097
rect 17472 -3473 17484 -3097
rect 17426 -3485 17484 -3473
rect 17544 -3097 17680 -3085
rect 17544 -3473 17556 -3097
rect 17590 -3273 17634 -3097
rect 17668 -3273 17680 -3097
rect 17590 -3285 17680 -3273
rect 17740 -3097 17798 -3085
rect 17740 -3273 17752 -3097
rect 17786 -3273 17798 -3097
rect 17740 -3285 17798 -3273
rect 20012 -3093 20070 -3081
rect 20012 -3269 20024 -3093
rect 20058 -3269 20070 -3093
rect 20012 -3281 20070 -3269
rect 20130 -3093 20262 -3081
rect 20130 -3269 20142 -3093
rect 20176 -3269 20216 -3093
rect 20130 -3281 20216 -3269
rect 17590 -3473 17602 -3285
rect 17544 -3485 17602 -3473
rect 20204 -3469 20216 -3281
rect 20250 -3469 20262 -3093
rect 20204 -3481 20262 -3469
rect 20322 -3093 20380 -3081
rect 20322 -3469 20334 -3093
rect 20368 -3469 20380 -3093
rect 20322 -3481 20380 -3469
rect 20440 -3093 20498 -3081
rect 20440 -3469 20452 -3093
rect 20486 -3469 20498 -3093
rect 20440 -3481 20498 -3469
rect 20558 -3093 20616 -3081
rect 20558 -3469 20570 -3093
rect 20604 -3469 20616 -3093
rect 20558 -3481 20616 -3469
rect 20676 -3093 20812 -3081
rect 20676 -3469 20688 -3093
rect 20722 -3269 20766 -3093
rect 20800 -3269 20812 -3093
rect 20722 -3281 20812 -3269
rect 20872 -3093 20930 -3081
rect 20872 -3269 20884 -3093
rect 20918 -3269 20930 -3093
rect 20872 -3281 20930 -3269
rect 23156 -3093 23214 -3081
rect 23156 -3269 23168 -3093
rect 23202 -3269 23214 -3093
rect 23156 -3281 23214 -3269
rect 23274 -3093 23406 -3081
rect 23274 -3269 23286 -3093
rect 23320 -3269 23360 -3093
rect 23274 -3281 23360 -3269
rect 20722 -3469 20734 -3281
rect 20676 -3481 20734 -3469
rect 23348 -3469 23360 -3281
rect 23394 -3469 23406 -3093
rect 23348 -3481 23406 -3469
rect 23466 -3093 23524 -3081
rect 23466 -3469 23478 -3093
rect 23512 -3469 23524 -3093
rect 23466 -3481 23524 -3469
rect 23584 -3093 23642 -3081
rect 23584 -3469 23596 -3093
rect 23630 -3469 23642 -3093
rect 23584 -3481 23642 -3469
rect 23702 -3093 23760 -3081
rect 23702 -3469 23714 -3093
rect 23748 -3469 23760 -3093
rect 23702 -3481 23760 -3469
rect 23820 -3093 23956 -3081
rect 23820 -3469 23832 -3093
rect 23866 -3269 23910 -3093
rect 23944 -3269 23956 -3093
rect 23866 -3281 23956 -3269
rect 24016 -3093 24074 -3081
rect 24016 -3269 24028 -3093
rect 24062 -3269 24074 -3093
rect 24016 -3281 24074 -3269
rect 23866 -3469 23878 -3281
rect 23820 -3481 23878 -3469
<< pdiff >>
rect 895 21980 953 21992
rect 895 21792 907 21980
rect 454 21780 512 21792
rect 454 21604 466 21780
rect 500 21604 512 21780
rect 454 21592 512 21604
rect 572 21780 630 21792
rect 572 21604 584 21780
rect 618 21604 630 21780
rect 572 21592 630 21604
rect 690 21780 748 21792
rect 690 21604 702 21780
rect 736 21604 748 21780
rect 690 21592 748 21604
rect 808 21780 907 21792
rect 808 21604 820 21780
rect 854 21604 907 21780
rect 941 21604 953 21980
rect 808 21592 953 21604
rect 1013 21980 1071 21992
rect 1013 21604 1025 21980
rect 1059 21604 1071 21980
rect 1013 21592 1071 21604
rect 1131 21980 1189 21992
rect 1131 21604 1143 21980
rect 1177 21604 1189 21980
rect 1131 21592 1189 21604
rect 1249 21980 1307 21992
rect 1249 21604 1261 21980
rect 1295 21604 1307 21980
rect 1249 21592 1307 21604
rect 1362 21980 1420 21992
rect 1362 21604 1374 21980
rect 1408 21604 1420 21980
rect 1362 21592 1420 21604
rect 1480 21980 1538 21992
rect 1480 21604 1492 21980
rect 1526 21604 1538 21980
rect 1480 21592 1538 21604
rect 1598 21980 1656 21992
rect 1598 21604 1610 21980
rect 1644 21604 1656 21980
rect 1598 21592 1656 21604
rect 1716 21980 1774 21992
rect 1716 21604 1728 21980
rect 1762 21604 1774 21980
rect 1716 21592 1774 21604
rect 1834 21980 1892 21992
rect 1834 21604 1846 21980
rect 1880 21604 1892 21980
rect 1834 21592 1892 21604
rect 1952 21980 2010 21992
rect 1952 21604 1964 21980
rect 1998 21604 2010 21980
rect 1952 21592 2010 21604
rect 2070 21980 2128 21992
rect 2070 21604 2082 21980
rect 2116 21604 2128 21980
rect 2070 21592 2128 21604
rect 2189 21980 2247 21992
rect 2189 21604 2201 21980
rect 2235 21604 2247 21980
rect 2189 21592 2247 21604
rect 2307 21980 2365 21992
rect 2307 21604 2319 21980
rect 2353 21604 2365 21980
rect 2307 21592 2365 21604
rect 2425 21980 2483 21992
rect 2425 21604 2437 21980
rect 2471 21604 2483 21980
rect 2425 21592 2483 21604
rect 2543 21980 2601 21992
rect 2543 21604 2555 21980
rect 2589 21604 2601 21980
rect 4039 21980 4097 21992
rect 4039 21792 4051 21980
rect 2543 21592 2601 21604
rect 2662 21780 2720 21792
rect 2662 21604 2674 21780
rect 2708 21604 2720 21780
rect 2662 21592 2720 21604
rect 2780 21780 2838 21792
rect 2780 21604 2792 21780
rect 2826 21604 2838 21780
rect 2780 21592 2838 21604
rect 2898 21780 2956 21792
rect 2898 21604 2910 21780
rect 2944 21604 2956 21780
rect 2898 21592 2956 21604
rect 3016 21780 3074 21792
rect 3016 21604 3028 21780
rect 3062 21604 3074 21780
rect 3016 21592 3074 21604
rect 3598 21780 3656 21792
rect 3598 21604 3610 21780
rect 3644 21604 3656 21780
rect 3598 21592 3656 21604
rect 3716 21780 3774 21792
rect 3716 21604 3728 21780
rect 3762 21604 3774 21780
rect 3716 21592 3774 21604
rect 3834 21780 3892 21792
rect 3834 21604 3846 21780
rect 3880 21604 3892 21780
rect 3834 21592 3892 21604
rect 3952 21780 4051 21792
rect 3952 21604 3964 21780
rect 3998 21604 4051 21780
rect 4085 21604 4097 21980
rect 3952 21592 4097 21604
rect 4157 21980 4215 21992
rect 4157 21604 4169 21980
rect 4203 21604 4215 21980
rect 4157 21592 4215 21604
rect 4275 21980 4333 21992
rect 4275 21604 4287 21980
rect 4321 21604 4333 21980
rect 4275 21592 4333 21604
rect 4393 21980 4451 21992
rect 4393 21604 4405 21980
rect 4439 21604 4451 21980
rect 4393 21592 4451 21604
rect 4506 21980 4564 21992
rect 4506 21604 4518 21980
rect 4552 21604 4564 21980
rect 4506 21592 4564 21604
rect 4624 21980 4682 21992
rect 4624 21604 4636 21980
rect 4670 21604 4682 21980
rect 4624 21592 4682 21604
rect 4742 21980 4800 21992
rect 4742 21604 4754 21980
rect 4788 21604 4800 21980
rect 4742 21592 4800 21604
rect 4860 21980 4918 21992
rect 4860 21604 4872 21980
rect 4906 21604 4918 21980
rect 4860 21592 4918 21604
rect 4978 21980 5036 21992
rect 4978 21604 4990 21980
rect 5024 21604 5036 21980
rect 4978 21592 5036 21604
rect 5096 21980 5154 21992
rect 5096 21604 5108 21980
rect 5142 21604 5154 21980
rect 5096 21592 5154 21604
rect 5214 21980 5272 21992
rect 5214 21604 5226 21980
rect 5260 21604 5272 21980
rect 5214 21592 5272 21604
rect 5333 21980 5391 21992
rect 5333 21604 5345 21980
rect 5379 21604 5391 21980
rect 5333 21592 5391 21604
rect 5451 21980 5509 21992
rect 5451 21604 5463 21980
rect 5497 21604 5509 21980
rect 5451 21592 5509 21604
rect 5569 21980 5627 21992
rect 5569 21604 5581 21980
rect 5615 21604 5627 21980
rect 5569 21592 5627 21604
rect 5687 21980 5745 21992
rect 5687 21604 5699 21980
rect 5733 21604 5745 21980
rect 7171 21984 7229 21996
rect 7171 21796 7183 21984
rect 5687 21592 5745 21604
rect 5806 21780 5864 21792
rect 5806 21604 5818 21780
rect 5852 21604 5864 21780
rect 5806 21592 5864 21604
rect 5924 21780 5982 21792
rect 5924 21604 5936 21780
rect 5970 21604 5982 21780
rect 5924 21592 5982 21604
rect 6042 21780 6100 21792
rect 6042 21604 6054 21780
rect 6088 21604 6100 21780
rect 6042 21592 6100 21604
rect 6160 21780 6218 21792
rect 6160 21604 6172 21780
rect 6206 21604 6218 21780
rect 6160 21592 6218 21604
rect 6730 21784 6788 21796
rect 6730 21608 6742 21784
rect 6776 21608 6788 21784
rect 6730 21596 6788 21608
rect 6848 21784 6906 21796
rect 6848 21608 6860 21784
rect 6894 21608 6906 21784
rect 6848 21596 6906 21608
rect 6966 21784 7024 21796
rect 6966 21608 6978 21784
rect 7012 21608 7024 21784
rect 6966 21596 7024 21608
rect 7084 21784 7183 21796
rect 7084 21608 7096 21784
rect 7130 21608 7183 21784
rect 7217 21608 7229 21984
rect 7084 21596 7229 21608
rect 7289 21984 7347 21996
rect 7289 21608 7301 21984
rect 7335 21608 7347 21984
rect 7289 21596 7347 21608
rect 7407 21984 7465 21996
rect 7407 21608 7419 21984
rect 7453 21608 7465 21984
rect 7407 21596 7465 21608
rect 7525 21984 7583 21996
rect 7525 21608 7537 21984
rect 7571 21608 7583 21984
rect 7525 21596 7583 21608
rect 7638 21984 7696 21996
rect 7638 21608 7650 21984
rect 7684 21608 7696 21984
rect 7638 21596 7696 21608
rect 7756 21984 7814 21996
rect 7756 21608 7768 21984
rect 7802 21608 7814 21984
rect 7756 21596 7814 21608
rect 7874 21984 7932 21996
rect 7874 21608 7886 21984
rect 7920 21608 7932 21984
rect 7874 21596 7932 21608
rect 7992 21984 8050 21996
rect 7992 21608 8004 21984
rect 8038 21608 8050 21984
rect 7992 21596 8050 21608
rect 8110 21984 8168 21996
rect 8110 21608 8122 21984
rect 8156 21608 8168 21984
rect 8110 21596 8168 21608
rect 8228 21984 8286 21996
rect 8228 21608 8240 21984
rect 8274 21608 8286 21984
rect 8228 21596 8286 21608
rect 8346 21984 8404 21996
rect 8346 21608 8358 21984
rect 8392 21608 8404 21984
rect 8346 21596 8404 21608
rect 8465 21984 8523 21996
rect 8465 21608 8477 21984
rect 8511 21608 8523 21984
rect 8465 21596 8523 21608
rect 8583 21984 8641 21996
rect 8583 21608 8595 21984
rect 8629 21608 8641 21984
rect 8583 21596 8641 21608
rect 8701 21984 8759 21996
rect 8701 21608 8713 21984
rect 8747 21608 8759 21984
rect 8701 21596 8759 21608
rect 8819 21984 8877 21996
rect 8819 21608 8831 21984
rect 8865 21608 8877 21984
rect 10315 21984 10373 21996
rect 10315 21796 10327 21984
rect 8819 21596 8877 21608
rect 8938 21784 8996 21796
rect 8938 21608 8950 21784
rect 8984 21608 8996 21784
rect 8938 21596 8996 21608
rect 9056 21784 9114 21796
rect 9056 21608 9068 21784
rect 9102 21608 9114 21784
rect 9056 21596 9114 21608
rect 9174 21784 9232 21796
rect 9174 21608 9186 21784
rect 9220 21608 9232 21784
rect 9174 21596 9232 21608
rect 9292 21784 9350 21796
rect 9292 21608 9304 21784
rect 9338 21608 9350 21784
rect 9292 21596 9350 21608
rect 9874 21784 9932 21796
rect 9874 21608 9886 21784
rect 9920 21608 9932 21784
rect 9874 21596 9932 21608
rect 9992 21784 10050 21796
rect 9992 21608 10004 21784
rect 10038 21608 10050 21784
rect 9992 21596 10050 21608
rect 10110 21784 10168 21796
rect 10110 21608 10122 21784
rect 10156 21608 10168 21784
rect 10110 21596 10168 21608
rect 10228 21784 10327 21796
rect 10228 21608 10240 21784
rect 10274 21608 10327 21784
rect 10361 21608 10373 21984
rect 10228 21596 10373 21608
rect 10433 21984 10491 21996
rect 10433 21608 10445 21984
rect 10479 21608 10491 21984
rect 10433 21596 10491 21608
rect 10551 21984 10609 21996
rect 10551 21608 10563 21984
rect 10597 21608 10609 21984
rect 10551 21596 10609 21608
rect 10669 21984 10727 21996
rect 10669 21608 10681 21984
rect 10715 21608 10727 21984
rect 10669 21596 10727 21608
rect 10782 21984 10840 21996
rect 10782 21608 10794 21984
rect 10828 21608 10840 21984
rect 10782 21596 10840 21608
rect 10900 21984 10958 21996
rect 10900 21608 10912 21984
rect 10946 21608 10958 21984
rect 10900 21596 10958 21608
rect 11018 21984 11076 21996
rect 11018 21608 11030 21984
rect 11064 21608 11076 21984
rect 11018 21596 11076 21608
rect 11136 21984 11194 21996
rect 11136 21608 11148 21984
rect 11182 21608 11194 21984
rect 11136 21596 11194 21608
rect 11254 21984 11312 21996
rect 11254 21608 11266 21984
rect 11300 21608 11312 21984
rect 11254 21596 11312 21608
rect 11372 21984 11430 21996
rect 11372 21608 11384 21984
rect 11418 21608 11430 21984
rect 11372 21596 11430 21608
rect 11490 21984 11548 21996
rect 11490 21608 11502 21984
rect 11536 21608 11548 21984
rect 11490 21596 11548 21608
rect 11609 21984 11667 21996
rect 11609 21608 11621 21984
rect 11655 21608 11667 21984
rect 11609 21596 11667 21608
rect 11727 21984 11785 21996
rect 11727 21608 11739 21984
rect 11773 21608 11785 21984
rect 11727 21596 11785 21608
rect 11845 21984 11903 21996
rect 11845 21608 11857 21984
rect 11891 21608 11903 21984
rect 11845 21596 11903 21608
rect 11963 21984 12021 21996
rect 11963 21608 11975 21984
rect 12009 21608 12021 21984
rect 13517 21980 13575 21992
rect 11963 21596 12021 21608
rect 12082 21784 12140 21796
rect 12082 21608 12094 21784
rect 12128 21608 12140 21784
rect 12082 21596 12140 21608
rect 12200 21784 12258 21796
rect 12200 21608 12212 21784
rect 12246 21608 12258 21784
rect 12200 21596 12258 21608
rect 12318 21784 12376 21796
rect 12318 21608 12330 21784
rect 12364 21608 12376 21784
rect 12318 21596 12376 21608
rect 12436 21784 12494 21796
rect 13517 21792 13529 21980
rect 12436 21608 12448 21784
rect 12482 21608 12494 21784
rect 12436 21596 12494 21608
rect 13076 21780 13134 21792
rect 13076 21604 13088 21780
rect 13122 21604 13134 21780
rect 13076 21592 13134 21604
rect 13194 21780 13252 21792
rect 13194 21604 13206 21780
rect 13240 21604 13252 21780
rect 13194 21592 13252 21604
rect 13312 21780 13370 21792
rect 13312 21604 13324 21780
rect 13358 21604 13370 21780
rect 13312 21592 13370 21604
rect 13430 21780 13529 21792
rect 13430 21604 13442 21780
rect 13476 21604 13529 21780
rect 13563 21604 13575 21980
rect 13430 21592 13575 21604
rect 13635 21980 13693 21992
rect 13635 21604 13647 21980
rect 13681 21604 13693 21980
rect 13635 21592 13693 21604
rect 13753 21980 13811 21992
rect 13753 21604 13765 21980
rect 13799 21604 13811 21980
rect 13753 21592 13811 21604
rect 13871 21980 13929 21992
rect 13871 21604 13883 21980
rect 13917 21604 13929 21980
rect 13871 21592 13929 21604
rect 13984 21980 14042 21992
rect 13984 21604 13996 21980
rect 14030 21604 14042 21980
rect 13984 21592 14042 21604
rect 14102 21980 14160 21992
rect 14102 21604 14114 21980
rect 14148 21604 14160 21980
rect 14102 21592 14160 21604
rect 14220 21980 14278 21992
rect 14220 21604 14232 21980
rect 14266 21604 14278 21980
rect 14220 21592 14278 21604
rect 14338 21980 14396 21992
rect 14338 21604 14350 21980
rect 14384 21604 14396 21980
rect 14338 21592 14396 21604
rect 14456 21980 14514 21992
rect 14456 21604 14468 21980
rect 14502 21604 14514 21980
rect 14456 21592 14514 21604
rect 14574 21980 14632 21992
rect 14574 21604 14586 21980
rect 14620 21604 14632 21980
rect 14574 21592 14632 21604
rect 14692 21980 14750 21992
rect 14692 21604 14704 21980
rect 14738 21604 14750 21980
rect 14692 21592 14750 21604
rect 14811 21980 14869 21992
rect 14811 21604 14823 21980
rect 14857 21604 14869 21980
rect 14811 21592 14869 21604
rect 14929 21980 14987 21992
rect 14929 21604 14941 21980
rect 14975 21604 14987 21980
rect 14929 21592 14987 21604
rect 15047 21980 15105 21992
rect 15047 21604 15059 21980
rect 15093 21604 15105 21980
rect 15047 21592 15105 21604
rect 15165 21980 15223 21992
rect 15165 21604 15177 21980
rect 15211 21604 15223 21980
rect 16661 21980 16719 21992
rect 16661 21792 16673 21980
rect 15165 21592 15223 21604
rect 15284 21780 15342 21792
rect 15284 21604 15296 21780
rect 15330 21604 15342 21780
rect 15284 21592 15342 21604
rect 15402 21780 15460 21792
rect 15402 21604 15414 21780
rect 15448 21604 15460 21780
rect 15402 21592 15460 21604
rect 15520 21780 15578 21792
rect 15520 21604 15532 21780
rect 15566 21604 15578 21780
rect 15520 21592 15578 21604
rect 15638 21780 15696 21792
rect 15638 21604 15650 21780
rect 15684 21604 15696 21780
rect 15638 21592 15696 21604
rect 16220 21780 16278 21792
rect 16220 21604 16232 21780
rect 16266 21604 16278 21780
rect 16220 21592 16278 21604
rect 16338 21780 16396 21792
rect 16338 21604 16350 21780
rect 16384 21604 16396 21780
rect 16338 21592 16396 21604
rect 16456 21780 16514 21792
rect 16456 21604 16468 21780
rect 16502 21604 16514 21780
rect 16456 21592 16514 21604
rect 16574 21780 16673 21792
rect 16574 21604 16586 21780
rect 16620 21604 16673 21780
rect 16707 21604 16719 21980
rect 16574 21592 16719 21604
rect 16779 21980 16837 21992
rect 16779 21604 16791 21980
rect 16825 21604 16837 21980
rect 16779 21592 16837 21604
rect 16897 21980 16955 21992
rect 16897 21604 16909 21980
rect 16943 21604 16955 21980
rect 16897 21592 16955 21604
rect 17015 21980 17073 21992
rect 17015 21604 17027 21980
rect 17061 21604 17073 21980
rect 17015 21592 17073 21604
rect 17128 21980 17186 21992
rect 17128 21604 17140 21980
rect 17174 21604 17186 21980
rect 17128 21592 17186 21604
rect 17246 21980 17304 21992
rect 17246 21604 17258 21980
rect 17292 21604 17304 21980
rect 17246 21592 17304 21604
rect 17364 21980 17422 21992
rect 17364 21604 17376 21980
rect 17410 21604 17422 21980
rect 17364 21592 17422 21604
rect 17482 21980 17540 21992
rect 17482 21604 17494 21980
rect 17528 21604 17540 21980
rect 17482 21592 17540 21604
rect 17600 21980 17658 21992
rect 17600 21604 17612 21980
rect 17646 21604 17658 21980
rect 17600 21592 17658 21604
rect 17718 21980 17776 21992
rect 17718 21604 17730 21980
rect 17764 21604 17776 21980
rect 17718 21592 17776 21604
rect 17836 21980 17894 21992
rect 17836 21604 17848 21980
rect 17882 21604 17894 21980
rect 17836 21592 17894 21604
rect 17955 21980 18013 21992
rect 17955 21604 17967 21980
rect 18001 21604 18013 21980
rect 17955 21592 18013 21604
rect 18073 21980 18131 21992
rect 18073 21604 18085 21980
rect 18119 21604 18131 21980
rect 18073 21592 18131 21604
rect 18191 21980 18249 21992
rect 18191 21604 18203 21980
rect 18237 21604 18249 21980
rect 18191 21592 18249 21604
rect 18309 21980 18367 21992
rect 18309 21604 18321 21980
rect 18355 21604 18367 21980
rect 19793 21984 19851 21996
rect 19793 21796 19805 21984
rect 18309 21592 18367 21604
rect 18428 21780 18486 21792
rect 18428 21604 18440 21780
rect 18474 21604 18486 21780
rect 18428 21592 18486 21604
rect 18546 21780 18604 21792
rect 18546 21604 18558 21780
rect 18592 21604 18604 21780
rect 18546 21592 18604 21604
rect 18664 21780 18722 21792
rect 18664 21604 18676 21780
rect 18710 21604 18722 21780
rect 18664 21592 18722 21604
rect 18782 21780 18840 21792
rect 18782 21604 18794 21780
rect 18828 21604 18840 21780
rect 18782 21592 18840 21604
rect 19352 21784 19410 21796
rect 19352 21608 19364 21784
rect 19398 21608 19410 21784
rect 19352 21596 19410 21608
rect 19470 21784 19528 21796
rect 19470 21608 19482 21784
rect 19516 21608 19528 21784
rect 19470 21596 19528 21608
rect 19588 21784 19646 21796
rect 19588 21608 19600 21784
rect 19634 21608 19646 21784
rect 19588 21596 19646 21608
rect 19706 21784 19805 21796
rect 19706 21608 19718 21784
rect 19752 21608 19805 21784
rect 19839 21608 19851 21984
rect 19706 21596 19851 21608
rect 19911 21984 19969 21996
rect 19911 21608 19923 21984
rect 19957 21608 19969 21984
rect 19911 21596 19969 21608
rect 20029 21984 20087 21996
rect 20029 21608 20041 21984
rect 20075 21608 20087 21984
rect 20029 21596 20087 21608
rect 20147 21984 20205 21996
rect 20147 21608 20159 21984
rect 20193 21608 20205 21984
rect 20147 21596 20205 21608
rect 20260 21984 20318 21996
rect 20260 21608 20272 21984
rect 20306 21608 20318 21984
rect 20260 21596 20318 21608
rect 20378 21984 20436 21996
rect 20378 21608 20390 21984
rect 20424 21608 20436 21984
rect 20378 21596 20436 21608
rect 20496 21984 20554 21996
rect 20496 21608 20508 21984
rect 20542 21608 20554 21984
rect 20496 21596 20554 21608
rect 20614 21984 20672 21996
rect 20614 21608 20626 21984
rect 20660 21608 20672 21984
rect 20614 21596 20672 21608
rect 20732 21984 20790 21996
rect 20732 21608 20744 21984
rect 20778 21608 20790 21984
rect 20732 21596 20790 21608
rect 20850 21984 20908 21996
rect 20850 21608 20862 21984
rect 20896 21608 20908 21984
rect 20850 21596 20908 21608
rect 20968 21984 21026 21996
rect 20968 21608 20980 21984
rect 21014 21608 21026 21984
rect 20968 21596 21026 21608
rect 21087 21984 21145 21996
rect 21087 21608 21099 21984
rect 21133 21608 21145 21984
rect 21087 21596 21145 21608
rect 21205 21984 21263 21996
rect 21205 21608 21217 21984
rect 21251 21608 21263 21984
rect 21205 21596 21263 21608
rect 21323 21984 21381 21996
rect 21323 21608 21335 21984
rect 21369 21608 21381 21984
rect 21323 21596 21381 21608
rect 21441 21984 21499 21996
rect 21441 21608 21453 21984
rect 21487 21608 21499 21984
rect 22937 21984 22995 21996
rect 22937 21796 22949 21984
rect 21441 21596 21499 21608
rect 21560 21784 21618 21796
rect 21560 21608 21572 21784
rect 21606 21608 21618 21784
rect 21560 21596 21618 21608
rect 21678 21784 21736 21796
rect 21678 21608 21690 21784
rect 21724 21608 21736 21784
rect 21678 21596 21736 21608
rect 21796 21784 21854 21796
rect 21796 21608 21808 21784
rect 21842 21608 21854 21784
rect 21796 21596 21854 21608
rect 21914 21784 21972 21796
rect 21914 21608 21926 21784
rect 21960 21608 21972 21784
rect 21914 21596 21972 21608
rect 22496 21784 22554 21796
rect 22496 21608 22508 21784
rect 22542 21608 22554 21784
rect 22496 21596 22554 21608
rect 22614 21784 22672 21796
rect 22614 21608 22626 21784
rect 22660 21608 22672 21784
rect 22614 21596 22672 21608
rect 22732 21784 22790 21796
rect 22732 21608 22744 21784
rect 22778 21608 22790 21784
rect 22732 21596 22790 21608
rect 22850 21784 22949 21796
rect 22850 21608 22862 21784
rect 22896 21608 22949 21784
rect 22983 21608 22995 21984
rect 22850 21596 22995 21608
rect 23055 21984 23113 21996
rect 23055 21608 23067 21984
rect 23101 21608 23113 21984
rect 23055 21596 23113 21608
rect 23173 21984 23231 21996
rect 23173 21608 23185 21984
rect 23219 21608 23231 21984
rect 23173 21596 23231 21608
rect 23291 21984 23349 21996
rect 23291 21608 23303 21984
rect 23337 21608 23349 21984
rect 23291 21596 23349 21608
rect 23404 21984 23462 21996
rect 23404 21608 23416 21984
rect 23450 21608 23462 21984
rect 23404 21596 23462 21608
rect 23522 21984 23580 21996
rect 23522 21608 23534 21984
rect 23568 21608 23580 21984
rect 23522 21596 23580 21608
rect 23640 21984 23698 21996
rect 23640 21608 23652 21984
rect 23686 21608 23698 21984
rect 23640 21596 23698 21608
rect 23758 21984 23816 21996
rect 23758 21608 23770 21984
rect 23804 21608 23816 21984
rect 23758 21596 23816 21608
rect 23876 21984 23934 21996
rect 23876 21608 23888 21984
rect 23922 21608 23934 21984
rect 23876 21596 23934 21608
rect 23994 21984 24052 21996
rect 23994 21608 24006 21984
rect 24040 21608 24052 21984
rect 23994 21596 24052 21608
rect 24112 21984 24170 21996
rect 24112 21608 24124 21984
rect 24158 21608 24170 21984
rect 24112 21596 24170 21608
rect 24231 21984 24289 21996
rect 24231 21608 24243 21984
rect 24277 21608 24289 21984
rect 24231 21596 24289 21608
rect 24349 21984 24407 21996
rect 24349 21608 24361 21984
rect 24395 21608 24407 21984
rect 24349 21596 24407 21608
rect 24467 21984 24525 21996
rect 24467 21608 24479 21984
rect 24513 21608 24525 21984
rect 24467 21596 24525 21608
rect 24585 21984 24643 21996
rect 24585 21608 24597 21984
rect 24631 21608 24643 21984
rect 24585 21596 24643 21608
rect 24704 21784 24762 21796
rect 24704 21608 24716 21784
rect 24750 21608 24762 21784
rect 24704 21596 24762 21608
rect 24822 21784 24880 21796
rect 24822 21608 24834 21784
rect 24868 21608 24880 21784
rect 24822 21596 24880 21608
rect 24940 21784 24998 21796
rect 24940 21608 24952 21784
rect 24986 21608 24998 21784
rect 24940 21596 24998 21608
rect 25058 21784 25116 21796
rect 25058 21608 25070 21784
rect 25104 21608 25116 21784
rect 25058 21596 25116 21608
rect 14660 16796 14718 16808
rect 2897 16599 2955 16611
rect 2897 16423 2909 16599
rect 2943 16423 2955 16599
rect 2897 16411 2955 16423
rect 3015 16599 3073 16611
rect 3015 16423 3027 16599
rect 3061 16423 3073 16599
rect 3015 16411 3073 16423
rect 3133 16599 3191 16611
rect 3133 16423 3145 16599
rect 3179 16423 3191 16599
rect 3133 16411 3191 16423
rect 3251 16599 3309 16611
rect 3251 16423 3263 16599
rect 3297 16423 3309 16599
rect 3251 16411 3309 16423
rect 3369 16599 3427 16611
rect 3369 16423 3381 16599
rect 3415 16423 3427 16599
rect 3369 16411 3427 16423
rect 3487 16599 3545 16611
rect 3487 16423 3499 16599
rect 3533 16423 3545 16599
rect 3487 16411 3545 16423
rect 3605 16599 3663 16611
rect 3605 16423 3617 16599
rect 3651 16423 3663 16599
rect 3605 16411 3663 16423
rect 3723 16599 3781 16611
rect 3723 16423 3735 16599
rect 3769 16423 3781 16599
rect 3723 16411 3781 16423
rect 3841 16599 3899 16611
rect 3841 16423 3853 16599
rect 3887 16423 3899 16599
rect 3841 16411 3899 16423
rect 3959 16599 4017 16611
rect 3959 16423 3971 16599
rect 4005 16423 4017 16599
rect 3959 16411 4017 16423
rect 4345 16599 4403 16611
rect 4345 16423 4357 16599
rect 4391 16423 4403 16599
rect 4345 16411 4403 16423
rect 4463 16599 4521 16611
rect 4463 16423 4475 16599
rect 4509 16423 4521 16599
rect 4463 16411 4521 16423
rect 4581 16599 4639 16611
rect 4581 16423 4593 16599
rect 4627 16423 4639 16599
rect 4581 16411 4639 16423
rect 4699 16599 4757 16611
rect 4699 16423 4711 16599
rect 4745 16423 4757 16599
rect 4699 16411 4757 16423
rect 4817 16599 4875 16611
rect 4817 16423 4829 16599
rect 4863 16423 4875 16599
rect 4817 16411 4875 16423
rect 4935 16599 4993 16611
rect 4935 16423 4947 16599
rect 4981 16423 4993 16599
rect 4935 16411 4993 16423
rect 5053 16599 5111 16611
rect 5053 16423 5065 16599
rect 5099 16423 5111 16599
rect 5053 16411 5111 16423
rect 5171 16599 5229 16611
rect 5171 16423 5183 16599
rect 5217 16423 5229 16599
rect 5171 16411 5229 16423
rect 5289 16599 5347 16611
rect 5289 16423 5301 16599
rect 5335 16423 5347 16599
rect 5289 16411 5347 16423
rect 5407 16599 5465 16611
rect 5407 16423 5419 16599
rect 5453 16423 5465 16599
rect 5407 16411 5465 16423
rect 5843 16601 5901 16613
rect 5843 16425 5855 16601
rect 5889 16425 5901 16601
rect 5843 16413 5901 16425
rect 5961 16601 6019 16613
rect 5961 16425 5973 16601
rect 6007 16425 6019 16601
rect 5961 16413 6019 16425
rect 6079 16601 6137 16613
rect 6079 16425 6091 16601
rect 6125 16425 6137 16601
rect 6079 16413 6137 16425
rect 6197 16601 6255 16613
rect 6197 16425 6209 16601
rect 6243 16425 6255 16601
rect 6197 16413 6255 16425
rect 6315 16601 6373 16613
rect 6315 16425 6327 16601
rect 6361 16425 6373 16601
rect 6315 16413 6373 16425
rect 6433 16601 6491 16613
rect 6433 16425 6445 16601
rect 6479 16425 6491 16601
rect 6433 16413 6491 16425
rect 6551 16601 6609 16613
rect 6551 16425 6563 16601
rect 6597 16425 6609 16601
rect 6551 16413 6609 16425
rect 6669 16601 6727 16613
rect 6669 16425 6681 16601
rect 6715 16425 6727 16601
rect 6669 16413 6727 16425
rect 6787 16601 6845 16613
rect 6787 16425 6799 16601
rect 6833 16425 6845 16601
rect 6787 16413 6845 16425
rect 6905 16601 6963 16613
rect 6905 16425 6917 16601
rect 6951 16425 6963 16601
rect 6905 16413 6963 16425
rect 7291 16601 7349 16613
rect 7291 16425 7303 16601
rect 7337 16425 7349 16601
rect 7291 16413 7349 16425
rect 7409 16601 7467 16613
rect 7409 16425 7421 16601
rect 7455 16425 7467 16601
rect 7409 16413 7467 16425
rect 7527 16601 7585 16613
rect 7527 16425 7539 16601
rect 7573 16425 7585 16601
rect 7527 16413 7585 16425
rect 7645 16601 7703 16613
rect 7645 16425 7657 16601
rect 7691 16425 7703 16601
rect 7645 16413 7703 16425
rect 7763 16601 7821 16613
rect 7763 16425 7775 16601
rect 7809 16425 7821 16601
rect 7763 16413 7821 16425
rect 7881 16601 7939 16613
rect 7881 16425 7893 16601
rect 7927 16425 7939 16601
rect 7881 16413 7939 16425
rect 7999 16601 8057 16613
rect 7999 16425 8011 16601
rect 8045 16425 8057 16601
rect 7999 16413 8057 16425
rect 8117 16601 8175 16613
rect 8117 16425 8129 16601
rect 8163 16425 8175 16601
rect 8117 16413 8175 16425
rect 8235 16601 8293 16613
rect 8235 16425 8247 16601
rect 8281 16425 8293 16601
rect 8235 16413 8293 16425
rect 8353 16601 8411 16613
rect 8353 16425 8365 16601
rect 8399 16425 8411 16601
rect 8353 16413 8411 16425
rect 8811 16599 8869 16611
rect 8811 16423 8823 16599
rect 8857 16423 8869 16599
rect 8811 16411 8869 16423
rect 8929 16599 8987 16611
rect 8929 16423 8941 16599
rect 8975 16423 8987 16599
rect 8929 16411 8987 16423
rect 9047 16599 9105 16611
rect 9047 16423 9059 16599
rect 9093 16423 9105 16599
rect 9047 16411 9105 16423
rect 9165 16599 9223 16611
rect 9165 16423 9177 16599
rect 9211 16423 9223 16599
rect 9165 16411 9223 16423
rect 9283 16599 9341 16611
rect 9283 16423 9295 16599
rect 9329 16423 9341 16599
rect 9283 16411 9341 16423
rect 9401 16599 9459 16611
rect 9401 16423 9413 16599
rect 9447 16423 9459 16599
rect 9401 16411 9459 16423
rect 9519 16599 9577 16611
rect 9519 16423 9531 16599
rect 9565 16423 9577 16599
rect 9519 16411 9577 16423
rect 9637 16599 9695 16611
rect 9637 16423 9649 16599
rect 9683 16423 9695 16599
rect 9637 16411 9695 16423
rect 9755 16599 9813 16611
rect 9755 16423 9767 16599
rect 9801 16423 9813 16599
rect 9755 16411 9813 16423
rect 9873 16599 9931 16611
rect 9873 16423 9885 16599
rect 9919 16423 9931 16599
rect 9873 16411 9931 16423
rect 10259 16599 10317 16611
rect 10259 16423 10271 16599
rect 10305 16423 10317 16599
rect 10259 16411 10317 16423
rect 10377 16599 10435 16611
rect 10377 16423 10389 16599
rect 10423 16423 10435 16599
rect 10377 16411 10435 16423
rect 10495 16599 10553 16611
rect 10495 16423 10507 16599
rect 10541 16423 10553 16599
rect 10495 16411 10553 16423
rect 10613 16599 10671 16611
rect 10613 16423 10625 16599
rect 10659 16423 10671 16599
rect 10613 16411 10671 16423
rect 10731 16599 10789 16611
rect 10731 16423 10743 16599
rect 10777 16423 10789 16599
rect 10731 16411 10789 16423
rect 10849 16599 10907 16611
rect 10849 16423 10861 16599
rect 10895 16423 10907 16599
rect 10849 16411 10907 16423
rect 10967 16599 11025 16611
rect 10967 16423 10979 16599
rect 11013 16423 11025 16599
rect 10967 16411 11025 16423
rect 11085 16599 11143 16611
rect 11085 16423 11097 16599
rect 11131 16423 11143 16599
rect 11085 16411 11143 16423
rect 11203 16599 11261 16611
rect 11203 16423 11215 16599
rect 11249 16423 11261 16599
rect 11203 16411 11261 16423
rect 11321 16599 11379 16611
rect 11321 16423 11333 16599
rect 11367 16423 11379 16599
rect 11321 16411 11379 16423
rect 11757 16601 11815 16613
rect 11757 16425 11769 16601
rect 11803 16425 11815 16601
rect 11757 16413 11815 16425
rect 11875 16601 11933 16613
rect 11875 16425 11887 16601
rect 11921 16425 11933 16601
rect 11875 16413 11933 16425
rect 11993 16601 12051 16613
rect 11993 16425 12005 16601
rect 12039 16425 12051 16601
rect 11993 16413 12051 16425
rect 12111 16601 12169 16613
rect 12111 16425 12123 16601
rect 12157 16425 12169 16601
rect 12111 16413 12169 16425
rect 12229 16601 12287 16613
rect 12229 16425 12241 16601
rect 12275 16425 12287 16601
rect 12229 16413 12287 16425
rect 12347 16601 12405 16613
rect 12347 16425 12359 16601
rect 12393 16425 12405 16601
rect 12347 16413 12405 16425
rect 12465 16601 12523 16613
rect 12465 16425 12477 16601
rect 12511 16425 12523 16601
rect 12465 16413 12523 16425
rect 12583 16601 12641 16613
rect 12583 16425 12595 16601
rect 12629 16425 12641 16601
rect 12583 16413 12641 16425
rect 12701 16601 12759 16613
rect 12701 16425 12713 16601
rect 12747 16425 12759 16601
rect 12701 16413 12759 16425
rect 12819 16601 12877 16613
rect 12819 16425 12831 16601
rect 12865 16425 12877 16601
rect 12819 16413 12877 16425
rect 13205 16601 13263 16613
rect 13205 16425 13217 16601
rect 13251 16425 13263 16601
rect 13205 16413 13263 16425
rect 13323 16601 13381 16613
rect 13323 16425 13335 16601
rect 13369 16425 13381 16601
rect 13323 16413 13381 16425
rect 13441 16601 13499 16613
rect 13441 16425 13453 16601
rect 13487 16425 13499 16601
rect 13441 16413 13499 16425
rect 13559 16601 13617 16613
rect 13559 16425 13571 16601
rect 13605 16425 13617 16601
rect 13559 16413 13617 16425
rect 13677 16601 13735 16613
rect 13677 16425 13689 16601
rect 13723 16425 13735 16601
rect 13677 16413 13735 16425
rect 13795 16601 13853 16613
rect 13795 16425 13807 16601
rect 13841 16425 13853 16601
rect 13795 16413 13853 16425
rect 13913 16601 13971 16613
rect 13913 16425 13925 16601
rect 13959 16425 13971 16601
rect 13913 16413 13971 16425
rect 14031 16601 14089 16613
rect 14031 16425 14043 16601
rect 14077 16425 14089 16601
rect 14031 16413 14089 16425
rect 14149 16601 14207 16613
rect 14149 16425 14161 16601
rect 14195 16425 14207 16601
rect 14149 16413 14207 16425
rect 14267 16601 14325 16613
rect 14267 16425 14279 16601
rect 14313 16425 14325 16601
rect 14267 16413 14325 16425
rect 14660 16420 14672 16796
rect 14706 16420 14718 16796
rect 14660 16408 14718 16420
rect 14778 16796 14836 16808
rect 14778 16420 14790 16796
rect 14824 16420 14836 16796
rect 14778 16408 14836 16420
rect 14896 16796 14954 16808
rect 14896 16420 14908 16796
rect 14942 16420 14954 16796
rect 14896 16408 14954 16420
rect 15014 16796 15072 16808
rect 15014 16420 15026 16796
rect 15060 16420 15072 16796
rect 15014 16408 15072 16420
rect 15132 16796 15190 16808
rect 15132 16420 15144 16796
rect 15178 16420 15190 16796
rect 15132 16408 15190 16420
rect 15250 16796 15308 16808
rect 15250 16420 15262 16796
rect 15296 16420 15308 16796
rect 15250 16408 15308 16420
rect 15368 16796 15426 16808
rect 15368 16420 15380 16796
rect 15414 16420 15426 16796
rect 15368 16408 15426 16420
rect 15828 16796 15886 16808
rect 15828 16420 15840 16796
rect 15874 16420 15886 16796
rect 15828 16408 15886 16420
rect 15946 16796 16004 16808
rect 15946 16420 15958 16796
rect 15992 16420 16004 16796
rect 15946 16408 16004 16420
rect 16064 16796 16122 16808
rect 16064 16420 16076 16796
rect 16110 16420 16122 16796
rect 16064 16408 16122 16420
rect 16182 16796 16240 16808
rect 16182 16420 16194 16796
rect 16228 16420 16240 16796
rect 16182 16408 16240 16420
rect 16300 16796 16358 16808
rect 16300 16420 16312 16796
rect 16346 16420 16358 16796
rect 16300 16408 16358 16420
rect 16418 16796 16476 16808
rect 16418 16420 16430 16796
rect 16464 16420 16476 16796
rect 16418 16408 16476 16420
rect 16536 16796 16594 16808
rect 16536 16420 16548 16796
rect 16582 16420 16594 16796
rect 16536 16408 16594 16420
rect 16996 16794 17054 16806
rect 16996 16418 17008 16794
rect 17042 16418 17054 16794
rect 16996 16406 17054 16418
rect 17114 16794 17172 16806
rect 17114 16418 17126 16794
rect 17160 16418 17172 16794
rect 17114 16406 17172 16418
rect 17232 16794 17290 16806
rect 17232 16418 17244 16794
rect 17278 16418 17290 16794
rect 17232 16406 17290 16418
rect 17350 16794 17408 16806
rect 17350 16418 17362 16794
rect 17396 16418 17408 16794
rect 17350 16406 17408 16418
rect 17468 16794 17526 16806
rect 17468 16418 17480 16794
rect 17514 16418 17526 16794
rect 17468 16406 17526 16418
rect 17586 16794 17644 16806
rect 17586 16418 17598 16794
rect 17632 16418 17644 16794
rect 17586 16406 17644 16418
rect 17704 16794 17762 16806
rect 17704 16418 17716 16794
rect 17750 16418 17762 16794
rect 17704 16406 17762 16418
rect 18164 16796 18222 16808
rect 18164 16420 18176 16796
rect 18210 16420 18222 16796
rect 18164 16408 18222 16420
rect 18282 16796 18340 16808
rect 18282 16420 18294 16796
rect 18328 16420 18340 16796
rect 18282 16408 18340 16420
rect 18400 16796 18458 16808
rect 18400 16420 18412 16796
rect 18446 16420 18458 16796
rect 18400 16408 18458 16420
rect 18518 16796 18576 16808
rect 18518 16420 18530 16796
rect 18564 16420 18576 16796
rect 18518 16408 18576 16420
rect 18636 16796 18694 16808
rect 18636 16420 18648 16796
rect 18682 16420 18694 16796
rect 18636 16408 18694 16420
rect 18754 16796 18812 16808
rect 18754 16420 18766 16796
rect 18800 16420 18812 16796
rect 18754 16408 18812 16420
rect 18872 16796 18930 16808
rect 18872 16420 18884 16796
rect 18918 16420 18930 16796
rect 18872 16408 18930 16420
rect 19338 16798 19396 16810
rect 19338 16422 19350 16798
rect 19384 16422 19396 16798
rect 19338 16410 19396 16422
rect 19456 16798 19514 16810
rect 19456 16422 19468 16798
rect 19502 16422 19514 16798
rect 19456 16410 19514 16422
rect 19574 16798 19632 16810
rect 19574 16422 19586 16798
rect 19620 16422 19632 16798
rect 19574 16410 19632 16422
rect 19692 16798 19750 16810
rect 19692 16422 19704 16798
rect 19738 16422 19750 16798
rect 19692 16410 19750 16422
rect 19810 16798 19868 16810
rect 19810 16422 19822 16798
rect 19856 16422 19868 16798
rect 19810 16410 19868 16422
rect 19928 16798 19986 16810
rect 19928 16422 19940 16798
rect 19974 16422 19986 16798
rect 19928 16410 19986 16422
rect 20046 16798 20104 16810
rect 20046 16422 20058 16798
rect 20092 16422 20104 16798
rect 20046 16410 20104 16422
rect 20506 16796 20564 16808
rect 20506 16420 20518 16796
rect 20552 16420 20564 16796
rect 20506 16408 20564 16420
rect 20624 16796 20682 16808
rect 20624 16420 20636 16796
rect 20670 16420 20682 16796
rect 20624 16408 20682 16420
rect 20742 16796 20800 16808
rect 20742 16420 20754 16796
rect 20788 16420 20800 16796
rect 20742 16408 20800 16420
rect 20860 16796 20918 16808
rect 20860 16420 20872 16796
rect 20906 16420 20918 16796
rect 20860 16408 20918 16420
rect 20978 16796 21036 16808
rect 20978 16420 20990 16796
rect 21024 16420 21036 16796
rect 20978 16408 21036 16420
rect 21096 16796 21154 16808
rect 21096 16420 21108 16796
rect 21142 16420 21154 16796
rect 21096 16408 21154 16420
rect 21214 16796 21272 16808
rect 21214 16420 21226 16796
rect 21260 16420 21272 16796
rect 21214 16408 21272 16420
rect 21674 16798 21732 16810
rect 21674 16422 21686 16798
rect 21720 16422 21732 16798
rect 21674 16410 21732 16422
rect 21792 16798 21850 16810
rect 21792 16422 21804 16798
rect 21838 16422 21850 16798
rect 21792 16410 21850 16422
rect 21910 16798 21968 16810
rect 21910 16422 21922 16798
rect 21956 16422 21968 16798
rect 21910 16410 21968 16422
rect 22028 16798 22086 16810
rect 22028 16422 22040 16798
rect 22074 16422 22086 16798
rect 22028 16410 22086 16422
rect 22146 16798 22204 16810
rect 22146 16422 22158 16798
rect 22192 16422 22204 16798
rect 22146 16410 22204 16422
rect 22264 16798 22322 16810
rect 22264 16422 22276 16798
rect 22310 16422 22322 16798
rect 22264 16410 22322 16422
rect 22382 16798 22440 16810
rect 22382 16422 22394 16798
rect 22428 16422 22440 16798
rect 22382 16410 22440 16422
rect 22842 16796 22900 16808
rect 22842 16420 22854 16796
rect 22888 16420 22900 16796
rect 15090 16006 15148 16018
rect 15090 15830 15102 16006
rect 15136 15830 15148 16006
rect 15090 15818 15148 15830
rect 15208 16006 15266 16018
rect 15208 15830 15220 16006
rect 15254 15830 15266 16006
rect 15208 15818 15266 15830
rect 15326 16006 15384 16018
rect 15326 15830 15338 16006
rect 15372 15830 15384 16006
rect 15326 15818 15384 15830
rect 15444 16006 15502 16018
rect 15444 15830 15456 16006
rect 15490 15830 15502 16006
rect 15444 15818 15502 15830
rect 16257 16012 16315 16024
rect 16257 15836 16269 16012
rect 16303 15836 16315 16012
rect 16257 15824 16315 15836
rect 16375 16012 16433 16024
rect 16375 15836 16387 16012
rect 16421 15836 16433 16012
rect 16375 15824 16433 15836
rect 16493 16012 16551 16024
rect 16493 15836 16505 16012
rect 16539 15836 16551 16012
rect 16493 15824 16551 15836
rect 16611 16012 16669 16024
rect 16611 15836 16623 16012
rect 16657 15836 16669 16012
rect 16611 15824 16669 15836
rect 17425 16012 17483 16024
rect 17425 15836 17437 16012
rect 17471 15836 17483 16012
rect 17425 15824 17483 15836
rect 17543 16012 17601 16024
rect 17543 15836 17555 16012
rect 17589 15836 17601 16012
rect 17543 15824 17601 15836
rect 17661 16012 17719 16024
rect 17661 15836 17673 16012
rect 17707 15836 17719 16012
rect 17661 15824 17719 15836
rect 17779 16012 17837 16024
rect 17779 15836 17791 16012
rect 17825 15836 17837 16012
rect 17779 15824 17837 15836
rect 18594 16012 18652 16024
rect 18594 15836 18606 16012
rect 18640 15836 18652 16012
rect 18594 15824 18652 15836
rect 18712 16012 18770 16024
rect 18712 15836 18724 16012
rect 18758 15836 18770 16012
rect 18712 15824 18770 15836
rect 18830 16012 18888 16024
rect 18830 15836 18842 16012
rect 18876 15836 18888 16012
rect 18830 15824 18888 15836
rect 18948 16012 19006 16024
rect 18948 15836 18960 16012
rect 18994 15836 19006 16012
rect 18948 15824 19006 15836
rect 19766 16008 19824 16020
rect 19766 15832 19778 16008
rect 19812 15832 19824 16008
rect 19766 15820 19824 15832
rect 19884 16008 19942 16020
rect 19884 15832 19896 16008
rect 19930 15832 19942 16008
rect 19884 15820 19942 15832
rect 20002 16008 20060 16020
rect 20002 15832 20014 16008
rect 20048 15832 20060 16008
rect 20002 15820 20060 15832
rect 20120 16008 20178 16020
rect 20120 15832 20132 16008
rect 20166 15832 20178 16008
rect 20120 15820 20178 15832
rect 22842 16408 22900 16420
rect 22960 16796 23018 16808
rect 22960 16420 22972 16796
rect 23006 16420 23018 16796
rect 22960 16408 23018 16420
rect 23078 16796 23136 16808
rect 23078 16420 23090 16796
rect 23124 16420 23136 16796
rect 23078 16408 23136 16420
rect 23196 16796 23254 16808
rect 23196 16420 23208 16796
rect 23242 16420 23254 16796
rect 23196 16408 23254 16420
rect 23314 16796 23372 16808
rect 23314 16420 23326 16796
rect 23360 16420 23372 16796
rect 23314 16408 23372 16420
rect 23432 16796 23490 16808
rect 23432 16420 23444 16796
rect 23478 16420 23490 16796
rect 23432 16408 23490 16420
rect 23550 16796 23608 16808
rect 23550 16420 23562 16796
rect 23596 16420 23608 16796
rect 23550 16408 23608 16420
rect 20935 16007 20993 16019
rect 20935 15831 20947 16007
rect 20981 15831 20993 16007
rect 20935 15819 20993 15831
rect 21053 16007 21111 16019
rect 21053 15831 21065 16007
rect 21099 15831 21111 16007
rect 21053 15819 21111 15831
rect 21171 16007 21229 16019
rect 21171 15831 21183 16007
rect 21217 15831 21229 16007
rect 21171 15819 21229 15831
rect 21289 16007 21347 16019
rect 21289 15831 21301 16007
rect 21335 15831 21347 16007
rect 21289 15819 21347 15831
rect 22103 16007 22161 16019
rect 22103 15831 22115 16007
rect 22149 15831 22161 16007
rect 22103 15819 22161 15831
rect 22221 16007 22279 16019
rect 22221 15831 22233 16007
rect 22267 15831 22279 16007
rect 22221 15819 22279 15831
rect 22339 16007 22397 16019
rect 22339 15831 22351 16007
rect 22385 15831 22397 16007
rect 22339 15819 22397 15831
rect 22457 16007 22515 16019
rect 22457 15831 22469 16007
rect 22503 15831 22515 16007
rect 22457 15819 22515 15831
rect 23271 16008 23329 16020
rect 23271 15832 23283 16008
rect 23317 15832 23329 16008
rect 23271 15820 23329 15832
rect 23389 16008 23447 16020
rect 23389 15832 23401 16008
rect 23435 15832 23447 16008
rect 23389 15820 23447 15832
rect 23507 16008 23565 16020
rect 23507 15832 23519 16008
rect 23553 15832 23565 16008
rect 23507 15820 23565 15832
rect 23625 16008 23683 16020
rect 23625 15832 23637 16008
rect 23671 15832 23683 16008
rect 23625 15820 23683 15832
rect 3397 14842 3455 14854
rect 3397 14654 3409 14842
rect 2956 14642 3014 14654
rect 2956 14466 2968 14642
rect 3002 14466 3014 14642
rect 2956 14454 3014 14466
rect 3074 14642 3132 14654
rect 3074 14466 3086 14642
rect 3120 14466 3132 14642
rect 3074 14454 3132 14466
rect 3192 14642 3250 14654
rect 3192 14466 3204 14642
rect 3238 14466 3250 14642
rect 3192 14454 3250 14466
rect 3310 14642 3409 14654
rect 3310 14466 3322 14642
rect 3356 14466 3409 14642
rect 3443 14466 3455 14842
rect 3310 14454 3455 14466
rect 3515 14842 3573 14854
rect 3515 14466 3527 14842
rect 3561 14466 3573 14842
rect 3515 14454 3573 14466
rect 3633 14842 3691 14854
rect 3633 14466 3645 14842
rect 3679 14466 3691 14842
rect 3633 14454 3691 14466
rect 3751 14842 3809 14854
rect 3751 14466 3763 14842
rect 3797 14466 3809 14842
rect 3751 14454 3809 14466
rect 3864 14842 3922 14854
rect 3864 14466 3876 14842
rect 3910 14466 3922 14842
rect 3864 14454 3922 14466
rect 3982 14842 4040 14854
rect 3982 14466 3994 14842
rect 4028 14466 4040 14842
rect 3982 14454 4040 14466
rect 4100 14842 4158 14854
rect 4100 14466 4112 14842
rect 4146 14466 4158 14842
rect 4100 14454 4158 14466
rect 4218 14842 4276 14854
rect 4218 14466 4230 14842
rect 4264 14466 4276 14842
rect 4218 14454 4276 14466
rect 4336 14842 4394 14854
rect 4336 14466 4348 14842
rect 4382 14466 4394 14842
rect 4336 14454 4394 14466
rect 4454 14842 4512 14854
rect 4454 14466 4466 14842
rect 4500 14466 4512 14842
rect 4454 14454 4512 14466
rect 4572 14842 4630 14854
rect 4572 14466 4584 14842
rect 4618 14466 4630 14842
rect 4572 14454 4630 14466
rect 4691 14842 4749 14854
rect 4691 14466 4703 14842
rect 4737 14466 4749 14842
rect 4691 14454 4749 14466
rect 4809 14842 4867 14854
rect 4809 14466 4821 14842
rect 4855 14466 4867 14842
rect 4809 14454 4867 14466
rect 4927 14842 4985 14854
rect 4927 14466 4939 14842
rect 4973 14466 4985 14842
rect 4927 14454 4985 14466
rect 5045 14842 5103 14854
rect 5045 14466 5057 14842
rect 5091 14466 5103 14842
rect 6541 14842 6599 14854
rect 6541 14654 6553 14842
rect 5045 14454 5103 14466
rect 5164 14642 5222 14654
rect 5164 14466 5176 14642
rect 5210 14466 5222 14642
rect 5164 14454 5222 14466
rect 5282 14642 5340 14654
rect 5282 14466 5294 14642
rect 5328 14466 5340 14642
rect 5282 14454 5340 14466
rect 5400 14642 5458 14654
rect 5400 14466 5412 14642
rect 5446 14466 5458 14642
rect 5400 14454 5458 14466
rect 5518 14642 5576 14654
rect 5518 14466 5530 14642
rect 5564 14466 5576 14642
rect 5518 14454 5576 14466
rect 6100 14642 6158 14654
rect 6100 14466 6112 14642
rect 6146 14466 6158 14642
rect 6100 14454 6158 14466
rect 6218 14642 6276 14654
rect 6218 14466 6230 14642
rect 6264 14466 6276 14642
rect 6218 14454 6276 14466
rect 6336 14642 6394 14654
rect 6336 14466 6348 14642
rect 6382 14466 6394 14642
rect 6336 14454 6394 14466
rect 6454 14642 6553 14654
rect 6454 14466 6466 14642
rect 6500 14466 6553 14642
rect 6587 14466 6599 14842
rect 6454 14454 6599 14466
rect 6659 14842 6717 14854
rect 6659 14466 6671 14842
rect 6705 14466 6717 14842
rect 6659 14454 6717 14466
rect 6777 14842 6835 14854
rect 6777 14466 6789 14842
rect 6823 14466 6835 14842
rect 6777 14454 6835 14466
rect 6895 14842 6953 14854
rect 6895 14466 6907 14842
rect 6941 14466 6953 14842
rect 6895 14454 6953 14466
rect 7008 14842 7066 14854
rect 7008 14466 7020 14842
rect 7054 14466 7066 14842
rect 7008 14454 7066 14466
rect 7126 14842 7184 14854
rect 7126 14466 7138 14842
rect 7172 14466 7184 14842
rect 7126 14454 7184 14466
rect 7244 14842 7302 14854
rect 7244 14466 7256 14842
rect 7290 14466 7302 14842
rect 7244 14454 7302 14466
rect 7362 14842 7420 14854
rect 7362 14466 7374 14842
rect 7408 14466 7420 14842
rect 7362 14454 7420 14466
rect 7480 14842 7538 14854
rect 7480 14466 7492 14842
rect 7526 14466 7538 14842
rect 7480 14454 7538 14466
rect 7598 14842 7656 14854
rect 7598 14466 7610 14842
rect 7644 14466 7656 14842
rect 7598 14454 7656 14466
rect 7716 14842 7774 14854
rect 7716 14466 7728 14842
rect 7762 14466 7774 14842
rect 7716 14454 7774 14466
rect 7835 14842 7893 14854
rect 7835 14466 7847 14842
rect 7881 14466 7893 14842
rect 7835 14454 7893 14466
rect 7953 14842 8011 14854
rect 7953 14466 7965 14842
rect 7999 14466 8011 14842
rect 7953 14454 8011 14466
rect 8071 14842 8129 14854
rect 8071 14466 8083 14842
rect 8117 14466 8129 14842
rect 8071 14454 8129 14466
rect 8189 14842 8247 14854
rect 8189 14466 8201 14842
rect 8235 14466 8247 14842
rect 9673 14846 9731 14858
rect 9673 14658 9685 14846
rect 8189 14454 8247 14466
rect 8308 14642 8366 14654
rect 8308 14466 8320 14642
rect 8354 14466 8366 14642
rect 8308 14454 8366 14466
rect 8426 14642 8484 14654
rect 8426 14466 8438 14642
rect 8472 14466 8484 14642
rect 8426 14454 8484 14466
rect 8544 14642 8602 14654
rect 8544 14466 8556 14642
rect 8590 14466 8602 14642
rect 8544 14454 8602 14466
rect 8662 14642 8720 14654
rect 8662 14466 8674 14642
rect 8708 14466 8720 14642
rect 8662 14454 8720 14466
rect 9232 14646 9290 14658
rect 9232 14470 9244 14646
rect 9278 14470 9290 14646
rect 9232 14458 9290 14470
rect 9350 14646 9408 14658
rect 9350 14470 9362 14646
rect 9396 14470 9408 14646
rect 9350 14458 9408 14470
rect 9468 14646 9526 14658
rect 9468 14470 9480 14646
rect 9514 14470 9526 14646
rect 9468 14458 9526 14470
rect 9586 14646 9685 14658
rect 9586 14470 9598 14646
rect 9632 14470 9685 14646
rect 9719 14470 9731 14846
rect 9586 14458 9731 14470
rect 9791 14846 9849 14858
rect 9791 14470 9803 14846
rect 9837 14470 9849 14846
rect 9791 14458 9849 14470
rect 9909 14846 9967 14858
rect 9909 14470 9921 14846
rect 9955 14470 9967 14846
rect 9909 14458 9967 14470
rect 10027 14846 10085 14858
rect 10027 14470 10039 14846
rect 10073 14470 10085 14846
rect 10027 14458 10085 14470
rect 10140 14846 10198 14858
rect 10140 14470 10152 14846
rect 10186 14470 10198 14846
rect 10140 14458 10198 14470
rect 10258 14846 10316 14858
rect 10258 14470 10270 14846
rect 10304 14470 10316 14846
rect 10258 14458 10316 14470
rect 10376 14846 10434 14858
rect 10376 14470 10388 14846
rect 10422 14470 10434 14846
rect 10376 14458 10434 14470
rect 10494 14846 10552 14858
rect 10494 14470 10506 14846
rect 10540 14470 10552 14846
rect 10494 14458 10552 14470
rect 10612 14846 10670 14858
rect 10612 14470 10624 14846
rect 10658 14470 10670 14846
rect 10612 14458 10670 14470
rect 10730 14846 10788 14858
rect 10730 14470 10742 14846
rect 10776 14470 10788 14846
rect 10730 14458 10788 14470
rect 10848 14846 10906 14858
rect 10848 14470 10860 14846
rect 10894 14470 10906 14846
rect 10848 14458 10906 14470
rect 10967 14846 11025 14858
rect 10967 14470 10979 14846
rect 11013 14470 11025 14846
rect 10967 14458 11025 14470
rect 11085 14846 11143 14858
rect 11085 14470 11097 14846
rect 11131 14470 11143 14846
rect 11085 14458 11143 14470
rect 11203 14846 11261 14858
rect 11203 14470 11215 14846
rect 11249 14470 11261 14846
rect 11203 14458 11261 14470
rect 11321 14846 11379 14858
rect 11321 14470 11333 14846
rect 11367 14470 11379 14846
rect 12817 14846 12875 14858
rect 12817 14658 12829 14846
rect 11321 14458 11379 14470
rect 11440 14646 11498 14658
rect 11440 14470 11452 14646
rect 11486 14470 11498 14646
rect 11440 14458 11498 14470
rect 11558 14646 11616 14658
rect 11558 14470 11570 14646
rect 11604 14470 11616 14646
rect 11558 14458 11616 14470
rect 11676 14646 11734 14658
rect 11676 14470 11688 14646
rect 11722 14470 11734 14646
rect 11676 14458 11734 14470
rect 11794 14646 11852 14658
rect 11794 14470 11806 14646
rect 11840 14470 11852 14646
rect 11794 14458 11852 14470
rect 12376 14646 12434 14658
rect 12376 14470 12388 14646
rect 12422 14470 12434 14646
rect 12376 14458 12434 14470
rect 12494 14646 12552 14658
rect 12494 14470 12506 14646
rect 12540 14470 12552 14646
rect 12494 14458 12552 14470
rect 12612 14646 12670 14658
rect 12612 14470 12624 14646
rect 12658 14470 12670 14646
rect 12612 14458 12670 14470
rect 12730 14646 12829 14658
rect 12730 14470 12742 14646
rect 12776 14470 12829 14646
rect 12863 14470 12875 14846
rect 12730 14458 12875 14470
rect 12935 14846 12993 14858
rect 12935 14470 12947 14846
rect 12981 14470 12993 14846
rect 12935 14458 12993 14470
rect 13053 14846 13111 14858
rect 13053 14470 13065 14846
rect 13099 14470 13111 14846
rect 13053 14458 13111 14470
rect 13171 14846 13229 14858
rect 13171 14470 13183 14846
rect 13217 14470 13229 14846
rect 13171 14458 13229 14470
rect 13284 14846 13342 14858
rect 13284 14470 13296 14846
rect 13330 14470 13342 14846
rect 13284 14458 13342 14470
rect 13402 14846 13460 14858
rect 13402 14470 13414 14846
rect 13448 14470 13460 14846
rect 13402 14458 13460 14470
rect 13520 14846 13578 14858
rect 13520 14470 13532 14846
rect 13566 14470 13578 14846
rect 13520 14458 13578 14470
rect 13638 14846 13696 14858
rect 13638 14470 13650 14846
rect 13684 14470 13696 14846
rect 13638 14458 13696 14470
rect 13756 14846 13814 14858
rect 13756 14470 13768 14846
rect 13802 14470 13814 14846
rect 13756 14458 13814 14470
rect 13874 14846 13932 14858
rect 13874 14470 13886 14846
rect 13920 14470 13932 14846
rect 13874 14458 13932 14470
rect 13992 14846 14050 14858
rect 13992 14470 14004 14846
rect 14038 14470 14050 14846
rect 13992 14458 14050 14470
rect 14111 14846 14169 14858
rect 14111 14470 14123 14846
rect 14157 14470 14169 14846
rect 14111 14458 14169 14470
rect 14229 14846 14287 14858
rect 14229 14470 14241 14846
rect 14275 14470 14287 14846
rect 14229 14458 14287 14470
rect 14347 14846 14405 14858
rect 14347 14470 14359 14846
rect 14393 14470 14405 14846
rect 14347 14458 14405 14470
rect 14465 14846 14523 14858
rect 14465 14470 14477 14846
rect 14511 14470 14523 14846
rect 16019 14842 16077 14854
rect 14465 14458 14523 14470
rect 14584 14646 14642 14658
rect 14584 14470 14596 14646
rect 14630 14470 14642 14646
rect 14584 14458 14642 14470
rect 14702 14646 14760 14658
rect 14702 14470 14714 14646
rect 14748 14470 14760 14646
rect 14702 14458 14760 14470
rect 14820 14646 14878 14658
rect 14820 14470 14832 14646
rect 14866 14470 14878 14646
rect 14820 14458 14878 14470
rect 14938 14646 14996 14658
rect 16019 14654 16031 14842
rect 14938 14470 14950 14646
rect 14984 14470 14996 14646
rect 14938 14458 14996 14470
rect 15578 14642 15636 14654
rect 15578 14466 15590 14642
rect 15624 14466 15636 14642
rect 15578 14454 15636 14466
rect 15696 14642 15754 14654
rect 15696 14466 15708 14642
rect 15742 14466 15754 14642
rect 15696 14454 15754 14466
rect 15814 14642 15872 14654
rect 15814 14466 15826 14642
rect 15860 14466 15872 14642
rect 15814 14454 15872 14466
rect 15932 14642 16031 14654
rect 15932 14466 15944 14642
rect 15978 14466 16031 14642
rect 16065 14466 16077 14842
rect 15932 14454 16077 14466
rect 16137 14842 16195 14854
rect 16137 14466 16149 14842
rect 16183 14466 16195 14842
rect 16137 14454 16195 14466
rect 16255 14842 16313 14854
rect 16255 14466 16267 14842
rect 16301 14466 16313 14842
rect 16255 14454 16313 14466
rect 16373 14842 16431 14854
rect 16373 14466 16385 14842
rect 16419 14466 16431 14842
rect 16373 14454 16431 14466
rect 16486 14842 16544 14854
rect 16486 14466 16498 14842
rect 16532 14466 16544 14842
rect 16486 14454 16544 14466
rect 16604 14842 16662 14854
rect 16604 14466 16616 14842
rect 16650 14466 16662 14842
rect 16604 14454 16662 14466
rect 16722 14842 16780 14854
rect 16722 14466 16734 14842
rect 16768 14466 16780 14842
rect 16722 14454 16780 14466
rect 16840 14842 16898 14854
rect 16840 14466 16852 14842
rect 16886 14466 16898 14842
rect 16840 14454 16898 14466
rect 16958 14842 17016 14854
rect 16958 14466 16970 14842
rect 17004 14466 17016 14842
rect 16958 14454 17016 14466
rect 17076 14842 17134 14854
rect 17076 14466 17088 14842
rect 17122 14466 17134 14842
rect 17076 14454 17134 14466
rect 17194 14842 17252 14854
rect 17194 14466 17206 14842
rect 17240 14466 17252 14842
rect 17194 14454 17252 14466
rect 17313 14842 17371 14854
rect 17313 14466 17325 14842
rect 17359 14466 17371 14842
rect 17313 14454 17371 14466
rect 17431 14842 17489 14854
rect 17431 14466 17443 14842
rect 17477 14466 17489 14842
rect 17431 14454 17489 14466
rect 17549 14842 17607 14854
rect 17549 14466 17561 14842
rect 17595 14466 17607 14842
rect 17549 14454 17607 14466
rect 17667 14842 17725 14854
rect 17667 14466 17679 14842
rect 17713 14466 17725 14842
rect 19163 14842 19221 14854
rect 19163 14654 19175 14842
rect 17667 14454 17725 14466
rect 17786 14642 17844 14654
rect 17786 14466 17798 14642
rect 17832 14466 17844 14642
rect 17786 14454 17844 14466
rect 17904 14642 17962 14654
rect 17904 14466 17916 14642
rect 17950 14466 17962 14642
rect 17904 14454 17962 14466
rect 18022 14642 18080 14654
rect 18022 14466 18034 14642
rect 18068 14466 18080 14642
rect 18022 14454 18080 14466
rect 18140 14642 18198 14654
rect 18140 14466 18152 14642
rect 18186 14466 18198 14642
rect 18140 14454 18198 14466
rect 18722 14642 18780 14654
rect 18722 14466 18734 14642
rect 18768 14466 18780 14642
rect 18722 14454 18780 14466
rect 18840 14642 18898 14654
rect 18840 14466 18852 14642
rect 18886 14466 18898 14642
rect 18840 14454 18898 14466
rect 18958 14642 19016 14654
rect 18958 14466 18970 14642
rect 19004 14466 19016 14642
rect 18958 14454 19016 14466
rect 19076 14642 19175 14654
rect 19076 14466 19088 14642
rect 19122 14466 19175 14642
rect 19209 14466 19221 14842
rect 19076 14454 19221 14466
rect 19281 14842 19339 14854
rect 19281 14466 19293 14842
rect 19327 14466 19339 14842
rect 19281 14454 19339 14466
rect 19399 14842 19457 14854
rect 19399 14466 19411 14842
rect 19445 14466 19457 14842
rect 19399 14454 19457 14466
rect 19517 14842 19575 14854
rect 19517 14466 19529 14842
rect 19563 14466 19575 14842
rect 19517 14454 19575 14466
rect 19630 14842 19688 14854
rect 19630 14466 19642 14842
rect 19676 14466 19688 14842
rect 19630 14454 19688 14466
rect 19748 14842 19806 14854
rect 19748 14466 19760 14842
rect 19794 14466 19806 14842
rect 19748 14454 19806 14466
rect 19866 14842 19924 14854
rect 19866 14466 19878 14842
rect 19912 14466 19924 14842
rect 19866 14454 19924 14466
rect 19984 14842 20042 14854
rect 19984 14466 19996 14842
rect 20030 14466 20042 14842
rect 19984 14454 20042 14466
rect 20102 14842 20160 14854
rect 20102 14466 20114 14842
rect 20148 14466 20160 14842
rect 20102 14454 20160 14466
rect 20220 14842 20278 14854
rect 20220 14466 20232 14842
rect 20266 14466 20278 14842
rect 20220 14454 20278 14466
rect 20338 14842 20396 14854
rect 20338 14466 20350 14842
rect 20384 14466 20396 14842
rect 20338 14454 20396 14466
rect 20457 14842 20515 14854
rect 20457 14466 20469 14842
rect 20503 14466 20515 14842
rect 20457 14454 20515 14466
rect 20575 14842 20633 14854
rect 20575 14466 20587 14842
rect 20621 14466 20633 14842
rect 20575 14454 20633 14466
rect 20693 14842 20751 14854
rect 20693 14466 20705 14842
rect 20739 14466 20751 14842
rect 20693 14454 20751 14466
rect 20811 14842 20869 14854
rect 20811 14466 20823 14842
rect 20857 14466 20869 14842
rect 22295 14846 22353 14858
rect 22295 14658 22307 14846
rect 20811 14454 20869 14466
rect 20930 14642 20988 14654
rect 20930 14466 20942 14642
rect 20976 14466 20988 14642
rect 20930 14454 20988 14466
rect 21048 14642 21106 14654
rect 21048 14466 21060 14642
rect 21094 14466 21106 14642
rect 21048 14454 21106 14466
rect 21166 14642 21224 14654
rect 21166 14466 21178 14642
rect 21212 14466 21224 14642
rect 21166 14454 21224 14466
rect 21284 14642 21342 14654
rect 21284 14466 21296 14642
rect 21330 14466 21342 14642
rect 21284 14454 21342 14466
rect 21854 14646 21912 14658
rect 21854 14470 21866 14646
rect 21900 14470 21912 14646
rect 21854 14458 21912 14470
rect 21972 14646 22030 14658
rect 21972 14470 21984 14646
rect 22018 14470 22030 14646
rect 21972 14458 22030 14470
rect 22090 14646 22148 14658
rect 22090 14470 22102 14646
rect 22136 14470 22148 14646
rect 22090 14458 22148 14470
rect 22208 14646 22307 14658
rect 22208 14470 22220 14646
rect 22254 14470 22307 14646
rect 22341 14470 22353 14846
rect 22208 14458 22353 14470
rect 22413 14846 22471 14858
rect 22413 14470 22425 14846
rect 22459 14470 22471 14846
rect 22413 14458 22471 14470
rect 22531 14846 22589 14858
rect 22531 14470 22543 14846
rect 22577 14470 22589 14846
rect 22531 14458 22589 14470
rect 22649 14846 22707 14858
rect 22649 14470 22661 14846
rect 22695 14470 22707 14846
rect 22649 14458 22707 14470
rect 22762 14846 22820 14858
rect 22762 14470 22774 14846
rect 22808 14470 22820 14846
rect 22762 14458 22820 14470
rect 22880 14846 22938 14858
rect 22880 14470 22892 14846
rect 22926 14470 22938 14846
rect 22880 14458 22938 14470
rect 22998 14846 23056 14858
rect 22998 14470 23010 14846
rect 23044 14470 23056 14846
rect 22998 14458 23056 14470
rect 23116 14846 23174 14858
rect 23116 14470 23128 14846
rect 23162 14470 23174 14846
rect 23116 14458 23174 14470
rect 23234 14846 23292 14858
rect 23234 14470 23246 14846
rect 23280 14470 23292 14846
rect 23234 14458 23292 14470
rect 23352 14846 23410 14858
rect 23352 14470 23364 14846
rect 23398 14470 23410 14846
rect 23352 14458 23410 14470
rect 23470 14846 23528 14858
rect 23470 14470 23482 14846
rect 23516 14470 23528 14846
rect 23470 14458 23528 14470
rect 23589 14846 23647 14858
rect 23589 14470 23601 14846
rect 23635 14470 23647 14846
rect 23589 14458 23647 14470
rect 23707 14846 23765 14858
rect 23707 14470 23719 14846
rect 23753 14470 23765 14846
rect 23707 14458 23765 14470
rect 23825 14846 23883 14858
rect 23825 14470 23837 14846
rect 23871 14470 23883 14846
rect 23825 14458 23883 14470
rect 23943 14846 24001 14858
rect 23943 14470 23955 14846
rect 23989 14470 24001 14846
rect 25439 14846 25497 14858
rect 25439 14658 25451 14846
rect 23943 14458 24001 14470
rect 24062 14646 24120 14658
rect 24062 14470 24074 14646
rect 24108 14470 24120 14646
rect 24062 14458 24120 14470
rect 24180 14646 24238 14658
rect 24180 14470 24192 14646
rect 24226 14470 24238 14646
rect 24180 14458 24238 14470
rect 24298 14646 24356 14658
rect 24298 14470 24310 14646
rect 24344 14470 24356 14646
rect 24298 14458 24356 14470
rect 24416 14646 24474 14658
rect 24416 14470 24428 14646
rect 24462 14470 24474 14646
rect 24416 14458 24474 14470
rect 24998 14646 25056 14658
rect 24998 14470 25010 14646
rect 25044 14470 25056 14646
rect 24998 14458 25056 14470
rect 25116 14646 25174 14658
rect 25116 14470 25128 14646
rect 25162 14470 25174 14646
rect 25116 14458 25174 14470
rect 25234 14646 25292 14658
rect 25234 14470 25246 14646
rect 25280 14470 25292 14646
rect 25234 14458 25292 14470
rect 25352 14646 25451 14658
rect 25352 14470 25364 14646
rect 25398 14470 25451 14646
rect 25485 14470 25497 14846
rect 25352 14458 25497 14470
rect 25557 14846 25615 14858
rect 25557 14470 25569 14846
rect 25603 14470 25615 14846
rect 25557 14458 25615 14470
rect 25675 14846 25733 14858
rect 25675 14470 25687 14846
rect 25721 14470 25733 14846
rect 25675 14458 25733 14470
rect 25793 14846 25851 14858
rect 25793 14470 25805 14846
rect 25839 14470 25851 14846
rect 25793 14458 25851 14470
rect 25906 14846 25964 14858
rect 25906 14470 25918 14846
rect 25952 14470 25964 14846
rect 25906 14458 25964 14470
rect 26024 14846 26082 14858
rect 26024 14470 26036 14846
rect 26070 14470 26082 14846
rect 26024 14458 26082 14470
rect 26142 14846 26200 14858
rect 26142 14470 26154 14846
rect 26188 14470 26200 14846
rect 26142 14458 26200 14470
rect 26260 14846 26318 14858
rect 26260 14470 26272 14846
rect 26306 14470 26318 14846
rect 26260 14458 26318 14470
rect 26378 14846 26436 14858
rect 26378 14470 26390 14846
rect 26424 14470 26436 14846
rect 26378 14458 26436 14470
rect 26496 14846 26554 14858
rect 26496 14470 26508 14846
rect 26542 14470 26554 14846
rect 26496 14458 26554 14470
rect 26614 14846 26672 14858
rect 26614 14470 26626 14846
rect 26660 14470 26672 14846
rect 26614 14458 26672 14470
rect 26733 14846 26791 14858
rect 26733 14470 26745 14846
rect 26779 14470 26791 14846
rect 26733 14458 26791 14470
rect 26851 14846 26909 14858
rect 26851 14470 26863 14846
rect 26897 14470 26909 14846
rect 26851 14458 26909 14470
rect 26969 14846 27027 14858
rect 26969 14470 26981 14846
rect 27015 14470 27027 14846
rect 26969 14458 27027 14470
rect 27087 14846 27145 14858
rect 27087 14470 27099 14846
rect 27133 14470 27145 14846
rect 27087 14458 27145 14470
rect 27206 14646 27264 14658
rect 27206 14470 27218 14646
rect 27252 14470 27264 14646
rect 27206 14458 27264 14470
rect 27324 14646 27382 14658
rect 27324 14470 27336 14646
rect 27370 14470 27382 14646
rect 27324 14458 27382 14470
rect 27442 14646 27500 14658
rect 27442 14470 27454 14646
rect 27488 14470 27500 14646
rect 27442 14458 27500 14470
rect 27560 14646 27618 14658
rect 27560 14470 27572 14646
rect 27606 14470 27618 14646
rect 27560 14458 27618 14470
rect 3397 12108 3455 12120
rect 3397 11920 3409 12108
rect 2956 11908 3014 11920
rect 2956 11732 2968 11908
rect 3002 11732 3014 11908
rect 2956 11720 3014 11732
rect 3074 11908 3132 11920
rect 3074 11732 3086 11908
rect 3120 11732 3132 11908
rect 3074 11720 3132 11732
rect 3192 11908 3250 11920
rect 3192 11732 3204 11908
rect 3238 11732 3250 11908
rect 3192 11720 3250 11732
rect 3310 11908 3409 11920
rect 3310 11732 3322 11908
rect 3356 11732 3409 11908
rect 3443 11732 3455 12108
rect 3310 11720 3455 11732
rect 3515 12108 3573 12120
rect 3515 11732 3527 12108
rect 3561 11732 3573 12108
rect 3515 11720 3573 11732
rect 3633 12108 3691 12120
rect 3633 11732 3645 12108
rect 3679 11732 3691 12108
rect 3633 11720 3691 11732
rect 3751 12108 3809 12120
rect 3751 11732 3763 12108
rect 3797 11732 3809 12108
rect 3751 11720 3809 11732
rect 3864 12108 3922 12120
rect 3864 11732 3876 12108
rect 3910 11732 3922 12108
rect 3864 11720 3922 11732
rect 3982 12108 4040 12120
rect 3982 11732 3994 12108
rect 4028 11732 4040 12108
rect 3982 11720 4040 11732
rect 4100 12108 4158 12120
rect 4100 11732 4112 12108
rect 4146 11732 4158 12108
rect 4100 11720 4158 11732
rect 4218 12108 4276 12120
rect 4218 11732 4230 12108
rect 4264 11732 4276 12108
rect 4218 11720 4276 11732
rect 4336 12108 4394 12120
rect 4336 11732 4348 12108
rect 4382 11732 4394 12108
rect 4336 11720 4394 11732
rect 4454 12108 4512 12120
rect 4454 11732 4466 12108
rect 4500 11732 4512 12108
rect 4454 11720 4512 11732
rect 4572 12108 4630 12120
rect 4572 11732 4584 12108
rect 4618 11732 4630 12108
rect 4572 11720 4630 11732
rect 4691 12108 4749 12120
rect 4691 11732 4703 12108
rect 4737 11732 4749 12108
rect 4691 11720 4749 11732
rect 4809 12108 4867 12120
rect 4809 11732 4821 12108
rect 4855 11732 4867 12108
rect 4809 11720 4867 11732
rect 4927 12108 4985 12120
rect 4927 11732 4939 12108
rect 4973 11732 4985 12108
rect 4927 11720 4985 11732
rect 5045 12108 5103 12120
rect 5045 11732 5057 12108
rect 5091 11732 5103 12108
rect 6541 12108 6599 12120
rect 6541 11920 6553 12108
rect 5045 11720 5103 11732
rect 5164 11908 5222 11920
rect 5164 11732 5176 11908
rect 5210 11732 5222 11908
rect 5164 11720 5222 11732
rect 5282 11908 5340 11920
rect 5282 11732 5294 11908
rect 5328 11732 5340 11908
rect 5282 11720 5340 11732
rect 5400 11908 5458 11920
rect 5400 11732 5412 11908
rect 5446 11732 5458 11908
rect 5400 11720 5458 11732
rect 5518 11908 5576 11920
rect 5518 11732 5530 11908
rect 5564 11732 5576 11908
rect 5518 11720 5576 11732
rect 6100 11908 6158 11920
rect 6100 11732 6112 11908
rect 6146 11732 6158 11908
rect 6100 11720 6158 11732
rect 6218 11908 6276 11920
rect 6218 11732 6230 11908
rect 6264 11732 6276 11908
rect 6218 11720 6276 11732
rect 6336 11908 6394 11920
rect 6336 11732 6348 11908
rect 6382 11732 6394 11908
rect 6336 11720 6394 11732
rect 6454 11908 6553 11920
rect 6454 11732 6466 11908
rect 6500 11732 6553 11908
rect 6587 11732 6599 12108
rect 6454 11720 6599 11732
rect 6659 12108 6717 12120
rect 6659 11732 6671 12108
rect 6705 11732 6717 12108
rect 6659 11720 6717 11732
rect 6777 12108 6835 12120
rect 6777 11732 6789 12108
rect 6823 11732 6835 12108
rect 6777 11720 6835 11732
rect 6895 12108 6953 12120
rect 6895 11732 6907 12108
rect 6941 11732 6953 12108
rect 6895 11720 6953 11732
rect 7008 12108 7066 12120
rect 7008 11732 7020 12108
rect 7054 11732 7066 12108
rect 7008 11720 7066 11732
rect 7126 12108 7184 12120
rect 7126 11732 7138 12108
rect 7172 11732 7184 12108
rect 7126 11720 7184 11732
rect 7244 12108 7302 12120
rect 7244 11732 7256 12108
rect 7290 11732 7302 12108
rect 7244 11720 7302 11732
rect 7362 12108 7420 12120
rect 7362 11732 7374 12108
rect 7408 11732 7420 12108
rect 7362 11720 7420 11732
rect 7480 12108 7538 12120
rect 7480 11732 7492 12108
rect 7526 11732 7538 12108
rect 7480 11720 7538 11732
rect 7598 12108 7656 12120
rect 7598 11732 7610 12108
rect 7644 11732 7656 12108
rect 7598 11720 7656 11732
rect 7716 12108 7774 12120
rect 7716 11732 7728 12108
rect 7762 11732 7774 12108
rect 7716 11720 7774 11732
rect 7835 12108 7893 12120
rect 7835 11732 7847 12108
rect 7881 11732 7893 12108
rect 7835 11720 7893 11732
rect 7953 12108 8011 12120
rect 7953 11732 7965 12108
rect 7999 11732 8011 12108
rect 7953 11720 8011 11732
rect 8071 12108 8129 12120
rect 8071 11732 8083 12108
rect 8117 11732 8129 12108
rect 8071 11720 8129 11732
rect 8189 12108 8247 12120
rect 8189 11732 8201 12108
rect 8235 11732 8247 12108
rect 9673 12112 9731 12124
rect 9673 11924 9685 12112
rect 8189 11720 8247 11732
rect 8308 11908 8366 11920
rect 8308 11732 8320 11908
rect 8354 11732 8366 11908
rect 8308 11720 8366 11732
rect 8426 11908 8484 11920
rect 8426 11732 8438 11908
rect 8472 11732 8484 11908
rect 8426 11720 8484 11732
rect 8544 11908 8602 11920
rect 8544 11732 8556 11908
rect 8590 11732 8602 11908
rect 8544 11720 8602 11732
rect 8662 11908 8720 11920
rect 8662 11732 8674 11908
rect 8708 11732 8720 11908
rect 8662 11720 8720 11732
rect 9232 11912 9290 11924
rect 9232 11736 9244 11912
rect 9278 11736 9290 11912
rect 9232 11724 9290 11736
rect 9350 11912 9408 11924
rect 9350 11736 9362 11912
rect 9396 11736 9408 11912
rect 9350 11724 9408 11736
rect 9468 11912 9526 11924
rect 9468 11736 9480 11912
rect 9514 11736 9526 11912
rect 9468 11724 9526 11736
rect 9586 11912 9685 11924
rect 9586 11736 9598 11912
rect 9632 11736 9685 11912
rect 9719 11736 9731 12112
rect 9586 11724 9731 11736
rect 9791 12112 9849 12124
rect 9791 11736 9803 12112
rect 9837 11736 9849 12112
rect 9791 11724 9849 11736
rect 9909 12112 9967 12124
rect 9909 11736 9921 12112
rect 9955 11736 9967 12112
rect 9909 11724 9967 11736
rect 10027 12112 10085 12124
rect 10027 11736 10039 12112
rect 10073 11736 10085 12112
rect 10027 11724 10085 11736
rect 10140 12112 10198 12124
rect 10140 11736 10152 12112
rect 10186 11736 10198 12112
rect 10140 11724 10198 11736
rect 10258 12112 10316 12124
rect 10258 11736 10270 12112
rect 10304 11736 10316 12112
rect 10258 11724 10316 11736
rect 10376 12112 10434 12124
rect 10376 11736 10388 12112
rect 10422 11736 10434 12112
rect 10376 11724 10434 11736
rect 10494 12112 10552 12124
rect 10494 11736 10506 12112
rect 10540 11736 10552 12112
rect 10494 11724 10552 11736
rect 10612 12112 10670 12124
rect 10612 11736 10624 12112
rect 10658 11736 10670 12112
rect 10612 11724 10670 11736
rect 10730 12112 10788 12124
rect 10730 11736 10742 12112
rect 10776 11736 10788 12112
rect 10730 11724 10788 11736
rect 10848 12112 10906 12124
rect 10848 11736 10860 12112
rect 10894 11736 10906 12112
rect 10848 11724 10906 11736
rect 10967 12112 11025 12124
rect 10967 11736 10979 12112
rect 11013 11736 11025 12112
rect 10967 11724 11025 11736
rect 11085 12112 11143 12124
rect 11085 11736 11097 12112
rect 11131 11736 11143 12112
rect 11085 11724 11143 11736
rect 11203 12112 11261 12124
rect 11203 11736 11215 12112
rect 11249 11736 11261 12112
rect 11203 11724 11261 11736
rect 11321 12112 11379 12124
rect 11321 11736 11333 12112
rect 11367 11736 11379 12112
rect 12817 12112 12875 12124
rect 12817 11924 12829 12112
rect 11321 11724 11379 11736
rect 11440 11912 11498 11924
rect 11440 11736 11452 11912
rect 11486 11736 11498 11912
rect 11440 11724 11498 11736
rect 11558 11912 11616 11924
rect 11558 11736 11570 11912
rect 11604 11736 11616 11912
rect 11558 11724 11616 11736
rect 11676 11912 11734 11924
rect 11676 11736 11688 11912
rect 11722 11736 11734 11912
rect 11676 11724 11734 11736
rect 11794 11912 11852 11924
rect 11794 11736 11806 11912
rect 11840 11736 11852 11912
rect 11794 11724 11852 11736
rect 12376 11912 12434 11924
rect 12376 11736 12388 11912
rect 12422 11736 12434 11912
rect 12376 11724 12434 11736
rect 12494 11912 12552 11924
rect 12494 11736 12506 11912
rect 12540 11736 12552 11912
rect 12494 11724 12552 11736
rect 12612 11912 12670 11924
rect 12612 11736 12624 11912
rect 12658 11736 12670 11912
rect 12612 11724 12670 11736
rect 12730 11912 12829 11924
rect 12730 11736 12742 11912
rect 12776 11736 12829 11912
rect 12863 11736 12875 12112
rect 12730 11724 12875 11736
rect 12935 12112 12993 12124
rect 12935 11736 12947 12112
rect 12981 11736 12993 12112
rect 12935 11724 12993 11736
rect 13053 12112 13111 12124
rect 13053 11736 13065 12112
rect 13099 11736 13111 12112
rect 13053 11724 13111 11736
rect 13171 12112 13229 12124
rect 13171 11736 13183 12112
rect 13217 11736 13229 12112
rect 13171 11724 13229 11736
rect 13284 12112 13342 12124
rect 13284 11736 13296 12112
rect 13330 11736 13342 12112
rect 13284 11724 13342 11736
rect 13402 12112 13460 12124
rect 13402 11736 13414 12112
rect 13448 11736 13460 12112
rect 13402 11724 13460 11736
rect 13520 12112 13578 12124
rect 13520 11736 13532 12112
rect 13566 11736 13578 12112
rect 13520 11724 13578 11736
rect 13638 12112 13696 12124
rect 13638 11736 13650 12112
rect 13684 11736 13696 12112
rect 13638 11724 13696 11736
rect 13756 12112 13814 12124
rect 13756 11736 13768 12112
rect 13802 11736 13814 12112
rect 13756 11724 13814 11736
rect 13874 12112 13932 12124
rect 13874 11736 13886 12112
rect 13920 11736 13932 12112
rect 13874 11724 13932 11736
rect 13992 12112 14050 12124
rect 13992 11736 14004 12112
rect 14038 11736 14050 12112
rect 13992 11724 14050 11736
rect 14111 12112 14169 12124
rect 14111 11736 14123 12112
rect 14157 11736 14169 12112
rect 14111 11724 14169 11736
rect 14229 12112 14287 12124
rect 14229 11736 14241 12112
rect 14275 11736 14287 12112
rect 14229 11724 14287 11736
rect 14347 12112 14405 12124
rect 14347 11736 14359 12112
rect 14393 11736 14405 12112
rect 14347 11724 14405 11736
rect 14465 12112 14523 12124
rect 14465 11736 14477 12112
rect 14511 11736 14523 12112
rect 16019 12108 16077 12120
rect 14465 11724 14523 11736
rect 14584 11912 14642 11924
rect 14584 11736 14596 11912
rect 14630 11736 14642 11912
rect 14584 11724 14642 11736
rect 14702 11912 14760 11924
rect 14702 11736 14714 11912
rect 14748 11736 14760 11912
rect 14702 11724 14760 11736
rect 14820 11912 14878 11924
rect 14820 11736 14832 11912
rect 14866 11736 14878 11912
rect 14820 11724 14878 11736
rect 14938 11912 14996 11924
rect 16019 11920 16031 12108
rect 14938 11736 14950 11912
rect 14984 11736 14996 11912
rect 14938 11724 14996 11736
rect 15578 11908 15636 11920
rect 15578 11732 15590 11908
rect 15624 11732 15636 11908
rect 15578 11720 15636 11732
rect 15696 11908 15754 11920
rect 15696 11732 15708 11908
rect 15742 11732 15754 11908
rect 15696 11720 15754 11732
rect 15814 11908 15872 11920
rect 15814 11732 15826 11908
rect 15860 11732 15872 11908
rect 15814 11720 15872 11732
rect 15932 11908 16031 11920
rect 15932 11732 15944 11908
rect 15978 11732 16031 11908
rect 16065 11732 16077 12108
rect 15932 11720 16077 11732
rect 16137 12108 16195 12120
rect 16137 11732 16149 12108
rect 16183 11732 16195 12108
rect 16137 11720 16195 11732
rect 16255 12108 16313 12120
rect 16255 11732 16267 12108
rect 16301 11732 16313 12108
rect 16255 11720 16313 11732
rect 16373 12108 16431 12120
rect 16373 11732 16385 12108
rect 16419 11732 16431 12108
rect 16373 11720 16431 11732
rect 16486 12108 16544 12120
rect 16486 11732 16498 12108
rect 16532 11732 16544 12108
rect 16486 11720 16544 11732
rect 16604 12108 16662 12120
rect 16604 11732 16616 12108
rect 16650 11732 16662 12108
rect 16604 11720 16662 11732
rect 16722 12108 16780 12120
rect 16722 11732 16734 12108
rect 16768 11732 16780 12108
rect 16722 11720 16780 11732
rect 16840 12108 16898 12120
rect 16840 11732 16852 12108
rect 16886 11732 16898 12108
rect 16840 11720 16898 11732
rect 16958 12108 17016 12120
rect 16958 11732 16970 12108
rect 17004 11732 17016 12108
rect 16958 11720 17016 11732
rect 17076 12108 17134 12120
rect 17076 11732 17088 12108
rect 17122 11732 17134 12108
rect 17076 11720 17134 11732
rect 17194 12108 17252 12120
rect 17194 11732 17206 12108
rect 17240 11732 17252 12108
rect 17194 11720 17252 11732
rect 17313 12108 17371 12120
rect 17313 11732 17325 12108
rect 17359 11732 17371 12108
rect 17313 11720 17371 11732
rect 17431 12108 17489 12120
rect 17431 11732 17443 12108
rect 17477 11732 17489 12108
rect 17431 11720 17489 11732
rect 17549 12108 17607 12120
rect 17549 11732 17561 12108
rect 17595 11732 17607 12108
rect 17549 11720 17607 11732
rect 17667 12108 17725 12120
rect 17667 11732 17679 12108
rect 17713 11732 17725 12108
rect 19163 12108 19221 12120
rect 19163 11920 19175 12108
rect 17667 11720 17725 11732
rect 17786 11908 17844 11920
rect 17786 11732 17798 11908
rect 17832 11732 17844 11908
rect 17786 11720 17844 11732
rect 17904 11908 17962 11920
rect 17904 11732 17916 11908
rect 17950 11732 17962 11908
rect 17904 11720 17962 11732
rect 18022 11908 18080 11920
rect 18022 11732 18034 11908
rect 18068 11732 18080 11908
rect 18022 11720 18080 11732
rect 18140 11908 18198 11920
rect 18140 11732 18152 11908
rect 18186 11732 18198 11908
rect 18140 11720 18198 11732
rect 18722 11908 18780 11920
rect 18722 11732 18734 11908
rect 18768 11732 18780 11908
rect 18722 11720 18780 11732
rect 18840 11908 18898 11920
rect 18840 11732 18852 11908
rect 18886 11732 18898 11908
rect 18840 11720 18898 11732
rect 18958 11908 19016 11920
rect 18958 11732 18970 11908
rect 19004 11732 19016 11908
rect 18958 11720 19016 11732
rect 19076 11908 19175 11920
rect 19076 11732 19088 11908
rect 19122 11732 19175 11908
rect 19209 11732 19221 12108
rect 19076 11720 19221 11732
rect 19281 12108 19339 12120
rect 19281 11732 19293 12108
rect 19327 11732 19339 12108
rect 19281 11720 19339 11732
rect 19399 12108 19457 12120
rect 19399 11732 19411 12108
rect 19445 11732 19457 12108
rect 19399 11720 19457 11732
rect 19517 12108 19575 12120
rect 19517 11732 19529 12108
rect 19563 11732 19575 12108
rect 19517 11720 19575 11732
rect 19630 12108 19688 12120
rect 19630 11732 19642 12108
rect 19676 11732 19688 12108
rect 19630 11720 19688 11732
rect 19748 12108 19806 12120
rect 19748 11732 19760 12108
rect 19794 11732 19806 12108
rect 19748 11720 19806 11732
rect 19866 12108 19924 12120
rect 19866 11732 19878 12108
rect 19912 11732 19924 12108
rect 19866 11720 19924 11732
rect 19984 12108 20042 12120
rect 19984 11732 19996 12108
rect 20030 11732 20042 12108
rect 19984 11720 20042 11732
rect 20102 12108 20160 12120
rect 20102 11732 20114 12108
rect 20148 11732 20160 12108
rect 20102 11720 20160 11732
rect 20220 12108 20278 12120
rect 20220 11732 20232 12108
rect 20266 11732 20278 12108
rect 20220 11720 20278 11732
rect 20338 12108 20396 12120
rect 20338 11732 20350 12108
rect 20384 11732 20396 12108
rect 20338 11720 20396 11732
rect 20457 12108 20515 12120
rect 20457 11732 20469 12108
rect 20503 11732 20515 12108
rect 20457 11720 20515 11732
rect 20575 12108 20633 12120
rect 20575 11732 20587 12108
rect 20621 11732 20633 12108
rect 20575 11720 20633 11732
rect 20693 12108 20751 12120
rect 20693 11732 20705 12108
rect 20739 11732 20751 12108
rect 20693 11720 20751 11732
rect 20811 12108 20869 12120
rect 20811 11732 20823 12108
rect 20857 11732 20869 12108
rect 22295 12112 22353 12124
rect 22295 11924 22307 12112
rect 20811 11720 20869 11732
rect 20930 11908 20988 11920
rect 20930 11732 20942 11908
rect 20976 11732 20988 11908
rect 20930 11720 20988 11732
rect 21048 11908 21106 11920
rect 21048 11732 21060 11908
rect 21094 11732 21106 11908
rect 21048 11720 21106 11732
rect 21166 11908 21224 11920
rect 21166 11732 21178 11908
rect 21212 11732 21224 11908
rect 21166 11720 21224 11732
rect 21284 11908 21342 11920
rect 21284 11732 21296 11908
rect 21330 11732 21342 11908
rect 21284 11720 21342 11732
rect 21854 11912 21912 11924
rect 21854 11736 21866 11912
rect 21900 11736 21912 11912
rect 21854 11724 21912 11736
rect 21972 11912 22030 11924
rect 21972 11736 21984 11912
rect 22018 11736 22030 11912
rect 21972 11724 22030 11736
rect 22090 11912 22148 11924
rect 22090 11736 22102 11912
rect 22136 11736 22148 11912
rect 22090 11724 22148 11736
rect 22208 11912 22307 11924
rect 22208 11736 22220 11912
rect 22254 11736 22307 11912
rect 22341 11736 22353 12112
rect 22208 11724 22353 11736
rect 22413 12112 22471 12124
rect 22413 11736 22425 12112
rect 22459 11736 22471 12112
rect 22413 11724 22471 11736
rect 22531 12112 22589 12124
rect 22531 11736 22543 12112
rect 22577 11736 22589 12112
rect 22531 11724 22589 11736
rect 22649 12112 22707 12124
rect 22649 11736 22661 12112
rect 22695 11736 22707 12112
rect 22649 11724 22707 11736
rect 22762 12112 22820 12124
rect 22762 11736 22774 12112
rect 22808 11736 22820 12112
rect 22762 11724 22820 11736
rect 22880 12112 22938 12124
rect 22880 11736 22892 12112
rect 22926 11736 22938 12112
rect 22880 11724 22938 11736
rect 22998 12112 23056 12124
rect 22998 11736 23010 12112
rect 23044 11736 23056 12112
rect 22998 11724 23056 11736
rect 23116 12112 23174 12124
rect 23116 11736 23128 12112
rect 23162 11736 23174 12112
rect 23116 11724 23174 11736
rect 23234 12112 23292 12124
rect 23234 11736 23246 12112
rect 23280 11736 23292 12112
rect 23234 11724 23292 11736
rect 23352 12112 23410 12124
rect 23352 11736 23364 12112
rect 23398 11736 23410 12112
rect 23352 11724 23410 11736
rect 23470 12112 23528 12124
rect 23470 11736 23482 12112
rect 23516 11736 23528 12112
rect 23470 11724 23528 11736
rect 23589 12112 23647 12124
rect 23589 11736 23601 12112
rect 23635 11736 23647 12112
rect 23589 11724 23647 11736
rect 23707 12112 23765 12124
rect 23707 11736 23719 12112
rect 23753 11736 23765 12112
rect 23707 11724 23765 11736
rect 23825 12112 23883 12124
rect 23825 11736 23837 12112
rect 23871 11736 23883 12112
rect 23825 11724 23883 11736
rect 23943 12112 24001 12124
rect 23943 11736 23955 12112
rect 23989 11736 24001 12112
rect 25439 12112 25497 12124
rect 25439 11924 25451 12112
rect 23943 11724 24001 11736
rect 24062 11912 24120 11924
rect 24062 11736 24074 11912
rect 24108 11736 24120 11912
rect 24062 11724 24120 11736
rect 24180 11912 24238 11924
rect 24180 11736 24192 11912
rect 24226 11736 24238 11912
rect 24180 11724 24238 11736
rect 24298 11912 24356 11924
rect 24298 11736 24310 11912
rect 24344 11736 24356 11912
rect 24298 11724 24356 11736
rect 24416 11912 24474 11924
rect 24416 11736 24428 11912
rect 24462 11736 24474 11912
rect 24416 11724 24474 11736
rect 24998 11912 25056 11924
rect 24998 11736 25010 11912
rect 25044 11736 25056 11912
rect 24998 11724 25056 11736
rect 25116 11912 25174 11924
rect 25116 11736 25128 11912
rect 25162 11736 25174 11912
rect 25116 11724 25174 11736
rect 25234 11912 25292 11924
rect 25234 11736 25246 11912
rect 25280 11736 25292 11912
rect 25234 11724 25292 11736
rect 25352 11912 25451 11924
rect 25352 11736 25364 11912
rect 25398 11736 25451 11912
rect 25485 11736 25497 12112
rect 25352 11724 25497 11736
rect 25557 12112 25615 12124
rect 25557 11736 25569 12112
rect 25603 11736 25615 12112
rect 25557 11724 25615 11736
rect 25675 12112 25733 12124
rect 25675 11736 25687 12112
rect 25721 11736 25733 12112
rect 25675 11724 25733 11736
rect 25793 12112 25851 12124
rect 25793 11736 25805 12112
rect 25839 11736 25851 12112
rect 25793 11724 25851 11736
rect 25906 12112 25964 12124
rect 25906 11736 25918 12112
rect 25952 11736 25964 12112
rect 25906 11724 25964 11736
rect 26024 12112 26082 12124
rect 26024 11736 26036 12112
rect 26070 11736 26082 12112
rect 26024 11724 26082 11736
rect 26142 12112 26200 12124
rect 26142 11736 26154 12112
rect 26188 11736 26200 12112
rect 26142 11724 26200 11736
rect 26260 12112 26318 12124
rect 26260 11736 26272 12112
rect 26306 11736 26318 12112
rect 26260 11724 26318 11736
rect 26378 12112 26436 12124
rect 26378 11736 26390 12112
rect 26424 11736 26436 12112
rect 26378 11724 26436 11736
rect 26496 12112 26554 12124
rect 26496 11736 26508 12112
rect 26542 11736 26554 12112
rect 26496 11724 26554 11736
rect 26614 12112 26672 12124
rect 26614 11736 26626 12112
rect 26660 11736 26672 12112
rect 26614 11724 26672 11736
rect 26733 12112 26791 12124
rect 26733 11736 26745 12112
rect 26779 11736 26791 12112
rect 26733 11724 26791 11736
rect 26851 12112 26909 12124
rect 26851 11736 26863 12112
rect 26897 11736 26909 12112
rect 26851 11724 26909 11736
rect 26969 12112 27027 12124
rect 26969 11736 26981 12112
rect 27015 11736 27027 12112
rect 26969 11724 27027 11736
rect 27087 12112 27145 12124
rect 27087 11736 27099 12112
rect 27133 11736 27145 12112
rect 27087 11724 27145 11736
rect 27206 11912 27264 11924
rect 27206 11736 27218 11912
rect 27252 11736 27264 11912
rect 27206 11724 27264 11736
rect 27324 11912 27382 11924
rect 27324 11736 27336 11912
rect 27370 11736 27382 11912
rect 27324 11724 27382 11736
rect 27442 11912 27500 11924
rect 27442 11736 27454 11912
rect 27488 11736 27500 11912
rect 27442 11724 27500 11736
rect 27560 11912 27618 11924
rect 27560 11736 27572 11912
rect 27606 11736 27618 11912
rect 27560 11724 27618 11736
rect 3387 9376 3445 9388
rect 3387 9188 3399 9376
rect 2946 9176 3004 9188
rect 2946 9000 2958 9176
rect 2992 9000 3004 9176
rect 2946 8988 3004 9000
rect 3064 9176 3122 9188
rect 3064 9000 3076 9176
rect 3110 9000 3122 9176
rect 3064 8988 3122 9000
rect 3182 9176 3240 9188
rect 3182 9000 3194 9176
rect 3228 9000 3240 9176
rect 3182 8988 3240 9000
rect 3300 9176 3399 9188
rect 3300 9000 3312 9176
rect 3346 9000 3399 9176
rect 3433 9000 3445 9376
rect 3300 8988 3445 9000
rect 3505 9376 3563 9388
rect 3505 9000 3517 9376
rect 3551 9000 3563 9376
rect 3505 8988 3563 9000
rect 3623 9376 3681 9388
rect 3623 9000 3635 9376
rect 3669 9000 3681 9376
rect 3623 8988 3681 9000
rect 3741 9376 3799 9388
rect 3741 9000 3753 9376
rect 3787 9000 3799 9376
rect 3741 8988 3799 9000
rect 3854 9376 3912 9388
rect 3854 9000 3866 9376
rect 3900 9000 3912 9376
rect 3854 8988 3912 9000
rect 3972 9376 4030 9388
rect 3972 9000 3984 9376
rect 4018 9000 4030 9376
rect 3972 8988 4030 9000
rect 4090 9376 4148 9388
rect 4090 9000 4102 9376
rect 4136 9000 4148 9376
rect 4090 8988 4148 9000
rect 4208 9376 4266 9388
rect 4208 9000 4220 9376
rect 4254 9000 4266 9376
rect 4208 8988 4266 9000
rect 4326 9376 4384 9388
rect 4326 9000 4338 9376
rect 4372 9000 4384 9376
rect 4326 8988 4384 9000
rect 4444 9376 4502 9388
rect 4444 9000 4456 9376
rect 4490 9000 4502 9376
rect 4444 8988 4502 9000
rect 4562 9376 4620 9388
rect 4562 9000 4574 9376
rect 4608 9000 4620 9376
rect 4562 8988 4620 9000
rect 4681 9376 4739 9388
rect 4681 9000 4693 9376
rect 4727 9000 4739 9376
rect 4681 8988 4739 9000
rect 4799 9376 4857 9388
rect 4799 9000 4811 9376
rect 4845 9000 4857 9376
rect 4799 8988 4857 9000
rect 4917 9376 4975 9388
rect 4917 9000 4929 9376
rect 4963 9000 4975 9376
rect 4917 8988 4975 9000
rect 5035 9376 5093 9388
rect 5035 9000 5047 9376
rect 5081 9000 5093 9376
rect 6531 9376 6589 9388
rect 6531 9188 6543 9376
rect 5035 8988 5093 9000
rect 5154 9176 5212 9188
rect 5154 9000 5166 9176
rect 5200 9000 5212 9176
rect 5154 8988 5212 9000
rect 5272 9176 5330 9188
rect 5272 9000 5284 9176
rect 5318 9000 5330 9176
rect 5272 8988 5330 9000
rect 5390 9176 5448 9188
rect 5390 9000 5402 9176
rect 5436 9000 5448 9176
rect 5390 8988 5448 9000
rect 5508 9176 5566 9188
rect 5508 9000 5520 9176
rect 5554 9000 5566 9176
rect 5508 8988 5566 9000
rect 6090 9176 6148 9188
rect 6090 9000 6102 9176
rect 6136 9000 6148 9176
rect 6090 8988 6148 9000
rect 6208 9176 6266 9188
rect 6208 9000 6220 9176
rect 6254 9000 6266 9176
rect 6208 8988 6266 9000
rect 6326 9176 6384 9188
rect 6326 9000 6338 9176
rect 6372 9000 6384 9176
rect 6326 8988 6384 9000
rect 6444 9176 6543 9188
rect 6444 9000 6456 9176
rect 6490 9000 6543 9176
rect 6577 9000 6589 9376
rect 6444 8988 6589 9000
rect 6649 9376 6707 9388
rect 6649 9000 6661 9376
rect 6695 9000 6707 9376
rect 6649 8988 6707 9000
rect 6767 9376 6825 9388
rect 6767 9000 6779 9376
rect 6813 9000 6825 9376
rect 6767 8988 6825 9000
rect 6885 9376 6943 9388
rect 6885 9000 6897 9376
rect 6931 9000 6943 9376
rect 6885 8988 6943 9000
rect 6998 9376 7056 9388
rect 6998 9000 7010 9376
rect 7044 9000 7056 9376
rect 6998 8988 7056 9000
rect 7116 9376 7174 9388
rect 7116 9000 7128 9376
rect 7162 9000 7174 9376
rect 7116 8988 7174 9000
rect 7234 9376 7292 9388
rect 7234 9000 7246 9376
rect 7280 9000 7292 9376
rect 7234 8988 7292 9000
rect 7352 9376 7410 9388
rect 7352 9000 7364 9376
rect 7398 9000 7410 9376
rect 7352 8988 7410 9000
rect 7470 9376 7528 9388
rect 7470 9000 7482 9376
rect 7516 9000 7528 9376
rect 7470 8988 7528 9000
rect 7588 9376 7646 9388
rect 7588 9000 7600 9376
rect 7634 9000 7646 9376
rect 7588 8988 7646 9000
rect 7706 9376 7764 9388
rect 7706 9000 7718 9376
rect 7752 9000 7764 9376
rect 7706 8988 7764 9000
rect 7825 9376 7883 9388
rect 7825 9000 7837 9376
rect 7871 9000 7883 9376
rect 7825 8988 7883 9000
rect 7943 9376 8001 9388
rect 7943 9000 7955 9376
rect 7989 9000 8001 9376
rect 7943 8988 8001 9000
rect 8061 9376 8119 9388
rect 8061 9000 8073 9376
rect 8107 9000 8119 9376
rect 8061 8988 8119 9000
rect 8179 9376 8237 9388
rect 8179 9000 8191 9376
rect 8225 9000 8237 9376
rect 9663 9380 9721 9392
rect 9663 9192 9675 9380
rect 8179 8988 8237 9000
rect 8298 9176 8356 9188
rect 8298 9000 8310 9176
rect 8344 9000 8356 9176
rect 8298 8988 8356 9000
rect 8416 9176 8474 9188
rect 8416 9000 8428 9176
rect 8462 9000 8474 9176
rect 8416 8988 8474 9000
rect 8534 9176 8592 9188
rect 8534 9000 8546 9176
rect 8580 9000 8592 9176
rect 8534 8988 8592 9000
rect 8652 9176 8710 9188
rect 8652 9000 8664 9176
rect 8698 9000 8710 9176
rect 8652 8988 8710 9000
rect 9222 9180 9280 9192
rect 9222 9004 9234 9180
rect 9268 9004 9280 9180
rect 9222 8992 9280 9004
rect 9340 9180 9398 9192
rect 9340 9004 9352 9180
rect 9386 9004 9398 9180
rect 9340 8992 9398 9004
rect 9458 9180 9516 9192
rect 9458 9004 9470 9180
rect 9504 9004 9516 9180
rect 9458 8992 9516 9004
rect 9576 9180 9675 9192
rect 9576 9004 9588 9180
rect 9622 9004 9675 9180
rect 9709 9004 9721 9380
rect 9576 8992 9721 9004
rect 9781 9380 9839 9392
rect 9781 9004 9793 9380
rect 9827 9004 9839 9380
rect 9781 8992 9839 9004
rect 9899 9380 9957 9392
rect 9899 9004 9911 9380
rect 9945 9004 9957 9380
rect 9899 8992 9957 9004
rect 10017 9380 10075 9392
rect 10017 9004 10029 9380
rect 10063 9004 10075 9380
rect 10017 8992 10075 9004
rect 10130 9380 10188 9392
rect 10130 9004 10142 9380
rect 10176 9004 10188 9380
rect 10130 8992 10188 9004
rect 10248 9380 10306 9392
rect 10248 9004 10260 9380
rect 10294 9004 10306 9380
rect 10248 8992 10306 9004
rect 10366 9380 10424 9392
rect 10366 9004 10378 9380
rect 10412 9004 10424 9380
rect 10366 8992 10424 9004
rect 10484 9380 10542 9392
rect 10484 9004 10496 9380
rect 10530 9004 10542 9380
rect 10484 8992 10542 9004
rect 10602 9380 10660 9392
rect 10602 9004 10614 9380
rect 10648 9004 10660 9380
rect 10602 8992 10660 9004
rect 10720 9380 10778 9392
rect 10720 9004 10732 9380
rect 10766 9004 10778 9380
rect 10720 8992 10778 9004
rect 10838 9380 10896 9392
rect 10838 9004 10850 9380
rect 10884 9004 10896 9380
rect 10838 8992 10896 9004
rect 10957 9380 11015 9392
rect 10957 9004 10969 9380
rect 11003 9004 11015 9380
rect 10957 8992 11015 9004
rect 11075 9380 11133 9392
rect 11075 9004 11087 9380
rect 11121 9004 11133 9380
rect 11075 8992 11133 9004
rect 11193 9380 11251 9392
rect 11193 9004 11205 9380
rect 11239 9004 11251 9380
rect 11193 8992 11251 9004
rect 11311 9380 11369 9392
rect 11311 9004 11323 9380
rect 11357 9004 11369 9380
rect 12807 9380 12865 9392
rect 12807 9192 12819 9380
rect 11311 8992 11369 9004
rect 11430 9180 11488 9192
rect 11430 9004 11442 9180
rect 11476 9004 11488 9180
rect 11430 8992 11488 9004
rect 11548 9180 11606 9192
rect 11548 9004 11560 9180
rect 11594 9004 11606 9180
rect 11548 8992 11606 9004
rect 11666 9180 11724 9192
rect 11666 9004 11678 9180
rect 11712 9004 11724 9180
rect 11666 8992 11724 9004
rect 11784 9180 11842 9192
rect 11784 9004 11796 9180
rect 11830 9004 11842 9180
rect 11784 8992 11842 9004
rect 12366 9180 12424 9192
rect 12366 9004 12378 9180
rect 12412 9004 12424 9180
rect 12366 8992 12424 9004
rect 12484 9180 12542 9192
rect 12484 9004 12496 9180
rect 12530 9004 12542 9180
rect 12484 8992 12542 9004
rect 12602 9180 12660 9192
rect 12602 9004 12614 9180
rect 12648 9004 12660 9180
rect 12602 8992 12660 9004
rect 12720 9180 12819 9192
rect 12720 9004 12732 9180
rect 12766 9004 12819 9180
rect 12853 9004 12865 9380
rect 12720 8992 12865 9004
rect 12925 9380 12983 9392
rect 12925 9004 12937 9380
rect 12971 9004 12983 9380
rect 12925 8992 12983 9004
rect 13043 9380 13101 9392
rect 13043 9004 13055 9380
rect 13089 9004 13101 9380
rect 13043 8992 13101 9004
rect 13161 9380 13219 9392
rect 13161 9004 13173 9380
rect 13207 9004 13219 9380
rect 13161 8992 13219 9004
rect 13274 9380 13332 9392
rect 13274 9004 13286 9380
rect 13320 9004 13332 9380
rect 13274 8992 13332 9004
rect 13392 9380 13450 9392
rect 13392 9004 13404 9380
rect 13438 9004 13450 9380
rect 13392 8992 13450 9004
rect 13510 9380 13568 9392
rect 13510 9004 13522 9380
rect 13556 9004 13568 9380
rect 13510 8992 13568 9004
rect 13628 9380 13686 9392
rect 13628 9004 13640 9380
rect 13674 9004 13686 9380
rect 13628 8992 13686 9004
rect 13746 9380 13804 9392
rect 13746 9004 13758 9380
rect 13792 9004 13804 9380
rect 13746 8992 13804 9004
rect 13864 9380 13922 9392
rect 13864 9004 13876 9380
rect 13910 9004 13922 9380
rect 13864 8992 13922 9004
rect 13982 9380 14040 9392
rect 13982 9004 13994 9380
rect 14028 9004 14040 9380
rect 13982 8992 14040 9004
rect 14101 9380 14159 9392
rect 14101 9004 14113 9380
rect 14147 9004 14159 9380
rect 14101 8992 14159 9004
rect 14219 9380 14277 9392
rect 14219 9004 14231 9380
rect 14265 9004 14277 9380
rect 14219 8992 14277 9004
rect 14337 9380 14395 9392
rect 14337 9004 14349 9380
rect 14383 9004 14395 9380
rect 14337 8992 14395 9004
rect 14455 9380 14513 9392
rect 14455 9004 14467 9380
rect 14501 9004 14513 9380
rect 16009 9376 16067 9388
rect 14455 8992 14513 9004
rect 14574 9180 14632 9192
rect 14574 9004 14586 9180
rect 14620 9004 14632 9180
rect 14574 8992 14632 9004
rect 14692 9180 14750 9192
rect 14692 9004 14704 9180
rect 14738 9004 14750 9180
rect 14692 8992 14750 9004
rect 14810 9180 14868 9192
rect 14810 9004 14822 9180
rect 14856 9004 14868 9180
rect 14810 8992 14868 9004
rect 14928 9180 14986 9192
rect 16009 9188 16021 9376
rect 14928 9004 14940 9180
rect 14974 9004 14986 9180
rect 14928 8992 14986 9004
rect 15568 9176 15626 9188
rect 15568 9000 15580 9176
rect 15614 9000 15626 9176
rect 15568 8988 15626 9000
rect 15686 9176 15744 9188
rect 15686 9000 15698 9176
rect 15732 9000 15744 9176
rect 15686 8988 15744 9000
rect 15804 9176 15862 9188
rect 15804 9000 15816 9176
rect 15850 9000 15862 9176
rect 15804 8988 15862 9000
rect 15922 9176 16021 9188
rect 15922 9000 15934 9176
rect 15968 9000 16021 9176
rect 16055 9000 16067 9376
rect 15922 8988 16067 9000
rect 16127 9376 16185 9388
rect 16127 9000 16139 9376
rect 16173 9000 16185 9376
rect 16127 8988 16185 9000
rect 16245 9376 16303 9388
rect 16245 9000 16257 9376
rect 16291 9000 16303 9376
rect 16245 8988 16303 9000
rect 16363 9376 16421 9388
rect 16363 9000 16375 9376
rect 16409 9000 16421 9376
rect 16363 8988 16421 9000
rect 16476 9376 16534 9388
rect 16476 9000 16488 9376
rect 16522 9000 16534 9376
rect 16476 8988 16534 9000
rect 16594 9376 16652 9388
rect 16594 9000 16606 9376
rect 16640 9000 16652 9376
rect 16594 8988 16652 9000
rect 16712 9376 16770 9388
rect 16712 9000 16724 9376
rect 16758 9000 16770 9376
rect 16712 8988 16770 9000
rect 16830 9376 16888 9388
rect 16830 9000 16842 9376
rect 16876 9000 16888 9376
rect 16830 8988 16888 9000
rect 16948 9376 17006 9388
rect 16948 9000 16960 9376
rect 16994 9000 17006 9376
rect 16948 8988 17006 9000
rect 17066 9376 17124 9388
rect 17066 9000 17078 9376
rect 17112 9000 17124 9376
rect 17066 8988 17124 9000
rect 17184 9376 17242 9388
rect 17184 9000 17196 9376
rect 17230 9000 17242 9376
rect 17184 8988 17242 9000
rect 17303 9376 17361 9388
rect 17303 9000 17315 9376
rect 17349 9000 17361 9376
rect 17303 8988 17361 9000
rect 17421 9376 17479 9388
rect 17421 9000 17433 9376
rect 17467 9000 17479 9376
rect 17421 8988 17479 9000
rect 17539 9376 17597 9388
rect 17539 9000 17551 9376
rect 17585 9000 17597 9376
rect 17539 8988 17597 9000
rect 17657 9376 17715 9388
rect 17657 9000 17669 9376
rect 17703 9000 17715 9376
rect 19153 9376 19211 9388
rect 19153 9188 19165 9376
rect 17657 8988 17715 9000
rect 17776 9176 17834 9188
rect 17776 9000 17788 9176
rect 17822 9000 17834 9176
rect 17776 8988 17834 9000
rect 17894 9176 17952 9188
rect 17894 9000 17906 9176
rect 17940 9000 17952 9176
rect 17894 8988 17952 9000
rect 18012 9176 18070 9188
rect 18012 9000 18024 9176
rect 18058 9000 18070 9176
rect 18012 8988 18070 9000
rect 18130 9176 18188 9188
rect 18130 9000 18142 9176
rect 18176 9000 18188 9176
rect 18130 8988 18188 9000
rect 18712 9176 18770 9188
rect 18712 9000 18724 9176
rect 18758 9000 18770 9176
rect 18712 8988 18770 9000
rect 18830 9176 18888 9188
rect 18830 9000 18842 9176
rect 18876 9000 18888 9176
rect 18830 8988 18888 9000
rect 18948 9176 19006 9188
rect 18948 9000 18960 9176
rect 18994 9000 19006 9176
rect 18948 8988 19006 9000
rect 19066 9176 19165 9188
rect 19066 9000 19078 9176
rect 19112 9000 19165 9176
rect 19199 9000 19211 9376
rect 19066 8988 19211 9000
rect 19271 9376 19329 9388
rect 19271 9000 19283 9376
rect 19317 9000 19329 9376
rect 19271 8988 19329 9000
rect 19389 9376 19447 9388
rect 19389 9000 19401 9376
rect 19435 9000 19447 9376
rect 19389 8988 19447 9000
rect 19507 9376 19565 9388
rect 19507 9000 19519 9376
rect 19553 9000 19565 9376
rect 19507 8988 19565 9000
rect 19620 9376 19678 9388
rect 19620 9000 19632 9376
rect 19666 9000 19678 9376
rect 19620 8988 19678 9000
rect 19738 9376 19796 9388
rect 19738 9000 19750 9376
rect 19784 9000 19796 9376
rect 19738 8988 19796 9000
rect 19856 9376 19914 9388
rect 19856 9000 19868 9376
rect 19902 9000 19914 9376
rect 19856 8988 19914 9000
rect 19974 9376 20032 9388
rect 19974 9000 19986 9376
rect 20020 9000 20032 9376
rect 19974 8988 20032 9000
rect 20092 9376 20150 9388
rect 20092 9000 20104 9376
rect 20138 9000 20150 9376
rect 20092 8988 20150 9000
rect 20210 9376 20268 9388
rect 20210 9000 20222 9376
rect 20256 9000 20268 9376
rect 20210 8988 20268 9000
rect 20328 9376 20386 9388
rect 20328 9000 20340 9376
rect 20374 9000 20386 9376
rect 20328 8988 20386 9000
rect 20447 9376 20505 9388
rect 20447 9000 20459 9376
rect 20493 9000 20505 9376
rect 20447 8988 20505 9000
rect 20565 9376 20623 9388
rect 20565 9000 20577 9376
rect 20611 9000 20623 9376
rect 20565 8988 20623 9000
rect 20683 9376 20741 9388
rect 20683 9000 20695 9376
rect 20729 9000 20741 9376
rect 20683 8988 20741 9000
rect 20801 9376 20859 9388
rect 20801 9000 20813 9376
rect 20847 9000 20859 9376
rect 22285 9380 22343 9392
rect 22285 9192 22297 9380
rect 20801 8988 20859 9000
rect 20920 9176 20978 9188
rect 20920 9000 20932 9176
rect 20966 9000 20978 9176
rect 20920 8988 20978 9000
rect 21038 9176 21096 9188
rect 21038 9000 21050 9176
rect 21084 9000 21096 9176
rect 21038 8988 21096 9000
rect 21156 9176 21214 9188
rect 21156 9000 21168 9176
rect 21202 9000 21214 9176
rect 21156 8988 21214 9000
rect 21274 9176 21332 9188
rect 21274 9000 21286 9176
rect 21320 9000 21332 9176
rect 21274 8988 21332 9000
rect 21844 9180 21902 9192
rect 21844 9004 21856 9180
rect 21890 9004 21902 9180
rect 21844 8992 21902 9004
rect 21962 9180 22020 9192
rect 21962 9004 21974 9180
rect 22008 9004 22020 9180
rect 21962 8992 22020 9004
rect 22080 9180 22138 9192
rect 22080 9004 22092 9180
rect 22126 9004 22138 9180
rect 22080 8992 22138 9004
rect 22198 9180 22297 9192
rect 22198 9004 22210 9180
rect 22244 9004 22297 9180
rect 22331 9004 22343 9380
rect 22198 8992 22343 9004
rect 22403 9380 22461 9392
rect 22403 9004 22415 9380
rect 22449 9004 22461 9380
rect 22403 8992 22461 9004
rect 22521 9380 22579 9392
rect 22521 9004 22533 9380
rect 22567 9004 22579 9380
rect 22521 8992 22579 9004
rect 22639 9380 22697 9392
rect 22639 9004 22651 9380
rect 22685 9004 22697 9380
rect 22639 8992 22697 9004
rect 22752 9380 22810 9392
rect 22752 9004 22764 9380
rect 22798 9004 22810 9380
rect 22752 8992 22810 9004
rect 22870 9380 22928 9392
rect 22870 9004 22882 9380
rect 22916 9004 22928 9380
rect 22870 8992 22928 9004
rect 22988 9380 23046 9392
rect 22988 9004 23000 9380
rect 23034 9004 23046 9380
rect 22988 8992 23046 9004
rect 23106 9380 23164 9392
rect 23106 9004 23118 9380
rect 23152 9004 23164 9380
rect 23106 8992 23164 9004
rect 23224 9380 23282 9392
rect 23224 9004 23236 9380
rect 23270 9004 23282 9380
rect 23224 8992 23282 9004
rect 23342 9380 23400 9392
rect 23342 9004 23354 9380
rect 23388 9004 23400 9380
rect 23342 8992 23400 9004
rect 23460 9380 23518 9392
rect 23460 9004 23472 9380
rect 23506 9004 23518 9380
rect 23460 8992 23518 9004
rect 23579 9380 23637 9392
rect 23579 9004 23591 9380
rect 23625 9004 23637 9380
rect 23579 8992 23637 9004
rect 23697 9380 23755 9392
rect 23697 9004 23709 9380
rect 23743 9004 23755 9380
rect 23697 8992 23755 9004
rect 23815 9380 23873 9392
rect 23815 9004 23827 9380
rect 23861 9004 23873 9380
rect 23815 8992 23873 9004
rect 23933 9380 23991 9392
rect 23933 9004 23945 9380
rect 23979 9004 23991 9380
rect 25429 9380 25487 9392
rect 25429 9192 25441 9380
rect 23933 8992 23991 9004
rect 24052 9180 24110 9192
rect 24052 9004 24064 9180
rect 24098 9004 24110 9180
rect 24052 8992 24110 9004
rect 24170 9180 24228 9192
rect 24170 9004 24182 9180
rect 24216 9004 24228 9180
rect 24170 8992 24228 9004
rect 24288 9180 24346 9192
rect 24288 9004 24300 9180
rect 24334 9004 24346 9180
rect 24288 8992 24346 9004
rect 24406 9180 24464 9192
rect 24406 9004 24418 9180
rect 24452 9004 24464 9180
rect 24406 8992 24464 9004
rect 24988 9180 25046 9192
rect 24988 9004 25000 9180
rect 25034 9004 25046 9180
rect 24988 8992 25046 9004
rect 25106 9180 25164 9192
rect 25106 9004 25118 9180
rect 25152 9004 25164 9180
rect 25106 8992 25164 9004
rect 25224 9180 25282 9192
rect 25224 9004 25236 9180
rect 25270 9004 25282 9180
rect 25224 8992 25282 9004
rect 25342 9180 25441 9192
rect 25342 9004 25354 9180
rect 25388 9004 25441 9180
rect 25475 9004 25487 9380
rect 25342 8992 25487 9004
rect 25547 9380 25605 9392
rect 25547 9004 25559 9380
rect 25593 9004 25605 9380
rect 25547 8992 25605 9004
rect 25665 9380 25723 9392
rect 25665 9004 25677 9380
rect 25711 9004 25723 9380
rect 25665 8992 25723 9004
rect 25783 9380 25841 9392
rect 25783 9004 25795 9380
rect 25829 9004 25841 9380
rect 25783 8992 25841 9004
rect 25896 9380 25954 9392
rect 25896 9004 25908 9380
rect 25942 9004 25954 9380
rect 25896 8992 25954 9004
rect 26014 9380 26072 9392
rect 26014 9004 26026 9380
rect 26060 9004 26072 9380
rect 26014 8992 26072 9004
rect 26132 9380 26190 9392
rect 26132 9004 26144 9380
rect 26178 9004 26190 9380
rect 26132 8992 26190 9004
rect 26250 9380 26308 9392
rect 26250 9004 26262 9380
rect 26296 9004 26308 9380
rect 26250 8992 26308 9004
rect 26368 9380 26426 9392
rect 26368 9004 26380 9380
rect 26414 9004 26426 9380
rect 26368 8992 26426 9004
rect 26486 9380 26544 9392
rect 26486 9004 26498 9380
rect 26532 9004 26544 9380
rect 26486 8992 26544 9004
rect 26604 9380 26662 9392
rect 26604 9004 26616 9380
rect 26650 9004 26662 9380
rect 26604 8992 26662 9004
rect 26723 9380 26781 9392
rect 26723 9004 26735 9380
rect 26769 9004 26781 9380
rect 26723 8992 26781 9004
rect 26841 9380 26899 9392
rect 26841 9004 26853 9380
rect 26887 9004 26899 9380
rect 26841 8992 26899 9004
rect 26959 9380 27017 9392
rect 26959 9004 26971 9380
rect 27005 9004 27017 9380
rect 26959 8992 27017 9004
rect 27077 9380 27135 9392
rect 27077 9004 27089 9380
rect 27123 9004 27135 9380
rect 27077 8992 27135 9004
rect 27196 9180 27254 9192
rect 27196 9004 27208 9180
rect 27242 9004 27254 9180
rect 27196 8992 27254 9004
rect 27314 9180 27372 9192
rect 27314 9004 27326 9180
rect 27360 9004 27372 9180
rect 27314 8992 27372 9004
rect 27432 9180 27490 9192
rect 27432 9004 27444 9180
rect 27478 9004 27490 9180
rect 27432 8992 27490 9004
rect 27550 9180 27608 9192
rect 27550 9004 27562 9180
rect 27596 9004 27608 9180
rect 27550 8992 27608 9004
rect 19415 6547 19473 6559
rect 3167 6431 3225 6443
rect 2683 6231 2741 6243
rect 2683 6055 2695 6231
rect 2729 6055 2741 6231
rect 2683 6043 2741 6055
rect 2801 6231 2859 6243
rect 2801 6055 2813 6231
rect 2847 6055 2859 6231
rect 2801 6043 2859 6055
rect 2919 6231 2977 6243
rect 2919 6055 2931 6231
rect 2965 6055 2977 6231
rect 2919 6043 2977 6055
rect 3037 6231 3095 6243
rect 3037 6055 3049 6231
rect 3083 6055 3095 6231
rect 3037 6043 3095 6055
rect 3167 6055 3179 6431
rect 3213 6055 3225 6431
rect 3167 6043 3225 6055
rect 3285 6431 3343 6443
rect 3285 6055 3297 6431
rect 3331 6055 3343 6431
rect 3285 6043 3343 6055
rect 3403 6431 3461 6443
rect 3403 6055 3415 6431
rect 3449 6055 3461 6431
rect 3403 6043 3461 6055
rect 3521 6431 3579 6443
rect 3521 6055 3533 6431
rect 3567 6055 3579 6431
rect 3521 6043 3579 6055
rect 3639 6431 3697 6443
rect 3639 6055 3651 6431
rect 3685 6055 3697 6431
rect 3639 6043 3697 6055
rect 3757 6431 3815 6443
rect 3757 6055 3769 6431
rect 3803 6055 3815 6431
rect 3757 6043 3815 6055
rect 3875 6431 3933 6443
rect 3875 6055 3887 6431
rect 3921 6055 3933 6431
rect 5235 6433 5293 6445
rect 3875 6043 3933 6055
rect 4004 6231 4062 6243
rect 4004 6055 4016 6231
rect 4050 6055 4062 6231
rect 4004 6043 4062 6055
rect 4122 6231 4180 6243
rect 4122 6055 4134 6231
rect 4168 6055 4180 6231
rect 4122 6043 4180 6055
rect 4240 6231 4298 6243
rect 4240 6055 4252 6231
rect 4286 6055 4298 6231
rect 4240 6043 4298 6055
rect 4358 6231 4416 6243
rect 4358 6055 4370 6231
rect 4404 6055 4416 6231
rect 4358 6043 4416 6055
rect 4751 6233 4809 6245
rect 4751 6057 4763 6233
rect 4797 6057 4809 6233
rect 4751 6045 4809 6057
rect 4869 6233 4927 6245
rect 4869 6057 4881 6233
rect 4915 6057 4927 6233
rect 4869 6045 4927 6057
rect 4987 6233 5045 6245
rect 4987 6057 4999 6233
rect 5033 6057 5045 6233
rect 4987 6045 5045 6057
rect 5105 6233 5163 6245
rect 5105 6057 5117 6233
rect 5151 6057 5163 6233
rect 5105 6045 5163 6057
rect 5235 6057 5247 6433
rect 5281 6057 5293 6433
rect 5235 6045 5293 6057
rect 5353 6433 5411 6445
rect 5353 6057 5365 6433
rect 5399 6057 5411 6433
rect 5353 6045 5411 6057
rect 5471 6433 5529 6445
rect 5471 6057 5483 6433
rect 5517 6057 5529 6433
rect 5471 6045 5529 6057
rect 5589 6433 5647 6445
rect 5589 6057 5601 6433
rect 5635 6057 5647 6433
rect 5589 6045 5647 6057
rect 5707 6433 5765 6445
rect 5707 6057 5719 6433
rect 5753 6057 5765 6433
rect 5707 6045 5765 6057
rect 5825 6433 5883 6445
rect 5825 6057 5837 6433
rect 5871 6057 5883 6433
rect 5825 6045 5883 6057
rect 5943 6433 6001 6445
rect 5943 6057 5955 6433
rect 5989 6057 6001 6433
rect 7304 6431 7362 6443
rect 5943 6045 6001 6057
rect 6072 6233 6130 6245
rect 6072 6057 6084 6233
rect 6118 6057 6130 6233
rect 6072 6045 6130 6057
rect 6190 6233 6248 6245
rect 6190 6057 6202 6233
rect 6236 6057 6248 6233
rect 6190 6045 6248 6057
rect 6308 6233 6366 6245
rect 6308 6057 6320 6233
rect 6354 6057 6366 6233
rect 6308 6045 6366 6057
rect 6426 6233 6484 6245
rect 6426 6057 6438 6233
rect 6472 6057 6484 6233
rect 6426 6045 6484 6057
rect 6820 6231 6878 6243
rect 6820 6055 6832 6231
rect 6866 6055 6878 6231
rect 3110 5738 3168 5750
rect 3110 5362 3122 5738
rect 3156 5362 3168 5738
rect 3110 5350 3168 5362
rect 3228 5738 3286 5750
rect 3228 5362 3240 5738
rect 3274 5362 3286 5738
rect 3228 5350 3286 5362
rect 3346 5738 3404 5750
rect 3346 5362 3358 5738
rect 3392 5362 3404 5738
rect 3346 5350 3404 5362
rect 3464 5738 3522 5750
rect 3464 5362 3476 5738
rect 3510 5362 3522 5738
rect 3464 5350 3522 5362
rect 3582 5738 3640 5750
rect 3582 5362 3594 5738
rect 3628 5362 3640 5738
rect 3582 5350 3640 5362
rect 3700 5738 3758 5750
rect 3700 5362 3712 5738
rect 3746 5362 3758 5738
rect 3700 5350 3758 5362
rect 3818 5738 3876 5750
rect 3818 5362 3830 5738
rect 3864 5362 3876 5738
rect 3818 5350 3876 5362
rect 6820 6043 6878 6055
rect 6938 6231 6996 6243
rect 6938 6055 6950 6231
rect 6984 6055 6996 6231
rect 6938 6043 6996 6055
rect 7056 6231 7114 6243
rect 7056 6055 7068 6231
rect 7102 6055 7114 6231
rect 7056 6043 7114 6055
rect 7174 6231 7232 6243
rect 7174 6055 7186 6231
rect 7220 6055 7232 6231
rect 7174 6043 7232 6055
rect 7304 6055 7316 6431
rect 7350 6055 7362 6431
rect 7304 6043 7362 6055
rect 7422 6431 7480 6443
rect 7422 6055 7434 6431
rect 7468 6055 7480 6431
rect 7422 6043 7480 6055
rect 7540 6431 7598 6443
rect 7540 6055 7552 6431
rect 7586 6055 7598 6431
rect 7540 6043 7598 6055
rect 7658 6431 7716 6443
rect 7658 6055 7670 6431
rect 7704 6055 7716 6431
rect 7658 6043 7716 6055
rect 7776 6431 7834 6443
rect 7776 6055 7788 6431
rect 7822 6055 7834 6431
rect 7776 6043 7834 6055
rect 7894 6431 7952 6443
rect 7894 6055 7906 6431
rect 7940 6055 7952 6431
rect 7894 6043 7952 6055
rect 8012 6431 8070 6443
rect 8012 6055 8024 6431
rect 8058 6055 8070 6431
rect 9372 6433 9430 6445
rect 8012 6043 8070 6055
rect 8141 6231 8199 6243
rect 8141 6055 8153 6231
rect 8187 6055 8199 6231
rect 8141 6043 8199 6055
rect 8259 6231 8317 6243
rect 8259 6055 8271 6231
rect 8305 6055 8317 6231
rect 8259 6043 8317 6055
rect 8377 6231 8435 6243
rect 8377 6055 8389 6231
rect 8423 6055 8435 6231
rect 8377 6043 8435 6055
rect 8495 6231 8553 6243
rect 8495 6055 8507 6231
rect 8541 6055 8553 6231
rect 8495 6043 8553 6055
rect 8888 6233 8946 6245
rect 8888 6057 8900 6233
rect 8934 6057 8946 6233
rect 8888 6045 8946 6057
rect 9006 6233 9064 6245
rect 9006 6057 9018 6233
rect 9052 6057 9064 6233
rect 9006 6045 9064 6057
rect 9124 6233 9182 6245
rect 9124 6057 9136 6233
rect 9170 6057 9182 6233
rect 9124 6045 9182 6057
rect 9242 6233 9300 6245
rect 9242 6057 9254 6233
rect 9288 6057 9300 6233
rect 9242 6045 9300 6057
rect 9372 6057 9384 6433
rect 9418 6057 9430 6433
rect 9372 6045 9430 6057
rect 9490 6433 9548 6445
rect 9490 6057 9502 6433
rect 9536 6057 9548 6433
rect 9490 6045 9548 6057
rect 9608 6433 9666 6445
rect 9608 6057 9620 6433
rect 9654 6057 9666 6433
rect 9608 6045 9666 6057
rect 9726 6433 9784 6445
rect 9726 6057 9738 6433
rect 9772 6057 9784 6433
rect 9726 6045 9784 6057
rect 9844 6433 9902 6445
rect 9844 6057 9856 6433
rect 9890 6057 9902 6433
rect 9844 6045 9902 6057
rect 9962 6433 10020 6445
rect 9962 6057 9974 6433
rect 10008 6057 10020 6433
rect 9962 6045 10020 6057
rect 10080 6433 10138 6445
rect 10080 6057 10092 6433
rect 10126 6057 10138 6433
rect 11441 6433 11499 6445
rect 10080 6045 10138 6057
rect 10209 6233 10267 6245
rect 10209 6057 10221 6233
rect 10255 6057 10267 6233
rect 10209 6045 10267 6057
rect 10327 6233 10385 6245
rect 10327 6057 10339 6233
rect 10373 6057 10385 6233
rect 10327 6045 10385 6057
rect 10445 6233 10503 6245
rect 10445 6057 10457 6233
rect 10491 6057 10503 6233
rect 10445 6045 10503 6057
rect 10563 6233 10621 6245
rect 10563 6057 10575 6233
rect 10609 6057 10621 6233
rect 10563 6045 10621 6057
rect 10957 6233 11015 6245
rect 10957 6057 10969 6233
rect 11003 6057 11015 6233
rect 10957 6045 11015 6057
rect 11075 6233 11133 6245
rect 11075 6057 11087 6233
rect 11121 6057 11133 6233
rect 11075 6045 11133 6057
rect 11193 6233 11251 6245
rect 11193 6057 11205 6233
rect 11239 6057 11251 6233
rect 11193 6045 11251 6057
rect 11311 6233 11369 6245
rect 11311 6057 11323 6233
rect 11357 6057 11369 6233
rect 11311 6045 11369 6057
rect 11441 6057 11453 6433
rect 11487 6057 11499 6433
rect 11441 6045 11499 6057
rect 11559 6433 11617 6445
rect 11559 6057 11571 6433
rect 11605 6057 11617 6433
rect 11559 6045 11617 6057
rect 11677 6433 11735 6445
rect 11677 6057 11689 6433
rect 11723 6057 11735 6433
rect 11677 6045 11735 6057
rect 11795 6433 11853 6445
rect 11795 6057 11807 6433
rect 11841 6057 11853 6433
rect 11795 6045 11853 6057
rect 11913 6433 11971 6445
rect 11913 6057 11925 6433
rect 11959 6057 11971 6433
rect 11913 6045 11971 6057
rect 12031 6433 12089 6445
rect 12031 6057 12043 6433
rect 12077 6057 12089 6433
rect 12031 6045 12089 6057
rect 12149 6433 12207 6445
rect 12149 6057 12161 6433
rect 12195 6057 12207 6433
rect 13509 6435 13567 6447
rect 12149 6045 12207 6057
rect 12278 6233 12336 6245
rect 12278 6057 12290 6233
rect 12324 6057 12336 6233
rect 12278 6045 12336 6057
rect 12396 6233 12454 6245
rect 12396 6057 12408 6233
rect 12442 6057 12454 6233
rect 12396 6045 12454 6057
rect 12514 6233 12572 6245
rect 12514 6057 12526 6233
rect 12560 6057 12572 6233
rect 12514 6045 12572 6057
rect 12632 6233 12690 6245
rect 12632 6057 12644 6233
rect 12678 6057 12690 6233
rect 12632 6045 12690 6057
rect 13025 6235 13083 6247
rect 13025 6059 13037 6235
rect 13071 6059 13083 6235
rect 13025 6047 13083 6059
rect 13143 6235 13201 6247
rect 13143 6059 13155 6235
rect 13189 6059 13201 6235
rect 13143 6047 13201 6059
rect 13261 6235 13319 6247
rect 13261 6059 13273 6235
rect 13307 6059 13319 6235
rect 13261 6047 13319 6059
rect 13379 6235 13437 6247
rect 13379 6059 13391 6235
rect 13425 6059 13437 6235
rect 13379 6047 13437 6059
rect 13509 6059 13521 6435
rect 13555 6059 13567 6435
rect 13509 6047 13567 6059
rect 13627 6435 13685 6447
rect 13627 6059 13639 6435
rect 13673 6059 13685 6435
rect 13627 6047 13685 6059
rect 13745 6435 13803 6447
rect 13745 6059 13757 6435
rect 13791 6059 13803 6435
rect 13745 6047 13803 6059
rect 13863 6435 13921 6447
rect 13863 6059 13875 6435
rect 13909 6059 13921 6435
rect 13863 6047 13921 6059
rect 13981 6435 14039 6447
rect 13981 6059 13993 6435
rect 14027 6059 14039 6435
rect 13981 6047 14039 6059
rect 14099 6435 14157 6447
rect 14099 6059 14111 6435
rect 14145 6059 14157 6435
rect 14099 6047 14157 6059
rect 14217 6435 14275 6447
rect 14217 6059 14229 6435
rect 14263 6059 14275 6435
rect 15578 6433 15636 6445
rect 14217 6047 14275 6059
rect 14346 6235 14404 6247
rect 14346 6059 14358 6235
rect 14392 6059 14404 6235
rect 14346 6047 14404 6059
rect 14464 6235 14522 6247
rect 14464 6059 14476 6235
rect 14510 6059 14522 6235
rect 14464 6047 14522 6059
rect 14582 6235 14640 6247
rect 14582 6059 14594 6235
rect 14628 6059 14640 6235
rect 14582 6047 14640 6059
rect 14700 6235 14758 6247
rect 14700 6059 14712 6235
rect 14746 6059 14758 6235
rect 14700 6047 14758 6059
rect 15094 6233 15152 6245
rect 15094 6057 15106 6233
rect 15140 6057 15152 6233
rect 5178 5740 5236 5752
rect 5178 5364 5190 5740
rect 5224 5364 5236 5740
rect 5178 5352 5236 5364
rect 5296 5740 5354 5752
rect 5296 5364 5308 5740
rect 5342 5364 5354 5740
rect 5296 5352 5354 5364
rect 5414 5740 5472 5752
rect 5414 5364 5426 5740
rect 5460 5364 5472 5740
rect 5414 5352 5472 5364
rect 5532 5740 5590 5752
rect 5532 5364 5544 5740
rect 5578 5364 5590 5740
rect 5532 5352 5590 5364
rect 5650 5740 5708 5752
rect 5650 5364 5662 5740
rect 5696 5364 5708 5740
rect 5650 5352 5708 5364
rect 5768 5740 5826 5752
rect 5768 5364 5780 5740
rect 5814 5364 5826 5740
rect 5768 5352 5826 5364
rect 5886 5740 5944 5752
rect 5886 5364 5898 5740
rect 5932 5364 5944 5740
rect 5886 5352 5944 5364
rect 7247 5738 7305 5750
rect 7247 5362 7259 5738
rect 7293 5362 7305 5738
rect 7247 5350 7305 5362
rect 7365 5738 7423 5750
rect 7365 5362 7377 5738
rect 7411 5362 7423 5738
rect 7365 5350 7423 5362
rect 7483 5738 7541 5750
rect 7483 5362 7495 5738
rect 7529 5362 7541 5738
rect 7483 5350 7541 5362
rect 7601 5738 7659 5750
rect 7601 5362 7613 5738
rect 7647 5362 7659 5738
rect 7601 5350 7659 5362
rect 7719 5738 7777 5750
rect 7719 5362 7731 5738
rect 7765 5362 7777 5738
rect 7719 5350 7777 5362
rect 7837 5738 7895 5750
rect 7837 5362 7849 5738
rect 7883 5362 7895 5738
rect 7837 5350 7895 5362
rect 7955 5738 8013 5750
rect 7955 5362 7967 5738
rect 8001 5362 8013 5738
rect 7955 5350 8013 5362
rect 9315 5740 9373 5752
rect 9315 5364 9327 5740
rect 9361 5364 9373 5740
rect 9315 5352 9373 5364
rect 9433 5740 9491 5752
rect 9433 5364 9445 5740
rect 9479 5364 9491 5740
rect 9433 5352 9491 5364
rect 9551 5740 9609 5752
rect 9551 5364 9563 5740
rect 9597 5364 9609 5740
rect 9551 5352 9609 5364
rect 9669 5740 9727 5752
rect 9669 5364 9681 5740
rect 9715 5364 9727 5740
rect 9669 5352 9727 5364
rect 9787 5740 9845 5752
rect 9787 5364 9799 5740
rect 9833 5364 9845 5740
rect 9787 5352 9845 5364
rect 9905 5740 9963 5752
rect 9905 5364 9917 5740
rect 9951 5364 9963 5740
rect 9905 5352 9963 5364
rect 10023 5740 10081 5752
rect 10023 5364 10035 5740
rect 10069 5364 10081 5740
rect 10023 5352 10081 5364
rect 11384 5740 11442 5752
rect 11384 5364 11396 5740
rect 11430 5364 11442 5740
rect 11384 5352 11442 5364
rect 11502 5740 11560 5752
rect 11502 5364 11514 5740
rect 11548 5364 11560 5740
rect 11502 5352 11560 5364
rect 11620 5740 11678 5752
rect 11620 5364 11632 5740
rect 11666 5364 11678 5740
rect 11620 5352 11678 5364
rect 11738 5740 11796 5752
rect 11738 5364 11750 5740
rect 11784 5364 11796 5740
rect 11738 5352 11796 5364
rect 11856 5740 11914 5752
rect 11856 5364 11868 5740
rect 11902 5364 11914 5740
rect 11856 5352 11914 5364
rect 11974 5740 12032 5752
rect 11974 5364 11986 5740
rect 12020 5364 12032 5740
rect 11974 5352 12032 5364
rect 12092 5740 12150 5752
rect 12092 5364 12104 5740
rect 12138 5364 12150 5740
rect 12092 5352 12150 5364
rect 15094 6045 15152 6057
rect 15212 6233 15270 6245
rect 15212 6057 15224 6233
rect 15258 6057 15270 6233
rect 15212 6045 15270 6057
rect 15330 6233 15388 6245
rect 15330 6057 15342 6233
rect 15376 6057 15388 6233
rect 15330 6045 15388 6057
rect 15448 6233 15506 6245
rect 15448 6057 15460 6233
rect 15494 6057 15506 6233
rect 15448 6045 15506 6057
rect 15578 6057 15590 6433
rect 15624 6057 15636 6433
rect 15578 6045 15636 6057
rect 15696 6433 15754 6445
rect 15696 6057 15708 6433
rect 15742 6057 15754 6433
rect 15696 6045 15754 6057
rect 15814 6433 15872 6445
rect 15814 6057 15826 6433
rect 15860 6057 15872 6433
rect 15814 6045 15872 6057
rect 15932 6433 15990 6445
rect 15932 6057 15944 6433
rect 15978 6057 15990 6433
rect 15932 6045 15990 6057
rect 16050 6433 16108 6445
rect 16050 6057 16062 6433
rect 16096 6057 16108 6433
rect 16050 6045 16108 6057
rect 16168 6433 16226 6445
rect 16168 6057 16180 6433
rect 16214 6057 16226 6433
rect 16168 6045 16226 6057
rect 16286 6433 16344 6445
rect 16286 6057 16298 6433
rect 16332 6057 16344 6433
rect 17646 6435 17704 6447
rect 16286 6045 16344 6057
rect 16415 6233 16473 6245
rect 16415 6057 16427 6233
rect 16461 6057 16473 6233
rect 16415 6045 16473 6057
rect 16533 6233 16591 6245
rect 16533 6057 16545 6233
rect 16579 6057 16591 6233
rect 16533 6045 16591 6057
rect 16651 6233 16709 6245
rect 16651 6057 16663 6233
rect 16697 6057 16709 6233
rect 16651 6045 16709 6057
rect 16769 6233 16827 6245
rect 16769 6057 16781 6233
rect 16815 6057 16827 6233
rect 16769 6045 16827 6057
rect 17162 6235 17220 6247
rect 17162 6059 17174 6235
rect 17208 6059 17220 6235
rect 17162 6047 17220 6059
rect 17280 6235 17338 6247
rect 17280 6059 17292 6235
rect 17326 6059 17338 6235
rect 17280 6047 17338 6059
rect 17398 6235 17456 6247
rect 17398 6059 17410 6235
rect 17444 6059 17456 6235
rect 17398 6047 17456 6059
rect 17516 6235 17574 6247
rect 17516 6059 17528 6235
rect 17562 6059 17574 6235
rect 17516 6047 17574 6059
rect 17646 6059 17658 6435
rect 17692 6059 17704 6435
rect 17646 6047 17704 6059
rect 17764 6435 17822 6447
rect 17764 6059 17776 6435
rect 17810 6059 17822 6435
rect 17764 6047 17822 6059
rect 17882 6435 17940 6447
rect 17882 6059 17894 6435
rect 17928 6059 17940 6435
rect 17882 6047 17940 6059
rect 18000 6435 18058 6447
rect 18000 6059 18012 6435
rect 18046 6059 18058 6435
rect 18000 6047 18058 6059
rect 18118 6435 18176 6447
rect 18118 6059 18130 6435
rect 18164 6059 18176 6435
rect 18118 6047 18176 6059
rect 18236 6435 18294 6447
rect 18236 6059 18248 6435
rect 18282 6059 18294 6435
rect 18236 6047 18294 6059
rect 18354 6435 18412 6447
rect 18354 6059 18366 6435
rect 18400 6059 18412 6435
rect 19415 6371 19427 6547
rect 19461 6371 19473 6547
rect 19415 6359 19473 6371
rect 19533 6547 19591 6559
rect 19533 6371 19545 6547
rect 19579 6371 19591 6547
rect 19533 6359 19591 6371
rect 19651 6547 19709 6559
rect 19651 6371 19663 6547
rect 19697 6371 19709 6547
rect 19651 6359 19709 6371
rect 19769 6547 19827 6559
rect 19769 6371 19781 6547
rect 19815 6371 19827 6547
rect 19769 6359 19827 6371
rect 20153 6551 20211 6563
rect 20153 6375 20165 6551
rect 20199 6375 20211 6551
rect 20153 6363 20211 6375
rect 20271 6551 20329 6563
rect 20271 6375 20283 6551
rect 20317 6375 20329 6551
rect 20271 6363 20329 6375
rect 20389 6551 20447 6563
rect 20389 6375 20401 6551
rect 20435 6375 20447 6551
rect 20389 6363 20447 6375
rect 20507 6551 20565 6563
rect 20507 6375 20519 6551
rect 20553 6375 20565 6551
rect 20507 6363 20565 6375
rect 20891 6547 20949 6559
rect 20891 6371 20903 6547
rect 20937 6371 20949 6547
rect 20891 6359 20949 6371
rect 21009 6547 21067 6559
rect 21009 6371 21021 6547
rect 21055 6371 21067 6547
rect 21009 6359 21067 6371
rect 21127 6547 21185 6559
rect 21127 6371 21139 6547
rect 21173 6371 21185 6547
rect 21127 6359 21185 6371
rect 21245 6547 21303 6559
rect 21245 6371 21257 6547
rect 21291 6371 21303 6547
rect 21245 6359 21303 6371
rect 21633 6545 21691 6557
rect 21633 6369 21645 6545
rect 21679 6369 21691 6545
rect 21633 6357 21691 6369
rect 21751 6545 21809 6557
rect 21751 6369 21763 6545
rect 21797 6369 21809 6545
rect 21751 6357 21809 6369
rect 21869 6545 21927 6557
rect 21869 6369 21881 6545
rect 21915 6369 21927 6545
rect 21869 6357 21927 6369
rect 21987 6545 22045 6557
rect 21987 6369 21999 6545
rect 22033 6369 22045 6545
rect 21987 6357 22045 6369
rect 22373 6545 22431 6557
rect 22373 6369 22385 6545
rect 22419 6369 22431 6545
rect 22373 6357 22431 6369
rect 22491 6545 22549 6557
rect 22491 6369 22503 6545
rect 22537 6369 22549 6545
rect 22491 6357 22549 6369
rect 22609 6545 22667 6557
rect 22609 6369 22621 6545
rect 22655 6369 22667 6545
rect 22609 6357 22667 6369
rect 22727 6545 22785 6557
rect 22727 6369 22739 6545
rect 22773 6369 22785 6545
rect 22727 6357 22785 6369
rect 23111 6545 23169 6557
rect 23111 6369 23123 6545
rect 23157 6369 23169 6545
rect 23111 6357 23169 6369
rect 23229 6545 23287 6557
rect 23229 6369 23241 6545
rect 23275 6369 23287 6545
rect 23229 6357 23287 6369
rect 23347 6545 23405 6557
rect 23347 6369 23359 6545
rect 23393 6369 23405 6545
rect 23347 6357 23405 6369
rect 23465 6545 23523 6557
rect 23465 6369 23477 6545
rect 23511 6369 23523 6545
rect 23465 6357 23523 6369
rect 23849 6545 23907 6557
rect 23849 6369 23861 6545
rect 23895 6369 23907 6545
rect 23849 6357 23907 6369
rect 23967 6545 24025 6557
rect 23967 6369 23979 6545
rect 24013 6369 24025 6545
rect 23967 6357 24025 6369
rect 24085 6545 24143 6557
rect 24085 6369 24097 6545
rect 24131 6369 24143 6545
rect 24085 6357 24143 6369
rect 24203 6545 24261 6557
rect 24203 6369 24215 6545
rect 24249 6369 24261 6545
rect 24203 6357 24261 6369
rect 24587 6545 24645 6557
rect 24587 6369 24599 6545
rect 24633 6369 24645 6545
rect 24587 6357 24645 6369
rect 24705 6545 24763 6557
rect 24705 6369 24717 6545
rect 24751 6369 24763 6545
rect 24705 6357 24763 6369
rect 24823 6545 24881 6557
rect 24823 6369 24835 6545
rect 24869 6369 24881 6545
rect 24823 6357 24881 6369
rect 24941 6545 24999 6557
rect 24941 6369 24953 6545
rect 24987 6369 24999 6545
rect 24941 6357 24999 6369
rect 18354 6047 18412 6059
rect 18483 6235 18541 6247
rect 18483 6059 18495 6235
rect 18529 6059 18541 6235
rect 18483 6047 18541 6059
rect 18601 6235 18659 6247
rect 18601 6059 18613 6235
rect 18647 6059 18659 6235
rect 18601 6047 18659 6059
rect 18719 6235 18777 6247
rect 18719 6059 18731 6235
rect 18765 6059 18777 6235
rect 18719 6047 18777 6059
rect 18837 6235 18895 6247
rect 18837 6059 18849 6235
rect 18883 6059 18895 6235
rect 18837 6047 18895 6059
rect 13452 5742 13510 5754
rect 13452 5366 13464 5742
rect 13498 5366 13510 5742
rect 13452 5354 13510 5366
rect 13570 5742 13628 5754
rect 13570 5366 13582 5742
rect 13616 5366 13628 5742
rect 13570 5354 13628 5366
rect 13688 5742 13746 5754
rect 13688 5366 13700 5742
rect 13734 5366 13746 5742
rect 13688 5354 13746 5366
rect 13806 5742 13864 5754
rect 13806 5366 13818 5742
rect 13852 5366 13864 5742
rect 13806 5354 13864 5366
rect 13924 5742 13982 5754
rect 13924 5366 13936 5742
rect 13970 5366 13982 5742
rect 13924 5354 13982 5366
rect 14042 5742 14100 5754
rect 14042 5366 14054 5742
rect 14088 5366 14100 5742
rect 14042 5354 14100 5366
rect 14160 5742 14218 5754
rect 14160 5366 14172 5742
rect 14206 5366 14218 5742
rect 14160 5354 14218 5366
rect 15521 5740 15579 5752
rect 15521 5364 15533 5740
rect 15567 5364 15579 5740
rect 15521 5352 15579 5364
rect 15639 5740 15697 5752
rect 15639 5364 15651 5740
rect 15685 5364 15697 5740
rect 15639 5352 15697 5364
rect 15757 5740 15815 5752
rect 15757 5364 15769 5740
rect 15803 5364 15815 5740
rect 15757 5352 15815 5364
rect 15875 5740 15933 5752
rect 15875 5364 15887 5740
rect 15921 5364 15933 5740
rect 15875 5352 15933 5364
rect 15993 5740 16051 5752
rect 15993 5364 16005 5740
rect 16039 5364 16051 5740
rect 15993 5352 16051 5364
rect 16111 5740 16169 5752
rect 16111 5364 16123 5740
rect 16157 5364 16169 5740
rect 16111 5352 16169 5364
rect 16229 5740 16287 5752
rect 16229 5364 16241 5740
rect 16275 5364 16287 5740
rect 16229 5352 16287 5364
rect 17589 5742 17647 5754
rect 17589 5366 17601 5742
rect 17635 5366 17647 5742
rect 17589 5354 17647 5366
rect 17707 5742 17765 5754
rect 17707 5366 17719 5742
rect 17753 5366 17765 5742
rect 17707 5354 17765 5366
rect 17825 5742 17883 5754
rect 17825 5366 17837 5742
rect 17871 5366 17883 5742
rect 17825 5354 17883 5366
rect 17943 5742 18001 5754
rect 17943 5366 17955 5742
rect 17989 5366 18001 5742
rect 17943 5354 18001 5366
rect 18061 5742 18119 5754
rect 18061 5366 18073 5742
rect 18107 5366 18119 5742
rect 18061 5354 18119 5366
rect 18179 5742 18237 5754
rect 18179 5366 18191 5742
rect 18225 5366 18237 5742
rect 18179 5354 18237 5366
rect 18297 5742 18355 5754
rect 18297 5366 18309 5742
rect 18343 5366 18355 5742
rect 18297 5354 18355 5366
rect 689 2128 747 2140
rect 689 1940 701 2128
rect 248 1928 306 1940
rect 248 1752 260 1928
rect 294 1752 306 1928
rect 248 1740 306 1752
rect 366 1928 424 1940
rect 366 1752 378 1928
rect 412 1752 424 1928
rect 366 1740 424 1752
rect 484 1928 542 1940
rect 484 1752 496 1928
rect 530 1752 542 1928
rect 484 1740 542 1752
rect 602 1928 701 1940
rect 602 1752 614 1928
rect 648 1752 701 1928
rect 735 1752 747 2128
rect 602 1740 747 1752
rect 807 2128 865 2140
rect 807 1752 819 2128
rect 853 1752 865 2128
rect 807 1740 865 1752
rect 925 2128 983 2140
rect 925 1752 937 2128
rect 971 1752 983 2128
rect 925 1740 983 1752
rect 1043 2128 1101 2140
rect 1043 1752 1055 2128
rect 1089 1752 1101 2128
rect 1043 1740 1101 1752
rect 1156 2128 1214 2140
rect 1156 1752 1168 2128
rect 1202 1752 1214 2128
rect 1156 1740 1214 1752
rect 1274 2128 1332 2140
rect 1274 1752 1286 2128
rect 1320 1752 1332 2128
rect 1274 1740 1332 1752
rect 1392 2128 1450 2140
rect 1392 1752 1404 2128
rect 1438 1752 1450 2128
rect 1392 1740 1450 1752
rect 1510 2128 1568 2140
rect 1510 1752 1522 2128
rect 1556 1752 1568 2128
rect 1510 1740 1568 1752
rect 1628 2128 1686 2140
rect 1628 1752 1640 2128
rect 1674 1752 1686 2128
rect 1628 1740 1686 1752
rect 1746 2128 1804 2140
rect 1746 1752 1758 2128
rect 1792 1752 1804 2128
rect 1746 1740 1804 1752
rect 1864 2128 1922 2140
rect 1864 1752 1876 2128
rect 1910 1752 1922 2128
rect 1864 1740 1922 1752
rect 1983 2128 2041 2140
rect 1983 1752 1995 2128
rect 2029 1752 2041 2128
rect 1983 1740 2041 1752
rect 2101 2128 2159 2140
rect 2101 1752 2113 2128
rect 2147 1752 2159 2128
rect 2101 1740 2159 1752
rect 2219 2128 2277 2140
rect 2219 1752 2231 2128
rect 2265 1752 2277 2128
rect 2219 1740 2277 1752
rect 2337 2128 2395 2140
rect 2337 1752 2349 2128
rect 2383 1752 2395 2128
rect 3833 2128 3891 2140
rect 3833 1940 3845 2128
rect 2337 1740 2395 1752
rect 2456 1928 2514 1940
rect 2456 1752 2468 1928
rect 2502 1752 2514 1928
rect 2456 1740 2514 1752
rect 2574 1928 2632 1940
rect 2574 1752 2586 1928
rect 2620 1752 2632 1928
rect 2574 1740 2632 1752
rect 2692 1928 2750 1940
rect 2692 1752 2704 1928
rect 2738 1752 2750 1928
rect 2692 1740 2750 1752
rect 2810 1928 2868 1940
rect 2810 1752 2822 1928
rect 2856 1752 2868 1928
rect 2810 1740 2868 1752
rect 3392 1928 3450 1940
rect 3392 1752 3404 1928
rect 3438 1752 3450 1928
rect 3392 1740 3450 1752
rect 3510 1928 3568 1940
rect 3510 1752 3522 1928
rect 3556 1752 3568 1928
rect 3510 1740 3568 1752
rect 3628 1928 3686 1940
rect 3628 1752 3640 1928
rect 3674 1752 3686 1928
rect 3628 1740 3686 1752
rect 3746 1928 3845 1940
rect 3746 1752 3758 1928
rect 3792 1752 3845 1928
rect 3879 1752 3891 2128
rect 3746 1740 3891 1752
rect 3951 2128 4009 2140
rect 3951 1752 3963 2128
rect 3997 1752 4009 2128
rect 3951 1740 4009 1752
rect 4069 2128 4127 2140
rect 4069 1752 4081 2128
rect 4115 1752 4127 2128
rect 4069 1740 4127 1752
rect 4187 2128 4245 2140
rect 4187 1752 4199 2128
rect 4233 1752 4245 2128
rect 4187 1740 4245 1752
rect 4300 2128 4358 2140
rect 4300 1752 4312 2128
rect 4346 1752 4358 2128
rect 4300 1740 4358 1752
rect 4418 2128 4476 2140
rect 4418 1752 4430 2128
rect 4464 1752 4476 2128
rect 4418 1740 4476 1752
rect 4536 2128 4594 2140
rect 4536 1752 4548 2128
rect 4582 1752 4594 2128
rect 4536 1740 4594 1752
rect 4654 2128 4712 2140
rect 4654 1752 4666 2128
rect 4700 1752 4712 2128
rect 4654 1740 4712 1752
rect 4772 2128 4830 2140
rect 4772 1752 4784 2128
rect 4818 1752 4830 2128
rect 4772 1740 4830 1752
rect 4890 2128 4948 2140
rect 4890 1752 4902 2128
rect 4936 1752 4948 2128
rect 4890 1740 4948 1752
rect 5008 2128 5066 2140
rect 5008 1752 5020 2128
rect 5054 1752 5066 2128
rect 5008 1740 5066 1752
rect 5127 2128 5185 2140
rect 5127 1752 5139 2128
rect 5173 1752 5185 2128
rect 5127 1740 5185 1752
rect 5245 2128 5303 2140
rect 5245 1752 5257 2128
rect 5291 1752 5303 2128
rect 5245 1740 5303 1752
rect 5363 2128 5421 2140
rect 5363 1752 5375 2128
rect 5409 1752 5421 2128
rect 5363 1740 5421 1752
rect 5481 2128 5539 2140
rect 5481 1752 5493 2128
rect 5527 1752 5539 2128
rect 6965 2132 7023 2144
rect 6965 1944 6977 2132
rect 5481 1740 5539 1752
rect 5600 1928 5658 1940
rect 5600 1752 5612 1928
rect 5646 1752 5658 1928
rect 5600 1740 5658 1752
rect 5718 1928 5776 1940
rect 5718 1752 5730 1928
rect 5764 1752 5776 1928
rect 5718 1740 5776 1752
rect 5836 1928 5894 1940
rect 5836 1752 5848 1928
rect 5882 1752 5894 1928
rect 5836 1740 5894 1752
rect 5954 1928 6012 1940
rect 5954 1752 5966 1928
rect 6000 1752 6012 1928
rect 5954 1740 6012 1752
rect 6524 1932 6582 1944
rect 6524 1756 6536 1932
rect 6570 1756 6582 1932
rect 6524 1744 6582 1756
rect 6642 1932 6700 1944
rect 6642 1756 6654 1932
rect 6688 1756 6700 1932
rect 6642 1744 6700 1756
rect 6760 1932 6818 1944
rect 6760 1756 6772 1932
rect 6806 1756 6818 1932
rect 6760 1744 6818 1756
rect 6878 1932 6977 1944
rect 6878 1756 6890 1932
rect 6924 1756 6977 1932
rect 7011 1756 7023 2132
rect 6878 1744 7023 1756
rect 7083 2132 7141 2144
rect 7083 1756 7095 2132
rect 7129 1756 7141 2132
rect 7083 1744 7141 1756
rect 7201 2132 7259 2144
rect 7201 1756 7213 2132
rect 7247 1756 7259 2132
rect 7201 1744 7259 1756
rect 7319 2132 7377 2144
rect 7319 1756 7331 2132
rect 7365 1756 7377 2132
rect 7319 1744 7377 1756
rect 7432 2132 7490 2144
rect 7432 1756 7444 2132
rect 7478 1756 7490 2132
rect 7432 1744 7490 1756
rect 7550 2132 7608 2144
rect 7550 1756 7562 2132
rect 7596 1756 7608 2132
rect 7550 1744 7608 1756
rect 7668 2132 7726 2144
rect 7668 1756 7680 2132
rect 7714 1756 7726 2132
rect 7668 1744 7726 1756
rect 7786 2132 7844 2144
rect 7786 1756 7798 2132
rect 7832 1756 7844 2132
rect 7786 1744 7844 1756
rect 7904 2132 7962 2144
rect 7904 1756 7916 2132
rect 7950 1756 7962 2132
rect 7904 1744 7962 1756
rect 8022 2132 8080 2144
rect 8022 1756 8034 2132
rect 8068 1756 8080 2132
rect 8022 1744 8080 1756
rect 8140 2132 8198 2144
rect 8140 1756 8152 2132
rect 8186 1756 8198 2132
rect 8140 1744 8198 1756
rect 8259 2132 8317 2144
rect 8259 1756 8271 2132
rect 8305 1756 8317 2132
rect 8259 1744 8317 1756
rect 8377 2132 8435 2144
rect 8377 1756 8389 2132
rect 8423 1756 8435 2132
rect 8377 1744 8435 1756
rect 8495 2132 8553 2144
rect 8495 1756 8507 2132
rect 8541 1756 8553 2132
rect 8495 1744 8553 1756
rect 8613 2132 8671 2144
rect 8613 1756 8625 2132
rect 8659 1756 8671 2132
rect 10109 2132 10167 2144
rect 10109 1944 10121 2132
rect 8613 1744 8671 1756
rect 8732 1932 8790 1944
rect 8732 1756 8744 1932
rect 8778 1756 8790 1932
rect 8732 1744 8790 1756
rect 8850 1932 8908 1944
rect 8850 1756 8862 1932
rect 8896 1756 8908 1932
rect 8850 1744 8908 1756
rect 8968 1932 9026 1944
rect 8968 1756 8980 1932
rect 9014 1756 9026 1932
rect 8968 1744 9026 1756
rect 9086 1932 9144 1944
rect 9086 1756 9098 1932
rect 9132 1756 9144 1932
rect 9086 1744 9144 1756
rect 9668 1932 9726 1944
rect 9668 1756 9680 1932
rect 9714 1756 9726 1932
rect 9668 1744 9726 1756
rect 9786 1932 9844 1944
rect 9786 1756 9798 1932
rect 9832 1756 9844 1932
rect 9786 1744 9844 1756
rect 9904 1932 9962 1944
rect 9904 1756 9916 1932
rect 9950 1756 9962 1932
rect 9904 1744 9962 1756
rect 10022 1932 10121 1944
rect 10022 1756 10034 1932
rect 10068 1756 10121 1932
rect 10155 1756 10167 2132
rect 10022 1744 10167 1756
rect 10227 2132 10285 2144
rect 10227 1756 10239 2132
rect 10273 1756 10285 2132
rect 10227 1744 10285 1756
rect 10345 2132 10403 2144
rect 10345 1756 10357 2132
rect 10391 1756 10403 2132
rect 10345 1744 10403 1756
rect 10463 2132 10521 2144
rect 10463 1756 10475 2132
rect 10509 1756 10521 2132
rect 10463 1744 10521 1756
rect 10576 2132 10634 2144
rect 10576 1756 10588 2132
rect 10622 1756 10634 2132
rect 10576 1744 10634 1756
rect 10694 2132 10752 2144
rect 10694 1756 10706 2132
rect 10740 1756 10752 2132
rect 10694 1744 10752 1756
rect 10812 2132 10870 2144
rect 10812 1756 10824 2132
rect 10858 1756 10870 2132
rect 10812 1744 10870 1756
rect 10930 2132 10988 2144
rect 10930 1756 10942 2132
rect 10976 1756 10988 2132
rect 10930 1744 10988 1756
rect 11048 2132 11106 2144
rect 11048 1756 11060 2132
rect 11094 1756 11106 2132
rect 11048 1744 11106 1756
rect 11166 2132 11224 2144
rect 11166 1756 11178 2132
rect 11212 1756 11224 2132
rect 11166 1744 11224 1756
rect 11284 2132 11342 2144
rect 11284 1756 11296 2132
rect 11330 1756 11342 2132
rect 11284 1744 11342 1756
rect 11403 2132 11461 2144
rect 11403 1756 11415 2132
rect 11449 1756 11461 2132
rect 11403 1744 11461 1756
rect 11521 2132 11579 2144
rect 11521 1756 11533 2132
rect 11567 1756 11579 2132
rect 11521 1744 11579 1756
rect 11639 2132 11697 2144
rect 11639 1756 11651 2132
rect 11685 1756 11697 2132
rect 11639 1744 11697 1756
rect 11757 2132 11815 2144
rect 11757 1756 11769 2132
rect 11803 1756 11815 2132
rect 13311 2128 13369 2140
rect 11757 1744 11815 1756
rect 11876 1932 11934 1944
rect 11876 1756 11888 1932
rect 11922 1756 11934 1932
rect 11876 1744 11934 1756
rect 11994 1932 12052 1944
rect 11994 1756 12006 1932
rect 12040 1756 12052 1932
rect 11994 1744 12052 1756
rect 12112 1932 12170 1944
rect 12112 1756 12124 1932
rect 12158 1756 12170 1932
rect 12112 1744 12170 1756
rect 12230 1932 12288 1944
rect 13311 1940 13323 2128
rect 12230 1756 12242 1932
rect 12276 1756 12288 1932
rect 12230 1744 12288 1756
rect 12870 1928 12928 1940
rect 12870 1752 12882 1928
rect 12916 1752 12928 1928
rect 12870 1740 12928 1752
rect 12988 1928 13046 1940
rect 12988 1752 13000 1928
rect 13034 1752 13046 1928
rect 12988 1740 13046 1752
rect 13106 1928 13164 1940
rect 13106 1752 13118 1928
rect 13152 1752 13164 1928
rect 13106 1740 13164 1752
rect 13224 1928 13323 1940
rect 13224 1752 13236 1928
rect 13270 1752 13323 1928
rect 13357 1752 13369 2128
rect 13224 1740 13369 1752
rect 13429 2128 13487 2140
rect 13429 1752 13441 2128
rect 13475 1752 13487 2128
rect 13429 1740 13487 1752
rect 13547 2128 13605 2140
rect 13547 1752 13559 2128
rect 13593 1752 13605 2128
rect 13547 1740 13605 1752
rect 13665 2128 13723 2140
rect 13665 1752 13677 2128
rect 13711 1752 13723 2128
rect 13665 1740 13723 1752
rect 13778 2128 13836 2140
rect 13778 1752 13790 2128
rect 13824 1752 13836 2128
rect 13778 1740 13836 1752
rect 13896 2128 13954 2140
rect 13896 1752 13908 2128
rect 13942 1752 13954 2128
rect 13896 1740 13954 1752
rect 14014 2128 14072 2140
rect 14014 1752 14026 2128
rect 14060 1752 14072 2128
rect 14014 1740 14072 1752
rect 14132 2128 14190 2140
rect 14132 1752 14144 2128
rect 14178 1752 14190 2128
rect 14132 1740 14190 1752
rect 14250 2128 14308 2140
rect 14250 1752 14262 2128
rect 14296 1752 14308 2128
rect 14250 1740 14308 1752
rect 14368 2128 14426 2140
rect 14368 1752 14380 2128
rect 14414 1752 14426 2128
rect 14368 1740 14426 1752
rect 14486 2128 14544 2140
rect 14486 1752 14498 2128
rect 14532 1752 14544 2128
rect 14486 1740 14544 1752
rect 14605 2128 14663 2140
rect 14605 1752 14617 2128
rect 14651 1752 14663 2128
rect 14605 1740 14663 1752
rect 14723 2128 14781 2140
rect 14723 1752 14735 2128
rect 14769 1752 14781 2128
rect 14723 1740 14781 1752
rect 14841 2128 14899 2140
rect 14841 1752 14853 2128
rect 14887 1752 14899 2128
rect 14841 1740 14899 1752
rect 14959 2128 15017 2140
rect 14959 1752 14971 2128
rect 15005 1752 15017 2128
rect 16455 2128 16513 2140
rect 16455 1940 16467 2128
rect 14959 1740 15017 1752
rect 15078 1928 15136 1940
rect 15078 1752 15090 1928
rect 15124 1752 15136 1928
rect 15078 1740 15136 1752
rect 15196 1928 15254 1940
rect 15196 1752 15208 1928
rect 15242 1752 15254 1928
rect 15196 1740 15254 1752
rect 15314 1928 15372 1940
rect 15314 1752 15326 1928
rect 15360 1752 15372 1928
rect 15314 1740 15372 1752
rect 15432 1928 15490 1940
rect 15432 1752 15444 1928
rect 15478 1752 15490 1928
rect 15432 1740 15490 1752
rect 16014 1928 16072 1940
rect 16014 1752 16026 1928
rect 16060 1752 16072 1928
rect 16014 1740 16072 1752
rect 16132 1928 16190 1940
rect 16132 1752 16144 1928
rect 16178 1752 16190 1928
rect 16132 1740 16190 1752
rect 16250 1928 16308 1940
rect 16250 1752 16262 1928
rect 16296 1752 16308 1928
rect 16250 1740 16308 1752
rect 16368 1928 16467 1940
rect 16368 1752 16380 1928
rect 16414 1752 16467 1928
rect 16501 1752 16513 2128
rect 16368 1740 16513 1752
rect 16573 2128 16631 2140
rect 16573 1752 16585 2128
rect 16619 1752 16631 2128
rect 16573 1740 16631 1752
rect 16691 2128 16749 2140
rect 16691 1752 16703 2128
rect 16737 1752 16749 2128
rect 16691 1740 16749 1752
rect 16809 2128 16867 2140
rect 16809 1752 16821 2128
rect 16855 1752 16867 2128
rect 16809 1740 16867 1752
rect 16922 2128 16980 2140
rect 16922 1752 16934 2128
rect 16968 1752 16980 2128
rect 16922 1740 16980 1752
rect 17040 2128 17098 2140
rect 17040 1752 17052 2128
rect 17086 1752 17098 2128
rect 17040 1740 17098 1752
rect 17158 2128 17216 2140
rect 17158 1752 17170 2128
rect 17204 1752 17216 2128
rect 17158 1740 17216 1752
rect 17276 2128 17334 2140
rect 17276 1752 17288 2128
rect 17322 1752 17334 2128
rect 17276 1740 17334 1752
rect 17394 2128 17452 2140
rect 17394 1752 17406 2128
rect 17440 1752 17452 2128
rect 17394 1740 17452 1752
rect 17512 2128 17570 2140
rect 17512 1752 17524 2128
rect 17558 1752 17570 2128
rect 17512 1740 17570 1752
rect 17630 2128 17688 2140
rect 17630 1752 17642 2128
rect 17676 1752 17688 2128
rect 17630 1740 17688 1752
rect 17749 2128 17807 2140
rect 17749 1752 17761 2128
rect 17795 1752 17807 2128
rect 17749 1740 17807 1752
rect 17867 2128 17925 2140
rect 17867 1752 17879 2128
rect 17913 1752 17925 2128
rect 17867 1740 17925 1752
rect 17985 2128 18043 2140
rect 17985 1752 17997 2128
rect 18031 1752 18043 2128
rect 17985 1740 18043 1752
rect 18103 2128 18161 2140
rect 18103 1752 18115 2128
rect 18149 1752 18161 2128
rect 19587 2132 19645 2144
rect 19587 1944 19599 2132
rect 18103 1740 18161 1752
rect 18222 1928 18280 1940
rect 18222 1752 18234 1928
rect 18268 1752 18280 1928
rect 18222 1740 18280 1752
rect 18340 1928 18398 1940
rect 18340 1752 18352 1928
rect 18386 1752 18398 1928
rect 18340 1740 18398 1752
rect 18458 1928 18516 1940
rect 18458 1752 18470 1928
rect 18504 1752 18516 1928
rect 18458 1740 18516 1752
rect 18576 1928 18634 1940
rect 18576 1752 18588 1928
rect 18622 1752 18634 1928
rect 18576 1740 18634 1752
rect 19146 1932 19204 1944
rect 19146 1756 19158 1932
rect 19192 1756 19204 1932
rect 19146 1744 19204 1756
rect 19264 1932 19322 1944
rect 19264 1756 19276 1932
rect 19310 1756 19322 1932
rect 19264 1744 19322 1756
rect 19382 1932 19440 1944
rect 19382 1756 19394 1932
rect 19428 1756 19440 1932
rect 19382 1744 19440 1756
rect 19500 1932 19599 1944
rect 19500 1756 19512 1932
rect 19546 1756 19599 1932
rect 19633 1756 19645 2132
rect 19500 1744 19645 1756
rect 19705 2132 19763 2144
rect 19705 1756 19717 2132
rect 19751 1756 19763 2132
rect 19705 1744 19763 1756
rect 19823 2132 19881 2144
rect 19823 1756 19835 2132
rect 19869 1756 19881 2132
rect 19823 1744 19881 1756
rect 19941 2132 19999 2144
rect 19941 1756 19953 2132
rect 19987 1756 19999 2132
rect 19941 1744 19999 1756
rect 20054 2132 20112 2144
rect 20054 1756 20066 2132
rect 20100 1756 20112 2132
rect 20054 1744 20112 1756
rect 20172 2132 20230 2144
rect 20172 1756 20184 2132
rect 20218 1756 20230 2132
rect 20172 1744 20230 1756
rect 20290 2132 20348 2144
rect 20290 1756 20302 2132
rect 20336 1756 20348 2132
rect 20290 1744 20348 1756
rect 20408 2132 20466 2144
rect 20408 1756 20420 2132
rect 20454 1756 20466 2132
rect 20408 1744 20466 1756
rect 20526 2132 20584 2144
rect 20526 1756 20538 2132
rect 20572 1756 20584 2132
rect 20526 1744 20584 1756
rect 20644 2132 20702 2144
rect 20644 1756 20656 2132
rect 20690 1756 20702 2132
rect 20644 1744 20702 1756
rect 20762 2132 20820 2144
rect 20762 1756 20774 2132
rect 20808 1756 20820 2132
rect 20762 1744 20820 1756
rect 20881 2132 20939 2144
rect 20881 1756 20893 2132
rect 20927 1756 20939 2132
rect 20881 1744 20939 1756
rect 20999 2132 21057 2144
rect 20999 1756 21011 2132
rect 21045 1756 21057 2132
rect 20999 1744 21057 1756
rect 21117 2132 21175 2144
rect 21117 1756 21129 2132
rect 21163 1756 21175 2132
rect 21117 1744 21175 1756
rect 21235 2132 21293 2144
rect 21235 1756 21247 2132
rect 21281 1756 21293 2132
rect 22731 2132 22789 2144
rect 22731 1944 22743 2132
rect 21235 1744 21293 1756
rect 21354 1932 21412 1944
rect 21354 1756 21366 1932
rect 21400 1756 21412 1932
rect 21354 1744 21412 1756
rect 21472 1932 21530 1944
rect 21472 1756 21484 1932
rect 21518 1756 21530 1932
rect 21472 1744 21530 1756
rect 21590 1932 21648 1944
rect 21590 1756 21602 1932
rect 21636 1756 21648 1932
rect 21590 1744 21648 1756
rect 21708 1932 21766 1944
rect 21708 1756 21720 1932
rect 21754 1756 21766 1932
rect 21708 1744 21766 1756
rect 22290 1932 22348 1944
rect 22290 1756 22302 1932
rect 22336 1756 22348 1932
rect 22290 1744 22348 1756
rect 22408 1932 22466 1944
rect 22408 1756 22420 1932
rect 22454 1756 22466 1932
rect 22408 1744 22466 1756
rect 22526 1932 22584 1944
rect 22526 1756 22538 1932
rect 22572 1756 22584 1932
rect 22526 1744 22584 1756
rect 22644 1932 22743 1944
rect 22644 1756 22656 1932
rect 22690 1756 22743 1932
rect 22777 1756 22789 2132
rect 22644 1744 22789 1756
rect 22849 2132 22907 2144
rect 22849 1756 22861 2132
rect 22895 1756 22907 2132
rect 22849 1744 22907 1756
rect 22967 2132 23025 2144
rect 22967 1756 22979 2132
rect 23013 1756 23025 2132
rect 22967 1744 23025 1756
rect 23085 2132 23143 2144
rect 23085 1756 23097 2132
rect 23131 1756 23143 2132
rect 23085 1744 23143 1756
rect 23198 2132 23256 2144
rect 23198 1756 23210 2132
rect 23244 1756 23256 2132
rect 23198 1744 23256 1756
rect 23316 2132 23374 2144
rect 23316 1756 23328 2132
rect 23362 1756 23374 2132
rect 23316 1744 23374 1756
rect 23434 2132 23492 2144
rect 23434 1756 23446 2132
rect 23480 1756 23492 2132
rect 23434 1744 23492 1756
rect 23552 2132 23610 2144
rect 23552 1756 23564 2132
rect 23598 1756 23610 2132
rect 23552 1744 23610 1756
rect 23670 2132 23728 2144
rect 23670 1756 23682 2132
rect 23716 1756 23728 2132
rect 23670 1744 23728 1756
rect 23788 2132 23846 2144
rect 23788 1756 23800 2132
rect 23834 1756 23846 2132
rect 23788 1744 23846 1756
rect 23906 2132 23964 2144
rect 23906 1756 23918 2132
rect 23952 1756 23964 2132
rect 23906 1744 23964 1756
rect 24025 2132 24083 2144
rect 24025 1756 24037 2132
rect 24071 1756 24083 2132
rect 24025 1744 24083 1756
rect 24143 2132 24201 2144
rect 24143 1756 24155 2132
rect 24189 1756 24201 2132
rect 24143 1744 24201 1756
rect 24261 2132 24319 2144
rect 24261 1756 24273 2132
rect 24307 1756 24319 2132
rect 24261 1744 24319 1756
rect 24379 2132 24437 2144
rect 24379 1756 24391 2132
rect 24425 1756 24437 2132
rect 24379 1744 24437 1756
rect 24498 1932 24556 1944
rect 24498 1756 24510 1932
rect 24544 1756 24556 1932
rect 24498 1744 24556 1756
rect 24616 1932 24674 1944
rect 24616 1756 24628 1932
rect 24662 1756 24674 1932
rect 24616 1744 24674 1756
rect 24734 1932 24792 1944
rect 24734 1756 24746 1932
rect 24780 1756 24792 1932
rect 24734 1744 24792 1756
rect 24852 1932 24910 1944
rect 24852 1756 24864 1932
rect 24898 1756 24910 1932
rect 24852 1744 24910 1756
rect 721 -1764 779 -1752
rect 721 -1952 733 -1764
rect 280 -1964 338 -1952
rect 280 -2140 292 -1964
rect 326 -2140 338 -1964
rect 280 -2152 338 -2140
rect 398 -1964 456 -1952
rect 398 -2140 410 -1964
rect 444 -2140 456 -1964
rect 398 -2152 456 -2140
rect 516 -1964 574 -1952
rect 516 -2140 528 -1964
rect 562 -2140 574 -1964
rect 516 -2152 574 -2140
rect 634 -1964 733 -1952
rect 634 -2140 646 -1964
rect 680 -2140 733 -1964
rect 767 -2140 779 -1764
rect 634 -2152 779 -2140
rect 839 -1764 897 -1752
rect 839 -2140 851 -1764
rect 885 -2140 897 -1764
rect 839 -2152 897 -2140
rect 957 -1764 1015 -1752
rect 957 -2140 969 -1764
rect 1003 -2140 1015 -1764
rect 957 -2152 1015 -2140
rect 1075 -1764 1133 -1752
rect 1075 -2140 1087 -1764
rect 1121 -2140 1133 -1764
rect 1075 -2152 1133 -2140
rect 1188 -1764 1246 -1752
rect 1188 -2140 1200 -1764
rect 1234 -2140 1246 -1764
rect 1188 -2152 1246 -2140
rect 1306 -1764 1364 -1752
rect 1306 -2140 1318 -1764
rect 1352 -2140 1364 -1764
rect 1306 -2152 1364 -2140
rect 1424 -1764 1482 -1752
rect 1424 -2140 1436 -1764
rect 1470 -2140 1482 -1764
rect 1424 -2152 1482 -2140
rect 1542 -1764 1600 -1752
rect 1542 -2140 1554 -1764
rect 1588 -2140 1600 -1764
rect 1542 -2152 1600 -2140
rect 1660 -1764 1718 -1752
rect 1660 -2140 1672 -1764
rect 1706 -2140 1718 -1764
rect 1660 -2152 1718 -2140
rect 1778 -1764 1836 -1752
rect 1778 -2140 1790 -1764
rect 1824 -2140 1836 -1764
rect 1778 -2152 1836 -2140
rect 1896 -1764 1954 -1752
rect 1896 -2140 1908 -1764
rect 1942 -2140 1954 -1764
rect 1896 -2152 1954 -2140
rect 2015 -1764 2073 -1752
rect 2015 -2140 2027 -1764
rect 2061 -2140 2073 -1764
rect 2015 -2152 2073 -2140
rect 2133 -1764 2191 -1752
rect 2133 -2140 2145 -1764
rect 2179 -2140 2191 -1764
rect 2133 -2152 2191 -2140
rect 2251 -1764 2309 -1752
rect 2251 -2140 2263 -1764
rect 2297 -2140 2309 -1764
rect 2251 -2152 2309 -2140
rect 2369 -1764 2427 -1752
rect 2369 -2140 2381 -1764
rect 2415 -2140 2427 -1764
rect 3865 -1764 3923 -1752
rect 3865 -1952 3877 -1764
rect 2369 -2152 2427 -2140
rect 2488 -1964 2546 -1952
rect 2488 -2140 2500 -1964
rect 2534 -2140 2546 -1964
rect 2488 -2152 2546 -2140
rect 2606 -1964 2664 -1952
rect 2606 -2140 2618 -1964
rect 2652 -2140 2664 -1964
rect 2606 -2152 2664 -2140
rect 2724 -1964 2782 -1952
rect 2724 -2140 2736 -1964
rect 2770 -2140 2782 -1964
rect 2724 -2152 2782 -2140
rect 2842 -1964 2900 -1952
rect 2842 -2140 2854 -1964
rect 2888 -2140 2900 -1964
rect 2842 -2152 2900 -2140
rect 3424 -1964 3482 -1952
rect 3424 -2140 3436 -1964
rect 3470 -2140 3482 -1964
rect 3424 -2152 3482 -2140
rect 3542 -1964 3600 -1952
rect 3542 -2140 3554 -1964
rect 3588 -2140 3600 -1964
rect 3542 -2152 3600 -2140
rect 3660 -1964 3718 -1952
rect 3660 -2140 3672 -1964
rect 3706 -2140 3718 -1964
rect 3660 -2152 3718 -2140
rect 3778 -1964 3877 -1952
rect 3778 -2140 3790 -1964
rect 3824 -2140 3877 -1964
rect 3911 -2140 3923 -1764
rect 3778 -2152 3923 -2140
rect 3983 -1764 4041 -1752
rect 3983 -2140 3995 -1764
rect 4029 -2140 4041 -1764
rect 3983 -2152 4041 -2140
rect 4101 -1764 4159 -1752
rect 4101 -2140 4113 -1764
rect 4147 -2140 4159 -1764
rect 4101 -2152 4159 -2140
rect 4219 -1764 4277 -1752
rect 4219 -2140 4231 -1764
rect 4265 -2140 4277 -1764
rect 4219 -2152 4277 -2140
rect 4332 -1764 4390 -1752
rect 4332 -2140 4344 -1764
rect 4378 -2140 4390 -1764
rect 4332 -2152 4390 -2140
rect 4450 -1764 4508 -1752
rect 4450 -2140 4462 -1764
rect 4496 -2140 4508 -1764
rect 4450 -2152 4508 -2140
rect 4568 -1764 4626 -1752
rect 4568 -2140 4580 -1764
rect 4614 -2140 4626 -1764
rect 4568 -2152 4626 -2140
rect 4686 -1764 4744 -1752
rect 4686 -2140 4698 -1764
rect 4732 -2140 4744 -1764
rect 4686 -2152 4744 -2140
rect 4804 -1764 4862 -1752
rect 4804 -2140 4816 -1764
rect 4850 -2140 4862 -1764
rect 4804 -2152 4862 -2140
rect 4922 -1764 4980 -1752
rect 4922 -2140 4934 -1764
rect 4968 -2140 4980 -1764
rect 4922 -2152 4980 -2140
rect 5040 -1764 5098 -1752
rect 5040 -2140 5052 -1764
rect 5086 -2140 5098 -1764
rect 5040 -2152 5098 -2140
rect 5159 -1764 5217 -1752
rect 5159 -2140 5171 -1764
rect 5205 -2140 5217 -1764
rect 5159 -2152 5217 -2140
rect 5277 -1764 5335 -1752
rect 5277 -2140 5289 -1764
rect 5323 -2140 5335 -1764
rect 5277 -2152 5335 -2140
rect 5395 -1764 5453 -1752
rect 5395 -2140 5407 -1764
rect 5441 -2140 5453 -1764
rect 5395 -2152 5453 -2140
rect 5513 -1764 5571 -1752
rect 5513 -2140 5525 -1764
rect 5559 -2140 5571 -1764
rect 6997 -1760 7055 -1748
rect 6997 -1948 7009 -1760
rect 5513 -2152 5571 -2140
rect 5632 -1964 5690 -1952
rect 5632 -2140 5644 -1964
rect 5678 -2140 5690 -1964
rect 5632 -2152 5690 -2140
rect 5750 -1964 5808 -1952
rect 5750 -2140 5762 -1964
rect 5796 -2140 5808 -1964
rect 5750 -2152 5808 -2140
rect 5868 -1964 5926 -1952
rect 5868 -2140 5880 -1964
rect 5914 -2140 5926 -1964
rect 5868 -2152 5926 -2140
rect 5986 -1964 6044 -1952
rect 5986 -2140 5998 -1964
rect 6032 -2140 6044 -1964
rect 5986 -2152 6044 -2140
rect 6556 -1960 6614 -1948
rect 6556 -2136 6568 -1960
rect 6602 -2136 6614 -1960
rect 6556 -2148 6614 -2136
rect 6674 -1960 6732 -1948
rect 6674 -2136 6686 -1960
rect 6720 -2136 6732 -1960
rect 6674 -2148 6732 -2136
rect 6792 -1960 6850 -1948
rect 6792 -2136 6804 -1960
rect 6838 -2136 6850 -1960
rect 6792 -2148 6850 -2136
rect 6910 -1960 7009 -1948
rect 6910 -2136 6922 -1960
rect 6956 -2136 7009 -1960
rect 7043 -2136 7055 -1760
rect 6910 -2148 7055 -2136
rect 7115 -1760 7173 -1748
rect 7115 -2136 7127 -1760
rect 7161 -2136 7173 -1760
rect 7115 -2148 7173 -2136
rect 7233 -1760 7291 -1748
rect 7233 -2136 7245 -1760
rect 7279 -2136 7291 -1760
rect 7233 -2148 7291 -2136
rect 7351 -1760 7409 -1748
rect 7351 -2136 7363 -1760
rect 7397 -2136 7409 -1760
rect 7351 -2148 7409 -2136
rect 7464 -1760 7522 -1748
rect 7464 -2136 7476 -1760
rect 7510 -2136 7522 -1760
rect 7464 -2148 7522 -2136
rect 7582 -1760 7640 -1748
rect 7582 -2136 7594 -1760
rect 7628 -2136 7640 -1760
rect 7582 -2148 7640 -2136
rect 7700 -1760 7758 -1748
rect 7700 -2136 7712 -1760
rect 7746 -2136 7758 -1760
rect 7700 -2148 7758 -2136
rect 7818 -1760 7876 -1748
rect 7818 -2136 7830 -1760
rect 7864 -2136 7876 -1760
rect 7818 -2148 7876 -2136
rect 7936 -1760 7994 -1748
rect 7936 -2136 7948 -1760
rect 7982 -2136 7994 -1760
rect 7936 -2148 7994 -2136
rect 8054 -1760 8112 -1748
rect 8054 -2136 8066 -1760
rect 8100 -2136 8112 -1760
rect 8054 -2148 8112 -2136
rect 8172 -1760 8230 -1748
rect 8172 -2136 8184 -1760
rect 8218 -2136 8230 -1760
rect 8172 -2148 8230 -2136
rect 8291 -1760 8349 -1748
rect 8291 -2136 8303 -1760
rect 8337 -2136 8349 -1760
rect 8291 -2148 8349 -2136
rect 8409 -1760 8467 -1748
rect 8409 -2136 8421 -1760
rect 8455 -2136 8467 -1760
rect 8409 -2148 8467 -2136
rect 8527 -1760 8585 -1748
rect 8527 -2136 8539 -1760
rect 8573 -2136 8585 -1760
rect 8527 -2148 8585 -2136
rect 8645 -1760 8703 -1748
rect 8645 -2136 8657 -1760
rect 8691 -2136 8703 -1760
rect 10141 -1760 10199 -1748
rect 10141 -1948 10153 -1760
rect 8645 -2148 8703 -2136
rect 8764 -1960 8822 -1948
rect 8764 -2136 8776 -1960
rect 8810 -2136 8822 -1960
rect 8764 -2148 8822 -2136
rect 8882 -1960 8940 -1948
rect 8882 -2136 8894 -1960
rect 8928 -2136 8940 -1960
rect 8882 -2148 8940 -2136
rect 9000 -1960 9058 -1948
rect 9000 -2136 9012 -1960
rect 9046 -2136 9058 -1960
rect 9000 -2148 9058 -2136
rect 9118 -1960 9176 -1948
rect 9118 -2136 9130 -1960
rect 9164 -2136 9176 -1960
rect 9118 -2148 9176 -2136
rect 9700 -1960 9758 -1948
rect 9700 -2136 9712 -1960
rect 9746 -2136 9758 -1960
rect 9700 -2148 9758 -2136
rect 9818 -1960 9876 -1948
rect 9818 -2136 9830 -1960
rect 9864 -2136 9876 -1960
rect 9818 -2148 9876 -2136
rect 9936 -1960 9994 -1948
rect 9936 -2136 9948 -1960
rect 9982 -2136 9994 -1960
rect 9936 -2148 9994 -2136
rect 10054 -1960 10153 -1948
rect 10054 -2136 10066 -1960
rect 10100 -2136 10153 -1960
rect 10187 -2136 10199 -1760
rect 10054 -2148 10199 -2136
rect 10259 -1760 10317 -1748
rect 10259 -2136 10271 -1760
rect 10305 -2136 10317 -1760
rect 10259 -2148 10317 -2136
rect 10377 -1760 10435 -1748
rect 10377 -2136 10389 -1760
rect 10423 -2136 10435 -1760
rect 10377 -2148 10435 -2136
rect 10495 -1760 10553 -1748
rect 10495 -2136 10507 -1760
rect 10541 -2136 10553 -1760
rect 10495 -2148 10553 -2136
rect 10608 -1760 10666 -1748
rect 10608 -2136 10620 -1760
rect 10654 -2136 10666 -1760
rect 10608 -2148 10666 -2136
rect 10726 -1760 10784 -1748
rect 10726 -2136 10738 -1760
rect 10772 -2136 10784 -1760
rect 10726 -2148 10784 -2136
rect 10844 -1760 10902 -1748
rect 10844 -2136 10856 -1760
rect 10890 -2136 10902 -1760
rect 10844 -2148 10902 -2136
rect 10962 -1760 11020 -1748
rect 10962 -2136 10974 -1760
rect 11008 -2136 11020 -1760
rect 10962 -2148 11020 -2136
rect 11080 -1760 11138 -1748
rect 11080 -2136 11092 -1760
rect 11126 -2136 11138 -1760
rect 11080 -2148 11138 -2136
rect 11198 -1760 11256 -1748
rect 11198 -2136 11210 -1760
rect 11244 -2136 11256 -1760
rect 11198 -2148 11256 -2136
rect 11316 -1760 11374 -1748
rect 11316 -2136 11328 -1760
rect 11362 -2136 11374 -1760
rect 11316 -2148 11374 -2136
rect 11435 -1760 11493 -1748
rect 11435 -2136 11447 -1760
rect 11481 -2136 11493 -1760
rect 11435 -2148 11493 -2136
rect 11553 -1760 11611 -1748
rect 11553 -2136 11565 -1760
rect 11599 -2136 11611 -1760
rect 11553 -2148 11611 -2136
rect 11671 -1760 11729 -1748
rect 11671 -2136 11683 -1760
rect 11717 -2136 11729 -1760
rect 11671 -2148 11729 -2136
rect 11789 -1760 11847 -1748
rect 11789 -2136 11801 -1760
rect 11835 -2136 11847 -1760
rect 13343 -1764 13401 -1752
rect 11789 -2148 11847 -2136
rect 11908 -1960 11966 -1948
rect 11908 -2136 11920 -1960
rect 11954 -2136 11966 -1960
rect 11908 -2148 11966 -2136
rect 12026 -1960 12084 -1948
rect 12026 -2136 12038 -1960
rect 12072 -2136 12084 -1960
rect 12026 -2148 12084 -2136
rect 12144 -1960 12202 -1948
rect 12144 -2136 12156 -1960
rect 12190 -2136 12202 -1960
rect 12144 -2148 12202 -2136
rect 12262 -1960 12320 -1948
rect 13343 -1952 13355 -1764
rect 12262 -2136 12274 -1960
rect 12308 -2136 12320 -1960
rect 12262 -2148 12320 -2136
rect 12902 -1964 12960 -1952
rect 12902 -2140 12914 -1964
rect 12948 -2140 12960 -1964
rect 12902 -2152 12960 -2140
rect 13020 -1964 13078 -1952
rect 13020 -2140 13032 -1964
rect 13066 -2140 13078 -1964
rect 13020 -2152 13078 -2140
rect 13138 -1964 13196 -1952
rect 13138 -2140 13150 -1964
rect 13184 -2140 13196 -1964
rect 13138 -2152 13196 -2140
rect 13256 -1964 13355 -1952
rect 13256 -2140 13268 -1964
rect 13302 -2140 13355 -1964
rect 13389 -2140 13401 -1764
rect 13256 -2152 13401 -2140
rect 13461 -1764 13519 -1752
rect 13461 -2140 13473 -1764
rect 13507 -2140 13519 -1764
rect 13461 -2152 13519 -2140
rect 13579 -1764 13637 -1752
rect 13579 -2140 13591 -1764
rect 13625 -2140 13637 -1764
rect 13579 -2152 13637 -2140
rect 13697 -1764 13755 -1752
rect 13697 -2140 13709 -1764
rect 13743 -2140 13755 -1764
rect 13697 -2152 13755 -2140
rect 13810 -1764 13868 -1752
rect 13810 -2140 13822 -1764
rect 13856 -2140 13868 -1764
rect 13810 -2152 13868 -2140
rect 13928 -1764 13986 -1752
rect 13928 -2140 13940 -1764
rect 13974 -2140 13986 -1764
rect 13928 -2152 13986 -2140
rect 14046 -1764 14104 -1752
rect 14046 -2140 14058 -1764
rect 14092 -2140 14104 -1764
rect 14046 -2152 14104 -2140
rect 14164 -1764 14222 -1752
rect 14164 -2140 14176 -1764
rect 14210 -2140 14222 -1764
rect 14164 -2152 14222 -2140
rect 14282 -1764 14340 -1752
rect 14282 -2140 14294 -1764
rect 14328 -2140 14340 -1764
rect 14282 -2152 14340 -2140
rect 14400 -1764 14458 -1752
rect 14400 -2140 14412 -1764
rect 14446 -2140 14458 -1764
rect 14400 -2152 14458 -2140
rect 14518 -1764 14576 -1752
rect 14518 -2140 14530 -1764
rect 14564 -2140 14576 -1764
rect 14518 -2152 14576 -2140
rect 14637 -1764 14695 -1752
rect 14637 -2140 14649 -1764
rect 14683 -2140 14695 -1764
rect 14637 -2152 14695 -2140
rect 14755 -1764 14813 -1752
rect 14755 -2140 14767 -1764
rect 14801 -2140 14813 -1764
rect 14755 -2152 14813 -2140
rect 14873 -1764 14931 -1752
rect 14873 -2140 14885 -1764
rect 14919 -2140 14931 -1764
rect 14873 -2152 14931 -2140
rect 14991 -1764 15049 -1752
rect 14991 -2140 15003 -1764
rect 15037 -2140 15049 -1764
rect 16487 -1764 16545 -1752
rect 16487 -1952 16499 -1764
rect 14991 -2152 15049 -2140
rect 15110 -1964 15168 -1952
rect 15110 -2140 15122 -1964
rect 15156 -2140 15168 -1964
rect 15110 -2152 15168 -2140
rect 15228 -1964 15286 -1952
rect 15228 -2140 15240 -1964
rect 15274 -2140 15286 -1964
rect 15228 -2152 15286 -2140
rect 15346 -1964 15404 -1952
rect 15346 -2140 15358 -1964
rect 15392 -2140 15404 -1964
rect 15346 -2152 15404 -2140
rect 15464 -1964 15522 -1952
rect 15464 -2140 15476 -1964
rect 15510 -2140 15522 -1964
rect 15464 -2152 15522 -2140
rect 16046 -1964 16104 -1952
rect 16046 -2140 16058 -1964
rect 16092 -2140 16104 -1964
rect 16046 -2152 16104 -2140
rect 16164 -1964 16222 -1952
rect 16164 -2140 16176 -1964
rect 16210 -2140 16222 -1964
rect 16164 -2152 16222 -2140
rect 16282 -1964 16340 -1952
rect 16282 -2140 16294 -1964
rect 16328 -2140 16340 -1964
rect 16282 -2152 16340 -2140
rect 16400 -1964 16499 -1952
rect 16400 -2140 16412 -1964
rect 16446 -2140 16499 -1964
rect 16533 -2140 16545 -1764
rect 16400 -2152 16545 -2140
rect 16605 -1764 16663 -1752
rect 16605 -2140 16617 -1764
rect 16651 -2140 16663 -1764
rect 16605 -2152 16663 -2140
rect 16723 -1764 16781 -1752
rect 16723 -2140 16735 -1764
rect 16769 -2140 16781 -1764
rect 16723 -2152 16781 -2140
rect 16841 -1764 16899 -1752
rect 16841 -2140 16853 -1764
rect 16887 -2140 16899 -1764
rect 16841 -2152 16899 -2140
rect 16954 -1764 17012 -1752
rect 16954 -2140 16966 -1764
rect 17000 -2140 17012 -1764
rect 16954 -2152 17012 -2140
rect 17072 -1764 17130 -1752
rect 17072 -2140 17084 -1764
rect 17118 -2140 17130 -1764
rect 17072 -2152 17130 -2140
rect 17190 -1764 17248 -1752
rect 17190 -2140 17202 -1764
rect 17236 -2140 17248 -1764
rect 17190 -2152 17248 -2140
rect 17308 -1764 17366 -1752
rect 17308 -2140 17320 -1764
rect 17354 -2140 17366 -1764
rect 17308 -2152 17366 -2140
rect 17426 -1764 17484 -1752
rect 17426 -2140 17438 -1764
rect 17472 -2140 17484 -1764
rect 17426 -2152 17484 -2140
rect 17544 -1764 17602 -1752
rect 17544 -2140 17556 -1764
rect 17590 -2140 17602 -1764
rect 17544 -2152 17602 -2140
rect 17662 -1764 17720 -1752
rect 17662 -2140 17674 -1764
rect 17708 -2140 17720 -1764
rect 17662 -2152 17720 -2140
rect 17781 -1764 17839 -1752
rect 17781 -2140 17793 -1764
rect 17827 -2140 17839 -1764
rect 17781 -2152 17839 -2140
rect 17899 -1764 17957 -1752
rect 17899 -2140 17911 -1764
rect 17945 -2140 17957 -1764
rect 17899 -2152 17957 -2140
rect 18017 -1764 18075 -1752
rect 18017 -2140 18029 -1764
rect 18063 -2140 18075 -1764
rect 18017 -2152 18075 -2140
rect 18135 -1764 18193 -1752
rect 18135 -2140 18147 -1764
rect 18181 -2140 18193 -1764
rect 19619 -1760 19677 -1748
rect 19619 -1948 19631 -1760
rect 18135 -2152 18193 -2140
rect 18254 -1964 18312 -1952
rect 18254 -2140 18266 -1964
rect 18300 -2140 18312 -1964
rect 18254 -2152 18312 -2140
rect 18372 -1964 18430 -1952
rect 18372 -2140 18384 -1964
rect 18418 -2140 18430 -1964
rect 18372 -2152 18430 -2140
rect 18490 -1964 18548 -1952
rect 18490 -2140 18502 -1964
rect 18536 -2140 18548 -1964
rect 18490 -2152 18548 -2140
rect 18608 -1964 18666 -1952
rect 18608 -2140 18620 -1964
rect 18654 -2140 18666 -1964
rect 18608 -2152 18666 -2140
rect 19178 -1960 19236 -1948
rect 19178 -2136 19190 -1960
rect 19224 -2136 19236 -1960
rect 19178 -2148 19236 -2136
rect 19296 -1960 19354 -1948
rect 19296 -2136 19308 -1960
rect 19342 -2136 19354 -1960
rect 19296 -2148 19354 -2136
rect 19414 -1960 19472 -1948
rect 19414 -2136 19426 -1960
rect 19460 -2136 19472 -1960
rect 19414 -2148 19472 -2136
rect 19532 -1960 19631 -1948
rect 19532 -2136 19544 -1960
rect 19578 -2136 19631 -1960
rect 19665 -2136 19677 -1760
rect 19532 -2148 19677 -2136
rect 19737 -1760 19795 -1748
rect 19737 -2136 19749 -1760
rect 19783 -2136 19795 -1760
rect 19737 -2148 19795 -2136
rect 19855 -1760 19913 -1748
rect 19855 -2136 19867 -1760
rect 19901 -2136 19913 -1760
rect 19855 -2148 19913 -2136
rect 19973 -1760 20031 -1748
rect 19973 -2136 19985 -1760
rect 20019 -2136 20031 -1760
rect 19973 -2148 20031 -2136
rect 20086 -1760 20144 -1748
rect 20086 -2136 20098 -1760
rect 20132 -2136 20144 -1760
rect 20086 -2148 20144 -2136
rect 20204 -1760 20262 -1748
rect 20204 -2136 20216 -1760
rect 20250 -2136 20262 -1760
rect 20204 -2148 20262 -2136
rect 20322 -1760 20380 -1748
rect 20322 -2136 20334 -1760
rect 20368 -2136 20380 -1760
rect 20322 -2148 20380 -2136
rect 20440 -1760 20498 -1748
rect 20440 -2136 20452 -1760
rect 20486 -2136 20498 -1760
rect 20440 -2148 20498 -2136
rect 20558 -1760 20616 -1748
rect 20558 -2136 20570 -1760
rect 20604 -2136 20616 -1760
rect 20558 -2148 20616 -2136
rect 20676 -1760 20734 -1748
rect 20676 -2136 20688 -1760
rect 20722 -2136 20734 -1760
rect 20676 -2148 20734 -2136
rect 20794 -1760 20852 -1748
rect 20794 -2136 20806 -1760
rect 20840 -2136 20852 -1760
rect 20794 -2148 20852 -2136
rect 20913 -1760 20971 -1748
rect 20913 -2136 20925 -1760
rect 20959 -2136 20971 -1760
rect 20913 -2148 20971 -2136
rect 21031 -1760 21089 -1748
rect 21031 -2136 21043 -1760
rect 21077 -2136 21089 -1760
rect 21031 -2148 21089 -2136
rect 21149 -1760 21207 -1748
rect 21149 -2136 21161 -1760
rect 21195 -2136 21207 -1760
rect 21149 -2148 21207 -2136
rect 21267 -1760 21325 -1748
rect 21267 -2136 21279 -1760
rect 21313 -2136 21325 -1760
rect 22763 -1760 22821 -1748
rect 22763 -1948 22775 -1760
rect 21267 -2148 21325 -2136
rect 21386 -1960 21444 -1948
rect 21386 -2136 21398 -1960
rect 21432 -2136 21444 -1960
rect 21386 -2148 21444 -2136
rect 21504 -1960 21562 -1948
rect 21504 -2136 21516 -1960
rect 21550 -2136 21562 -1960
rect 21504 -2148 21562 -2136
rect 21622 -1960 21680 -1948
rect 21622 -2136 21634 -1960
rect 21668 -2136 21680 -1960
rect 21622 -2148 21680 -2136
rect 21740 -1960 21798 -1948
rect 21740 -2136 21752 -1960
rect 21786 -2136 21798 -1960
rect 21740 -2148 21798 -2136
rect 22322 -1960 22380 -1948
rect 22322 -2136 22334 -1960
rect 22368 -2136 22380 -1960
rect 22322 -2148 22380 -2136
rect 22440 -1960 22498 -1948
rect 22440 -2136 22452 -1960
rect 22486 -2136 22498 -1960
rect 22440 -2148 22498 -2136
rect 22558 -1960 22616 -1948
rect 22558 -2136 22570 -1960
rect 22604 -2136 22616 -1960
rect 22558 -2148 22616 -2136
rect 22676 -1960 22775 -1948
rect 22676 -2136 22688 -1960
rect 22722 -2136 22775 -1960
rect 22809 -2136 22821 -1760
rect 22676 -2148 22821 -2136
rect 22881 -1760 22939 -1748
rect 22881 -2136 22893 -1760
rect 22927 -2136 22939 -1760
rect 22881 -2148 22939 -2136
rect 22999 -1760 23057 -1748
rect 22999 -2136 23011 -1760
rect 23045 -2136 23057 -1760
rect 22999 -2148 23057 -2136
rect 23117 -1760 23175 -1748
rect 23117 -2136 23129 -1760
rect 23163 -2136 23175 -1760
rect 23117 -2148 23175 -2136
rect 23230 -1760 23288 -1748
rect 23230 -2136 23242 -1760
rect 23276 -2136 23288 -1760
rect 23230 -2148 23288 -2136
rect 23348 -1760 23406 -1748
rect 23348 -2136 23360 -1760
rect 23394 -2136 23406 -1760
rect 23348 -2148 23406 -2136
rect 23466 -1760 23524 -1748
rect 23466 -2136 23478 -1760
rect 23512 -2136 23524 -1760
rect 23466 -2148 23524 -2136
rect 23584 -1760 23642 -1748
rect 23584 -2136 23596 -1760
rect 23630 -2136 23642 -1760
rect 23584 -2148 23642 -2136
rect 23702 -1760 23760 -1748
rect 23702 -2136 23714 -1760
rect 23748 -2136 23760 -1760
rect 23702 -2148 23760 -2136
rect 23820 -1760 23878 -1748
rect 23820 -2136 23832 -1760
rect 23866 -2136 23878 -1760
rect 23820 -2148 23878 -2136
rect 23938 -1760 23996 -1748
rect 23938 -2136 23950 -1760
rect 23984 -2136 23996 -1760
rect 23938 -2148 23996 -2136
rect 24057 -1760 24115 -1748
rect 24057 -2136 24069 -1760
rect 24103 -2136 24115 -1760
rect 24057 -2148 24115 -2136
rect 24175 -1760 24233 -1748
rect 24175 -2136 24187 -1760
rect 24221 -2136 24233 -1760
rect 24175 -2148 24233 -2136
rect 24293 -1760 24351 -1748
rect 24293 -2136 24305 -1760
rect 24339 -2136 24351 -1760
rect 24293 -2148 24351 -2136
rect 24411 -1760 24469 -1748
rect 24411 -2136 24423 -1760
rect 24457 -2136 24469 -1760
rect 24411 -2148 24469 -2136
rect 24530 -1960 24588 -1948
rect 24530 -2136 24542 -1960
rect 24576 -2136 24588 -1960
rect 24530 -2148 24588 -2136
rect 24648 -1960 24706 -1948
rect 24648 -2136 24660 -1960
rect 24694 -2136 24706 -1960
rect 24648 -2148 24706 -2136
rect 24766 -1960 24824 -1948
rect 24766 -2136 24778 -1960
rect 24812 -2136 24824 -1960
rect 24766 -2148 24824 -2136
rect 24884 -1960 24942 -1948
rect 24884 -2136 24896 -1960
rect 24930 -2136 24942 -1960
rect 24884 -2148 24942 -2136
<< ndiffc >>
rect 1300 20471 1334 20647
rect 1418 20471 1452 20647
rect 1492 20271 1526 20647
rect 1610 20271 1644 20647
rect 1728 20271 1762 20647
rect 1846 20271 1880 20647
rect 1964 20271 1998 20647
rect 2042 20471 2076 20647
rect 2160 20471 2194 20647
rect 4444 20471 4478 20647
rect 4562 20471 4596 20647
rect 4636 20271 4670 20647
rect 4754 20271 4788 20647
rect 4872 20271 4906 20647
rect 4990 20271 5024 20647
rect 5108 20271 5142 20647
rect 5186 20471 5220 20647
rect 5304 20471 5338 20647
rect 7576 20475 7610 20651
rect 7694 20475 7728 20651
rect 7768 20275 7802 20651
rect 7886 20275 7920 20651
rect 8004 20275 8038 20651
rect 8122 20275 8156 20651
rect 8240 20275 8274 20651
rect 8318 20475 8352 20651
rect 8436 20475 8470 20651
rect 10720 20475 10754 20651
rect 10838 20475 10872 20651
rect 10912 20275 10946 20651
rect 11030 20275 11064 20651
rect 11148 20275 11182 20651
rect 11266 20275 11300 20651
rect 11384 20275 11418 20651
rect 11462 20475 11496 20651
rect 11580 20475 11614 20651
rect 13922 20471 13956 20647
rect 14040 20471 14074 20647
rect 14114 20271 14148 20647
rect 14232 20271 14266 20647
rect 14350 20271 14384 20647
rect 14468 20271 14502 20647
rect 14586 20271 14620 20647
rect 14664 20471 14698 20647
rect 14782 20471 14816 20647
rect 17066 20471 17100 20647
rect 17184 20471 17218 20647
rect 17258 20271 17292 20647
rect 17376 20271 17410 20647
rect 17494 20271 17528 20647
rect 17612 20271 17646 20647
rect 17730 20271 17764 20647
rect 17808 20471 17842 20647
rect 17926 20471 17960 20647
rect 20198 20475 20232 20651
rect 20316 20475 20350 20651
rect 20390 20275 20424 20651
rect 20508 20275 20542 20651
rect 20626 20275 20660 20651
rect 20744 20275 20778 20651
rect 20862 20275 20896 20651
rect 20940 20475 20974 20651
rect 21058 20475 21092 20651
rect 23342 20475 23376 20651
rect 23460 20475 23494 20651
rect 23534 20275 23568 20651
rect 23652 20275 23686 20651
rect 23770 20275 23804 20651
rect 23888 20275 23922 20651
rect 24006 20275 24040 20651
rect 24084 20475 24118 20651
rect 24202 20475 24236 20651
rect 3146 15786 3180 16162
rect 3264 15786 3298 16162
rect 3382 15786 3416 16162
rect 3499 15986 3533 16162
rect 3617 15986 3651 16162
rect 4594 15786 4628 16162
rect 4712 15786 4746 16162
rect 4830 15786 4864 16162
rect 4947 15986 4981 16162
rect 5065 15986 5099 16162
rect 6092 15788 6126 16164
rect 6210 15788 6244 16164
rect 6328 15788 6362 16164
rect 6445 15988 6479 16164
rect 6563 15988 6597 16164
rect 7540 15788 7574 16164
rect 7658 15788 7692 16164
rect 7776 15788 7810 16164
rect 7893 15988 7927 16164
rect 8011 15988 8045 16164
rect 9060 15786 9094 16162
rect 9178 15786 9212 16162
rect 9296 15786 9330 16162
rect 9413 15986 9447 16162
rect 9531 15986 9565 16162
rect 10508 15786 10542 16162
rect 10626 15786 10660 16162
rect 10744 15786 10778 16162
rect 10861 15986 10895 16162
rect 10979 15986 11013 16162
rect 12006 15788 12040 16164
rect 12124 15788 12158 16164
rect 12242 15788 12276 16164
rect 12359 15988 12393 16164
rect 12477 15988 12511 16164
rect 13454 15788 13488 16164
rect 13572 15788 13606 16164
rect 13690 15788 13724 16164
rect 13807 15988 13841 16164
rect 13925 15988 13959 16164
rect 14582 15834 14616 16010
rect 14700 15834 14734 16010
rect 14818 15834 14852 16010
rect 14936 15834 14970 16010
rect 15750 15836 15784 16012
rect 15868 15836 15902 16012
rect 15986 15836 16020 16012
rect 16104 15836 16138 16012
rect 16918 15836 16952 16012
rect 17036 15836 17070 16012
rect 17154 15836 17188 16012
rect 17272 15836 17306 16012
rect 18086 15836 18120 16012
rect 18204 15836 18238 16012
rect 18322 15836 18356 16012
rect 18440 15836 18474 16012
rect 19260 15836 19294 16012
rect 19378 15836 19412 16012
rect 19496 15836 19530 16012
rect 19614 15836 19648 16012
rect 20428 15836 20462 16012
rect 20546 15836 20580 16012
rect 20664 15836 20698 16012
rect 20782 15836 20816 16012
rect 21596 15838 21630 16014
rect 21714 15838 21748 16014
rect 21832 15838 21866 16014
rect 21950 15838 21984 16014
rect 22764 15838 22798 16014
rect 22882 15838 22916 16014
rect 23000 15838 23034 16014
rect 23118 15838 23152 16014
rect 3802 13333 3836 13509
rect 3920 13333 3954 13509
rect 3994 13133 4028 13509
rect 4112 13133 4146 13509
rect 4230 13133 4264 13509
rect 4348 13133 4382 13509
rect 4466 13133 4500 13509
rect 4544 13333 4578 13509
rect 4662 13333 4696 13509
rect 6946 13333 6980 13509
rect 7064 13333 7098 13509
rect 7138 13133 7172 13509
rect 7256 13133 7290 13509
rect 7374 13133 7408 13509
rect 7492 13133 7526 13509
rect 7610 13133 7644 13509
rect 7688 13333 7722 13509
rect 7806 13333 7840 13509
rect 10078 13337 10112 13513
rect 10196 13337 10230 13513
rect 10270 13137 10304 13513
rect 10388 13137 10422 13513
rect 10506 13137 10540 13513
rect 10624 13137 10658 13513
rect 10742 13137 10776 13513
rect 10820 13337 10854 13513
rect 10938 13337 10972 13513
rect 13222 13337 13256 13513
rect 13340 13337 13374 13513
rect 13414 13137 13448 13513
rect 13532 13137 13566 13513
rect 13650 13137 13684 13513
rect 13768 13137 13802 13513
rect 13886 13137 13920 13513
rect 13964 13337 13998 13513
rect 14082 13337 14116 13513
rect 16424 13333 16458 13509
rect 16542 13333 16576 13509
rect 16616 13133 16650 13509
rect 16734 13133 16768 13509
rect 16852 13133 16886 13509
rect 16970 13133 17004 13509
rect 17088 13133 17122 13509
rect 17166 13333 17200 13509
rect 17284 13333 17318 13509
rect 19568 13333 19602 13509
rect 19686 13333 19720 13509
rect 19760 13133 19794 13509
rect 19878 13133 19912 13509
rect 19996 13133 20030 13509
rect 20114 13133 20148 13509
rect 20232 13133 20266 13509
rect 20310 13333 20344 13509
rect 20428 13333 20462 13509
rect 22700 13337 22734 13513
rect 22818 13337 22852 13513
rect 22892 13137 22926 13513
rect 23010 13137 23044 13513
rect 23128 13137 23162 13513
rect 23246 13137 23280 13513
rect 23364 13137 23398 13513
rect 23442 13337 23476 13513
rect 23560 13337 23594 13513
rect 25844 13337 25878 13513
rect 25962 13337 25996 13513
rect 26036 13137 26070 13513
rect 26154 13137 26188 13513
rect 26272 13137 26306 13513
rect 26390 13137 26424 13513
rect 26508 13137 26542 13513
rect 26586 13337 26620 13513
rect 26704 13337 26738 13513
rect 3802 10599 3836 10775
rect 3920 10599 3954 10775
rect 3994 10399 4028 10775
rect 4112 10399 4146 10775
rect 4230 10399 4264 10775
rect 4348 10399 4382 10775
rect 4466 10399 4500 10775
rect 4544 10599 4578 10775
rect 4662 10599 4696 10775
rect 6946 10599 6980 10775
rect 7064 10599 7098 10775
rect 7138 10399 7172 10775
rect 7256 10399 7290 10775
rect 7374 10399 7408 10775
rect 7492 10399 7526 10775
rect 7610 10399 7644 10775
rect 7688 10599 7722 10775
rect 7806 10599 7840 10775
rect 10078 10603 10112 10779
rect 10196 10603 10230 10779
rect 10270 10403 10304 10779
rect 10388 10403 10422 10779
rect 10506 10403 10540 10779
rect 10624 10403 10658 10779
rect 10742 10403 10776 10779
rect 10820 10603 10854 10779
rect 10938 10603 10972 10779
rect 13222 10603 13256 10779
rect 13340 10603 13374 10779
rect 13414 10403 13448 10779
rect 13532 10403 13566 10779
rect 13650 10403 13684 10779
rect 13768 10403 13802 10779
rect 13886 10403 13920 10779
rect 13964 10603 13998 10779
rect 14082 10603 14116 10779
rect 16424 10599 16458 10775
rect 16542 10599 16576 10775
rect 16616 10399 16650 10775
rect 16734 10399 16768 10775
rect 16852 10399 16886 10775
rect 16970 10399 17004 10775
rect 17088 10399 17122 10775
rect 17166 10599 17200 10775
rect 17284 10599 17318 10775
rect 19568 10599 19602 10775
rect 19686 10599 19720 10775
rect 19760 10399 19794 10775
rect 19878 10399 19912 10775
rect 19996 10399 20030 10775
rect 20114 10399 20148 10775
rect 20232 10399 20266 10775
rect 20310 10599 20344 10775
rect 20428 10599 20462 10775
rect 22700 10603 22734 10779
rect 22818 10603 22852 10779
rect 22892 10403 22926 10779
rect 23010 10403 23044 10779
rect 23128 10403 23162 10779
rect 23246 10403 23280 10779
rect 23364 10403 23398 10779
rect 23442 10603 23476 10779
rect 23560 10603 23594 10779
rect 25844 10603 25878 10779
rect 25962 10603 25996 10779
rect 26036 10403 26070 10779
rect 26154 10403 26188 10779
rect 26272 10403 26306 10779
rect 26390 10403 26424 10779
rect 26508 10403 26542 10779
rect 26586 10603 26620 10779
rect 26704 10603 26738 10779
rect 3792 7867 3826 8043
rect 3910 7867 3944 8043
rect 3984 7667 4018 8043
rect 4102 7667 4136 8043
rect 4220 7667 4254 8043
rect 4338 7667 4372 8043
rect 4456 7667 4490 8043
rect 4534 7867 4568 8043
rect 4652 7867 4686 8043
rect 6936 7867 6970 8043
rect 7054 7867 7088 8043
rect 7128 7667 7162 8043
rect 7246 7667 7280 8043
rect 7364 7667 7398 8043
rect 7482 7667 7516 8043
rect 7600 7667 7634 8043
rect 7678 7867 7712 8043
rect 7796 7867 7830 8043
rect 10068 7871 10102 8047
rect 10186 7871 10220 8047
rect 10260 7671 10294 8047
rect 10378 7671 10412 8047
rect 10496 7671 10530 8047
rect 10614 7671 10648 8047
rect 10732 7671 10766 8047
rect 10810 7871 10844 8047
rect 10928 7871 10962 8047
rect 13212 7871 13246 8047
rect 13330 7871 13364 8047
rect 13404 7671 13438 8047
rect 13522 7671 13556 8047
rect 13640 7671 13674 8047
rect 13758 7671 13792 8047
rect 13876 7671 13910 8047
rect 13954 7871 13988 8047
rect 14072 7871 14106 8047
rect 16414 7867 16448 8043
rect 16532 7867 16566 8043
rect 16606 7667 16640 8043
rect 16724 7667 16758 8043
rect 16842 7667 16876 8043
rect 16960 7667 16994 8043
rect 17078 7667 17112 8043
rect 17156 7867 17190 8043
rect 17274 7867 17308 8043
rect 19558 7867 19592 8043
rect 19676 7867 19710 8043
rect 19750 7667 19784 8043
rect 19868 7667 19902 8043
rect 19986 7667 20020 8043
rect 20104 7667 20138 8043
rect 20222 7667 20256 8043
rect 20300 7867 20334 8043
rect 20418 7867 20452 8043
rect 22690 7871 22724 8047
rect 22808 7871 22842 8047
rect 22882 7671 22916 8047
rect 23000 7671 23034 8047
rect 23118 7671 23152 8047
rect 23236 7671 23270 8047
rect 23354 7671 23388 8047
rect 23432 7871 23466 8047
rect 23550 7871 23584 8047
rect 25834 7871 25868 8047
rect 25952 7871 25986 8047
rect 26026 7671 26060 8047
rect 26144 7671 26178 8047
rect 26262 7671 26296 8047
rect 26380 7671 26414 8047
rect 26498 7671 26532 8047
rect 26576 7871 26610 8047
rect 26694 7871 26728 8047
rect 2820 4830 2854 5006
rect 2938 4830 2972 5006
rect 3240 4630 3274 5006
rect 3358 4630 3392 5006
rect 3476 4630 3510 5006
rect 3594 4630 3628 5006
rect 3712 4630 3746 5006
rect 4118 4830 4152 5006
rect 4236 4830 4270 5006
rect 4888 4832 4922 5008
rect 5006 4832 5040 5008
rect 5308 4632 5342 5008
rect 5426 4632 5460 5008
rect 5544 4632 5578 5008
rect 5662 4632 5696 5008
rect 5780 4632 5814 5008
rect 6186 4832 6220 5008
rect 6304 4832 6338 5008
rect 6957 4830 6991 5006
rect 7075 4830 7109 5006
rect 7377 4630 7411 5006
rect 7495 4630 7529 5006
rect 7613 4630 7647 5006
rect 7731 4630 7765 5006
rect 7849 4630 7883 5006
rect 8255 4830 8289 5006
rect 8373 4830 8407 5006
rect 9025 4832 9059 5008
rect 9143 4832 9177 5008
rect 9445 4632 9479 5008
rect 9563 4632 9597 5008
rect 9681 4632 9715 5008
rect 9799 4632 9833 5008
rect 9917 4632 9951 5008
rect 10323 4832 10357 5008
rect 10441 4832 10475 5008
rect 11094 4832 11128 5008
rect 11212 4832 11246 5008
rect 11514 4632 11548 5008
rect 11632 4632 11666 5008
rect 11750 4632 11784 5008
rect 11868 4632 11902 5008
rect 11986 4632 12020 5008
rect 12392 4832 12426 5008
rect 12510 4832 12544 5008
rect 13162 4834 13196 5010
rect 13280 4834 13314 5010
rect 13582 4634 13616 5010
rect 13700 4634 13734 5010
rect 13818 4634 13852 5010
rect 13936 4634 13970 5010
rect 14054 4634 14088 5010
rect 14460 4834 14494 5010
rect 19545 5985 19579 6161
rect 19663 5985 19697 6161
rect 20283 5987 20317 6163
rect 20401 5987 20435 6163
rect 21021 5983 21055 6159
rect 21139 5983 21173 6159
rect 21763 5983 21797 6159
rect 21881 5983 21915 6159
rect 22503 5983 22537 6159
rect 22621 5983 22655 6159
rect 23241 5983 23275 6159
rect 23359 5983 23393 6159
rect 23979 5987 24013 6163
rect 24097 5987 24131 6163
rect 24717 5987 24751 6163
rect 24835 5987 24869 6163
rect 14578 4834 14612 5010
rect 15231 4832 15265 5008
rect 15349 4832 15383 5008
rect 15651 4632 15685 5008
rect 15769 4632 15803 5008
rect 15887 4632 15921 5008
rect 16005 4632 16039 5008
rect 16123 4632 16157 5008
rect 16529 4832 16563 5008
rect 16647 4832 16681 5008
rect 17299 4834 17333 5010
rect 17417 4834 17451 5010
rect 17719 4634 17753 5010
rect 17837 4634 17871 5010
rect 17955 4634 17989 5010
rect 18073 4634 18107 5010
rect 18191 4634 18225 5010
rect 18597 4834 18631 5010
rect 18715 4834 18749 5010
rect 1094 619 1128 795
rect 1212 619 1246 795
rect 1286 419 1320 795
rect 1404 419 1438 795
rect 1522 419 1556 795
rect 1640 419 1674 795
rect 1758 419 1792 795
rect 1836 619 1870 795
rect 1954 619 1988 795
rect 4238 619 4272 795
rect 4356 619 4390 795
rect 4430 419 4464 795
rect 4548 419 4582 795
rect 4666 419 4700 795
rect 4784 419 4818 795
rect 4902 419 4936 795
rect 4980 619 5014 795
rect 5098 619 5132 795
rect 7370 623 7404 799
rect 7488 623 7522 799
rect 7562 423 7596 799
rect 7680 423 7714 799
rect 7798 423 7832 799
rect 7916 423 7950 799
rect 8034 423 8068 799
rect 8112 623 8146 799
rect 8230 623 8264 799
rect 10514 623 10548 799
rect 10632 623 10666 799
rect 10706 423 10740 799
rect 10824 423 10858 799
rect 10942 423 10976 799
rect 11060 423 11094 799
rect 11178 423 11212 799
rect 11256 623 11290 799
rect 11374 623 11408 799
rect 13716 619 13750 795
rect 13834 619 13868 795
rect 13908 419 13942 795
rect 14026 419 14060 795
rect 14144 419 14178 795
rect 14262 419 14296 795
rect 14380 419 14414 795
rect 14458 619 14492 795
rect 14576 619 14610 795
rect 16860 619 16894 795
rect 16978 619 17012 795
rect 17052 419 17086 795
rect 17170 419 17204 795
rect 17288 419 17322 795
rect 17406 419 17440 795
rect 17524 419 17558 795
rect 17602 619 17636 795
rect 17720 619 17754 795
rect 19992 623 20026 799
rect 20110 623 20144 799
rect 20184 423 20218 799
rect 20302 423 20336 799
rect 20420 423 20454 799
rect 20538 423 20572 799
rect 20656 423 20690 799
rect 20734 623 20768 799
rect 20852 623 20886 799
rect 23136 623 23170 799
rect 23254 623 23288 799
rect 23328 423 23362 799
rect 23446 423 23480 799
rect 23564 423 23598 799
rect 23682 423 23716 799
rect 23800 423 23834 799
rect 23878 623 23912 799
rect 23996 623 24030 799
rect 1126 -3273 1160 -3097
rect 1244 -3273 1278 -3097
rect 1318 -3473 1352 -3097
rect 1436 -3473 1470 -3097
rect 1554 -3473 1588 -3097
rect 1672 -3473 1706 -3097
rect 1790 -3473 1824 -3097
rect 1868 -3273 1902 -3097
rect 1986 -3273 2020 -3097
rect 4270 -3273 4304 -3097
rect 4388 -3273 4422 -3097
rect 4462 -3473 4496 -3097
rect 4580 -3473 4614 -3097
rect 4698 -3473 4732 -3097
rect 4816 -3473 4850 -3097
rect 4934 -3473 4968 -3097
rect 5012 -3273 5046 -3097
rect 5130 -3273 5164 -3097
rect 7402 -3269 7436 -3093
rect 7520 -3269 7554 -3093
rect 7594 -3469 7628 -3093
rect 7712 -3469 7746 -3093
rect 7830 -3469 7864 -3093
rect 7948 -3469 7982 -3093
rect 8066 -3469 8100 -3093
rect 8144 -3269 8178 -3093
rect 8262 -3269 8296 -3093
rect 10546 -3269 10580 -3093
rect 10664 -3269 10698 -3093
rect 10738 -3469 10772 -3093
rect 10856 -3469 10890 -3093
rect 10974 -3469 11008 -3093
rect 11092 -3469 11126 -3093
rect 11210 -3469 11244 -3093
rect 11288 -3269 11322 -3093
rect 11406 -3269 11440 -3093
rect 13748 -3273 13782 -3097
rect 13866 -3273 13900 -3097
rect 13940 -3473 13974 -3097
rect 14058 -3473 14092 -3097
rect 14176 -3473 14210 -3097
rect 14294 -3473 14328 -3097
rect 14412 -3473 14446 -3097
rect 14490 -3273 14524 -3097
rect 14608 -3273 14642 -3097
rect 16892 -3273 16926 -3097
rect 17010 -3273 17044 -3097
rect 17084 -3473 17118 -3097
rect 17202 -3473 17236 -3097
rect 17320 -3473 17354 -3097
rect 17438 -3473 17472 -3097
rect 17556 -3473 17590 -3097
rect 17634 -3273 17668 -3097
rect 17752 -3273 17786 -3097
rect 20024 -3269 20058 -3093
rect 20142 -3269 20176 -3093
rect 20216 -3469 20250 -3093
rect 20334 -3469 20368 -3093
rect 20452 -3469 20486 -3093
rect 20570 -3469 20604 -3093
rect 20688 -3469 20722 -3093
rect 20766 -3269 20800 -3093
rect 20884 -3269 20918 -3093
rect 23168 -3269 23202 -3093
rect 23286 -3269 23320 -3093
rect 23360 -3469 23394 -3093
rect 23478 -3469 23512 -3093
rect 23596 -3469 23630 -3093
rect 23714 -3469 23748 -3093
rect 23832 -3469 23866 -3093
rect 23910 -3269 23944 -3093
rect 24028 -3269 24062 -3093
<< pdiffc >>
rect 466 21604 500 21780
rect 584 21604 618 21780
rect 702 21604 736 21780
rect 820 21604 854 21780
rect 907 21604 941 21980
rect 1025 21604 1059 21980
rect 1143 21604 1177 21980
rect 1261 21604 1295 21980
rect 1374 21604 1408 21980
rect 1492 21604 1526 21980
rect 1610 21604 1644 21980
rect 1728 21604 1762 21980
rect 1846 21604 1880 21980
rect 1964 21604 1998 21980
rect 2082 21604 2116 21980
rect 2201 21604 2235 21980
rect 2319 21604 2353 21980
rect 2437 21604 2471 21980
rect 2555 21604 2589 21980
rect 2674 21604 2708 21780
rect 2792 21604 2826 21780
rect 2910 21604 2944 21780
rect 3028 21604 3062 21780
rect 3610 21604 3644 21780
rect 3728 21604 3762 21780
rect 3846 21604 3880 21780
rect 3964 21604 3998 21780
rect 4051 21604 4085 21980
rect 4169 21604 4203 21980
rect 4287 21604 4321 21980
rect 4405 21604 4439 21980
rect 4518 21604 4552 21980
rect 4636 21604 4670 21980
rect 4754 21604 4788 21980
rect 4872 21604 4906 21980
rect 4990 21604 5024 21980
rect 5108 21604 5142 21980
rect 5226 21604 5260 21980
rect 5345 21604 5379 21980
rect 5463 21604 5497 21980
rect 5581 21604 5615 21980
rect 5699 21604 5733 21980
rect 5818 21604 5852 21780
rect 5936 21604 5970 21780
rect 6054 21604 6088 21780
rect 6172 21604 6206 21780
rect 6742 21608 6776 21784
rect 6860 21608 6894 21784
rect 6978 21608 7012 21784
rect 7096 21608 7130 21784
rect 7183 21608 7217 21984
rect 7301 21608 7335 21984
rect 7419 21608 7453 21984
rect 7537 21608 7571 21984
rect 7650 21608 7684 21984
rect 7768 21608 7802 21984
rect 7886 21608 7920 21984
rect 8004 21608 8038 21984
rect 8122 21608 8156 21984
rect 8240 21608 8274 21984
rect 8358 21608 8392 21984
rect 8477 21608 8511 21984
rect 8595 21608 8629 21984
rect 8713 21608 8747 21984
rect 8831 21608 8865 21984
rect 8950 21608 8984 21784
rect 9068 21608 9102 21784
rect 9186 21608 9220 21784
rect 9304 21608 9338 21784
rect 9886 21608 9920 21784
rect 10004 21608 10038 21784
rect 10122 21608 10156 21784
rect 10240 21608 10274 21784
rect 10327 21608 10361 21984
rect 10445 21608 10479 21984
rect 10563 21608 10597 21984
rect 10681 21608 10715 21984
rect 10794 21608 10828 21984
rect 10912 21608 10946 21984
rect 11030 21608 11064 21984
rect 11148 21608 11182 21984
rect 11266 21608 11300 21984
rect 11384 21608 11418 21984
rect 11502 21608 11536 21984
rect 11621 21608 11655 21984
rect 11739 21608 11773 21984
rect 11857 21608 11891 21984
rect 11975 21608 12009 21984
rect 12094 21608 12128 21784
rect 12212 21608 12246 21784
rect 12330 21608 12364 21784
rect 12448 21608 12482 21784
rect 13088 21604 13122 21780
rect 13206 21604 13240 21780
rect 13324 21604 13358 21780
rect 13442 21604 13476 21780
rect 13529 21604 13563 21980
rect 13647 21604 13681 21980
rect 13765 21604 13799 21980
rect 13883 21604 13917 21980
rect 13996 21604 14030 21980
rect 14114 21604 14148 21980
rect 14232 21604 14266 21980
rect 14350 21604 14384 21980
rect 14468 21604 14502 21980
rect 14586 21604 14620 21980
rect 14704 21604 14738 21980
rect 14823 21604 14857 21980
rect 14941 21604 14975 21980
rect 15059 21604 15093 21980
rect 15177 21604 15211 21980
rect 15296 21604 15330 21780
rect 15414 21604 15448 21780
rect 15532 21604 15566 21780
rect 15650 21604 15684 21780
rect 16232 21604 16266 21780
rect 16350 21604 16384 21780
rect 16468 21604 16502 21780
rect 16586 21604 16620 21780
rect 16673 21604 16707 21980
rect 16791 21604 16825 21980
rect 16909 21604 16943 21980
rect 17027 21604 17061 21980
rect 17140 21604 17174 21980
rect 17258 21604 17292 21980
rect 17376 21604 17410 21980
rect 17494 21604 17528 21980
rect 17612 21604 17646 21980
rect 17730 21604 17764 21980
rect 17848 21604 17882 21980
rect 17967 21604 18001 21980
rect 18085 21604 18119 21980
rect 18203 21604 18237 21980
rect 18321 21604 18355 21980
rect 18440 21604 18474 21780
rect 18558 21604 18592 21780
rect 18676 21604 18710 21780
rect 18794 21604 18828 21780
rect 19364 21608 19398 21784
rect 19482 21608 19516 21784
rect 19600 21608 19634 21784
rect 19718 21608 19752 21784
rect 19805 21608 19839 21984
rect 19923 21608 19957 21984
rect 20041 21608 20075 21984
rect 20159 21608 20193 21984
rect 20272 21608 20306 21984
rect 20390 21608 20424 21984
rect 20508 21608 20542 21984
rect 20626 21608 20660 21984
rect 20744 21608 20778 21984
rect 20862 21608 20896 21984
rect 20980 21608 21014 21984
rect 21099 21608 21133 21984
rect 21217 21608 21251 21984
rect 21335 21608 21369 21984
rect 21453 21608 21487 21984
rect 21572 21608 21606 21784
rect 21690 21608 21724 21784
rect 21808 21608 21842 21784
rect 21926 21608 21960 21784
rect 22508 21608 22542 21784
rect 22626 21608 22660 21784
rect 22744 21608 22778 21784
rect 22862 21608 22896 21784
rect 22949 21608 22983 21984
rect 23067 21608 23101 21984
rect 23185 21608 23219 21984
rect 23303 21608 23337 21984
rect 23416 21608 23450 21984
rect 23534 21608 23568 21984
rect 23652 21608 23686 21984
rect 23770 21608 23804 21984
rect 23888 21608 23922 21984
rect 24006 21608 24040 21984
rect 24124 21608 24158 21984
rect 24243 21608 24277 21984
rect 24361 21608 24395 21984
rect 24479 21608 24513 21984
rect 24597 21608 24631 21984
rect 24716 21608 24750 21784
rect 24834 21608 24868 21784
rect 24952 21608 24986 21784
rect 25070 21608 25104 21784
rect 2909 16423 2943 16599
rect 3027 16423 3061 16599
rect 3145 16423 3179 16599
rect 3263 16423 3297 16599
rect 3381 16423 3415 16599
rect 3499 16423 3533 16599
rect 3617 16423 3651 16599
rect 3735 16423 3769 16599
rect 3853 16423 3887 16599
rect 3971 16423 4005 16599
rect 4357 16423 4391 16599
rect 4475 16423 4509 16599
rect 4593 16423 4627 16599
rect 4711 16423 4745 16599
rect 4829 16423 4863 16599
rect 4947 16423 4981 16599
rect 5065 16423 5099 16599
rect 5183 16423 5217 16599
rect 5301 16423 5335 16599
rect 5419 16423 5453 16599
rect 5855 16425 5889 16601
rect 5973 16425 6007 16601
rect 6091 16425 6125 16601
rect 6209 16425 6243 16601
rect 6327 16425 6361 16601
rect 6445 16425 6479 16601
rect 6563 16425 6597 16601
rect 6681 16425 6715 16601
rect 6799 16425 6833 16601
rect 6917 16425 6951 16601
rect 7303 16425 7337 16601
rect 7421 16425 7455 16601
rect 7539 16425 7573 16601
rect 7657 16425 7691 16601
rect 7775 16425 7809 16601
rect 7893 16425 7927 16601
rect 8011 16425 8045 16601
rect 8129 16425 8163 16601
rect 8247 16425 8281 16601
rect 8365 16425 8399 16601
rect 8823 16423 8857 16599
rect 8941 16423 8975 16599
rect 9059 16423 9093 16599
rect 9177 16423 9211 16599
rect 9295 16423 9329 16599
rect 9413 16423 9447 16599
rect 9531 16423 9565 16599
rect 9649 16423 9683 16599
rect 9767 16423 9801 16599
rect 9885 16423 9919 16599
rect 10271 16423 10305 16599
rect 10389 16423 10423 16599
rect 10507 16423 10541 16599
rect 10625 16423 10659 16599
rect 10743 16423 10777 16599
rect 10861 16423 10895 16599
rect 10979 16423 11013 16599
rect 11097 16423 11131 16599
rect 11215 16423 11249 16599
rect 11333 16423 11367 16599
rect 11769 16425 11803 16601
rect 11887 16425 11921 16601
rect 12005 16425 12039 16601
rect 12123 16425 12157 16601
rect 12241 16425 12275 16601
rect 12359 16425 12393 16601
rect 12477 16425 12511 16601
rect 12595 16425 12629 16601
rect 12713 16425 12747 16601
rect 12831 16425 12865 16601
rect 13217 16425 13251 16601
rect 13335 16425 13369 16601
rect 13453 16425 13487 16601
rect 13571 16425 13605 16601
rect 13689 16425 13723 16601
rect 13807 16425 13841 16601
rect 13925 16425 13959 16601
rect 14043 16425 14077 16601
rect 14161 16425 14195 16601
rect 14279 16425 14313 16601
rect 14672 16420 14706 16796
rect 14790 16420 14824 16796
rect 14908 16420 14942 16796
rect 15026 16420 15060 16796
rect 15144 16420 15178 16796
rect 15262 16420 15296 16796
rect 15380 16420 15414 16796
rect 15840 16420 15874 16796
rect 15958 16420 15992 16796
rect 16076 16420 16110 16796
rect 16194 16420 16228 16796
rect 16312 16420 16346 16796
rect 16430 16420 16464 16796
rect 16548 16420 16582 16796
rect 17008 16418 17042 16794
rect 17126 16418 17160 16794
rect 17244 16418 17278 16794
rect 17362 16418 17396 16794
rect 17480 16418 17514 16794
rect 17598 16418 17632 16794
rect 17716 16418 17750 16794
rect 18176 16420 18210 16796
rect 18294 16420 18328 16796
rect 18412 16420 18446 16796
rect 18530 16420 18564 16796
rect 18648 16420 18682 16796
rect 18766 16420 18800 16796
rect 18884 16420 18918 16796
rect 19350 16422 19384 16798
rect 19468 16422 19502 16798
rect 19586 16422 19620 16798
rect 19704 16422 19738 16798
rect 19822 16422 19856 16798
rect 19940 16422 19974 16798
rect 20058 16422 20092 16798
rect 20518 16420 20552 16796
rect 20636 16420 20670 16796
rect 20754 16420 20788 16796
rect 20872 16420 20906 16796
rect 20990 16420 21024 16796
rect 21108 16420 21142 16796
rect 21226 16420 21260 16796
rect 21686 16422 21720 16798
rect 21804 16422 21838 16798
rect 21922 16422 21956 16798
rect 22040 16422 22074 16798
rect 22158 16422 22192 16798
rect 22276 16422 22310 16798
rect 22394 16422 22428 16798
rect 22854 16420 22888 16796
rect 15102 15830 15136 16006
rect 15220 15830 15254 16006
rect 15338 15830 15372 16006
rect 15456 15830 15490 16006
rect 16269 15836 16303 16012
rect 16387 15836 16421 16012
rect 16505 15836 16539 16012
rect 16623 15836 16657 16012
rect 17437 15836 17471 16012
rect 17555 15836 17589 16012
rect 17673 15836 17707 16012
rect 17791 15836 17825 16012
rect 18606 15836 18640 16012
rect 18724 15836 18758 16012
rect 18842 15836 18876 16012
rect 18960 15836 18994 16012
rect 19778 15832 19812 16008
rect 19896 15832 19930 16008
rect 20014 15832 20048 16008
rect 20132 15832 20166 16008
rect 22972 16420 23006 16796
rect 23090 16420 23124 16796
rect 23208 16420 23242 16796
rect 23326 16420 23360 16796
rect 23444 16420 23478 16796
rect 23562 16420 23596 16796
rect 20947 15831 20981 16007
rect 21065 15831 21099 16007
rect 21183 15831 21217 16007
rect 21301 15831 21335 16007
rect 22115 15831 22149 16007
rect 22233 15831 22267 16007
rect 22351 15831 22385 16007
rect 22469 15831 22503 16007
rect 23283 15832 23317 16008
rect 23401 15832 23435 16008
rect 23519 15832 23553 16008
rect 23637 15832 23671 16008
rect 2968 14466 3002 14642
rect 3086 14466 3120 14642
rect 3204 14466 3238 14642
rect 3322 14466 3356 14642
rect 3409 14466 3443 14842
rect 3527 14466 3561 14842
rect 3645 14466 3679 14842
rect 3763 14466 3797 14842
rect 3876 14466 3910 14842
rect 3994 14466 4028 14842
rect 4112 14466 4146 14842
rect 4230 14466 4264 14842
rect 4348 14466 4382 14842
rect 4466 14466 4500 14842
rect 4584 14466 4618 14842
rect 4703 14466 4737 14842
rect 4821 14466 4855 14842
rect 4939 14466 4973 14842
rect 5057 14466 5091 14842
rect 5176 14466 5210 14642
rect 5294 14466 5328 14642
rect 5412 14466 5446 14642
rect 5530 14466 5564 14642
rect 6112 14466 6146 14642
rect 6230 14466 6264 14642
rect 6348 14466 6382 14642
rect 6466 14466 6500 14642
rect 6553 14466 6587 14842
rect 6671 14466 6705 14842
rect 6789 14466 6823 14842
rect 6907 14466 6941 14842
rect 7020 14466 7054 14842
rect 7138 14466 7172 14842
rect 7256 14466 7290 14842
rect 7374 14466 7408 14842
rect 7492 14466 7526 14842
rect 7610 14466 7644 14842
rect 7728 14466 7762 14842
rect 7847 14466 7881 14842
rect 7965 14466 7999 14842
rect 8083 14466 8117 14842
rect 8201 14466 8235 14842
rect 8320 14466 8354 14642
rect 8438 14466 8472 14642
rect 8556 14466 8590 14642
rect 8674 14466 8708 14642
rect 9244 14470 9278 14646
rect 9362 14470 9396 14646
rect 9480 14470 9514 14646
rect 9598 14470 9632 14646
rect 9685 14470 9719 14846
rect 9803 14470 9837 14846
rect 9921 14470 9955 14846
rect 10039 14470 10073 14846
rect 10152 14470 10186 14846
rect 10270 14470 10304 14846
rect 10388 14470 10422 14846
rect 10506 14470 10540 14846
rect 10624 14470 10658 14846
rect 10742 14470 10776 14846
rect 10860 14470 10894 14846
rect 10979 14470 11013 14846
rect 11097 14470 11131 14846
rect 11215 14470 11249 14846
rect 11333 14470 11367 14846
rect 11452 14470 11486 14646
rect 11570 14470 11604 14646
rect 11688 14470 11722 14646
rect 11806 14470 11840 14646
rect 12388 14470 12422 14646
rect 12506 14470 12540 14646
rect 12624 14470 12658 14646
rect 12742 14470 12776 14646
rect 12829 14470 12863 14846
rect 12947 14470 12981 14846
rect 13065 14470 13099 14846
rect 13183 14470 13217 14846
rect 13296 14470 13330 14846
rect 13414 14470 13448 14846
rect 13532 14470 13566 14846
rect 13650 14470 13684 14846
rect 13768 14470 13802 14846
rect 13886 14470 13920 14846
rect 14004 14470 14038 14846
rect 14123 14470 14157 14846
rect 14241 14470 14275 14846
rect 14359 14470 14393 14846
rect 14477 14470 14511 14846
rect 14596 14470 14630 14646
rect 14714 14470 14748 14646
rect 14832 14470 14866 14646
rect 14950 14470 14984 14646
rect 15590 14466 15624 14642
rect 15708 14466 15742 14642
rect 15826 14466 15860 14642
rect 15944 14466 15978 14642
rect 16031 14466 16065 14842
rect 16149 14466 16183 14842
rect 16267 14466 16301 14842
rect 16385 14466 16419 14842
rect 16498 14466 16532 14842
rect 16616 14466 16650 14842
rect 16734 14466 16768 14842
rect 16852 14466 16886 14842
rect 16970 14466 17004 14842
rect 17088 14466 17122 14842
rect 17206 14466 17240 14842
rect 17325 14466 17359 14842
rect 17443 14466 17477 14842
rect 17561 14466 17595 14842
rect 17679 14466 17713 14842
rect 17798 14466 17832 14642
rect 17916 14466 17950 14642
rect 18034 14466 18068 14642
rect 18152 14466 18186 14642
rect 18734 14466 18768 14642
rect 18852 14466 18886 14642
rect 18970 14466 19004 14642
rect 19088 14466 19122 14642
rect 19175 14466 19209 14842
rect 19293 14466 19327 14842
rect 19411 14466 19445 14842
rect 19529 14466 19563 14842
rect 19642 14466 19676 14842
rect 19760 14466 19794 14842
rect 19878 14466 19912 14842
rect 19996 14466 20030 14842
rect 20114 14466 20148 14842
rect 20232 14466 20266 14842
rect 20350 14466 20384 14842
rect 20469 14466 20503 14842
rect 20587 14466 20621 14842
rect 20705 14466 20739 14842
rect 20823 14466 20857 14842
rect 20942 14466 20976 14642
rect 21060 14466 21094 14642
rect 21178 14466 21212 14642
rect 21296 14466 21330 14642
rect 21866 14470 21900 14646
rect 21984 14470 22018 14646
rect 22102 14470 22136 14646
rect 22220 14470 22254 14646
rect 22307 14470 22341 14846
rect 22425 14470 22459 14846
rect 22543 14470 22577 14846
rect 22661 14470 22695 14846
rect 22774 14470 22808 14846
rect 22892 14470 22926 14846
rect 23010 14470 23044 14846
rect 23128 14470 23162 14846
rect 23246 14470 23280 14846
rect 23364 14470 23398 14846
rect 23482 14470 23516 14846
rect 23601 14470 23635 14846
rect 23719 14470 23753 14846
rect 23837 14470 23871 14846
rect 23955 14470 23989 14846
rect 24074 14470 24108 14646
rect 24192 14470 24226 14646
rect 24310 14470 24344 14646
rect 24428 14470 24462 14646
rect 25010 14470 25044 14646
rect 25128 14470 25162 14646
rect 25246 14470 25280 14646
rect 25364 14470 25398 14646
rect 25451 14470 25485 14846
rect 25569 14470 25603 14846
rect 25687 14470 25721 14846
rect 25805 14470 25839 14846
rect 25918 14470 25952 14846
rect 26036 14470 26070 14846
rect 26154 14470 26188 14846
rect 26272 14470 26306 14846
rect 26390 14470 26424 14846
rect 26508 14470 26542 14846
rect 26626 14470 26660 14846
rect 26745 14470 26779 14846
rect 26863 14470 26897 14846
rect 26981 14470 27015 14846
rect 27099 14470 27133 14846
rect 27218 14470 27252 14646
rect 27336 14470 27370 14646
rect 27454 14470 27488 14646
rect 27572 14470 27606 14646
rect 2968 11732 3002 11908
rect 3086 11732 3120 11908
rect 3204 11732 3238 11908
rect 3322 11732 3356 11908
rect 3409 11732 3443 12108
rect 3527 11732 3561 12108
rect 3645 11732 3679 12108
rect 3763 11732 3797 12108
rect 3876 11732 3910 12108
rect 3994 11732 4028 12108
rect 4112 11732 4146 12108
rect 4230 11732 4264 12108
rect 4348 11732 4382 12108
rect 4466 11732 4500 12108
rect 4584 11732 4618 12108
rect 4703 11732 4737 12108
rect 4821 11732 4855 12108
rect 4939 11732 4973 12108
rect 5057 11732 5091 12108
rect 5176 11732 5210 11908
rect 5294 11732 5328 11908
rect 5412 11732 5446 11908
rect 5530 11732 5564 11908
rect 6112 11732 6146 11908
rect 6230 11732 6264 11908
rect 6348 11732 6382 11908
rect 6466 11732 6500 11908
rect 6553 11732 6587 12108
rect 6671 11732 6705 12108
rect 6789 11732 6823 12108
rect 6907 11732 6941 12108
rect 7020 11732 7054 12108
rect 7138 11732 7172 12108
rect 7256 11732 7290 12108
rect 7374 11732 7408 12108
rect 7492 11732 7526 12108
rect 7610 11732 7644 12108
rect 7728 11732 7762 12108
rect 7847 11732 7881 12108
rect 7965 11732 7999 12108
rect 8083 11732 8117 12108
rect 8201 11732 8235 12108
rect 8320 11732 8354 11908
rect 8438 11732 8472 11908
rect 8556 11732 8590 11908
rect 8674 11732 8708 11908
rect 9244 11736 9278 11912
rect 9362 11736 9396 11912
rect 9480 11736 9514 11912
rect 9598 11736 9632 11912
rect 9685 11736 9719 12112
rect 9803 11736 9837 12112
rect 9921 11736 9955 12112
rect 10039 11736 10073 12112
rect 10152 11736 10186 12112
rect 10270 11736 10304 12112
rect 10388 11736 10422 12112
rect 10506 11736 10540 12112
rect 10624 11736 10658 12112
rect 10742 11736 10776 12112
rect 10860 11736 10894 12112
rect 10979 11736 11013 12112
rect 11097 11736 11131 12112
rect 11215 11736 11249 12112
rect 11333 11736 11367 12112
rect 11452 11736 11486 11912
rect 11570 11736 11604 11912
rect 11688 11736 11722 11912
rect 11806 11736 11840 11912
rect 12388 11736 12422 11912
rect 12506 11736 12540 11912
rect 12624 11736 12658 11912
rect 12742 11736 12776 11912
rect 12829 11736 12863 12112
rect 12947 11736 12981 12112
rect 13065 11736 13099 12112
rect 13183 11736 13217 12112
rect 13296 11736 13330 12112
rect 13414 11736 13448 12112
rect 13532 11736 13566 12112
rect 13650 11736 13684 12112
rect 13768 11736 13802 12112
rect 13886 11736 13920 12112
rect 14004 11736 14038 12112
rect 14123 11736 14157 12112
rect 14241 11736 14275 12112
rect 14359 11736 14393 12112
rect 14477 11736 14511 12112
rect 14596 11736 14630 11912
rect 14714 11736 14748 11912
rect 14832 11736 14866 11912
rect 14950 11736 14984 11912
rect 15590 11732 15624 11908
rect 15708 11732 15742 11908
rect 15826 11732 15860 11908
rect 15944 11732 15978 11908
rect 16031 11732 16065 12108
rect 16149 11732 16183 12108
rect 16267 11732 16301 12108
rect 16385 11732 16419 12108
rect 16498 11732 16532 12108
rect 16616 11732 16650 12108
rect 16734 11732 16768 12108
rect 16852 11732 16886 12108
rect 16970 11732 17004 12108
rect 17088 11732 17122 12108
rect 17206 11732 17240 12108
rect 17325 11732 17359 12108
rect 17443 11732 17477 12108
rect 17561 11732 17595 12108
rect 17679 11732 17713 12108
rect 17798 11732 17832 11908
rect 17916 11732 17950 11908
rect 18034 11732 18068 11908
rect 18152 11732 18186 11908
rect 18734 11732 18768 11908
rect 18852 11732 18886 11908
rect 18970 11732 19004 11908
rect 19088 11732 19122 11908
rect 19175 11732 19209 12108
rect 19293 11732 19327 12108
rect 19411 11732 19445 12108
rect 19529 11732 19563 12108
rect 19642 11732 19676 12108
rect 19760 11732 19794 12108
rect 19878 11732 19912 12108
rect 19996 11732 20030 12108
rect 20114 11732 20148 12108
rect 20232 11732 20266 12108
rect 20350 11732 20384 12108
rect 20469 11732 20503 12108
rect 20587 11732 20621 12108
rect 20705 11732 20739 12108
rect 20823 11732 20857 12108
rect 20942 11732 20976 11908
rect 21060 11732 21094 11908
rect 21178 11732 21212 11908
rect 21296 11732 21330 11908
rect 21866 11736 21900 11912
rect 21984 11736 22018 11912
rect 22102 11736 22136 11912
rect 22220 11736 22254 11912
rect 22307 11736 22341 12112
rect 22425 11736 22459 12112
rect 22543 11736 22577 12112
rect 22661 11736 22695 12112
rect 22774 11736 22808 12112
rect 22892 11736 22926 12112
rect 23010 11736 23044 12112
rect 23128 11736 23162 12112
rect 23246 11736 23280 12112
rect 23364 11736 23398 12112
rect 23482 11736 23516 12112
rect 23601 11736 23635 12112
rect 23719 11736 23753 12112
rect 23837 11736 23871 12112
rect 23955 11736 23989 12112
rect 24074 11736 24108 11912
rect 24192 11736 24226 11912
rect 24310 11736 24344 11912
rect 24428 11736 24462 11912
rect 25010 11736 25044 11912
rect 25128 11736 25162 11912
rect 25246 11736 25280 11912
rect 25364 11736 25398 11912
rect 25451 11736 25485 12112
rect 25569 11736 25603 12112
rect 25687 11736 25721 12112
rect 25805 11736 25839 12112
rect 25918 11736 25952 12112
rect 26036 11736 26070 12112
rect 26154 11736 26188 12112
rect 26272 11736 26306 12112
rect 26390 11736 26424 12112
rect 26508 11736 26542 12112
rect 26626 11736 26660 12112
rect 26745 11736 26779 12112
rect 26863 11736 26897 12112
rect 26981 11736 27015 12112
rect 27099 11736 27133 12112
rect 27218 11736 27252 11912
rect 27336 11736 27370 11912
rect 27454 11736 27488 11912
rect 27572 11736 27606 11912
rect 2958 9000 2992 9176
rect 3076 9000 3110 9176
rect 3194 9000 3228 9176
rect 3312 9000 3346 9176
rect 3399 9000 3433 9376
rect 3517 9000 3551 9376
rect 3635 9000 3669 9376
rect 3753 9000 3787 9376
rect 3866 9000 3900 9376
rect 3984 9000 4018 9376
rect 4102 9000 4136 9376
rect 4220 9000 4254 9376
rect 4338 9000 4372 9376
rect 4456 9000 4490 9376
rect 4574 9000 4608 9376
rect 4693 9000 4727 9376
rect 4811 9000 4845 9376
rect 4929 9000 4963 9376
rect 5047 9000 5081 9376
rect 5166 9000 5200 9176
rect 5284 9000 5318 9176
rect 5402 9000 5436 9176
rect 5520 9000 5554 9176
rect 6102 9000 6136 9176
rect 6220 9000 6254 9176
rect 6338 9000 6372 9176
rect 6456 9000 6490 9176
rect 6543 9000 6577 9376
rect 6661 9000 6695 9376
rect 6779 9000 6813 9376
rect 6897 9000 6931 9376
rect 7010 9000 7044 9376
rect 7128 9000 7162 9376
rect 7246 9000 7280 9376
rect 7364 9000 7398 9376
rect 7482 9000 7516 9376
rect 7600 9000 7634 9376
rect 7718 9000 7752 9376
rect 7837 9000 7871 9376
rect 7955 9000 7989 9376
rect 8073 9000 8107 9376
rect 8191 9000 8225 9376
rect 8310 9000 8344 9176
rect 8428 9000 8462 9176
rect 8546 9000 8580 9176
rect 8664 9000 8698 9176
rect 9234 9004 9268 9180
rect 9352 9004 9386 9180
rect 9470 9004 9504 9180
rect 9588 9004 9622 9180
rect 9675 9004 9709 9380
rect 9793 9004 9827 9380
rect 9911 9004 9945 9380
rect 10029 9004 10063 9380
rect 10142 9004 10176 9380
rect 10260 9004 10294 9380
rect 10378 9004 10412 9380
rect 10496 9004 10530 9380
rect 10614 9004 10648 9380
rect 10732 9004 10766 9380
rect 10850 9004 10884 9380
rect 10969 9004 11003 9380
rect 11087 9004 11121 9380
rect 11205 9004 11239 9380
rect 11323 9004 11357 9380
rect 11442 9004 11476 9180
rect 11560 9004 11594 9180
rect 11678 9004 11712 9180
rect 11796 9004 11830 9180
rect 12378 9004 12412 9180
rect 12496 9004 12530 9180
rect 12614 9004 12648 9180
rect 12732 9004 12766 9180
rect 12819 9004 12853 9380
rect 12937 9004 12971 9380
rect 13055 9004 13089 9380
rect 13173 9004 13207 9380
rect 13286 9004 13320 9380
rect 13404 9004 13438 9380
rect 13522 9004 13556 9380
rect 13640 9004 13674 9380
rect 13758 9004 13792 9380
rect 13876 9004 13910 9380
rect 13994 9004 14028 9380
rect 14113 9004 14147 9380
rect 14231 9004 14265 9380
rect 14349 9004 14383 9380
rect 14467 9004 14501 9380
rect 14586 9004 14620 9180
rect 14704 9004 14738 9180
rect 14822 9004 14856 9180
rect 14940 9004 14974 9180
rect 15580 9000 15614 9176
rect 15698 9000 15732 9176
rect 15816 9000 15850 9176
rect 15934 9000 15968 9176
rect 16021 9000 16055 9376
rect 16139 9000 16173 9376
rect 16257 9000 16291 9376
rect 16375 9000 16409 9376
rect 16488 9000 16522 9376
rect 16606 9000 16640 9376
rect 16724 9000 16758 9376
rect 16842 9000 16876 9376
rect 16960 9000 16994 9376
rect 17078 9000 17112 9376
rect 17196 9000 17230 9376
rect 17315 9000 17349 9376
rect 17433 9000 17467 9376
rect 17551 9000 17585 9376
rect 17669 9000 17703 9376
rect 17788 9000 17822 9176
rect 17906 9000 17940 9176
rect 18024 9000 18058 9176
rect 18142 9000 18176 9176
rect 18724 9000 18758 9176
rect 18842 9000 18876 9176
rect 18960 9000 18994 9176
rect 19078 9000 19112 9176
rect 19165 9000 19199 9376
rect 19283 9000 19317 9376
rect 19401 9000 19435 9376
rect 19519 9000 19553 9376
rect 19632 9000 19666 9376
rect 19750 9000 19784 9376
rect 19868 9000 19902 9376
rect 19986 9000 20020 9376
rect 20104 9000 20138 9376
rect 20222 9000 20256 9376
rect 20340 9000 20374 9376
rect 20459 9000 20493 9376
rect 20577 9000 20611 9376
rect 20695 9000 20729 9376
rect 20813 9000 20847 9376
rect 20932 9000 20966 9176
rect 21050 9000 21084 9176
rect 21168 9000 21202 9176
rect 21286 9000 21320 9176
rect 21856 9004 21890 9180
rect 21974 9004 22008 9180
rect 22092 9004 22126 9180
rect 22210 9004 22244 9180
rect 22297 9004 22331 9380
rect 22415 9004 22449 9380
rect 22533 9004 22567 9380
rect 22651 9004 22685 9380
rect 22764 9004 22798 9380
rect 22882 9004 22916 9380
rect 23000 9004 23034 9380
rect 23118 9004 23152 9380
rect 23236 9004 23270 9380
rect 23354 9004 23388 9380
rect 23472 9004 23506 9380
rect 23591 9004 23625 9380
rect 23709 9004 23743 9380
rect 23827 9004 23861 9380
rect 23945 9004 23979 9380
rect 24064 9004 24098 9180
rect 24182 9004 24216 9180
rect 24300 9004 24334 9180
rect 24418 9004 24452 9180
rect 25000 9004 25034 9180
rect 25118 9004 25152 9180
rect 25236 9004 25270 9180
rect 25354 9004 25388 9180
rect 25441 9004 25475 9380
rect 25559 9004 25593 9380
rect 25677 9004 25711 9380
rect 25795 9004 25829 9380
rect 25908 9004 25942 9380
rect 26026 9004 26060 9380
rect 26144 9004 26178 9380
rect 26262 9004 26296 9380
rect 26380 9004 26414 9380
rect 26498 9004 26532 9380
rect 26616 9004 26650 9380
rect 26735 9004 26769 9380
rect 26853 9004 26887 9380
rect 26971 9004 27005 9380
rect 27089 9004 27123 9380
rect 27208 9004 27242 9180
rect 27326 9004 27360 9180
rect 27444 9004 27478 9180
rect 27562 9004 27596 9180
rect 2695 6055 2729 6231
rect 2813 6055 2847 6231
rect 2931 6055 2965 6231
rect 3049 6055 3083 6231
rect 3179 6055 3213 6431
rect 3297 6055 3331 6431
rect 3415 6055 3449 6431
rect 3533 6055 3567 6431
rect 3651 6055 3685 6431
rect 3769 6055 3803 6431
rect 3887 6055 3921 6431
rect 4016 6055 4050 6231
rect 4134 6055 4168 6231
rect 4252 6055 4286 6231
rect 4370 6055 4404 6231
rect 4763 6057 4797 6233
rect 4881 6057 4915 6233
rect 4999 6057 5033 6233
rect 5117 6057 5151 6233
rect 5247 6057 5281 6433
rect 5365 6057 5399 6433
rect 5483 6057 5517 6433
rect 5601 6057 5635 6433
rect 5719 6057 5753 6433
rect 5837 6057 5871 6433
rect 5955 6057 5989 6433
rect 6084 6057 6118 6233
rect 6202 6057 6236 6233
rect 6320 6057 6354 6233
rect 6438 6057 6472 6233
rect 6832 6055 6866 6231
rect 3122 5362 3156 5738
rect 3240 5362 3274 5738
rect 3358 5362 3392 5738
rect 3476 5362 3510 5738
rect 3594 5362 3628 5738
rect 3712 5362 3746 5738
rect 3830 5362 3864 5738
rect 6950 6055 6984 6231
rect 7068 6055 7102 6231
rect 7186 6055 7220 6231
rect 7316 6055 7350 6431
rect 7434 6055 7468 6431
rect 7552 6055 7586 6431
rect 7670 6055 7704 6431
rect 7788 6055 7822 6431
rect 7906 6055 7940 6431
rect 8024 6055 8058 6431
rect 8153 6055 8187 6231
rect 8271 6055 8305 6231
rect 8389 6055 8423 6231
rect 8507 6055 8541 6231
rect 8900 6057 8934 6233
rect 9018 6057 9052 6233
rect 9136 6057 9170 6233
rect 9254 6057 9288 6233
rect 9384 6057 9418 6433
rect 9502 6057 9536 6433
rect 9620 6057 9654 6433
rect 9738 6057 9772 6433
rect 9856 6057 9890 6433
rect 9974 6057 10008 6433
rect 10092 6057 10126 6433
rect 10221 6057 10255 6233
rect 10339 6057 10373 6233
rect 10457 6057 10491 6233
rect 10575 6057 10609 6233
rect 10969 6057 11003 6233
rect 11087 6057 11121 6233
rect 11205 6057 11239 6233
rect 11323 6057 11357 6233
rect 11453 6057 11487 6433
rect 11571 6057 11605 6433
rect 11689 6057 11723 6433
rect 11807 6057 11841 6433
rect 11925 6057 11959 6433
rect 12043 6057 12077 6433
rect 12161 6057 12195 6433
rect 12290 6057 12324 6233
rect 12408 6057 12442 6233
rect 12526 6057 12560 6233
rect 12644 6057 12678 6233
rect 13037 6059 13071 6235
rect 13155 6059 13189 6235
rect 13273 6059 13307 6235
rect 13391 6059 13425 6235
rect 13521 6059 13555 6435
rect 13639 6059 13673 6435
rect 13757 6059 13791 6435
rect 13875 6059 13909 6435
rect 13993 6059 14027 6435
rect 14111 6059 14145 6435
rect 14229 6059 14263 6435
rect 14358 6059 14392 6235
rect 14476 6059 14510 6235
rect 14594 6059 14628 6235
rect 14712 6059 14746 6235
rect 15106 6057 15140 6233
rect 5190 5364 5224 5740
rect 5308 5364 5342 5740
rect 5426 5364 5460 5740
rect 5544 5364 5578 5740
rect 5662 5364 5696 5740
rect 5780 5364 5814 5740
rect 5898 5364 5932 5740
rect 7259 5362 7293 5738
rect 7377 5362 7411 5738
rect 7495 5362 7529 5738
rect 7613 5362 7647 5738
rect 7731 5362 7765 5738
rect 7849 5362 7883 5738
rect 7967 5362 8001 5738
rect 9327 5364 9361 5740
rect 9445 5364 9479 5740
rect 9563 5364 9597 5740
rect 9681 5364 9715 5740
rect 9799 5364 9833 5740
rect 9917 5364 9951 5740
rect 10035 5364 10069 5740
rect 11396 5364 11430 5740
rect 11514 5364 11548 5740
rect 11632 5364 11666 5740
rect 11750 5364 11784 5740
rect 11868 5364 11902 5740
rect 11986 5364 12020 5740
rect 12104 5364 12138 5740
rect 15224 6057 15258 6233
rect 15342 6057 15376 6233
rect 15460 6057 15494 6233
rect 15590 6057 15624 6433
rect 15708 6057 15742 6433
rect 15826 6057 15860 6433
rect 15944 6057 15978 6433
rect 16062 6057 16096 6433
rect 16180 6057 16214 6433
rect 16298 6057 16332 6433
rect 16427 6057 16461 6233
rect 16545 6057 16579 6233
rect 16663 6057 16697 6233
rect 16781 6057 16815 6233
rect 17174 6059 17208 6235
rect 17292 6059 17326 6235
rect 17410 6059 17444 6235
rect 17528 6059 17562 6235
rect 17658 6059 17692 6435
rect 17776 6059 17810 6435
rect 17894 6059 17928 6435
rect 18012 6059 18046 6435
rect 18130 6059 18164 6435
rect 18248 6059 18282 6435
rect 18366 6059 18400 6435
rect 19427 6371 19461 6547
rect 19545 6371 19579 6547
rect 19663 6371 19697 6547
rect 19781 6371 19815 6547
rect 20165 6375 20199 6551
rect 20283 6375 20317 6551
rect 20401 6375 20435 6551
rect 20519 6375 20553 6551
rect 20903 6371 20937 6547
rect 21021 6371 21055 6547
rect 21139 6371 21173 6547
rect 21257 6371 21291 6547
rect 21645 6369 21679 6545
rect 21763 6369 21797 6545
rect 21881 6369 21915 6545
rect 21999 6369 22033 6545
rect 22385 6369 22419 6545
rect 22503 6369 22537 6545
rect 22621 6369 22655 6545
rect 22739 6369 22773 6545
rect 23123 6369 23157 6545
rect 23241 6369 23275 6545
rect 23359 6369 23393 6545
rect 23477 6369 23511 6545
rect 23861 6369 23895 6545
rect 23979 6369 24013 6545
rect 24097 6369 24131 6545
rect 24215 6369 24249 6545
rect 24599 6369 24633 6545
rect 24717 6369 24751 6545
rect 24835 6369 24869 6545
rect 24953 6369 24987 6545
rect 18495 6059 18529 6235
rect 18613 6059 18647 6235
rect 18731 6059 18765 6235
rect 18849 6059 18883 6235
rect 13464 5366 13498 5742
rect 13582 5366 13616 5742
rect 13700 5366 13734 5742
rect 13818 5366 13852 5742
rect 13936 5366 13970 5742
rect 14054 5366 14088 5742
rect 14172 5366 14206 5742
rect 15533 5364 15567 5740
rect 15651 5364 15685 5740
rect 15769 5364 15803 5740
rect 15887 5364 15921 5740
rect 16005 5364 16039 5740
rect 16123 5364 16157 5740
rect 16241 5364 16275 5740
rect 17601 5366 17635 5742
rect 17719 5366 17753 5742
rect 17837 5366 17871 5742
rect 17955 5366 17989 5742
rect 18073 5366 18107 5742
rect 18191 5366 18225 5742
rect 18309 5366 18343 5742
rect 260 1752 294 1928
rect 378 1752 412 1928
rect 496 1752 530 1928
rect 614 1752 648 1928
rect 701 1752 735 2128
rect 819 1752 853 2128
rect 937 1752 971 2128
rect 1055 1752 1089 2128
rect 1168 1752 1202 2128
rect 1286 1752 1320 2128
rect 1404 1752 1438 2128
rect 1522 1752 1556 2128
rect 1640 1752 1674 2128
rect 1758 1752 1792 2128
rect 1876 1752 1910 2128
rect 1995 1752 2029 2128
rect 2113 1752 2147 2128
rect 2231 1752 2265 2128
rect 2349 1752 2383 2128
rect 2468 1752 2502 1928
rect 2586 1752 2620 1928
rect 2704 1752 2738 1928
rect 2822 1752 2856 1928
rect 3404 1752 3438 1928
rect 3522 1752 3556 1928
rect 3640 1752 3674 1928
rect 3758 1752 3792 1928
rect 3845 1752 3879 2128
rect 3963 1752 3997 2128
rect 4081 1752 4115 2128
rect 4199 1752 4233 2128
rect 4312 1752 4346 2128
rect 4430 1752 4464 2128
rect 4548 1752 4582 2128
rect 4666 1752 4700 2128
rect 4784 1752 4818 2128
rect 4902 1752 4936 2128
rect 5020 1752 5054 2128
rect 5139 1752 5173 2128
rect 5257 1752 5291 2128
rect 5375 1752 5409 2128
rect 5493 1752 5527 2128
rect 5612 1752 5646 1928
rect 5730 1752 5764 1928
rect 5848 1752 5882 1928
rect 5966 1752 6000 1928
rect 6536 1756 6570 1932
rect 6654 1756 6688 1932
rect 6772 1756 6806 1932
rect 6890 1756 6924 1932
rect 6977 1756 7011 2132
rect 7095 1756 7129 2132
rect 7213 1756 7247 2132
rect 7331 1756 7365 2132
rect 7444 1756 7478 2132
rect 7562 1756 7596 2132
rect 7680 1756 7714 2132
rect 7798 1756 7832 2132
rect 7916 1756 7950 2132
rect 8034 1756 8068 2132
rect 8152 1756 8186 2132
rect 8271 1756 8305 2132
rect 8389 1756 8423 2132
rect 8507 1756 8541 2132
rect 8625 1756 8659 2132
rect 8744 1756 8778 1932
rect 8862 1756 8896 1932
rect 8980 1756 9014 1932
rect 9098 1756 9132 1932
rect 9680 1756 9714 1932
rect 9798 1756 9832 1932
rect 9916 1756 9950 1932
rect 10034 1756 10068 1932
rect 10121 1756 10155 2132
rect 10239 1756 10273 2132
rect 10357 1756 10391 2132
rect 10475 1756 10509 2132
rect 10588 1756 10622 2132
rect 10706 1756 10740 2132
rect 10824 1756 10858 2132
rect 10942 1756 10976 2132
rect 11060 1756 11094 2132
rect 11178 1756 11212 2132
rect 11296 1756 11330 2132
rect 11415 1756 11449 2132
rect 11533 1756 11567 2132
rect 11651 1756 11685 2132
rect 11769 1756 11803 2132
rect 11888 1756 11922 1932
rect 12006 1756 12040 1932
rect 12124 1756 12158 1932
rect 12242 1756 12276 1932
rect 12882 1752 12916 1928
rect 13000 1752 13034 1928
rect 13118 1752 13152 1928
rect 13236 1752 13270 1928
rect 13323 1752 13357 2128
rect 13441 1752 13475 2128
rect 13559 1752 13593 2128
rect 13677 1752 13711 2128
rect 13790 1752 13824 2128
rect 13908 1752 13942 2128
rect 14026 1752 14060 2128
rect 14144 1752 14178 2128
rect 14262 1752 14296 2128
rect 14380 1752 14414 2128
rect 14498 1752 14532 2128
rect 14617 1752 14651 2128
rect 14735 1752 14769 2128
rect 14853 1752 14887 2128
rect 14971 1752 15005 2128
rect 15090 1752 15124 1928
rect 15208 1752 15242 1928
rect 15326 1752 15360 1928
rect 15444 1752 15478 1928
rect 16026 1752 16060 1928
rect 16144 1752 16178 1928
rect 16262 1752 16296 1928
rect 16380 1752 16414 1928
rect 16467 1752 16501 2128
rect 16585 1752 16619 2128
rect 16703 1752 16737 2128
rect 16821 1752 16855 2128
rect 16934 1752 16968 2128
rect 17052 1752 17086 2128
rect 17170 1752 17204 2128
rect 17288 1752 17322 2128
rect 17406 1752 17440 2128
rect 17524 1752 17558 2128
rect 17642 1752 17676 2128
rect 17761 1752 17795 2128
rect 17879 1752 17913 2128
rect 17997 1752 18031 2128
rect 18115 1752 18149 2128
rect 18234 1752 18268 1928
rect 18352 1752 18386 1928
rect 18470 1752 18504 1928
rect 18588 1752 18622 1928
rect 19158 1756 19192 1932
rect 19276 1756 19310 1932
rect 19394 1756 19428 1932
rect 19512 1756 19546 1932
rect 19599 1756 19633 2132
rect 19717 1756 19751 2132
rect 19835 1756 19869 2132
rect 19953 1756 19987 2132
rect 20066 1756 20100 2132
rect 20184 1756 20218 2132
rect 20302 1756 20336 2132
rect 20420 1756 20454 2132
rect 20538 1756 20572 2132
rect 20656 1756 20690 2132
rect 20774 1756 20808 2132
rect 20893 1756 20927 2132
rect 21011 1756 21045 2132
rect 21129 1756 21163 2132
rect 21247 1756 21281 2132
rect 21366 1756 21400 1932
rect 21484 1756 21518 1932
rect 21602 1756 21636 1932
rect 21720 1756 21754 1932
rect 22302 1756 22336 1932
rect 22420 1756 22454 1932
rect 22538 1756 22572 1932
rect 22656 1756 22690 1932
rect 22743 1756 22777 2132
rect 22861 1756 22895 2132
rect 22979 1756 23013 2132
rect 23097 1756 23131 2132
rect 23210 1756 23244 2132
rect 23328 1756 23362 2132
rect 23446 1756 23480 2132
rect 23564 1756 23598 2132
rect 23682 1756 23716 2132
rect 23800 1756 23834 2132
rect 23918 1756 23952 2132
rect 24037 1756 24071 2132
rect 24155 1756 24189 2132
rect 24273 1756 24307 2132
rect 24391 1756 24425 2132
rect 24510 1756 24544 1932
rect 24628 1756 24662 1932
rect 24746 1756 24780 1932
rect 24864 1756 24898 1932
rect 292 -2140 326 -1964
rect 410 -2140 444 -1964
rect 528 -2140 562 -1964
rect 646 -2140 680 -1964
rect 733 -2140 767 -1764
rect 851 -2140 885 -1764
rect 969 -2140 1003 -1764
rect 1087 -2140 1121 -1764
rect 1200 -2140 1234 -1764
rect 1318 -2140 1352 -1764
rect 1436 -2140 1470 -1764
rect 1554 -2140 1588 -1764
rect 1672 -2140 1706 -1764
rect 1790 -2140 1824 -1764
rect 1908 -2140 1942 -1764
rect 2027 -2140 2061 -1764
rect 2145 -2140 2179 -1764
rect 2263 -2140 2297 -1764
rect 2381 -2140 2415 -1764
rect 2500 -2140 2534 -1964
rect 2618 -2140 2652 -1964
rect 2736 -2140 2770 -1964
rect 2854 -2140 2888 -1964
rect 3436 -2140 3470 -1964
rect 3554 -2140 3588 -1964
rect 3672 -2140 3706 -1964
rect 3790 -2140 3824 -1964
rect 3877 -2140 3911 -1764
rect 3995 -2140 4029 -1764
rect 4113 -2140 4147 -1764
rect 4231 -2140 4265 -1764
rect 4344 -2140 4378 -1764
rect 4462 -2140 4496 -1764
rect 4580 -2140 4614 -1764
rect 4698 -2140 4732 -1764
rect 4816 -2140 4850 -1764
rect 4934 -2140 4968 -1764
rect 5052 -2140 5086 -1764
rect 5171 -2140 5205 -1764
rect 5289 -2140 5323 -1764
rect 5407 -2140 5441 -1764
rect 5525 -2140 5559 -1764
rect 5644 -2140 5678 -1964
rect 5762 -2140 5796 -1964
rect 5880 -2140 5914 -1964
rect 5998 -2140 6032 -1964
rect 6568 -2136 6602 -1960
rect 6686 -2136 6720 -1960
rect 6804 -2136 6838 -1960
rect 6922 -2136 6956 -1960
rect 7009 -2136 7043 -1760
rect 7127 -2136 7161 -1760
rect 7245 -2136 7279 -1760
rect 7363 -2136 7397 -1760
rect 7476 -2136 7510 -1760
rect 7594 -2136 7628 -1760
rect 7712 -2136 7746 -1760
rect 7830 -2136 7864 -1760
rect 7948 -2136 7982 -1760
rect 8066 -2136 8100 -1760
rect 8184 -2136 8218 -1760
rect 8303 -2136 8337 -1760
rect 8421 -2136 8455 -1760
rect 8539 -2136 8573 -1760
rect 8657 -2136 8691 -1760
rect 8776 -2136 8810 -1960
rect 8894 -2136 8928 -1960
rect 9012 -2136 9046 -1960
rect 9130 -2136 9164 -1960
rect 9712 -2136 9746 -1960
rect 9830 -2136 9864 -1960
rect 9948 -2136 9982 -1960
rect 10066 -2136 10100 -1960
rect 10153 -2136 10187 -1760
rect 10271 -2136 10305 -1760
rect 10389 -2136 10423 -1760
rect 10507 -2136 10541 -1760
rect 10620 -2136 10654 -1760
rect 10738 -2136 10772 -1760
rect 10856 -2136 10890 -1760
rect 10974 -2136 11008 -1760
rect 11092 -2136 11126 -1760
rect 11210 -2136 11244 -1760
rect 11328 -2136 11362 -1760
rect 11447 -2136 11481 -1760
rect 11565 -2136 11599 -1760
rect 11683 -2136 11717 -1760
rect 11801 -2136 11835 -1760
rect 11920 -2136 11954 -1960
rect 12038 -2136 12072 -1960
rect 12156 -2136 12190 -1960
rect 12274 -2136 12308 -1960
rect 12914 -2140 12948 -1964
rect 13032 -2140 13066 -1964
rect 13150 -2140 13184 -1964
rect 13268 -2140 13302 -1964
rect 13355 -2140 13389 -1764
rect 13473 -2140 13507 -1764
rect 13591 -2140 13625 -1764
rect 13709 -2140 13743 -1764
rect 13822 -2140 13856 -1764
rect 13940 -2140 13974 -1764
rect 14058 -2140 14092 -1764
rect 14176 -2140 14210 -1764
rect 14294 -2140 14328 -1764
rect 14412 -2140 14446 -1764
rect 14530 -2140 14564 -1764
rect 14649 -2140 14683 -1764
rect 14767 -2140 14801 -1764
rect 14885 -2140 14919 -1764
rect 15003 -2140 15037 -1764
rect 15122 -2140 15156 -1964
rect 15240 -2140 15274 -1964
rect 15358 -2140 15392 -1964
rect 15476 -2140 15510 -1964
rect 16058 -2140 16092 -1964
rect 16176 -2140 16210 -1964
rect 16294 -2140 16328 -1964
rect 16412 -2140 16446 -1964
rect 16499 -2140 16533 -1764
rect 16617 -2140 16651 -1764
rect 16735 -2140 16769 -1764
rect 16853 -2140 16887 -1764
rect 16966 -2140 17000 -1764
rect 17084 -2140 17118 -1764
rect 17202 -2140 17236 -1764
rect 17320 -2140 17354 -1764
rect 17438 -2140 17472 -1764
rect 17556 -2140 17590 -1764
rect 17674 -2140 17708 -1764
rect 17793 -2140 17827 -1764
rect 17911 -2140 17945 -1764
rect 18029 -2140 18063 -1764
rect 18147 -2140 18181 -1764
rect 18266 -2140 18300 -1964
rect 18384 -2140 18418 -1964
rect 18502 -2140 18536 -1964
rect 18620 -2140 18654 -1964
rect 19190 -2136 19224 -1960
rect 19308 -2136 19342 -1960
rect 19426 -2136 19460 -1960
rect 19544 -2136 19578 -1960
rect 19631 -2136 19665 -1760
rect 19749 -2136 19783 -1760
rect 19867 -2136 19901 -1760
rect 19985 -2136 20019 -1760
rect 20098 -2136 20132 -1760
rect 20216 -2136 20250 -1760
rect 20334 -2136 20368 -1760
rect 20452 -2136 20486 -1760
rect 20570 -2136 20604 -1760
rect 20688 -2136 20722 -1760
rect 20806 -2136 20840 -1760
rect 20925 -2136 20959 -1760
rect 21043 -2136 21077 -1760
rect 21161 -2136 21195 -1760
rect 21279 -2136 21313 -1760
rect 21398 -2136 21432 -1960
rect 21516 -2136 21550 -1960
rect 21634 -2136 21668 -1960
rect 21752 -2136 21786 -1960
rect 22334 -2136 22368 -1960
rect 22452 -2136 22486 -1960
rect 22570 -2136 22604 -1960
rect 22688 -2136 22722 -1960
rect 22775 -2136 22809 -1760
rect 22893 -2136 22927 -1760
rect 23011 -2136 23045 -1760
rect 23129 -2136 23163 -1760
rect 23242 -2136 23276 -1760
rect 23360 -2136 23394 -1760
rect 23478 -2136 23512 -1760
rect 23596 -2136 23630 -1760
rect 23714 -2136 23748 -1760
rect 23832 -2136 23866 -1760
rect 23950 -2136 23984 -1760
rect 24069 -2136 24103 -1760
rect 24187 -2136 24221 -1760
rect 24305 -2136 24339 -1760
rect 24423 -2136 24457 -1760
rect 24542 -2136 24576 -1960
rect 24660 -2136 24694 -1960
rect 24778 -2136 24812 -1960
rect 24896 -2136 24930 -1960
<< psubdiff >>
rect 1668 20004 1854 20028
rect 1668 19958 1710 20004
rect 1814 19958 1854 20004
rect 1668 19922 1854 19958
rect 4812 20004 4998 20028
rect 4812 19958 4854 20004
rect 4958 19958 4998 20004
rect 4812 19922 4998 19958
rect 7944 20008 8130 20032
rect 7944 19962 7986 20008
rect 8090 19962 8130 20008
rect 7944 19926 8130 19962
rect 11088 20008 11274 20032
rect 11088 19962 11130 20008
rect 11234 19962 11274 20008
rect 11088 19926 11274 19962
rect 14290 20004 14476 20028
rect 14290 19958 14332 20004
rect 14436 19958 14476 20004
rect 14290 19922 14476 19958
rect 17434 20004 17620 20028
rect 17434 19958 17476 20004
rect 17580 19958 17620 20004
rect 17434 19922 17620 19958
rect 20566 20008 20752 20032
rect 20566 19962 20608 20008
rect 20712 19962 20752 20008
rect 20566 19926 20752 19962
rect 23710 20008 23896 20032
rect 23710 19962 23752 20008
rect 23856 19962 23896 20008
rect 23710 19926 23896 19962
rect 14704 15702 14900 15732
rect 3398 15631 3610 15661
rect 3398 15575 3438 15631
rect 3572 15575 3610 15631
rect 3398 15553 3610 15575
rect 4846 15631 5058 15661
rect 4846 15575 4886 15631
rect 5020 15575 5058 15631
rect 4846 15553 5058 15575
rect 6344 15633 6556 15663
rect 6344 15577 6384 15633
rect 6518 15577 6556 15633
rect 6344 15555 6556 15577
rect 7792 15633 8004 15663
rect 7792 15577 7832 15633
rect 7966 15577 8004 15633
rect 7792 15555 8004 15577
rect 9312 15631 9524 15661
rect 9312 15575 9352 15631
rect 9486 15575 9524 15631
rect 9312 15553 9524 15575
rect 10760 15631 10972 15661
rect 10760 15575 10800 15631
rect 10934 15575 10972 15631
rect 10760 15553 10972 15575
rect 12258 15633 12470 15663
rect 12258 15577 12298 15633
rect 12432 15577 12470 15633
rect 12258 15555 12470 15577
rect 13706 15633 13918 15663
rect 13706 15577 13746 15633
rect 13880 15577 13918 15633
rect 14704 15636 14744 15702
rect 14862 15636 14900 15702
rect 14704 15588 14900 15636
rect 15872 15702 16068 15732
rect 15872 15636 15912 15702
rect 16030 15636 16068 15702
rect 15872 15588 16068 15636
rect 17040 15702 17236 15732
rect 17040 15636 17080 15702
rect 17198 15636 17236 15702
rect 17040 15588 17236 15636
rect 18208 15702 18404 15732
rect 18208 15636 18248 15702
rect 18366 15636 18404 15702
rect 18208 15588 18404 15636
rect 19382 15704 19578 15734
rect 19382 15638 19422 15704
rect 19540 15638 19578 15704
rect 19382 15590 19578 15638
rect 20550 15704 20746 15734
rect 20550 15638 20590 15704
rect 20708 15638 20746 15704
rect 20550 15590 20746 15638
rect 21718 15704 21914 15734
rect 21718 15638 21758 15704
rect 21876 15638 21914 15704
rect 21718 15590 21914 15638
rect 22886 15704 23082 15734
rect 22886 15638 22926 15704
rect 23044 15638 23082 15704
rect 22886 15590 23082 15638
rect 13706 15555 13918 15577
rect 4170 12866 4356 12890
rect 4170 12820 4212 12866
rect 4316 12820 4356 12866
rect 4170 12784 4356 12820
rect 7314 12866 7500 12890
rect 7314 12820 7356 12866
rect 7460 12820 7500 12866
rect 7314 12784 7500 12820
rect 10446 12870 10632 12894
rect 10446 12824 10488 12870
rect 10592 12824 10632 12870
rect 10446 12788 10632 12824
rect 13590 12870 13776 12894
rect 13590 12824 13632 12870
rect 13736 12824 13776 12870
rect 13590 12788 13776 12824
rect 16792 12866 16978 12890
rect 16792 12820 16834 12866
rect 16938 12820 16978 12866
rect 16792 12784 16978 12820
rect 19936 12866 20122 12890
rect 19936 12820 19978 12866
rect 20082 12820 20122 12866
rect 19936 12784 20122 12820
rect 23068 12870 23254 12894
rect 23068 12824 23110 12870
rect 23214 12824 23254 12870
rect 23068 12788 23254 12824
rect 26212 12870 26398 12894
rect 26212 12824 26254 12870
rect 26358 12824 26398 12870
rect 26212 12788 26398 12824
rect 4170 10132 4356 10156
rect 4170 10086 4212 10132
rect 4316 10086 4356 10132
rect 4170 10050 4356 10086
rect 7314 10132 7500 10156
rect 7314 10086 7356 10132
rect 7460 10086 7500 10132
rect 7314 10050 7500 10086
rect 10446 10136 10632 10160
rect 10446 10090 10488 10136
rect 10592 10090 10632 10136
rect 10446 10054 10632 10090
rect 13590 10136 13776 10160
rect 13590 10090 13632 10136
rect 13736 10090 13776 10136
rect 13590 10054 13776 10090
rect 16792 10132 16978 10156
rect 16792 10086 16834 10132
rect 16938 10086 16978 10132
rect 16792 10050 16978 10086
rect 19936 10132 20122 10156
rect 19936 10086 19978 10132
rect 20082 10086 20122 10132
rect 19936 10050 20122 10086
rect 23068 10136 23254 10160
rect 23068 10090 23110 10136
rect 23214 10090 23254 10136
rect 23068 10054 23254 10090
rect 26212 10136 26398 10160
rect 26212 10090 26254 10136
rect 26358 10090 26398 10136
rect 26212 10054 26398 10090
rect 4160 7400 4346 7424
rect 4160 7354 4202 7400
rect 4306 7354 4346 7400
rect 4160 7318 4346 7354
rect 7304 7400 7490 7424
rect 7304 7354 7346 7400
rect 7450 7354 7490 7400
rect 7304 7318 7490 7354
rect 10436 7404 10622 7428
rect 10436 7358 10478 7404
rect 10582 7358 10622 7404
rect 10436 7322 10622 7358
rect 13580 7404 13766 7428
rect 13580 7358 13622 7404
rect 13726 7358 13766 7404
rect 13580 7322 13766 7358
rect 16782 7400 16968 7424
rect 16782 7354 16824 7400
rect 16928 7354 16968 7400
rect 16782 7318 16968 7354
rect 19926 7400 20112 7424
rect 19926 7354 19968 7400
rect 20072 7354 20112 7400
rect 19926 7318 20112 7354
rect 23058 7404 23244 7428
rect 23058 7358 23100 7404
rect 23204 7358 23244 7404
rect 23058 7322 23244 7358
rect 26202 7404 26388 7428
rect 26202 7358 26244 7404
rect 26348 7358 26388 7404
rect 26202 7322 26388 7358
rect 19423 5873 19683 5919
rect 19423 5803 19485 5873
rect 19629 5803 19683 5873
rect 19423 5769 19683 5803
rect 20161 5871 20421 5917
rect 20161 5801 20223 5871
rect 20367 5801 20421 5871
rect 20161 5767 20421 5801
rect 20899 5871 21159 5917
rect 20899 5801 20961 5871
rect 21105 5801 21159 5871
rect 20899 5767 21159 5801
rect 21641 5871 21901 5917
rect 21641 5801 21703 5871
rect 21847 5801 21901 5871
rect 21641 5767 21901 5801
rect 22381 5871 22641 5917
rect 22381 5801 22443 5871
rect 22587 5801 22641 5871
rect 22381 5767 22641 5801
rect 23119 5871 23379 5917
rect 23119 5801 23181 5871
rect 23325 5801 23379 5871
rect 23119 5767 23379 5801
rect 23857 5871 24117 5917
rect 23857 5801 23919 5871
rect 24063 5801 24117 5871
rect 23857 5767 24117 5801
rect 24595 5871 24855 5917
rect 24595 5801 24657 5871
rect 24801 5801 24855 5871
rect 24595 5767 24855 5801
rect 3372 4442 3624 4462
rect 3372 4386 3430 4442
rect 3562 4386 3624 4442
rect 3372 4364 3624 4386
rect 5440 4444 5692 4464
rect 5440 4388 5498 4444
rect 5630 4388 5692 4444
rect 5440 4366 5692 4388
rect 7509 4442 7761 4462
rect 7509 4386 7567 4442
rect 7699 4386 7761 4442
rect 7509 4364 7761 4386
rect 9577 4444 9829 4464
rect 9577 4388 9635 4444
rect 9767 4388 9829 4444
rect 9577 4366 9829 4388
rect 11646 4444 11898 4464
rect 11646 4388 11704 4444
rect 11836 4388 11898 4444
rect 11646 4366 11898 4388
rect 13714 4446 13966 4466
rect 13714 4390 13772 4446
rect 13904 4390 13966 4446
rect 13714 4368 13966 4390
rect 15783 4444 16035 4464
rect 15783 4388 15841 4444
rect 15973 4388 16035 4444
rect 15783 4366 16035 4388
rect 17851 4446 18103 4466
rect 17851 4390 17909 4446
rect 18041 4390 18103 4446
rect 17851 4368 18103 4390
rect 1462 152 1648 176
rect 1462 106 1504 152
rect 1608 106 1648 152
rect 1462 70 1648 106
rect 4606 152 4792 176
rect 4606 106 4648 152
rect 4752 106 4792 152
rect 4606 70 4792 106
rect 7738 156 7924 180
rect 7738 110 7780 156
rect 7884 110 7924 156
rect 7738 74 7924 110
rect 10882 156 11068 180
rect 10882 110 10924 156
rect 11028 110 11068 156
rect 10882 74 11068 110
rect 14084 152 14270 176
rect 14084 106 14126 152
rect 14230 106 14270 152
rect 14084 70 14270 106
rect 17228 152 17414 176
rect 17228 106 17270 152
rect 17374 106 17414 152
rect 17228 70 17414 106
rect 20360 156 20546 180
rect 20360 110 20402 156
rect 20506 110 20546 156
rect 20360 74 20546 110
rect 23504 156 23690 180
rect 23504 110 23546 156
rect 23650 110 23690 156
rect 23504 74 23690 110
rect 1494 -3740 1680 -3716
rect 1494 -3786 1536 -3740
rect 1640 -3786 1680 -3740
rect 1494 -3822 1680 -3786
rect 4638 -3740 4824 -3716
rect 4638 -3786 4680 -3740
rect 4784 -3786 4824 -3740
rect 4638 -3822 4824 -3786
rect 7770 -3736 7956 -3712
rect 7770 -3782 7812 -3736
rect 7916 -3782 7956 -3736
rect 7770 -3818 7956 -3782
rect 10914 -3736 11100 -3712
rect 10914 -3782 10956 -3736
rect 11060 -3782 11100 -3736
rect 10914 -3818 11100 -3782
rect 14116 -3740 14302 -3716
rect 14116 -3786 14158 -3740
rect 14262 -3786 14302 -3740
rect 14116 -3822 14302 -3786
rect 17260 -3740 17446 -3716
rect 17260 -3786 17302 -3740
rect 17406 -3786 17446 -3740
rect 17260 -3822 17446 -3786
rect 20392 -3736 20578 -3712
rect 20392 -3782 20434 -3736
rect 20538 -3782 20578 -3736
rect 20392 -3818 20578 -3782
rect 23536 -3736 23722 -3712
rect 23536 -3782 23578 -3736
rect 23682 -3782 23722 -3736
rect 23536 -3818 23722 -3782
<< nsubdiff >>
rect 1598 22250 1902 22306
rect 1598 22174 1652 22250
rect 1848 22174 1902 22250
rect 1598 22160 1902 22174
rect 4742 22250 5046 22306
rect 4742 22174 4796 22250
rect 4992 22174 5046 22250
rect 4742 22160 5046 22174
rect 7874 22254 8178 22310
rect 7874 22178 7928 22254
rect 8124 22178 8178 22254
rect 7874 22164 8178 22178
rect 11018 22254 11322 22310
rect 11018 22178 11072 22254
rect 11268 22178 11322 22254
rect 11018 22164 11322 22178
rect 14220 22250 14524 22306
rect 14220 22174 14274 22250
rect 14470 22174 14524 22250
rect 14220 22160 14524 22174
rect 17364 22250 17668 22306
rect 17364 22174 17418 22250
rect 17614 22174 17668 22250
rect 17364 22160 17668 22174
rect 20496 22254 20800 22310
rect 20496 22178 20550 22254
rect 20746 22178 20800 22254
rect 20496 22164 20800 22178
rect 23640 22254 23944 22310
rect 23640 22178 23694 22254
rect 23890 22178 23944 22254
rect 23640 22164 23944 22178
rect 15144 17046 15410 17084
rect 15144 16974 15200 17046
rect 15344 16974 15410 17046
rect 16312 17046 16578 17084
rect 15144 16944 15410 16974
rect 3158 16839 3402 16877
rect 3158 16769 3214 16839
rect 3350 16769 3402 16839
rect 3158 16747 3402 16769
rect 4606 16839 4850 16877
rect 4606 16769 4662 16839
rect 4798 16769 4850 16839
rect 4606 16747 4850 16769
rect 6104 16841 6348 16879
rect 6104 16771 6160 16841
rect 6296 16771 6348 16841
rect 6104 16749 6348 16771
rect 7552 16841 7796 16879
rect 7552 16771 7608 16841
rect 7744 16771 7796 16841
rect 7552 16749 7796 16771
rect 9072 16839 9316 16877
rect 9072 16769 9128 16839
rect 9264 16769 9316 16839
rect 9072 16747 9316 16769
rect 10520 16839 10764 16877
rect 10520 16769 10576 16839
rect 10712 16769 10764 16839
rect 10520 16747 10764 16769
rect 12018 16841 12262 16879
rect 12018 16771 12074 16841
rect 12210 16771 12262 16841
rect 12018 16749 12262 16771
rect 13466 16841 13710 16879
rect 13466 16771 13522 16841
rect 13658 16771 13710 16841
rect 16312 16974 16368 17046
rect 16512 16974 16578 17046
rect 17480 17046 17746 17084
rect 16312 16944 16578 16974
rect 17480 16974 17536 17046
rect 17680 16974 17746 17046
rect 18648 17046 18914 17084
rect 17480 16944 17746 16974
rect 18648 16974 18704 17046
rect 18848 16974 18914 17046
rect 19822 17048 20088 17086
rect 18648 16944 18914 16974
rect 19822 16976 19878 17048
rect 20022 16976 20088 17048
rect 20990 17048 21256 17086
rect 19822 16946 20088 16976
rect 20990 16976 21046 17048
rect 21190 16976 21256 17048
rect 22158 17048 22424 17086
rect 20990 16946 21256 16976
rect 22158 16976 22214 17048
rect 22358 16976 22424 17048
rect 23326 17048 23592 17086
rect 22158 16946 22424 16976
rect 23326 16976 23382 17048
rect 23526 16976 23592 17048
rect 23326 16946 23592 16976
rect 13466 16749 13710 16771
rect 4100 15112 4404 15168
rect 4100 15036 4154 15112
rect 4350 15036 4404 15112
rect 4100 15022 4404 15036
rect 7244 15112 7548 15168
rect 7244 15036 7298 15112
rect 7494 15036 7548 15112
rect 7244 15022 7548 15036
rect 10376 15116 10680 15172
rect 10376 15040 10430 15116
rect 10626 15040 10680 15116
rect 10376 15026 10680 15040
rect 13520 15116 13824 15172
rect 13520 15040 13574 15116
rect 13770 15040 13824 15116
rect 13520 15026 13824 15040
rect 16722 15112 17026 15168
rect 16722 15036 16776 15112
rect 16972 15036 17026 15112
rect 16722 15022 17026 15036
rect 19866 15112 20170 15168
rect 19866 15036 19920 15112
rect 20116 15036 20170 15112
rect 19866 15022 20170 15036
rect 22998 15116 23302 15172
rect 22998 15040 23052 15116
rect 23248 15040 23302 15116
rect 22998 15026 23302 15040
rect 26142 15116 26446 15172
rect 26142 15040 26196 15116
rect 26392 15040 26446 15116
rect 26142 15026 26446 15040
rect 4100 12378 4404 12434
rect 4100 12302 4154 12378
rect 4350 12302 4404 12378
rect 4100 12288 4404 12302
rect 7244 12378 7548 12434
rect 7244 12302 7298 12378
rect 7494 12302 7548 12378
rect 7244 12288 7548 12302
rect 10376 12382 10680 12438
rect 10376 12306 10430 12382
rect 10626 12306 10680 12382
rect 10376 12292 10680 12306
rect 13520 12382 13824 12438
rect 13520 12306 13574 12382
rect 13770 12306 13824 12382
rect 13520 12292 13824 12306
rect 16722 12378 17026 12434
rect 16722 12302 16776 12378
rect 16972 12302 17026 12378
rect 16722 12288 17026 12302
rect 19866 12378 20170 12434
rect 19866 12302 19920 12378
rect 20116 12302 20170 12378
rect 19866 12288 20170 12302
rect 22998 12382 23302 12438
rect 22998 12306 23052 12382
rect 23248 12306 23302 12382
rect 22998 12292 23302 12306
rect 26142 12382 26446 12438
rect 26142 12306 26196 12382
rect 26392 12306 26446 12382
rect 26142 12292 26446 12306
rect 4090 9646 4394 9702
rect 4090 9570 4144 9646
rect 4340 9570 4394 9646
rect 4090 9556 4394 9570
rect 7234 9646 7538 9702
rect 7234 9570 7288 9646
rect 7484 9570 7538 9646
rect 7234 9556 7538 9570
rect 10366 9650 10670 9706
rect 10366 9574 10420 9650
rect 10616 9574 10670 9650
rect 10366 9560 10670 9574
rect 13510 9650 13814 9706
rect 13510 9574 13564 9650
rect 13760 9574 13814 9650
rect 13510 9560 13814 9574
rect 16712 9646 17016 9702
rect 16712 9570 16766 9646
rect 16962 9570 17016 9646
rect 16712 9556 17016 9570
rect 19856 9646 20160 9702
rect 19856 9570 19910 9646
rect 20106 9570 20160 9646
rect 19856 9556 20160 9570
rect 22988 9650 23292 9706
rect 22988 9574 23042 9650
rect 23238 9574 23292 9650
rect 22988 9560 23292 9574
rect 26132 9650 26436 9706
rect 26132 9574 26186 9650
rect 26382 9574 26436 9650
rect 26132 9560 26436 9574
rect 3356 6702 3756 6754
rect 3356 6658 3480 6702
rect 3602 6658 3756 6702
rect 3356 6610 3756 6658
rect 5424 6704 5824 6756
rect 5424 6660 5548 6704
rect 5670 6660 5824 6704
rect 5424 6612 5824 6660
rect 7493 6702 7893 6754
rect 7493 6658 7617 6702
rect 7739 6658 7893 6702
rect 7493 6610 7893 6658
rect 9561 6704 9961 6756
rect 9561 6660 9685 6704
rect 9807 6660 9961 6704
rect 9561 6612 9961 6660
rect 11630 6704 12030 6756
rect 11630 6660 11754 6704
rect 11876 6660 12030 6704
rect 11630 6612 12030 6660
rect 13698 6706 14098 6758
rect 13698 6662 13822 6706
rect 13944 6662 14098 6706
rect 13698 6614 14098 6662
rect 15767 6704 16167 6756
rect 15767 6660 15891 6704
rect 16013 6660 16167 6704
rect 15767 6612 16167 6660
rect 17835 6706 18235 6758
rect 17835 6662 17959 6706
rect 18081 6662 18235 6706
rect 17835 6614 18235 6662
rect 19473 6753 19769 6767
rect 19473 6691 19551 6753
rect 19691 6691 19769 6753
rect 19473 6635 19769 6691
rect 20211 6751 20507 6765
rect 20211 6689 20289 6751
rect 20429 6689 20507 6751
rect 20211 6633 20507 6689
rect 20949 6751 21245 6765
rect 20949 6689 21027 6751
rect 21167 6689 21245 6751
rect 20949 6633 21245 6689
rect 21691 6751 21987 6765
rect 21691 6689 21769 6751
rect 21909 6689 21987 6751
rect 21691 6633 21987 6689
rect 22431 6751 22727 6765
rect 22431 6689 22509 6751
rect 22649 6689 22727 6751
rect 22431 6633 22727 6689
rect 23169 6751 23465 6765
rect 23169 6689 23247 6751
rect 23387 6689 23465 6751
rect 23169 6633 23465 6689
rect 23907 6751 24203 6765
rect 23907 6689 23985 6751
rect 24125 6689 24203 6751
rect 23907 6633 24203 6689
rect 24645 6751 24941 6765
rect 24645 6689 24723 6751
rect 24863 6689 24941 6751
rect 24645 6633 24941 6689
rect 1392 2398 1696 2454
rect 1392 2322 1446 2398
rect 1642 2322 1696 2398
rect 1392 2308 1696 2322
rect 4536 2398 4840 2454
rect 4536 2322 4590 2398
rect 4786 2322 4840 2398
rect 4536 2308 4840 2322
rect 7668 2402 7972 2458
rect 7668 2326 7722 2402
rect 7918 2326 7972 2402
rect 7668 2312 7972 2326
rect 10812 2402 11116 2458
rect 10812 2326 10866 2402
rect 11062 2326 11116 2402
rect 10812 2312 11116 2326
rect 14014 2398 14318 2454
rect 14014 2322 14068 2398
rect 14264 2322 14318 2398
rect 14014 2308 14318 2322
rect 17158 2398 17462 2454
rect 17158 2322 17212 2398
rect 17408 2322 17462 2398
rect 17158 2308 17462 2322
rect 20290 2402 20594 2458
rect 20290 2326 20344 2402
rect 20540 2326 20594 2402
rect 20290 2312 20594 2326
rect 23434 2402 23738 2458
rect 23434 2326 23488 2402
rect 23684 2326 23738 2402
rect 23434 2312 23738 2326
rect 1424 -1494 1728 -1438
rect 1424 -1570 1478 -1494
rect 1674 -1570 1728 -1494
rect 1424 -1584 1728 -1570
rect 4568 -1494 4872 -1438
rect 4568 -1570 4622 -1494
rect 4818 -1570 4872 -1494
rect 4568 -1584 4872 -1570
rect 7700 -1490 8004 -1434
rect 7700 -1566 7754 -1490
rect 7950 -1566 8004 -1490
rect 7700 -1580 8004 -1566
rect 10844 -1490 11148 -1434
rect 10844 -1566 10898 -1490
rect 11094 -1566 11148 -1490
rect 10844 -1580 11148 -1566
rect 14046 -1494 14350 -1438
rect 14046 -1570 14100 -1494
rect 14296 -1570 14350 -1494
rect 14046 -1584 14350 -1570
rect 17190 -1494 17494 -1438
rect 17190 -1570 17244 -1494
rect 17440 -1570 17494 -1494
rect 17190 -1584 17494 -1570
rect 20322 -1490 20626 -1434
rect 20322 -1566 20376 -1490
rect 20572 -1566 20626 -1490
rect 20322 -1580 20626 -1566
rect 23466 -1490 23770 -1434
rect 23466 -1566 23520 -1490
rect 23716 -1566 23770 -1490
rect 23466 -1580 23770 -1566
<< psubdiffcont >>
rect 1710 19958 1814 20004
rect 4854 19958 4958 20004
rect 7986 19962 8090 20008
rect 11130 19962 11234 20008
rect 14332 19958 14436 20004
rect 17476 19958 17580 20004
rect 20608 19962 20712 20008
rect 23752 19962 23856 20008
rect 3438 15575 3572 15631
rect 4886 15575 5020 15631
rect 6384 15577 6518 15633
rect 7832 15577 7966 15633
rect 9352 15575 9486 15631
rect 10800 15575 10934 15631
rect 12298 15577 12432 15633
rect 13746 15577 13880 15633
rect 14744 15636 14862 15702
rect 15912 15636 16030 15702
rect 17080 15636 17198 15702
rect 18248 15636 18366 15702
rect 19422 15638 19540 15704
rect 20590 15638 20708 15704
rect 21758 15638 21876 15704
rect 22926 15638 23044 15704
rect 4212 12820 4316 12866
rect 7356 12820 7460 12866
rect 10488 12824 10592 12870
rect 13632 12824 13736 12870
rect 16834 12820 16938 12866
rect 19978 12820 20082 12866
rect 23110 12824 23214 12870
rect 26254 12824 26358 12870
rect 4212 10086 4316 10132
rect 7356 10086 7460 10132
rect 10488 10090 10592 10136
rect 13632 10090 13736 10136
rect 16834 10086 16938 10132
rect 19978 10086 20082 10132
rect 23110 10090 23214 10136
rect 26254 10090 26358 10136
rect 4202 7354 4306 7400
rect 7346 7354 7450 7400
rect 10478 7358 10582 7404
rect 13622 7358 13726 7404
rect 16824 7354 16928 7400
rect 19968 7354 20072 7400
rect 23100 7358 23204 7404
rect 26244 7358 26348 7404
rect 19485 5803 19629 5873
rect 20223 5801 20367 5871
rect 20961 5801 21105 5871
rect 21703 5801 21847 5871
rect 22443 5801 22587 5871
rect 23181 5801 23325 5871
rect 23919 5801 24063 5871
rect 24657 5801 24801 5871
rect 3430 4386 3562 4442
rect 5498 4388 5630 4444
rect 7567 4386 7699 4442
rect 9635 4388 9767 4444
rect 11704 4388 11836 4444
rect 13772 4390 13904 4446
rect 15841 4388 15973 4444
rect 17909 4390 18041 4446
rect 1504 106 1608 152
rect 4648 106 4752 152
rect 7780 110 7884 156
rect 10924 110 11028 156
rect 14126 106 14230 152
rect 17270 106 17374 152
rect 20402 110 20506 156
rect 23546 110 23650 156
rect 1536 -3786 1640 -3740
rect 4680 -3786 4784 -3740
rect 7812 -3782 7916 -3736
rect 10956 -3782 11060 -3736
rect 14158 -3786 14262 -3740
rect 17302 -3786 17406 -3740
rect 20434 -3782 20538 -3736
rect 23578 -3782 23682 -3736
<< nsubdiffcont >>
rect 1652 22174 1848 22250
rect 4796 22174 4992 22250
rect 7928 22178 8124 22254
rect 11072 22178 11268 22254
rect 14274 22174 14470 22250
rect 17418 22174 17614 22250
rect 20550 22178 20746 22254
rect 23694 22178 23890 22254
rect 15200 16974 15344 17046
rect 3214 16769 3350 16839
rect 4662 16769 4798 16839
rect 6160 16771 6296 16841
rect 7608 16771 7744 16841
rect 9128 16769 9264 16839
rect 10576 16769 10712 16839
rect 12074 16771 12210 16841
rect 13522 16771 13658 16841
rect 16368 16974 16512 17046
rect 17536 16974 17680 17046
rect 18704 16974 18848 17046
rect 19878 16976 20022 17048
rect 21046 16976 21190 17048
rect 22214 16976 22358 17048
rect 23382 16976 23526 17048
rect 4154 15036 4350 15112
rect 7298 15036 7494 15112
rect 10430 15040 10626 15116
rect 13574 15040 13770 15116
rect 16776 15036 16972 15112
rect 19920 15036 20116 15112
rect 23052 15040 23248 15116
rect 26196 15040 26392 15116
rect 4154 12302 4350 12378
rect 7298 12302 7494 12378
rect 10430 12306 10626 12382
rect 13574 12306 13770 12382
rect 16776 12302 16972 12378
rect 19920 12302 20116 12378
rect 23052 12306 23248 12382
rect 26196 12306 26392 12382
rect 4144 9570 4340 9646
rect 7288 9570 7484 9646
rect 10420 9574 10616 9650
rect 13564 9574 13760 9650
rect 16766 9570 16962 9646
rect 19910 9570 20106 9646
rect 23042 9574 23238 9650
rect 26186 9574 26382 9650
rect 3480 6658 3602 6702
rect 5548 6660 5670 6704
rect 7617 6658 7739 6702
rect 9685 6660 9807 6704
rect 11754 6660 11876 6704
rect 13822 6662 13944 6706
rect 15891 6660 16013 6704
rect 17959 6662 18081 6706
rect 19551 6691 19691 6753
rect 20289 6689 20429 6751
rect 21027 6689 21167 6751
rect 21769 6689 21909 6751
rect 22509 6689 22649 6751
rect 23247 6689 23387 6751
rect 23985 6689 24125 6751
rect 24723 6689 24863 6751
rect 1446 2322 1642 2398
rect 4590 2322 4786 2398
rect 7722 2326 7918 2402
rect 10866 2326 11062 2402
rect 14068 2322 14264 2398
rect 17212 2322 17408 2398
rect 20344 2326 20540 2402
rect 23488 2326 23684 2402
rect 1478 -1570 1674 -1494
rect 4622 -1570 4818 -1494
rect 7754 -1566 7950 -1490
rect 10898 -1566 11094 -1490
rect 14100 -1570 14296 -1494
rect 17244 -1570 17440 -1494
rect 20376 -1566 20572 -1490
rect 23520 -1566 23716 -1490
<< poly >>
rect 953 22007 1249 22046
rect 953 21992 1013 22007
rect 1071 21992 1131 22007
rect 1189 21992 1249 22007
rect 1420 22007 1716 22046
rect 1420 21992 1480 22007
rect 1538 21992 1598 22007
rect 1656 21992 1716 22007
rect 1774 22007 2070 22046
rect 1774 21992 1834 22007
rect 1892 21992 1952 22007
rect 2010 21992 2070 22007
rect 2247 22007 2543 22046
rect 2247 21992 2307 22007
rect 2365 21992 2425 22007
rect 2483 21992 2543 22007
rect 4097 22007 4393 22046
rect 4097 21992 4157 22007
rect 4215 21992 4275 22007
rect 4333 21992 4393 22007
rect 4564 22007 4860 22046
rect 4564 21992 4624 22007
rect 4682 21992 4742 22007
rect 4800 21992 4860 22007
rect 4918 22007 5214 22046
rect 4918 21992 4978 22007
rect 5036 21992 5096 22007
rect 5154 21992 5214 22007
rect 5391 22007 5687 22046
rect 5391 21992 5451 22007
rect 5509 21992 5569 22007
rect 5627 21992 5687 22007
rect 7229 22011 7525 22050
rect 7229 21996 7289 22011
rect 7347 21996 7407 22011
rect 7465 21996 7525 22011
rect 7696 22011 7992 22050
rect 7696 21996 7756 22011
rect 7814 21996 7874 22011
rect 7932 21996 7992 22011
rect 8050 22011 8346 22050
rect 8050 21996 8110 22011
rect 8168 21996 8228 22011
rect 8286 21996 8346 22011
rect 8523 22011 8819 22050
rect 8523 21996 8583 22011
rect 8641 21996 8701 22011
rect 8759 21996 8819 22011
rect 10373 22011 10669 22050
rect 10373 21996 10433 22011
rect 10491 21996 10551 22011
rect 10609 21996 10669 22011
rect 10840 22011 11136 22050
rect 10840 21996 10900 22011
rect 10958 21996 11018 22011
rect 11076 21996 11136 22011
rect 11194 22011 11490 22050
rect 11194 21996 11254 22011
rect 11312 21996 11372 22011
rect 11430 21996 11490 22011
rect 11667 22011 11963 22050
rect 11667 21996 11727 22011
rect 11785 21996 11845 22011
rect 11903 21996 11963 22011
rect 13575 22007 13871 22046
rect 512 21808 808 21847
rect 512 21792 572 21808
rect 630 21792 690 21808
rect 748 21792 808 21808
rect 2720 21808 3016 21847
rect 2720 21792 2780 21808
rect 2838 21792 2898 21808
rect 2956 21792 3016 21808
rect 3656 21808 3952 21847
rect 3656 21792 3716 21808
rect 3774 21792 3834 21808
rect 3892 21792 3952 21808
rect 5864 21808 6160 21847
rect 5864 21792 5924 21808
rect 5982 21792 6042 21808
rect 6100 21792 6160 21808
rect 6788 21812 7084 21851
rect 6788 21796 6848 21812
rect 6906 21796 6966 21812
rect 7024 21796 7084 21812
rect 8996 21812 9292 21851
rect 8996 21796 9056 21812
rect 9114 21796 9174 21812
rect 9232 21796 9292 21812
rect 9932 21812 10228 21851
rect 9932 21796 9992 21812
rect 10050 21796 10110 21812
rect 10168 21796 10228 21812
rect 13575 21992 13635 22007
rect 13693 21992 13753 22007
rect 13811 21992 13871 22007
rect 14042 22007 14338 22046
rect 14042 21992 14102 22007
rect 14160 21992 14220 22007
rect 14278 21992 14338 22007
rect 14396 22007 14692 22046
rect 14396 21992 14456 22007
rect 14514 21992 14574 22007
rect 14632 21992 14692 22007
rect 14869 22007 15165 22046
rect 14869 21992 14929 22007
rect 14987 21992 15047 22007
rect 15105 21992 15165 22007
rect 16719 22007 17015 22046
rect 16719 21992 16779 22007
rect 16837 21992 16897 22007
rect 16955 21992 17015 22007
rect 17186 22007 17482 22046
rect 17186 21992 17246 22007
rect 17304 21992 17364 22007
rect 17422 21992 17482 22007
rect 17540 22007 17836 22046
rect 17540 21992 17600 22007
rect 17658 21992 17718 22007
rect 17776 21992 17836 22007
rect 18013 22007 18309 22046
rect 18013 21992 18073 22007
rect 18131 21992 18191 22007
rect 18249 21992 18309 22007
rect 19851 22011 20147 22050
rect 19851 21996 19911 22011
rect 19969 21996 20029 22011
rect 20087 21996 20147 22011
rect 20318 22011 20614 22050
rect 20318 21996 20378 22011
rect 20436 21996 20496 22011
rect 20554 21996 20614 22011
rect 20672 22011 20968 22050
rect 20672 21996 20732 22011
rect 20790 21996 20850 22011
rect 20908 21996 20968 22011
rect 21145 22011 21441 22050
rect 21145 21996 21205 22011
rect 21263 21996 21323 22011
rect 21381 21996 21441 22011
rect 22995 22011 23291 22050
rect 22995 21996 23055 22011
rect 23113 21996 23173 22011
rect 23231 21996 23291 22011
rect 23462 22011 23758 22050
rect 23462 21996 23522 22011
rect 23580 21996 23640 22011
rect 23698 21996 23758 22011
rect 23816 22011 24112 22050
rect 23816 21996 23876 22011
rect 23934 21996 23994 22011
rect 24052 21996 24112 22011
rect 24289 22011 24585 22050
rect 24289 21996 24349 22011
rect 24407 21996 24467 22011
rect 24525 21996 24585 22011
rect 12140 21812 12436 21851
rect 12140 21796 12200 21812
rect 12258 21796 12318 21812
rect 12376 21796 12436 21812
rect 13134 21808 13430 21847
rect 13134 21792 13194 21808
rect 13252 21792 13312 21808
rect 13370 21792 13430 21808
rect 512 21306 572 21592
rect 630 21566 690 21592
rect 748 21566 808 21592
rect 953 21566 1013 21592
rect 512 21289 648 21306
rect 512 21234 571 21289
rect 629 21234 648 21289
rect 512 21219 648 21234
rect 512 20907 572 21219
rect 1071 21174 1131 21592
rect 1189 21566 1249 21592
rect 1420 21566 1480 21592
rect 1538 21566 1598 21592
rect 1656 21566 1716 21592
rect 1774 21566 1834 21592
rect 1539 21406 1598 21566
rect 1539 21405 1602 21406
rect 1536 21389 1602 21405
rect 1536 21355 1552 21389
rect 1586 21355 1602 21389
rect 1536 21339 1602 21355
rect 1639 21290 1734 21305
rect 1639 21235 1658 21290
rect 1716 21267 1734 21290
rect 1892 21267 1952 21592
rect 2010 21566 2070 21592
rect 2247 21566 2307 21592
rect 1716 21235 1952 21267
rect 1639 21218 1952 21235
rect 1071 21117 1598 21174
rect 1538 21018 1598 21117
rect 1527 21005 1608 21018
rect 1527 20950 1540 21005
rect 1598 20950 1608 21005
rect 1527 20939 1608 20950
rect 512 20862 1406 20907
rect 1346 20659 1406 20862
rect 1538 20659 1598 20939
rect 1656 20659 1716 21218
rect 2365 21176 2425 21592
rect 2483 21566 2543 21592
rect 2720 21566 2780 21592
rect 2838 21566 2898 21592
rect 2846 21443 2912 21446
rect 2956 21443 3016 21592
rect 2846 21430 3016 21443
rect 2846 21396 2862 21430
rect 2896 21396 3016 21430
rect 2846 21383 3016 21396
rect 2846 21380 2912 21383
rect 1887 21159 2425 21176
rect 1887 21125 1906 21159
rect 1940 21125 2425 21159
rect 1887 21119 2425 21125
rect 1887 21109 1956 21119
rect 1887 21107 1952 21109
rect 1771 20769 1837 20785
rect 1771 20735 1787 20769
rect 1821 20735 1837 20769
rect 1771 20719 1837 20735
rect 1774 20659 1834 20719
rect 1892 20659 1952 21107
rect 2956 20907 3016 21383
rect 2088 20862 3016 20907
rect 3656 21306 3716 21592
rect 3774 21566 3834 21592
rect 3892 21566 3952 21592
rect 4097 21566 4157 21592
rect 3656 21289 3792 21306
rect 3656 21234 3715 21289
rect 3773 21234 3792 21289
rect 3656 21219 3792 21234
rect 3656 20907 3716 21219
rect 4215 21174 4275 21592
rect 4333 21566 4393 21592
rect 4564 21566 4624 21592
rect 4682 21566 4742 21592
rect 4800 21566 4860 21592
rect 4918 21566 4978 21592
rect 4683 21406 4742 21566
rect 4683 21405 4746 21406
rect 4680 21389 4746 21405
rect 4680 21355 4696 21389
rect 4730 21355 4746 21389
rect 4680 21339 4746 21355
rect 4783 21290 4878 21305
rect 4783 21235 4802 21290
rect 4860 21267 4878 21290
rect 5036 21267 5096 21592
rect 5154 21566 5214 21592
rect 5391 21566 5451 21592
rect 4860 21235 5096 21267
rect 4783 21218 5096 21235
rect 4215 21117 4742 21174
rect 4682 21018 4742 21117
rect 4671 21005 4752 21018
rect 4671 20950 4684 21005
rect 4742 20950 4752 21005
rect 4671 20939 4752 20950
rect 3656 20862 4550 20907
rect 2088 20659 2148 20862
rect 4490 20659 4550 20862
rect 4682 20659 4742 20939
rect 4800 20659 4860 21218
rect 5509 21176 5569 21592
rect 5627 21566 5687 21592
rect 5864 21566 5924 21592
rect 5982 21566 6042 21592
rect 5990 21443 6056 21446
rect 6100 21443 6160 21592
rect 5990 21430 6160 21443
rect 5990 21396 6006 21430
rect 6040 21396 6160 21430
rect 5990 21383 6160 21396
rect 5990 21380 6056 21383
rect 5031 21159 5569 21176
rect 5031 21125 5050 21159
rect 5084 21125 5569 21159
rect 5031 21119 5569 21125
rect 5031 21109 5100 21119
rect 5031 21107 5096 21109
rect 4915 20769 4981 20785
rect 4915 20735 4931 20769
rect 4965 20735 4981 20769
rect 4915 20719 4981 20735
rect 4918 20659 4978 20719
rect 5036 20659 5096 21107
rect 6100 20907 6160 21383
rect 5232 20862 6160 20907
rect 6788 21310 6848 21596
rect 6906 21570 6966 21596
rect 7024 21570 7084 21596
rect 7229 21570 7289 21596
rect 6788 21293 6924 21310
rect 6788 21238 6847 21293
rect 6905 21238 6924 21293
rect 6788 21223 6924 21238
rect 6788 20911 6848 21223
rect 7347 21178 7407 21596
rect 7465 21570 7525 21596
rect 7696 21570 7756 21596
rect 7814 21570 7874 21596
rect 7932 21570 7992 21596
rect 8050 21570 8110 21596
rect 7815 21410 7874 21570
rect 7815 21409 7878 21410
rect 7812 21393 7878 21409
rect 7812 21359 7828 21393
rect 7862 21359 7878 21393
rect 7812 21343 7878 21359
rect 7915 21294 8010 21309
rect 7915 21239 7934 21294
rect 7992 21271 8010 21294
rect 8168 21271 8228 21596
rect 8286 21570 8346 21596
rect 8523 21570 8583 21596
rect 7992 21239 8228 21271
rect 7915 21222 8228 21239
rect 7347 21121 7874 21178
rect 7814 21022 7874 21121
rect 7803 21009 7884 21022
rect 7803 20954 7816 21009
rect 7874 20954 7884 21009
rect 7803 20943 7884 20954
rect 6788 20866 7682 20911
rect 5232 20659 5292 20862
rect 7622 20663 7682 20866
rect 7814 20663 7874 20943
rect 7932 20663 7992 21222
rect 8641 21180 8701 21596
rect 8759 21570 8819 21596
rect 8996 21570 9056 21596
rect 9114 21570 9174 21596
rect 9122 21447 9188 21450
rect 9232 21447 9292 21596
rect 9122 21434 9292 21447
rect 9122 21400 9138 21434
rect 9172 21400 9292 21434
rect 9122 21387 9292 21400
rect 9122 21384 9188 21387
rect 8163 21163 8701 21180
rect 8163 21129 8182 21163
rect 8216 21129 8701 21163
rect 8163 21123 8701 21129
rect 8163 21113 8232 21123
rect 8163 21111 8228 21113
rect 8047 20773 8113 20789
rect 8047 20739 8063 20773
rect 8097 20739 8113 20773
rect 8047 20723 8113 20739
rect 8050 20663 8110 20723
rect 8168 20663 8228 21111
rect 9232 20911 9292 21387
rect 8364 20866 9292 20911
rect 9932 21310 9992 21596
rect 10050 21570 10110 21596
rect 10168 21570 10228 21596
rect 10373 21570 10433 21596
rect 9932 21293 10068 21310
rect 9932 21238 9991 21293
rect 10049 21238 10068 21293
rect 9932 21223 10068 21238
rect 9932 20911 9992 21223
rect 10491 21178 10551 21596
rect 10609 21570 10669 21596
rect 10840 21570 10900 21596
rect 10958 21570 11018 21596
rect 11076 21570 11136 21596
rect 11194 21570 11254 21596
rect 10959 21410 11018 21570
rect 10959 21409 11022 21410
rect 10956 21393 11022 21409
rect 10956 21359 10972 21393
rect 11006 21359 11022 21393
rect 10956 21343 11022 21359
rect 11059 21294 11154 21309
rect 11059 21239 11078 21294
rect 11136 21271 11154 21294
rect 11312 21271 11372 21596
rect 11430 21570 11490 21596
rect 11667 21570 11727 21596
rect 11136 21239 11372 21271
rect 11059 21222 11372 21239
rect 10491 21121 11018 21178
rect 10958 21022 11018 21121
rect 10947 21009 11028 21022
rect 10947 20954 10960 21009
rect 11018 20954 11028 21009
rect 10947 20943 11028 20954
rect 9932 20866 10826 20911
rect 8364 20663 8424 20866
rect 10766 20663 10826 20866
rect 10958 20663 11018 20943
rect 11076 20663 11136 21222
rect 11785 21180 11845 21596
rect 11903 21570 11963 21596
rect 12140 21570 12200 21596
rect 12258 21570 12318 21596
rect 12266 21447 12332 21450
rect 12376 21447 12436 21596
rect 15342 21808 15638 21847
rect 15342 21792 15402 21808
rect 15460 21792 15520 21808
rect 15578 21792 15638 21808
rect 16278 21808 16574 21847
rect 16278 21792 16338 21808
rect 16396 21792 16456 21808
rect 16514 21792 16574 21808
rect 18486 21808 18782 21847
rect 18486 21792 18546 21808
rect 18604 21792 18664 21808
rect 18722 21792 18782 21808
rect 19410 21812 19706 21851
rect 19410 21796 19470 21812
rect 19528 21796 19588 21812
rect 19646 21796 19706 21812
rect 21618 21812 21914 21851
rect 21618 21796 21678 21812
rect 21736 21796 21796 21812
rect 21854 21796 21914 21812
rect 22554 21812 22850 21851
rect 22554 21796 22614 21812
rect 22672 21796 22732 21812
rect 22790 21796 22850 21812
rect 24762 21812 25058 21851
rect 24762 21796 24822 21812
rect 24880 21796 24940 21812
rect 24998 21796 25058 21812
rect 12266 21434 12436 21447
rect 12266 21400 12282 21434
rect 12316 21400 12436 21434
rect 12266 21387 12436 21400
rect 12266 21384 12332 21387
rect 11307 21163 11845 21180
rect 11307 21129 11326 21163
rect 11360 21129 11845 21163
rect 11307 21123 11845 21129
rect 11307 21113 11376 21123
rect 11307 21111 11372 21113
rect 11191 20773 11257 20789
rect 11191 20739 11207 20773
rect 11241 20739 11257 20773
rect 11191 20723 11257 20739
rect 11194 20663 11254 20723
rect 11312 20663 11372 21111
rect 12376 20911 12436 21387
rect 11508 20866 12436 20911
rect 13134 21306 13194 21592
rect 13252 21566 13312 21592
rect 13370 21566 13430 21592
rect 13575 21566 13635 21592
rect 13134 21289 13270 21306
rect 13134 21234 13193 21289
rect 13251 21234 13270 21289
rect 13134 21219 13270 21234
rect 13134 20907 13194 21219
rect 13693 21174 13753 21592
rect 13811 21566 13871 21592
rect 14042 21566 14102 21592
rect 14160 21566 14220 21592
rect 14278 21566 14338 21592
rect 14396 21566 14456 21592
rect 14161 21406 14220 21566
rect 14161 21405 14224 21406
rect 14158 21389 14224 21405
rect 14158 21355 14174 21389
rect 14208 21355 14224 21389
rect 14158 21339 14224 21355
rect 14261 21290 14356 21305
rect 14261 21235 14280 21290
rect 14338 21267 14356 21290
rect 14514 21267 14574 21592
rect 14632 21566 14692 21592
rect 14869 21566 14929 21592
rect 14338 21235 14574 21267
rect 14261 21218 14574 21235
rect 13693 21117 14220 21174
rect 14160 21018 14220 21117
rect 14149 21005 14230 21018
rect 14149 20950 14162 21005
rect 14220 20950 14230 21005
rect 14149 20939 14230 20950
rect 11508 20663 11568 20866
rect 13134 20862 14028 20907
rect 1346 20433 1406 20459
rect 1538 20233 1598 20259
rect 1656 20233 1716 20259
rect 1774 20233 1834 20259
rect 1892 20233 1952 20259
rect 1713 20178 1779 20186
rect 2088 20178 2148 20459
rect 4490 20433 4550 20459
rect 4682 20233 4742 20259
rect 4800 20233 4860 20259
rect 4918 20233 4978 20259
rect 5036 20233 5096 20259
rect 1713 20170 2148 20178
rect 1713 20136 1729 20170
rect 1763 20136 2148 20170
rect 1713 20127 2148 20136
rect 4857 20178 4923 20186
rect 5232 20178 5292 20459
rect 7622 20437 7682 20463
rect 7814 20237 7874 20263
rect 7932 20237 7992 20263
rect 8050 20237 8110 20263
rect 8168 20237 8228 20263
rect 4857 20170 5292 20178
rect 4857 20136 4873 20170
rect 4907 20136 5292 20170
rect 4857 20127 5292 20136
rect 7989 20182 8055 20190
rect 8364 20182 8424 20463
rect 10766 20437 10826 20463
rect 13968 20659 14028 20862
rect 14160 20659 14220 20939
rect 14278 20659 14338 21218
rect 14987 21176 15047 21592
rect 15105 21566 15165 21592
rect 15342 21566 15402 21592
rect 15460 21566 15520 21592
rect 15468 21443 15534 21446
rect 15578 21443 15638 21592
rect 15468 21430 15638 21443
rect 15468 21396 15484 21430
rect 15518 21396 15638 21430
rect 15468 21383 15638 21396
rect 15468 21380 15534 21383
rect 14509 21159 15047 21176
rect 14509 21125 14528 21159
rect 14562 21125 15047 21159
rect 14509 21119 15047 21125
rect 14509 21109 14578 21119
rect 14509 21107 14574 21109
rect 14393 20769 14459 20785
rect 14393 20735 14409 20769
rect 14443 20735 14459 20769
rect 14393 20719 14459 20735
rect 14396 20659 14456 20719
rect 14514 20659 14574 21107
rect 15578 20907 15638 21383
rect 14710 20862 15638 20907
rect 16278 21306 16338 21592
rect 16396 21566 16456 21592
rect 16514 21566 16574 21592
rect 16719 21566 16779 21592
rect 16278 21289 16414 21306
rect 16278 21234 16337 21289
rect 16395 21234 16414 21289
rect 16278 21219 16414 21234
rect 16278 20907 16338 21219
rect 16837 21174 16897 21592
rect 16955 21566 17015 21592
rect 17186 21566 17246 21592
rect 17304 21566 17364 21592
rect 17422 21566 17482 21592
rect 17540 21566 17600 21592
rect 17305 21406 17364 21566
rect 17305 21405 17368 21406
rect 17302 21389 17368 21405
rect 17302 21355 17318 21389
rect 17352 21355 17368 21389
rect 17302 21339 17368 21355
rect 17405 21290 17500 21305
rect 17405 21235 17424 21290
rect 17482 21267 17500 21290
rect 17658 21267 17718 21592
rect 17776 21566 17836 21592
rect 18013 21566 18073 21592
rect 17482 21235 17718 21267
rect 17405 21218 17718 21235
rect 16837 21117 17364 21174
rect 17304 21018 17364 21117
rect 17293 21005 17374 21018
rect 17293 20950 17306 21005
rect 17364 20950 17374 21005
rect 17293 20939 17374 20950
rect 16278 20862 17172 20907
rect 14710 20659 14770 20862
rect 17112 20659 17172 20862
rect 17304 20659 17364 20939
rect 17422 20659 17482 21218
rect 18131 21176 18191 21592
rect 18249 21566 18309 21592
rect 18486 21566 18546 21592
rect 18604 21566 18664 21592
rect 18612 21443 18678 21446
rect 18722 21443 18782 21592
rect 18612 21430 18782 21443
rect 18612 21396 18628 21430
rect 18662 21396 18782 21430
rect 18612 21383 18782 21396
rect 18612 21380 18678 21383
rect 17653 21159 18191 21176
rect 17653 21125 17672 21159
rect 17706 21125 18191 21159
rect 17653 21119 18191 21125
rect 17653 21109 17722 21119
rect 17653 21107 17718 21109
rect 17537 20769 17603 20785
rect 17537 20735 17553 20769
rect 17587 20735 17603 20769
rect 17537 20719 17603 20735
rect 17540 20659 17600 20719
rect 17658 20659 17718 21107
rect 18722 20907 18782 21383
rect 17854 20862 18782 20907
rect 19410 21310 19470 21596
rect 19528 21570 19588 21596
rect 19646 21570 19706 21596
rect 19851 21570 19911 21596
rect 19410 21293 19546 21310
rect 19410 21238 19469 21293
rect 19527 21238 19546 21293
rect 19410 21223 19546 21238
rect 19410 20911 19470 21223
rect 19969 21178 20029 21596
rect 20087 21570 20147 21596
rect 20318 21570 20378 21596
rect 20436 21570 20496 21596
rect 20554 21570 20614 21596
rect 20672 21570 20732 21596
rect 20437 21410 20496 21570
rect 20437 21409 20500 21410
rect 20434 21393 20500 21409
rect 20434 21359 20450 21393
rect 20484 21359 20500 21393
rect 20434 21343 20500 21359
rect 20537 21294 20632 21309
rect 20537 21239 20556 21294
rect 20614 21271 20632 21294
rect 20790 21271 20850 21596
rect 20908 21570 20968 21596
rect 21145 21570 21205 21596
rect 20614 21239 20850 21271
rect 20537 21222 20850 21239
rect 19969 21121 20496 21178
rect 20436 21022 20496 21121
rect 20425 21009 20506 21022
rect 20425 20954 20438 21009
rect 20496 20954 20506 21009
rect 20425 20943 20506 20954
rect 19410 20866 20304 20911
rect 17854 20659 17914 20862
rect 20244 20663 20304 20866
rect 20436 20663 20496 20943
rect 20554 20663 20614 21222
rect 21263 21180 21323 21596
rect 21381 21570 21441 21596
rect 21618 21570 21678 21596
rect 21736 21570 21796 21596
rect 21744 21447 21810 21450
rect 21854 21447 21914 21596
rect 21744 21434 21914 21447
rect 21744 21400 21760 21434
rect 21794 21400 21914 21434
rect 21744 21387 21914 21400
rect 21744 21384 21810 21387
rect 20785 21163 21323 21180
rect 20785 21129 20804 21163
rect 20838 21129 21323 21163
rect 20785 21123 21323 21129
rect 20785 21113 20854 21123
rect 20785 21111 20850 21113
rect 20669 20773 20735 20789
rect 20669 20739 20685 20773
rect 20719 20739 20735 20773
rect 20669 20723 20735 20739
rect 20672 20663 20732 20723
rect 20790 20663 20850 21111
rect 21854 20911 21914 21387
rect 20986 20866 21914 20911
rect 22554 21310 22614 21596
rect 22672 21570 22732 21596
rect 22790 21570 22850 21596
rect 22995 21570 23055 21596
rect 22554 21293 22690 21310
rect 22554 21238 22613 21293
rect 22671 21238 22690 21293
rect 22554 21223 22690 21238
rect 22554 20911 22614 21223
rect 23113 21178 23173 21596
rect 23231 21570 23291 21596
rect 23462 21570 23522 21596
rect 23580 21570 23640 21596
rect 23698 21570 23758 21596
rect 23816 21570 23876 21596
rect 23581 21410 23640 21570
rect 23581 21409 23644 21410
rect 23578 21393 23644 21409
rect 23578 21359 23594 21393
rect 23628 21359 23644 21393
rect 23578 21343 23644 21359
rect 23681 21294 23776 21309
rect 23681 21239 23700 21294
rect 23758 21271 23776 21294
rect 23934 21271 23994 21596
rect 24052 21570 24112 21596
rect 24289 21570 24349 21596
rect 23758 21239 23994 21271
rect 23681 21222 23994 21239
rect 23113 21121 23640 21178
rect 23580 21022 23640 21121
rect 23569 21009 23650 21022
rect 23569 20954 23582 21009
rect 23640 20954 23650 21009
rect 23569 20943 23650 20954
rect 22554 20866 23448 20911
rect 20986 20663 21046 20866
rect 23388 20663 23448 20866
rect 23580 20663 23640 20943
rect 23698 20663 23758 21222
rect 24407 21180 24467 21596
rect 24525 21570 24585 21596
rect 24762 21570 24822 21596
rect 24880 21570 24940 21596
rect 24888 21447 24954 21450
rect 24998 21447 25058 21596
rect 24888 21434 25058 21447
rect 24888 21400 24904 21434
rect 24938 21400 25058 21434
rect 24888 21387 25058 21400
rect 24888 21384 24954 21387
rect 23929 21163 24467 21180
rect 23929 21129 23948 21163
rect 23982 21129 24467 21163
rect 23929 21123 24467 21129
rect 23929 21113 23998 21123
rect 23929 21111 23994 21113
rect 23813 20773 23879 20789
rect 23813 20739 23829 20773
rect 23863 20739 23879 20773
rect 23813 20723 23879 20739
rect 23816 20663 23876 20723
rect 23934 20663 23994 21111
rect 24998 20911 25058 21387
rect 24130 20866 25058 20911
rect 24130 20663 24190 20866
rect 10958 20237 11018 20263
rect 11076 20237 11136 20263
rect 11194 20237 11254 20263
rect 11312 20237 11372 20263
rect 7989 20174 8424 20182
rect 7989 20140 8005 20174
rect 8039 20140 8424 20174
rect 7989 20131 8424 20140
rect 11133 20182 11199 20190
rect 11508 20182 11568 20463
rect 13968 20433 14028 20459
rect 14160 20233 14220 20259
rect 14278 20233 14338 20259
rect 14396 20233 14456 20259
rect 14514 20233 14574 20259
rect 11133 20174 11568 20182
rect 11133 20140 11149 20174
rect 11183 20140 11568 20174
rect 11133 20131 11568 20140
rect 14335 20178 14401 20186
rect 14710 20178 14770 20459
rect 17112 20433 17172 20459
rect 17304 20233 17364 20259
rect 17422 20233 17482 20259
rect 17540 20233 17600 20259
rect 17658 20233 17718 20259
rect 14335 20170 14770 20178
rect 14335 20136 14351 20170
rect 14385 20136 14770 20170
rect 1713 20120 1779 20127
rect 4857 20120 4923 20127
rect 7989 20124 8055 20131
rect 11133 20124 11199 20131
rect 14335 20127 14770 20136
rect 17479 20178 17545 20186
rect 17854 20178 17914 20459
rect 20244 20437 20304 20463
rect 20436 20237 20496 20263
rect 20554 20237 20614 20263
rect 20672 20237 20732 20263
rect 20790 20237 20850 20263
rect 17479 20170 17914 20178
rect 17479 20136 17495 20170
rect 17529 20136 17914 20170
rect 17479 20127 17914 20136
rect 20611 20182 20677 20190
rect 20986 20182 21046 20463
rect 23388 20437 23448 20463
rect 23580 20237 23640 20263
rect 23698 20237 23758 20263
rect 23816 20237 23876 20263
rect 23934 20237 23994 20263
rect 20611 20174 21046 20182
rect 20611 20140 20627 20174
rect 20661 20140 21046 20174
rect 20611 20131 21046 20140
rect 23755 20182 23821 20190
rect 24130 20182 24190 20463
rect 23755 20174 24190 20182
rect 23755 20140 23771 20174
rect 23805 20140 24190 20174
rect 23755 20131 24190 20140
rect 14335 20120 14401 20127
rect 17479 20120 17545 20127
rect 20611 20124 20677 20131
rect 23755 20124 23821 20131
rect 14566 16968 14632 16984
rect 14566 16934 14582 16968
rect 14616 16964 14632 16968
rect 14616 16934 15116 16964
rect 15734 16968 15800 16984
rect 14566 16921 15116 16934
rect 14566 16918 14632 16921
rect 14566 16869 14632 16876
rect 15072 16869 15116 16921
rect 15734 16934 15750 16968
rect 15784 16964 15800 16968
rect 15784 16934 16284 16964
rect 16902 16968 16968 16984
rect 15734 16921 16284 16934
rect 15734 16918 15800 16921
rect 15734 16869 15800 16876
rect 16240 16869 16284 16921
rect 16902 16934 16918 16968
rect 16952 16964 16968 16968
rect 16952 16934 17452 16964
rect 18070 16968 18136 16984
rect 16902 16921 17452 16934
rect 16902 16918 16968 16921
rect 16902 16869 16968 16876
rect 17408 16869 17452 16921
rect 18070 16934 18086 16968
rect 18120 16964 18136 16968
rect 18120 16934 18620 16964
rect 19244 16970 19310 16986
rect 18070 16921 18620 16934
rect 18070 16918 18136 16921
rect 18070 16869 18136 16876
rect 18576 16869 18620 16921
rect 19244 16936 19260 16970
rect 19294 16966 19310 16970
rect 19294 16936 19794 16966
rect 20412 16970 20478 16986
rect 19244 16923 19794 16936
rect 19244 16920 19310 16923
rect 19244 16871 19310 16878
rect 19750 16871 19794 16923
rect 20412 16936 20428 16970
rect 20462 16966 20478 16970
rect 20462 16936 20962 16966
rect 21580 16970 21646 16986
rect 20412 16923 20962 16936
rect 20412 16920 20478 16923
rect 20412 16871 20478 16878
rect 20918 16871 20962 16923
rect 21580 16936 21596 16970
rect 21630 16966 21646 16970
rect 21630 16936 22130 16966
rect 22748 16970 22814 16986
rect 21580 16923 22130 16936
rect 21580 16920 21646 16923
rect 21580 16871 21646 16878
rect 22086 16871 22130 16923
rect 22748 16936 22764 16970
rect 22798 16966 22814 16970
rect 22798 16936 23298 16966
rect 22748 16923 23298 16936
rect 22748 16920 22814 16923
rect 22748 16871 22814 16878
rect 23254 16871 23298 16923
rect 14566 16860 15014 16869
rect 14566 16826 14582 16860
rect 14616 16828 15014 16860
rect 14616 16827 14778 16828
rect 14616 16826 14632 16827
rect 14566 16810 14632 16826
rect 14718 16808 14778 16827
rect 14836 16808 14896 16828
rect 14954 16808 15014 16828
rect 15072 16828 15368 16869
rect 15072 16808 15132 16828
rect 15190 16808 15250 16828
rect 15308 16808 15368 16828
rect 15734 16860 16182 16869
rect 15734 16826 15750 16860
rect 15784 16828 16182 16860
rect 15784 16827 15946 16828
rect 15784 16826 15800 16827
rect 15734 16810 15800 16826
rect 15886 16808 15946 16827
rect 16004 16808 16064 16828
rect 16122 16808 16182 16828
rect 16240 16828 16536 16869
rect 16240 16808 16300 16828
rect 16358 16808 16418 16828
rect 16476 16808 16536 16828
rect 16902 16860 17350 16869
rect 16902 16826 16918 16860
rect 16952 16828 17350 16860
rect 16952 16827 17114 16828
rect 16952 16826 16968 16827
rect 16902 16810 16968 16826
rect 2955 16632 3251 16668
rect 2955 16611 3015 16632
rect 3073 16611 3133 16632
rect 3191 16611 3251 16632
rect 3309 16631 3605 16667
rect 3309 16611 3369 16631
rect 3427 16611 3487 16631
rect 3545 16611 3605 16631
rect 3663 16631 3959 16667
rect 3663 16611 3723 16631
rect 3781 16611 3841 16631
rect 3899 16611 3959 16631
rect 4403 16632 4699 16668
rect 4403 16611 4463 16632
rect 4521 16611 4581 16632
rect 4639 16611 4699 16632
rect 4757 16631 5053 16667
rect 4757 16611 4817 16631
rect 4875 16611 4935 16631
rect 4993 16611 5053 16631
rect 5111 16631 5407 16667
rect 5111 16611 5171 16631
rect 5229 16611 5289 16631
rect 5347 16611 5407 16631
rect 5901 16634 6197 16670
rect 5901 16613 5961 16634
rect 6019 16613 6079 16634
rect 6137 16613 6197 16634
rect 6255 16633 6551 16669
rect 6255 16613 6315 16633
rect 6373 16613 6433 16633
rect 6491 16613 6551 16633
rect 6609 16633 6905 16669
rect 6609 16613 6669 16633
rect 6727 16613 6787 16633
rect 6845 16613 6905 16633
rect 7349 16634 7645 16670
rect 7349 16613 7409 16634
rect 7467 16613 7527 16634
rect 7585 16613 7645 16634
rect 7703 16633 7999 16669
rect 7703 16613 7763 16633
rect 7821 16613 7881 16633
rect 7939 16613 7999 16633
rect 8057 16633 8353 16669
rect 8057 16613 8117 16633
rect 8175 16613 8235 16633
rect 8293 16613 8353 16633
rect 8869 16632 9165 16668
rect 8869 16611 8929 16632
rect 8987 16611 9047 16632
rect 9105 16611 9165 16632
rect 9223 16631 9519 16667
rect 9223 16611 9283 16631
rect 9341 16611 9401 16631
rect 9459 16611 9519 16631
rect 9577 16631 9873 16667
rect 9577 16611 9637 16631
rect 9695 16611 9755 16631
rect 9813 16611 9873 16631
rect 10317 16632 10613 16668
rect 10317 16611 10377 16632
rect 10435 16611 10495 16632
rect 10553 16611 10613 16632
rect 10671 16631 10967 16667
rect 10671 16611 10731 16631
rect 10789 16611 10849 16631
rect 10907 16611 10967 16631
rect 11025 16631 11321 16667
rect 11025 16611 11085 16631
rect 11143 16611 11203 16631
rect 11261 16611 11321 16631
rect 11815 16634 12111 16670
rect 11815 16613 11875 16634
rect 11933 16613 11993 16634
rect 12051 16613 12111 16634
rect 12169 16633 12465 16669
rect 12169 16613 12229 16633
rect 12287 16613 12347 16633
rect 12405 16613 12465 16633
rect 12523 16633 12819 16669
rect 12523 16613 12583 16633
rect 12641 16613 12701 16633
rect 12759 16613 12819 16633
rect 13263 16634 13559 16670
rect 13263 16613 13323 16634
rect 13381 16613 13441 16634
rect 13499 16613 13559 16634
rect 13617 16633 13913 16669
rect 13617 16613 13677 16633
rect 13735 16613 13795 16633
rect 13853 16613 13913 16633
rect 13971 16633 14267 16669
rect 13971 16613 14031 16633
rect 14089 16613 14149 16633
rect 14207 16613 14267 16633
rect 2955 16385 3015 16411
rect 3073 16385 3133 16411
rect 3191 16385 3251 16411
rect 3309 16391 3369 16411
rect 3309 16385 3370 16391
rect 3427 16385 3487 16411
rect 3545 16385 3605 16411
rect 3192 16200 3250 16385
rect 3192 16174 3252 16200
rect 3310 16174 3370 16385
rect 3663 16379 3723 16411
rect 3781 16385 3841 16411
rect 3899 16385 3959 16411
rect 4403 16385 4463 16411
rect 4521 16385 4581 16411
rect 4639 16385 4699 16411
rect 4757 16391 4817 16411
rect 4757 16385 4818 16391
rect 4875 16385 4935 16411
rect 4993 16385 5053 16411
rect 3660 16363 3726 16379
rect 3660 16329 3676 16363
rect 3710 16329 3726 16363
rect 3660 16313 3726 16329
rect 3542 16246 3608 16262
rect 3542 16212 3558 16246
rect 3592 16212 3608 16246
rect 3542 16196 3608 16212
rect 4640 16200 4698 16385
rect 3545 16174 3605 16196
rect 4640 16174 4700 16200
rect 4758 16174 4818 16385
rect 5111 16379 5171 16411
rect 5229 16385 5289 16411
rect 5347 16385 5407 16411
rect 5901 16387 5961 16413
rect 6019 16387 6079 16413
rect 6137 16387 6197 16413
rect 6255 16393 6315 16413
rect 6255 16387 6316 16393
rect 6373 16387 6433 16413
rect 6491 16387 6551 16413
rect 5108 16363 5174 16379
rect 5108 16329 5124 16363
rect 5158 16329 5174 16363
rect 5108 16313 5174 16329
rect 4990 16246 5056 16262
rect 4990 16212 5006 16246
rect 5040 16212 5056 16246
rect 4990 16196 5056 16212
rect 6138 16202 6196 16387
rect 4993 16174 5053 16196
rect 6138 16176 6198 16202
rect 6256 16176 6316 16387
rect 6609 16381 6669 16413
rect 6727 16387 6787 16413
rect 6845 16387 6905 16413
rect 7349 16387 7409 16413
rect 7467 16387 7527 16413
rect 7585 16387 7645 16413
rect 7703 16393 7763 16413
rect 7703 16387 7764 16393
rect 7821 16387 7881 16413
rect 7939 16387 7999 16413
rect 6606 16365 6672 16381
rect 6606 16331 6622 16365
rect 6656 16331 6672 16365
rect 6606 16315 6672 16331
rect 6488 16248 6554 16264
rect 6488 16214 6504 16248
rect 6538 16214 6554 16248
rect 6488 16198 6554 16214
rect 7586 16202 7644 16387
rect 6491 16176 6551 16198
rect 7586 16176 7646 16202
rect 7704 16176 7764 16387
rect 8057 16381 8117 16413
rect 8175 16387 8235 16413
rect 8293 16387 8353 16413
rect 8869 16385 8929 16411
rect 8987 16385 9047 16411
rect 9105 16385 9165 16411
rect 9223 16391 9283 16411
rect 9223 16385 9284 16391
rect 9341 16385 9401 16411
rect 9459 16385 9519 16411
rect 8054 16365 8120 16381
rect 8054 16331 8070 16365
rect 8104 16331 8120 16365
rect 8054 16315 8120 16331
rect 7936 16248 8002 16264
rect 7936 16214 7952 16248
rect 7986 16214 8002 16248
rect 7936 16198 8002 16214
rect 9106 16200 9164 16385
rect 7939 16176 7999 16198
rect 3545 15948 3605 15974
rect 4993 15948 5053 15974
rect 6491 15950 6551 15976
rect 9106 16174 9166 16200
rect 9224 16174 9284 16385
rect 9577 16379 9637 16411
rect 9695 16385 9755 16411
rect 9813 16385 9873 16411
rect 10317 16385 10377 16411
rect 10435 16385 10495 16411
rect 10553 16385 10613 16411
rect 10671 16391 10731 16411
rect 10671 16385 10732 16391
rect 10789 16385 10849 16411
rect 10907 16385 10967 16411
rect 9574 16363 9640 16379
rect 9574 16329 9590 16363
rect 9624 16329 9640 16363
rect 9574 16313 9640 16329
rect 9456 16246 9522 16262
rect 9456 16212 9472 16246
rect 9506 16212 9522 16246
rect 9456 16196 9522 16212
rect 10554 16200 10612 16385
rect 9459 16174 9519 16196
rect 10554 16174 10614 16200
rect 10672 16174 10732 16385
rect 11025 16379 11085 16411
rect 11143 16385 11203 16411
rect 11261 16385 11321 16411
rect 11815 16387 11875 16413
rect 11933 16387 11993 16413
rect 12051 16387 12111 16413
rect 12169 16393 12229 16413
rect 12169 16387 12230 16393
rect 12287 16387 12347 16413
rect 12405 16387 12465 16413
rect 11022 16363 11088 16379
rect 11022 16329 11038 16363
rect 11072 16329 11088 16363
rect 11022 16313 11088 16329
rect 10904 16246 10970 16262
rect 10904 16212 10920 16246
rect 10954 16212 10970 16246
rect 10904 16196 10970 16212
rect 12052 16202 12110 16387
rect 10907 16174 10967 16196
rect 12052 16176 12112 16202
rect 12170 16176 12230 16387
rect 12523 16381 12583 16413
rect 12641 16387 12701 16413
rect 12759 16387 12819 16413
rect 13263 16387 13323 16413
rect 13381 16387 13441 16413
rect 13499 16387 13559 16413
rect 13617 16393 13677 16413
rect 13617 16387 13678 16393
rect 13735 16387 13795 16413
rect 13853 16387 13913 16413
rect 12520 16365 12586 16381
rect 12520 16331 12536 16365
rect 12570 16331 12586 16365
rect 12520 16315 12586 16331
rect 12402 16248 12468 16264
rect 12402 16214 12418 16248
rect 12452 16214 12468 16248
rect 12402 16198 12468 16214
rect 13500 16202 13558 16387
rect 12405 16176 12465 16198
rect 13500 16176 13560 16202
rect 13618 16176 13678 16387
rect 13971 16381 14031 16413
rect 14089 16387 14149 16413
rect 14207 16387 14267 16413
rect 17054 16806 17114 16827
rect 17172 16806 17232 16828
rect 17290 16806 17350 16828
rect 17408 16828 17704 16869
rect 17408 16806 17468 16828
rect 17526 16806 17586 16828
rect 17644 16806 17704 16828
rect 18070 16860 18518 16869
rect 18070 16826 18086 16860
rect 18120 16828 18518 16860
rect 18120 16827 18282 16828
rect 18120 16826 18136 16827
rect 18070 16810 18136 16826
rect 18222 16808 18282 16827
rect 18340 16808 18400 16828
rect 18458 16808 18518 16828
rect 18576 16828 18872 16869
rect 18576 16808 18636 16828
rect 18694 16808 18754 16828
rect 18812 16808 18872 16828
rect 19244 16862 19692 16871
rect 19244 16828 19260 16862
rect 19294 16830 19692 16862
rect 19294 16829 19456 16830
rect 19294 16828 19310 16829
rect 19244 16812 19310 16828
rect 19396 16810 19456 16829
rect 19514 16810 19574 16830
rect 19632 16810 19692 16830
rect 19750 16830 20046 16871
rect 19750 16810 19810 16830
rect 19868 16810 19928 16830
rect 19986 16810 20046 16830
rect 20412 16862 20860 16871
rect 20412 16828 20428 16862
rect 20462 16830 20860 16862
rect 20462 16829 20624 16830
rect 20462 16828 20478 16829
rect 20412 16812 20478 16828
rect 14718 16390 14778 16408
rect 13968 16365 14034 16381
rect 13968 16331 13984 16365
rect 14018 16331 14034 16365
rect 13968 16315 14034 16331
rect 14718 16301 14779 16390
rect 14836 16382 14896 16408
rect 14954 16382 15014 16408
rect 13850 16248 13916 16264
rect 13850 16214 13866 16248
rect 13900 16214 13916 16248
rect 13850 16198 13916 16214
rect 14628 16248 14779 16301
rect 13853 16176 13913 16198
rect 7939 15950 7999 15976
rect 3192 15752 3252 15774
rect 3310 15752 3370 15774
rect 4640 15752 4700 15774
rect 4758 15752 4818 15774
rect 6138 15754 6198 15776
rect 6256 15754 6316 15776
rect 7586 15754 7646 15776
rect 7704 15754 7764 15776
rect 9459 15948 9519 15974
rect 10907 15948 10967 15974
rect 12405 15950 12465 15976
rect 14628 16022 14688 16248
rect 15072 16206 15132 16408
rect 15190 16382 15250 16408
rect 15308 16382 15368 16408
rect 15886 16390 15946 16408
rect 15886 16301 15947 16390
rect 16004 16382 16064 16408
rect 16122 16382 16182 16408
rect 14746 16155 15132 16206
rect 15796 16248 15947 16301
rect 14746 16022 14806 16155
rect 14861 16097 14927 16113
rect 14861 16063 14877 16097
rect 14911 16063 14927 16097
rect 14861 16047 14927 16063
rect 14864 16022 14924 16047
rect 13853 15950 13913 15976
rect 15148 16018 15208 16044
rect 15266 16018 15326 16044
rect 15384 16018 15444 16044
rect 15796 16024 15856 16248
rect 16240 16206 16300 16408
rect 16358 16382 16418 16408
rect 16476 16382 16536 16408
rect 20564 16808 20624 16829
rect 20682 16808 20742 16830
rect 20800 16808 20860 16830
rect 20918 16830 21214 16871
rect 20918 16808 20978 16830
rect 21036 16808 21096 16830
rect 21154 16808 21214 16830
rect 21580 16862 22028 16871
rect 21580 16828 21596 16862
rect 21630 16830 22028 16862
rect 21630 16829 21792 16830
rect 21630 16828 21646 16829
rect 21580 16812 21646 16828
rect 21732 16810 21792 16829
rect 21850 16810 21910 16830
rect 21968 16810 22028 16830
rect 22086 16830 22382 16871
rect 22086 16810 22146 16830
rect 22204 16810 22264 16830
rect 22322 16810 22382 16830
rect 22748 16862 23196 16871
rect 22748 16828 22764 16862
rect 22798 16830 23196 16862
rect 22798 16829 22960 16830
rect 22798 16828 22814 16829
rect 22748 16812 22814 16828
rect 17054 16390 17114 16406
rect 17054 16301 17115 16390
rect 17172 16380 17232 16406
rect 17290 16380 17350 16406
rect 15914 16155 16300 16206
rect 16964 16248 17115 16301
rect 15914 16024 15974 16155
rect 16029 16097 16095 16113
rect 16029 16063 16045 16097
rect 16079 16063 16095 16097
rect 16029 16047 16095 16063
rect 16032 16024 16092 16047
rect 16315 16024 16375 16050
rect 16433 16024 16493 16050
rect 16551 16024 16611 16050
rect 16964 16024 17024 16248
rect 17408 16206 17468 16406
rect 17526 16380 17586 16406
rect 17644 16380 17704 16406
rect 18222 16390 18282 16408
rect 18222 16301 18283 16390
rect 18340 16382 18400 16408
rect 18458 16382 18518 16408
rect 17082 16155 17468 16206
rect 18132 16248 18283 16301
rect 17082 16024 17142 16155
rect 17197 16097 17263 16113
rect 17197 16063 17213 16097
rect 17247 16063 17263 16097
rect 17197 16047 17263 16063
rect 17200 16024 17260 16047
rect 17483 16024 17543 16050
rect 17601 16024 17661 16050
rect 17719 16024 17779 16050
rect 18132 16024 18192 16248
rect 18576 16206 18636 16408
rect 18694 16382 18754 16408
rect 18812 16382 18872 16408
rect 19396 16392 19456 16410
rect 19396 16303 19457 16392
rect 19514 16384 19574 16410
rect 19632 16384 19692 16410
rect 18250 16155 18636 16206
rect 19306 16250 19457 16303
rect 18250 16024 18310 16155
rect 18365 16097 18431 16113
rect 18365 16063 18381 16097
rect 18415 16063 18431 16097
rect 18365 16047 18431 16063
rect 18368 16024 18428 16047
rect 18652 16024 18712 16050
rect 18770 16024 18830 16050
rect 18888 16024 18948 16050
rect 19306 16024 19366 16250
rect 19750 16208 19810 16410
rect 19868 16384 19928 16410
rect 19986 16384 20046 16410
rect 22900 16808 22960 16829
rect 23018 16808 23078 16830
rect 23136 16808 23196 16830
rect 23254 16830 23550 16871
rect 23254 16808 23314 16830
rect 23372 16808 23432 16830
rect 23490 16808 23550 16830
rect 20564 16392 20624 16408
rect 20564 16303 20625 16392
rect 20682 16382 20742 16408
rect 20800 16382 20860 16408
rect 19424 16157 19810 16208
rect 20474 16250 20625 16303
rect 19424 16024 19484 16157
rect 19539 16099 19605 16115
rect 19539 16065 19555 16099
rect 19589 16065 19605 16099
rect 19539 16049 19605 16065
rect 19542 16024 19602 16049
rect 14628 15796 14688 15822
rect 14746 15796 14806 15822
rect 14864 15792 14924 15822
rect 19824 16020 19884 16046
rect 19942 16020 20002 16046
rect 20060 16020 20120 16046
rect 20474 16024 20534 16250
rect 20918 16208 20978 16408
rect 21036 16382 21096 16408
rect 21154 16382 21214 16408
rect 21732 16392 21792 16410
rect 21732 16303 21793 16392
rect 21850 16384 21910 16410
rect 21968 16384 22028 16410
rect 20592 16157 20978 16208
rect 21642 16250 21793 16303
rect 20592 16024 20652 16157
rect 20707 16099 20773 16115
rect 20707 16065 20723 16099
rect 20757 16065 20773 16099
rect 20707 16049 20773 16065
rect 20710 16024 20770 16049
rect 15148 15792 15208 15818
rect 15266 15792 15326 15818
rect 15384 15792 15444 15818
rect 15796 15798 15856 15824
rect 15914 15798 15974 15824
rect 16032 15792 16092 15824
rect 16315 15792 16375 15824
rect 16433 15792 16493 15824
rect 16551 15792 16611 15824
rect 16964 15798 17024 15824
rect 17082 15798 17142 15824
rect 3189 15736 3255 15752
rect 3189 15702 3205 15736
rect 3239 15702 3255 15736
rect 3189 15686 3255 15702
rect 3307 15736 3373 15752
rect 3307 15702 3323 15736
rect 3357 15702 3373 15736
rect 3307 15686 3373 15702
rect 4637 15736 4703 15752
rect 4637 15702 4653 15736
rect 4687 15702 4703 15736
rect 4637 15686 4703 15702
rect 4755 15736 4821 15752
rect 4755 15702 4771 15736
rect 4805 15702 4821 15736
rect 4755 15686 4821 15702
rect 6135 15738 6201 15754
rect 6135 15704 6151 15738
rect 6185 15704 6201 15738
rect 6135 15688 6201 15704
rect 6253 15738 6319 15754
rect 6253 15704 6269 15738
rect 6303 15704 6319 15738
rect 6253 15688 6319 15704
rect 7583 15738 7649 15754
rect 7583 15704 7599 15738
rect 7633 15704 7649 15738
rect 7583 15688 7649 15704
rect 7701 15738 7767 15754
rect 9106 15752 9166 15774
rect 9224 15752 9284 15774
rect 10554 15752 10614 15774
rect 10672 15752 10732 15774
rect 12052 15754 12112 15776
rect 12170 15754 12230 15776
rect 13500 15754 13560 15776
rect 13618 15754 13678 15776
rect 7701 15704 7717 15738
rect 7751 15704 7767 15738
rect 7701 15688 7767 15704
rect 9103 15736 9169 15752
rect 9103 15702 9119 15736
rect 9153 15702 9169 15736
rect 9103 15686 9169 15702
rect 9221 15736 9287 15752
rect 9221 15702 9237 15736
rect 9271 15702 9287 15736
rect 9221 15686 9287 15702
rect 10551 15736 10617 15752
rect 10551 15702 10567 15736
rect 10601 15702 10617 15736
rect 10551 15686 10617 15702
rect 10669 15736 10735 15752
rect 10669 15702 10685 15736
rect 10719 15702 10735 15736
rect 10669 15686 10735 15702
rect 12049 15738 12115 15754
rect 12049 15704 12065 15738
rect 12099 15704 12115 15738
rect 12049 15688 12115 15704
rect 12167 15738 12233 15754
rect 12167 15704 12183 15738
rect 12217 15704 12233 15738
rect 12167 15688 12233 15704
rect 13497 15738 13563 15754
rect 13497 15704 13513 15738
rect 13547 15704 13563 15738
rect 13497 15688 13563 15704
rect 13615 15738 13681 15754
rect 14864 15751 15443 15792
rect 16032 15751 16611 15792
rect 17200 15792 17260 15824
rect 17483 15792 17543 15824
rect 17601 15792 17661 15824
rect 17719 15792 17779 15824
rect 18132 15798 18192 15824
rect 18250 15798 18310 15824
rect 17200 15751 17779 15792
rect 18368 15792 18428 15824
rect 18652 15792 18712 15824
rect 18770 15792 18830 15824
rect 18888 15798 18948 15824
rect 19306 15798 19366 15824
rect 19424 15798 19484 15824
rect 18888 15792 18947 15798
rect 18368 15751 18947 15792
rect 19542 15794 19602 15824
rect 20993 16019 21053 16045
rect 21111 16019 21171 16045
rect 21229 16019 21289 16045
rect 21642 16026 21702 16250
rect 22086 16208 22146 16410
rect 22204 16384 22264 16410
rect 22322 16384 22382 16410
rect 22900 16392 22960 16408
rect 22900 16303 22961 16392
rect 23018 16382 23078 16408
rect 23136 16382 23196 16408
rect 21760 16157 22146 16208
rect 22810 16250 22961 16303
rect 21760 16026 21820 16157
rect 21875 16099 21941 16115
rect 21875 16065 21891 16099
rect 21925 16065 21941 16099
rect 21875 16049 21941 16065
rect 21878 16026 21938 16049
rect 19824 15794 19884 15820
rect 19942 15794 20002 15820
rect 20060 15794 20120 15820
rect 20474 15798 20534 15824
rect 20592 15798 20652 15824
rect 19542 15788 20120 15794
rect 20710 15794 20770 15824
rect 22161 16019 22221 16045
rect 22279 16019 22339 16045
rect 22397 16019 22457 16045
rect 22810 16026 22870 16250
rect 23254 16208 23314 16408
rect 23372 16382 23432 16408
rect 23490 16382 23550 16408
rect 22928 16157 23314 16208
rect 22928 16026 22988 16157
rect 23043 16099 23109 16115
rect 23043 16065 23059 16099
rect 23093 16065 23109 16099
rect 23043 16049 23109 16065
rect 23046 16026 23106 16049
rect 20993 15794 21053 15819
rect 21111 15794 21171 15819
rect 21229 15794 21289 15819
rect 21642 15800 21702 15826
rect 21760 15800 21820 15826
rect 19542 15753 20121 15788
rect 20710 15753 21289 15794
rect 21878 15794 21938 15826
rect 23329 16020 23389 16046
rect 23447 16020 23507 16046
rect 23565 16020 23625 16046
rect 22161 15794 22221 15819
rect 22279 15794 22339 15819
rect 22397 15794 22457 15819
rect 22810 15800 22870 15826
rect 22928 15800 22988 15826
rect 21878 15753 22457 15794
rect 23046 15794 23106 15826
rect 23329 15794 23389 15820
rect 23447 15794 23507 15820
rect 23565 15794 23625 15820
rect 23046 15753 23625 15794
rect 13615 15704 13631 15738
rect 13665 15704 13681 15738
rect 13615 15688 13681 15704
rect 3455 14869 3751 14908
rect 3455 14854 3515 14869
rect 3573 14854 3633 14869
rect 3691 14854 3751 14869
rect 3922 14869 4218 14908
rect 3922 14854 3982 14869
rect 4040 14854 4100 14869
rect 4158 14854 4218 14869
rect 4276 14869 4572 14908
rect 4276 14854 4336 14869
rect 4394 14854 4454 14869
rect 4512 14854 4572 14869
rect 4749 14869 5045 14908
rect 4749 14854 4809 14869
rect 4867 14854 4927 14869
rect 4985 14854 5045 14869
rect 6599 14869 6895 14908
rect 6599 14854 6659 14869
rect 6717 14854 6777 14869
rect 6835 14854 6895 14869
rect 7066 14869 7362 14908
rect 7066 14854 7126 14869
rect 7184 14854 7244 14869
rect 7302 14854 7362 14869
rect 7420 14869 7716 14908
rect 7420 14854 7480 14869
rect 7538 14854 7598 14869
rect 7656 14854 7716 14869
rect 7893 14869 8189 14908
rect 7893 14854 7953 14869
rect 8011 14854 8071 14869
rect 8129 14854 8189 14869
rect 9731 14873 10027 14912
rect 9731 14858 9791 14873
rect 9849 14858 9909 14873
rect 9967 14858 10027 14873
rect 10198 14873 10494 14912
rect 10198 14858 10258 14873
rect 10316 14858 10376 14873
rect 10434 14858 10494 14873
rect 10552 14873 10848 14912
rect 10552 14858 10612 14873
rect 10670 14858 10730 14873
rect 10788 14858 10848 14873
rect 11025 14873 11321 14912
rect 11025 14858 11085 14873
rect 11143 14858 11203 14873
rect 11261 14858 11321 14873
rect 12875 14873 13171 14912
rect 12875 14858 12935 14873
rect 12993 14858 13053 14873
rect 13111 14858 13171 14873
rect 13342 14873 13638 14912
rect 13342 14858 13402 14873
rect 13460 14858 13520 14873
rect 13578 14858 13638 14873
rect 13696 14873 13992 14912
rect 13696 14858 13756 14873
rect 13814 14858 13874 14873
rect 13932 14858 13992 14873
rect 14169 14873 14465 14912
rect 14169 14858 14229 14873
rect 14287 14858 14347 14873
rect 14405 14858 14465 14873
rect 16077 14869 16373 14908
rect 3014 14670 3310 14709
rect 3014 14654 3074 14670
rect 3132 14654 3192 14670
rect 3250 14654 3310 14670
rect 5222 14670 5518 14709
rect 5222 14654 5282 14670
rect 5340 14654 5400 14670
rect 5458 14654 5518 14670
rect 6158 14670 6454 14709
rect 6158 14654 6218 14670
rect 6276 14654 6336 14670
rect 6394 14654 6454 14670
rect 8366 14670 8662 14709
rect 8366 14654 8426 14670
rect 8484 14654 8544 14670
rect 8602 14654 8662 14670
rect 9290 14674 9586 14713
rect 9290 14658 9350 14674
rect 9408 14658 9468 14674
rect 9526 14658 9586 14674
rect 11498 14674 11794 14713
rect 11498 14658 11558 14674
rect 11616 14658 11676 14674
rect 11734 14658 11794 14674
rect 12434 14674 12730 14713
rect 12434 14658 12494 14674
rect 12552 14658 12612 14674
rect 12670 14658 12730 14674
rect 16077 14854 16137 14869
rect 16195 14854 16255 14869
rect 16313 14854 16373 14869
rect 16544 14869 16840 14908
rect 16544 14854 16604 14869
rect 16662 14854 16722 14869
rect 16780 14854 16840 14869
rect 16898 14869 17194 14908
rect 16898 14854 16958 14869
rect 17016 14854 17076 14869
rect 17134 14854 17194 14869
rect 17371 14869 17667 14908
rect 17371 14854 17431 14869
rect 17489 14854 17549 14869
rect 17607 14854 17667 14869
rect 19221 14869 19517 14908
rect 19221 14854 19281 14869
rect 19339 14854 19399 14869
rect 19457 14854 19517 14869
rect 19688 14869 19984 14908
rect 19688 14854 19748 14869
rect 19806 14854 19866 14869
rect 19924 14854 19984 14869
rect 20042 14869 20338 14908
rect 20042 14854 20102 14869
rect 20160 14854 20220 14869
rect 20278 14854 20338 14869
rect 20515 14869 20811 14908
rect 20515 14854 20575 14869
rect 20633 14854 20693 14869
rect 20751 14854 20811 14869
rect 22353 14873 22649 14912
rect 22353 14858 22413 14873
rect 22471 14858 22531 14873
rect 22589 14858 22649 14873
rect 22820 14873 23116 14912
rect 22820 14858 22880 14873
rect 22938 14858 22998 14873
rect 23056 14858 23116 14873
rect 23174 14873 23470 14912
rect 23174 14858 23234 14873
rect 23292 14858 23352 14873
rect 23410 14858 23470 14873
rect 23647 14873 23943 14912
rect 23647 14858 23707 14873
rect 23765 14858 23825 14873
rect 23883 14858 23943 14873
rect 25497 14873 25793 14912
rect 25497 14858 25557 14873
rect 25615 14858 25675 14873
rect 25733 14858 25793 14873
rect 25964 14873 26260 14912
rect 25964 14858 26024 14873
rect 26082 14858 26142 14873
rect 26200 14858 26260 14873
rect 26318 14873 26614 14912
rect 26318 14858 26378 14873
rect 26436 14858 26496 14873
rect 26554 14858 26614 14873
rect 26791 14873 27087 14912
rect 26791 14858 26851 14873
rect 26909 14858 26969 14873
rect 27027 14858 27087 14873
rect 14642 14674 14938 14713
rect 14642 14658 14702 14674
rect 14760 14658 14820 14674
rect 14878 14658 14938 14674
rect 15636 14670 15932 14709
rect 15636 14654 15696 14670
rect 15754 14654 15814 14670
rect 15872 14654 15932 14670
rect 3014 14168 3074 14454
rect 3132 14428 3192 14454
rect 3250 14428 3310 14454
rect 3455 14428 3515 14454
rect 3014 14151 3150 14168
rect 3014 14096 3073 14151
rect 3131 14096 3150 14151
rect 3014 14081 3150 14096
rect 3014 13769 3074 14081
rect 3573 14036 3633 14454
rect 3691 14428 3751 14454
rect 3922 14428 3982 14454
rect 4040 14428 4100 14454
rect 4158 14428 4218 14454
rect 4276 14428 4336 14454
rect 4041 14268 4100 14428
rect 4041 14267 4104 14268
rect 4038 14251 4104 14267
rect 4038 14217 4054 14251
rect 4088 14217 4104 14251
rect 4038 14201 4104 14217
rect 4141 14152 4236 14167
rect 4141 14097 4160 14152
rect 4218 14129 4236 14152
rect 4394 14129 4454 14454
rect 4512 14428 4572 14454
rect 4749 14428 4809 14454
rect 4218 14097 4454 14129
rect 4141 14080 4454 14097
rect 3573 13979 4100 14036
rect 4040 13880 4100 13979
rect 4029 13867 4110 13880
rect 4029 13812 4042 13867
rect 4100 13812 4110 13867
rect 4029 13801 4110 13812
rect 3014 13724 3908 13769
rect 3848 13521 3908 13724
rect 4040 13521 4100 13801
rect 4158 13521 4218 14080
rect 4867 14038 4927 14454
rect 4985 14428 5045 14454
rect 5222 14428 5282 14454
rect 5340 14428 5400 14454
rect 5348 14305 5414 14308
rect 5458 14305 5518 14454
rect 5348 14292 5518 14305
rect 5348 14258 5364 14292
rect 5398 14258 5518 14292
rect 5348 14245 5518 14258
rect 5348 14242 5414 14245
rect 4389 14021 4927 14038
rect 4389 13987 4408 14021
rect 4442 13987 4927 14021
rect 4389 13981 4927 13987
rect 4389 13971 4458 13981
rect 4389 13969 4454 13971
rect 4273 13631 4339 13647
rect 4273 13597 4289 13631
rect 4323 13597 4339 13631
rect 4273 13581 4339 13597
rect 4276 13521 4336 13581
rect 4394 13521 4454 13969
rect 5458 13769 5518 14245
rect 4590 13724 5518 13769
rect 6158 14168 6218 14454
rect 6276 14428 6336 14454
rect 6394 14428 6454 14454
rect 6599 14428 6659 14454
rect 6158 14151 6294 14168
rect 6158 14096 6217 14151
rect 6275 14096 6294 14151
rect 6158 14081 6294 14096
rect 6158 13769 6218 14081
rect 6717 14036 6777 14454
rect 6835 14428 6895 14454
rect 7066 14428 7126 14454
rect 7184 14428 7244 14454
rect 7302 14428 7362 14454
rect 7420 14428 7480 14454
rect 7185 14268 7244 14428
rect 7185 14267 7248 14268
rect 7182 14251 7248 14267
rect 7182 14217 7198 14251
rect 7232 14217 7248 14251
rect 7182 14201 7248 14217
rect 7285 14152 7380 14167
rect 7285 14097 7304 14152
rect 7362 14129 7380 14152
rect 7538 14129 7598 14454
rect 7656 14428 7716 14454
rect 7893 14428 7953 14454
rect 7362 14097 7598 14129
rect 7285 14080 7598 14097
rect 6717 13979 7244 14036
rect 7184 13880 7244 13979
rect 7173 13867 7254 13880
rect 7173 13812 7186 13867
rect 7244 13812 7254 13867
rect 7173 13801 7254 13812
rect 6158 13724 7052 13769
rect 4590 13521 4650 13724
rect 6992 13521 7052 13724
rect 7184 13521 7244 13801
rect 7302 13521 7362 14080
rect 8011 14038 8071 14454
rect 8129 14428 8189 14454
rect 8366 14428 8426 14454
rect 8484 14428 8544 14454
rect 8492 14305 8558 14308
rect 8602 14305 8662 14454
rect 8492 14292 8662 14305
rect 8492 14258 8508 14292
rect 8542 14258 8662 14292
rect 8492 14245 8662 14258
rect 8492 14242 8558 14245
rect 7533 14021 8071 14038
rect 7533 13987 7552 14021
rect 7586 13987 8071 14021
rect 7533 13981 8071 13987
rect 7533 13971 7602 13981
rect 7533 13969 7598 13971
rect 7417 13631 7483 13647
rect 7417 13597 7433 13631
rect 7467 13597 7483 13631
rect 7417 13581 7483 13597
rect 7420 13521 7480 13581
rect 7538 13521 7598 13969
rect 8602 13769 8662 14245
rect 7734 13724 8662 13769
rect 9290 14172 9350 14458
rect 9408 14432 9468 14458
rect 9526 14432 9586 14458
rect 9731 14432 9791 14458
rect 9290 14155 9426 14172
rect 9290 14100 9349 14155
rect 9407 14100 9426 14155
rect 9290 14085 9426 14100
rect 9290 13773 9350 14085
rect 9849 14040 9909 14458
rect 9967 14432 10027 14458
rect 10198 14432 10258 14458
rect 10316 14432 10376 14458
rect 10434 14432 10494 14458
rect 10552 14432 10612 14458
rect 10317 14272 10376 14432
rect 10317 14271 10380 14272
rect 10314 14255 10380 14271
rect 10314 14221 10330 14255
rect 10364 14221 10380 14255
rect 10314 14205 10380 14221
rect 10417 14156 10512 14171
rect 10417 14101 10436 14156
rect 10494 14133 10512 14156
rect 10670 14133 10730 14458
rect 10788 14432 10848 14458
rect 11025 14432 11085 14458
rect 10494 14101 10730 14133
rect 10417 14084 10730 14101
rect 9849 13983 10376 14040
rect 10316 13884 10376 13983
rect 10305 13871 10386 13884
rect 10305 13816 10318 13871
rect 10376 13816 10386 13871
rect 10305 13805 10386 13816
rect 9290 13728 10184 13773
rect 7734 13521 7794 13724
rect 10124 13525 10184 13728
rect 10316 13525 10376 13805
rect 10434 13525 10494 14084
rect 11143 14042 11203 14458
rect 11261 14432 11321 14458
rect 11498 14432 11558 14458
rect 11616 14432 11676 14458
rect 11624 14309 11690 14312
rect 11734 14309 11794 14458
rect 11624 14296 11794 14309
rect 11624 14262 11640 14296
rect 11674 14262 11794 14296
rect 11624 14249 11794 14262
rect 11624 14246 11690 14249
rect 10665 14025 11203 14042
rect 10665 13991 10684 14025
rect 10718 13991 11203 14025
rect 10665 13985 11203 13991
rect 10665 13975 10734 13985
rect 10665 13973 10730 13975
rect 10549 13635 10615 13651
rect 10549 13601 10565 13635
rect 10599 13601 10615 13635
rect 10549 13585 10615 13601
rect 10552 13525 10612 13585
rect 10670 13525 10730 13973
rect 11734 13773 11794 14249
rect 10866 13728 11794 13773
rect 12434 14172 12494 14458
rect 12552 14432 12612 14458
rect 12670 14432 12730 14458
rect 12875 14432 12935 14458
rect 12434 14155 12570 14172
rect 12434 14100 12493 14155
rect 12551 14100 12570 14155
rect 12434 14085 12570 14100
rect 12434 13773 12494 14085
rect 12993 14040 13053 14458
rect 13111 14432 13171 14458
rect 13342 14432 13402 14458
rect 13460 14432 13520 14458
rect 13578 14432 13638 14458
rect 13696 14432 13756 14458
rect 13461 14272 13520 14432
rect 13461 14271 13524 14272
rect 13458 14255 13524 14271
rect 13458 14221 13474 14255
rect 13508 14221 13524 14255
rect 13458 14205 13524 14221
rect 13561 14156 13656 14171
rect 13561 14101 13580 14156
rect 13638 14133 13656 14156
rect 13814 14133 13874 14458
rect 13932 14432 13992 14458
rect 14169 14432 14229 14458
rect 13638 14101 13874 14133
rect 13561 14084 13874 14101
rect 12993 13983 13520 14040
rect 13460 13884 13520 13983
rect 13449 13871 13530 13884
rect 13449 13816 13462 13871
rect 13520 13816 13530 13871
rect 13449 13805 13530 13816
rect 12434 13728 13328 13773
rect 10866 13525 10926 13728
rect 13268 13525 13328 13728
rect 13460 13525 13520 13805
rect 13578 13525 13638 14084
rect 14287 14042 14347 14458
rect 14405 14432 14465 14458
rect 14642 14432 14702 14458
rect 14760 14432 14820 14458
rect 14768 14309 14834 14312
rect 14878 14309 14938 14458
rect 17844 14670 18140 14709
rect 17844 14654 17904 14670
rect 17962 14654 18022 14670
rect 18080 14654 18140 14670
rect 18780 14670 19076 14709
rect 18780 14654 18840 14670
rect 18898 14654 18958 14670
rect 19016 14654 19076 14670
rect 20988 14670 21284 14709
rect 20988 14654 21048 14670
rect 21106 14654 21166 14670
rect 21224 14654 21284 14670
rect 21912 14674 22208 14713
rect 21912 14658 21972 14674
rect 22030 14658 22090 14674
rect 22148 14658 22208 14674
rect 24120 14674 24416 14713
rect 24120 14658 24180 14674
rect 24238 14658 24298 14674
rect 24356 14658 24416 14674
rect 25056 14674 25352 14713
rect 25056 14658 25116 14674
rect 25174 14658 25234 14674
rect 25292 14658 25352 14674
rect 27264 14674 27560 14713
rect 27264 14658 27324 14674
rect 27382 14658 27442 14674
rect 27500 14658 27560 14674
rect 14768 14296 14938 14309
rect 14768 14262 14784 14296
rect 14818 14262 14938 14296
rect 14768 14249 14938 14262
rect 14768 14246 14834 14249
rect 13809 14025 14347 14042
rect 13809 13991 13828 14025
rect 13862 13991 14347 14025
rect 13809 13985 14347 13991
rect 13809 13975 13878 13985
rect 13809 13973 13874 13975
rect 13693 13635 13759 13651
rect 13693 13601 13709 13635
rect 13743 13601 13759 13635
rect 13693 13585 13759 13601
rect 13696 13525 13756 13585
rect 13814 13525 13874 13973
rect 14878 13773 14938 14249
rect 14010 13728 14938 13773
rect 15636 14168 15696 14454
rect 15754 14428 15814 14454
rect 15872 14428 15932 14454
rect 16077 14428 16137 14454
rect 15636 14151 15772 14168
rect 15636 14096 15695 14151
rect 15753 14096 15772 14151
rect 15636 14081 15772 14096
rect 15636 13769 15696 14081
rect 16195 14036 16255 14454
rect 16313 14428 16373 14454
rect 16544 14428 16604 14454
rect 16662 14428 16722 14454
rect 16780 14428 16840 14454
rect 16898 14428 16958 14454
rect 16663 14268 16722 14428
rect 16663 14267 16726 14268
rect 16660 14251 16726 14267
rect 16660 14217 16676 14251
rect 16710 14217 16726 14251
rect 16660 14201 16726 14217
rect 16763 14152 16858 14167
rect 16763 14097 16782 14152
rect 16840 14129 16858 14152
rect 17016 14129 17076 14454
rect 17134 14428 17194 14454
rect 17371 14428 17431 14454
rect 16840 14097 17076 14129
rect 16763 14080 17076 14097
rect 16195 13979 16722 14036
rect 16662 13880 16722 13979
rect 16651 13867 16732 13880
rect 16651 13812 16664 13867
rect 16722 13812 16732 13867
rect 16651 13801 16732 13812
rect 14010 13525 14070 13728
rect 15636 13724 16530 13769
rect 3848 13295 3908 13321
rect 4040 13095 4100 13121
rect 4158 13095 4218 13121
rect 4276 13095 4336 13121
rect 4394 13095 4454 13121
rect 4215 13040 4281 13048
rect 4590 13040 4650 13321
rect 6992 13295 7052 13321
rect 7184 13095 7244 13121
rect 7302 13095 7362 13121
rect 7420 13095 7480 13121
rect 7538 13095 7598 13121
rect 4215 13032 4650 13040
rect 4215 12998 4231 13032
rect 4265 12998 4650 13032
rect 4215 12989 4650 12998
rect 7359 13040 7425 13048
rect 7734 13040 7794 13321
rect 10124 13299 10184 13325
rect 10316 13099 10376 13125
rect 10434 13099 10494 13125
rect 10552 13099 10612 13125
rect 10670 13099 10730 13125
rect 7359 13032 7794 13040
rect 7359 12998 7375 13032
rect 7409 12998 7794 13032
rect 7359 12989 7794 12998
rect 10491 13044 10557 13052
rect 10866 13044 10926 13325
rect 13268 13299 13328 13325
rect 16470 13521 16530 13724
rect 16662 13521 16722 13801
rect 16780 13521 16840 14080
rect 17489 14038 17549 14454
rect 17607 14428 17667 14454
rect 17844 14428 17904 14454
rect 17962 14428 18022 14454
rect 17970 14305 18036 14308
rect 18080 14305 18140 14454
rect 17970 14292 18140 14305
rect 17970 14258 17986 14292
rect 18020 14258 18140 14292
rect 17970 14245 18140 14258
rect 17970 14242 18036 14245
rect 17011 14021 17549 14038
rect 17011 13987 17030 14021
rect 17064 13987 17549 14021
rect 17011 13981 17549 13987
rect 17011 13971 17080 13981
rect 17011 13969 17076 13971
rect 16895 13631 16961 13647
rect 16895 13597 16911 13631
rect 16945 13597 16961 13631
rect 16895 13581 16961 13597
rect 16898 13521 16958 13581
rect 17016 13521 17076 13969
rect 18080 13769 18140 14245
rect 17212 13724 18140 13769
rect 18780 14168 18840 14454
rect 18898 14428 18958 14454
rect 19016 14428 19076 14454
rect 19221 14428 19281 14454
rect 18780 14151 18916 14168
rect 18780 14096 18839 14151
rect 18897 14096 18916 14151
rect 18780 14081 18916 14096
rect 18780 13769 18840 14081
rect 19339 14036 19399 14454
rect 19457 14428 19517 14454
rect 19688 14428 19748 14454
rect 19806 14428 19866 14454
rect 19924 14428 19984 14454
rect 20042 14428 20102 14454
rect 19807 14268 19866 14428
rect 19807 14267 19870 14268
rect 19804 14251 19870 14267
rect 19804 14217 19820 14251
rect 19854 14217 19870 14251
rect 19804 14201 19870 14217
rect 19907 14152 20002 14167
rect 19907 14097 19926 14152
rect 19984 14129 20002 14152
rect 20160 14129 20220 14454
rect 20278 14428 20338 14454
rect 20515 14428 20575 14454
rect 19984 14097 20220 14129
rect 19907 14080 20220 14097
rect 19339 13979 19866 14036
rect 19806 13880 19866 13979
rect 19795 13867 19876 13880
rect 19795 13812 19808 13867
rect 19866 13812 19876 13867
rect 19795 13801 19876 13812
rect 18780 13724 19674 13769
rect 17212 13521 17272 13724
rect 19614 13521 19674 13724
rect 19806 13521 19866 13801
rect 19924 13521 19984 14080
rect 20633 14038 20693 14454
rect 20751 14428 20811 14454
rect 20988 14428 21048 14454
rect 21106 14428 21166 14454
rect 21114 14305 21180 14308
rect 21224 14305 21284 14454
rect 21114 14292 21284 14305
rect 21114 14258 21130 14292
rect 21164 14258 21284 14292
rect 21114 14245 21284 14258
rect 21114 14242 21180 14245
rect 20155 14021 20693 14038
rect 20155 13987 20174 14021
rect 20208 13987 20693 14021
rect 20155 13981 20693 13987
rect 20155 13971 20224 13981
rect 20155 13969 20220 13971
rect 20039 13631 20105 13647
rect 20039 13597 20055 13631
rect 20089 13597 20105 13631
rect 20039 13581 20105 13597
rect 20042 13521 20102 13581
rect 20160 13521 20220 13969
rect 21224 13769 21284 14245
rect 20356 13724 21284 13769
rect 21912 14172 21972 14458
rect 22030 14432 22090 14458
rect 22148 14432 22208 14458
rect 22353 14432 22413 14458
rect 21912 14155 22048 14172
rect 21912 14100 21971 14155
rect 22029 14100 22048 14155
rect 21912 14085 22048 14100
rect 21912 13773 21972 14085
rect 22471 14040 22531 14458
rect 22589 14432 22649 14458
rect 22820 14432 22880 14458
rect 22938 14432 22998 14458
rect 23056 14432 23116 14458
rect 23174 14432 23234 14458
rect 22939 14272 22998 14432
rect 22939 14271 23002 14272
rect 22936 14255 23002 14271
rect 22936 14221 22952 14255
rect 22986 14221 23002 14255
rect 22936 14205 23002 14221
rect 23039 14156 23134 14171
rect 23039 14101 23058 14156
rect 23116 14133 23134 14156
rect 23292 14133 23352 14458
rect 23410 14432 23470 14458
rect 23647 14432 23707 14458
rect 23116 14101 23352 14133
rect 23039 14084 23352 14101
rect 22471 13983 22998 14040
rect 22938 13884 22998 13983
rect 22927 13871 23008 13884
rect 22927 13816 22940 13871
rect 22998 13816 23008 13871
rect 22927 13805 23008 13816
rect 21912 13728 22806 13773
rect 20356 13521 20416 13724
rect 22746 13525 22806 13728
rect 22938 13525 22998 13805
rect 23056 13525 23116 14084
rect 23765 14042 23825 14458
rect 23883 14432 23943 14458
rect 24120 14432 24180 14458
rect 24238 14432 24298 14458
rect 24246 14309 24312 14312
rect 24356 14309 24416 14458
rect 24246 14296 24416 14309
rect 24246 14262 24262 14296
rect 24296 14262 24416 14296
rect 24246 14249 24416 14262
rect 24246 14246 24312 14249
rect 23287 14025 23825 14042
rect 23287 13991 23306 14025
rect 23340 13991 23825 14025
rect 23287 13985 23825 13991
rect 23287 13975 23356 13985
rect 23287 13973 23352 13975
rect 23171 13635 23237 13651
rect 23171 13601 23187 13635
rect 23221 13601 23237 13635
rect 23171 13585 23237 13601
rect 23174 13525 23234 13585
rect 23292 13525 23352 13973
rect 24356 13773 24416 14249
rect 23488 13728 24416 13773
rect 25056 14172 25116 14458
rect 25174 14432 25234 14458
rect 25292 14432 25352 14458
rect 25497 14432 25557 14458
rect 25056 14155 25192 14172
rect 25056 14100 25115 14155
rect 25173 14100 25192 14155
rect 25056 14085 25192 14100
rect 25056 13773 25116 14085
rect 25615 14040 25675 14458
rect 25733 14432 25793 14458
rect 25964 14432 26024 14458
rect 26082 14432 26142 14458
rect 26200 14432 26260 14458
rect 26318 14432 26378 14458
rect 26083 14272 26142 14432
rect 26083 14271 26146 14272
rect 26080 14255 26146 14271
rect 26080 14221 26096 14255
rect 26130 14221 26146 14255
rect 26080 14205 26146 14221
rect 26183 14156 26278 14171
rect 26183 14101 26202 14156
rect 26260 14133 26278 14156
rect 26436 14133 26496 14458
rect 26554 14432 26614 14458
rect 26791 14432 26851 14458
rect 26260 14101 26496 14133
rect 26183 14084 26496 14101
rect 25615 13983 26142 14040
rect 26082 13884 26142 13983
rect 26071 13871 26152 13884
rect 26071 13816 26084 13871
rect 26142 13816 26152 13871
rect 26071 13805 26152 13816
rect 25056 13728 25950 13773
rect 23488 13525 23548 13728
rect 25890 13525 25950 13728
rect 26082 13525 26142 13805
rect 26200 13525 26260 14084
rect 26909 14042 26969 14458
rect 27027 14432 27087 14458
rect 27264 14432 27324 14458
rect 27382 14432 27442 14458
rect 27390 14309 27456 14312
rect 27500 14309 27560 14458
rect 27390 14296 27560 14309
rect 27390 14262 27406 14296
rect 27440 14262 27560 14296
rect 27390 14249 27560 14262
rect 27390 14246 27456 14249
rect 26431 14025 26969 14042
rect 26431 13991 26450 14025
rect 26484 13991 26969 14025
rect 26431 13985 26969 13991
rect 26431 13975 26500 13985
rect 26431 13973 26496 13975
rect 26315 13635 26381 13651
rect 26315 13601 26331 13635
rect 26365 13601 26381 13635
rect 26315 13585 26381 13601
rect 26318 13525 26378 13585
rect 26436 13525 26496 13973
rect 27500 13773 27560 14249
rect 26632 13728 27560 13773
rect 26632 13525 26692 13728
rect 13460 13099 13520 13125
rect 13578 13099 13638 13125
rect 13696 13099 13756 13125
rect 13814 13099 13874 13125
rect 10491 13036 10926 13044
rect 10491 13002 10507 13036
rect 10541 13002 10926 13036
rect 10491 12993 10926 13002
rect 13635 13044 13701 13052
rect 14010 13044 14070 13325
rect 16470 13295 16530 13321
rect 16662 13095 16722 13121
rect 16780 13095 16840 13121
rect 16898 13095 16958 13121
rect 17016 13095 17076 13121
rect 13635 13036 14070 13044
rect 13635 13002 13651 13036
rect 13685 13002 14070 13036
rect 13635 12993 14070 13002
rect 16837 13040 16903 13048
rect 17212 13040 17272 13321
rect 19614 13295 19674 13321
rect 19806 13095 19866 13121
rect 19924 13095 19984 13121
rect 20042 13095 20102 13121
rect 20160 13095 20220 13121
rect 16837 13032 17272 13040
rect 16837 12998 16853 13032
rect 16887 12998 17272 13032
rect 4215 12982 4281 12989
rect 7359 12982 7425 12989
rect 10491 12986 10557 12993
rect 13635 12986 13701 12993
rect 16837 12989 17272 12998
rect 19981 13040 20047 13048
rect 20356 13040 20416 13321
rect 22746 13299 22806 13325
rect 22938 13099 22998 13125
rect 23056 13099 23116 13125
rect 23174 13099 23234 13125
rect 23292 13099 23352 13125
rect 19981 13032 20416 13040
rect 19981 12998 19997 13032
rect 20031 12998 20416 13032
rect 19981 12989 20416 12998
rect 23113 13044 23179 13052
rect 23488 13044 23548 13325
rect 25890 13299 25950 13325
rect 26082 13099 26142 13125
rect 26200 13099 26260 13125
rect 26318 13099 26378 13125
rect 26436 13099 26496 13125
rect 23113 13036 23548 13044
rect 23113 13002 23129 13036
rect 23163 13002 23548 13036
rect 23113 12993 23548 13002
rect 26257 13044 26323 13052
rect 26632 13044 26692 13325
rect 26257 13036 26692 13044
rect 26257 13002 26273 13036
rect 26307 13002 26692 13036
rect 26257 12993 26692 13002
rect 16837 12982 16903 12989
rect 19981 12982 20047 12989
rect 23113 12986 23179 12993
rect 26257 12986 26323 12993
rect 3455 12135 3751 12174
rect 3455 12120 3515 12135
rect 3573 12120 3633 12135
rect 3691 12120 3751 12135
rect 3922 12135 4218 12174
rect 3922 12120 3982 12135
rect 4040 12120 4100 12135
rect 4158 12120 4218 12135
rect 4276 12135 4572 12174
rect 4276 12120 4336 12135
rect 4394 12120 4454 12135
rect 4512 12120 4572 12135
rect 4749 12135 5045 12174
rect 4749 12120 4809 12135
rect 4867 12120 4927 12135
rect 4985 12120 5045 12135
rect 6599 12135 6895 12174
rect 6599 12120 6659 12135
rect 6717 12120 6777 12135
rect 6835 12120 6895 12135
rect 7066 12135 7362 12174
rect 7066 12120 7126 12135
rect 7184 12120 7244 12135
rect 7302 12120 7362 12135
rect 7420 12135 7716 12174
rect 7420 12120 7480 12135
rect 7538 12120 7598 12135
rect 7656 12120 7716 12135
rect 7893 12135 8189 12174
rect 7893 12120 7953 12135
rect 8011 12120 8071 12135
rect 8129 12120 8189 12135
rect 9731 12139 10027 12178
rect 9731 12124 9791 12139
rect 9849 12124 9909 12139
rect 9967 12124 10027 12139
rect 10198 12139 10494 12178
rect 10198 12124 10258 12139
rect 10316 12124 10376 12139
rect 10434 12124 10494 12139
rect 10552 12139 10848 12178
rect 10552 12124 10612 12139
rect 10670 12124 10730 12139
rect 10788 12124 10848 12139
rect 11025 12139 11321 12178
rect 11025 12124 11085 12139
rect 11143 12124 11203 12139
rect 11261 12124 11321 12139
rect 12875 12139 13171 12178
rect 12875 12124 12935 12139
rect 12993 12124 13053 12139
rect 13111 12124 13171 12139
rect 13342 12139 13638 12178
rect 13342 12124 13402 12139
rect 13460 12124 13520 12139
rect 13578 12124 13638 12139
rect 13696 12139 13992 12178
rect 13696 12124 13756 12139
rect 13814 12124 13874 12139
rect 13932 12124 13992 12139
rect 14169 12139 14465 12178
rect 14169 12124 14229 12139
rect 14287 12124 14347 12139
rect 14405 12124 14465 12139
rect 16077 12135 16373 12174
rect 3014 11936 3310 11975
rect 3014 11920 3074 11936
rect 3132 11920 3192 11936
rect 3250 11920 3310 11936
rect 5222 11936 5518 11975
rect 5222 11920 5282 11936
rect 5340 11920 5400 11936
rect 5458 11920 5518 11936
rect 6158 11936 6454 11975
rect 6158 11920 6218 11936
rect 6276 11920 6336 11936
rect 6394 11920 6454 11936
rect 8366 11936 8662 11975
rect 8366 11920 8426 11936
rect 8484 11920 8544 11936
rect 8602 11920 8662 11936
rect 9290 11940 9586 11979
rect 9290 11924 9350 11940
rect 9408 11924 9468 11940
rect 9526 11924 9586 11940
rect 11498 11940 11794 11979
rect 11498 11924 11558 11940
rect 11616 11924 11676 11940
rect 11734 11924 11794 11940
rect 12434 11940 12730 11979
rect 12434 11924 12494 11940
rect 12552 11924 12612 11940
rect 12670 11924 12730 11940
rect 16077 12120 16137 12135
rect 16195 12120 16255 12135
rect 16313 12120 16373 12135
rect 16544 12135 16840 12174
rect 16544 12120 16604 12135
rect 16662 12120 16722 12135
rect 16780 12120 16840 12135
rect 16898 12135 17194 12174
rect 16898 12120 16958 12135
rect 17016 12120 17076 12135
rect 17134 12120 17194 12135
rect 17371 12135 17667 12174
rect 17371 12120 17431 12135
rect 17489 12120 17549 12135
rect 17607 12120 17667 12135
rect 19221 12135 19517 12174
rect 19221 12120 19281 12135
rect 19339 12120 19399 12135
rect 19457 12120 19517 12135
rect 19688 12135 19984 12174
rect 19688 12120 19748 12135
rect 19806 12120 19866 12135
rect 19924 12120 19984 12135
rect 20042 12135 20338 12174
rect 20042 12120 20102 12135
rect 20160 12120 20220 12135
rect 20278 12120 20338 12135
rect 20515 12135 20811 12174
rect 20515 12120 20575 12135
rect 20633 12120 20693 12135
rect 20751 12120 20811 12135
rect 22353 12139 22649 12178
rect 22353 12124 22413 12139
rect 22471 12124 22531 12139
rect 22589 12124 22649 12139
rect 22820 12139 23116 12178
rect 22820 12124 22880 12139
rect 22938 12124 22998 12139
rect 23056 12124 23116 12139
rect 23174 12139 23470 12178
rect 23174 12124 23234 12139
rect 23292 12124 23352 12139
rect 23410 12124 23470 12139
rect 23647 12139 23943 12178
rect 23647 12124 23707 12139
rect 23765 12124 23825 12139
rect 23883 12124 23943 12139
rect 25497 12139 25793 12178
rect 25497 12124 25557 12139
rect 25615 12124 25675 12139
rect 25733 12124 25793 12139
rect 25964 12139 26260 12178
rect 25964 12124 26024 12139
rect 26082 12124 26142 12139
rect 26200 12124 26260 12139
rect 26318 12139 26614 12178
rect 26318 12124 26378 12139
rect 26436 12124 26496 12139
rect 26554 12124 26614 12139
rect 26791 12139 27087 12178
rect 26791 12124 26851 12139
rect 26909 12124 26969 12139
rect 27027 12124 27087 12139
rect 14642 11940 14938 11979
rect 14642 11924 14702 11940
rect 14760 11924 14820 11940
rect 14878 11924 14938 11940
rect 15636 11936 15932 11975
rect 15636 11920 15696 11936
rect 15754 11920 15814 11936
rect 15872 11920 15932 11936
rect 3014 11434 3074 11720
rect 3132 11694 3192 11720
rect 3250 11694 3310 11720
rect 3455 11694 3515 11720
rect 3014 11417 3150 11434
rect 3014 11362 3073 11417
rect 3131 11362 3150 11417
rect 3014 11347 3150 11362
rect 3014 11035 3074 11347
rect 3573 11302 3633 11720
rect 3691 11694 3751 11720
rect 3922 11694 3982 11720
rect 4040 11694 4100 11720
rect 4158 11694 4218 11720
rect 4276 11694 4336 11720
rect 4041 11534 4100 11694
rect 4041 11533 4104 11534
rect 4038 11517 4104 11533
rect 4038 11483 4054 11517
rect 4088 11483 4104 11517
rect 4038 11467 4104 11483
rect 4141 11418 4236 11433
rect 4141 11363 4160 11418
rect 4218 11395 4236 11418
rect 4394 11395 4454 11720
rect 4512 11694 4572 11720
rect 4749 11694 4809 11720
rect 4218 11363 4454 11395
rect 4141 11346 4454 11363
rect 3573 11245 4100 11302
rect 4040 11146 4100 11245
rect 4029 11133 4110 11146
rect 4029 11078 4042 11133
rect 4100 11078 4110 11133
rect 4029 11067 4110 11078
rect 3014 10990 3908 11035
rect 3848 10787 3908 10990
rect 4040 10787 4100 11067
rect 4158 10787 4218 11346
rect 4867 11304 4927 11720
rect 4985 11694 5045 11720
rect 5222 11694 5282 11720
rect 5340 11694 5400 11720
rect 5348 11571 5414 11574
rect 5458 11571 5518 11720
rect 5348 11558 5518 11571
rect 5348 11524 5364 11558
rect 5398 11524 5518 11558
rect 5348 11511 5518 11524
rect 5348 11508 5414 11511
rect 4389 11287 4927 11304
rect 4389 11253 4408 11287
rect 4442 11253 4927 11287
rect 4389 11247 4927 11253
rect 4389 11237 4458 11247
rect 4389 11235 4454 11237
rect 4273 10897 4339 10913
rect 4273 10863 4289 10897
rect 4323 10863 4339 10897
rect 4273 10847 4339 10863
rect 4276 10787 4336 10847
rect 4394 10787 4454 11235
rect 5458 11035 5518 11511
rect 4590 10990 5518 11035
rect 6158 11434 6218 11720
rect 6276 11694 6336 11720
rect 6394 11694 6454 11720
rect 6599 11694 6659 11720
rect 6158 11417 6294 11434
rect 6158 11362 6217 11417
rect 6275 11362 6294 11417
rect 6158 11347 6294 11362
rect 6158 11035 6218 11347
rect 6717 11302 6777 11720
rect 6835 11694 6895 11720
rect 7066 11694 7126 11720
rect 7184 11694 7244 11720
rect 7302 11694 7362 11720
rect 7420 11694 7480 11720
rect 7185 11534 7244 11694
rect 7185 11533 7248 11534
rect 7182 11517 7248 11533
rect 7182 11483 7198 11517
rect 7232 11483 7248 11517
rect 7182 11467 7248 11483
rect 7285 11418 7380 11433
rect 7285 11363 7304 11418
rect 7362 11395 7380 11418
rect 7538 11395 7598 11720
rect 7656 11694 7716 11720
rect 7893 11694 7953 11720
rect 7362 11363 7598 11395
rect 7285 11346 7598 11363
rect 6717 11245 7244 11302
rect 7184 11146 7244 11245
rect 7173 11133 7254 11146
rect 7173 11078 7186 11133
rect 7244 11078 7254 11133
rect 7173 11067 7254 11078
rect 6158 10990 7052 11035
rect 4590 10787 4650 10990
rect 6992 10787 7052 10990
rect 7184 10787 7244 11067
rect 7302 10787 7362 11346
rect 8011 11304 8071 11720
rect 8129 11694 8189 11720
rect 8366 11694 8426 11720
rect 8484 11694 8544 11720
rect 8492 11571 8558 11574
rect 8602 11571 8662 11720
rect 8492 11558 8662 11571
rect 8492 11524 8508 11558
rect 8542 11524 8662 11558
rect 8492 11511 8662 11524
rect 8492 11508 8558 11511
rect 7533 11287 8071 11304
rect 7533 11253 7552 11287
rect 7586 11253 8071 11287
rect 7533 11247 8071 11253
rect 7533 11237 7602 11247
rect 7533 11235 7598 11237
rect 7417 10897 7483 10913
rect 7417 10863 7433 10897
rect 7467 10863 7483 10897
rect 7417 10847 7483 10863
rect 7420 10787 7480 10847
rect 7538 10787 7598 11235
rect 8602 11035 8662 11511
rect 7734 10990 8662 11035
rect 9290 11438 9350 11724
rect 9408 11698 9468 11724
rect 9526 11698 9586 11724
rect 9731 11698 9791 11724
rect 9290 11421 9426 11438
rect 9290 11366 9349 11421
rect 9407 11366 9426 11421
rect 9290 11351 9426 11366
rect 9290 11039 9350 11351
rect 9849 11306 9909 11724
rect 9967 11698 10027 11724
rect 10198 11698 10258 11724
rect 10316 11698 10376 11724
rect 10434 11698 10494 11724
rect 10552 11698 10612 11724
rect 10317 11538 10376 11698
rect 10317 11537 10380 11538
rect 10314 11521 10380 11537
rect 10314 11487 10330 11521
rect 10364 11487 10380 11521
rect 10314 11471 10380 11487
rect 10417 11422 10512 11437
rect 10417 11367 10436 11422
rect 10494 11399 10512 11422
rect 10670 11399 10730 11724
rect 10788 11698 10848 11724
rect 11025 11698 11085 11724
rect 10494 11367 10730 11399
rect 10417 11350 10730 11367
rect 9849 11249 10376 11306
rect 10316 11150 10376 11249
rect 10305 11137 10386 11150
rect 10305 11082 10318 11137
rect 10376 11082 10386 11137
rect 10305 11071 10386 11082
rect 9290 10994 10184 11039
rect 7734 10787 7794 10990
rect 10124 10791 10184 10994
rect 10316 10791 10376 11071
rect 10434 10791 10494 11350
rect 11143 11308 11203 11724
rect 11261 11698 11321 11724
rect 11498 11698 11558 11724
rect 11616 11698 11676 11724
rect 11624 11575 11690 11578
rect 11734 11575 11794 11724
rect 11624 11562 11794 11575
rect 11624 11528 11640 11562
rect 11674 11528 11794 11562
rect 11624 11515 11794 11528
rect 11624 11512 11690 11515
rect 10665 11291 11203 11308
rect 10665 11257 10684 11291
rect 10718 11257 11203 11291
rect 10665 11251 11203 11257
rect 10665 11241 10734 11251
rect 10665 11239 10730 11241
rect 10549 10901 10615 10917
rect 10549 10867 10565 10901
rect 10599 10867 10615 10901
rect 10549 10851 10615 10867
rect 10552 10791 10612 10851
rect 10670 10791 10730 11239
rect 11734 11039 11794 11515
rect 10866 10994 11794 11039
rect 12434 11438 12494 11724
rect 12552 11698 12612 11724
rect 12670 11698 12730 11724
rect 12875 11698 12935 11724
rect 12434 11421 12570 11438
rect 12434 11366 12493 11421
rect 12551 11366 12570 11421
rect 12434 11351 12570 11366
rect 12434 11039 12494 11351
rect 12993 11306 13053 11724
rect 13111 11698 13171 11724
rect 13342 11698 13402 11724
rect 13460 11698 13520 11724
rect 13578 11698 13638 11724
rect 13696 11698 13756 11724
rect 13461 11538 13520 11698
rect 13461 11537 13524 11538
rect 13458 11521 13524 11537
rect 13458 11487 13474 11521
rect 13508 11487 13524 11521
rect 13458 11471 13524 11487
rect 13561 11422 13656 11437
rect 13561 11367 13580 11422
rect 13638 11399 13656 11422
rect 13814 11399 13874 11724
rect 13932 11698 13992 11724
rect 14169 11698 14229 11724
rect 13638 11367 13874 11399
rect 13561 11350 13874 11367
rect 12993 11249 13520 11306
rect 13460 11150 13520 11249
rect 13449 11137 13530 11150
rect 13449 11082 13462 11137
rect 13520 11082 13530 11137
rect 13449 11071 13530 11082
rect 12434 10994 13328 11039
rect 10866 10791 10926 10994
rect 13268 10791 13328 10994
rect 13460 10791 13520 11071
rect 13578 10791 13638 11350
rect 14287 11308 14347 11724
rect 14405 11698 14465 11724
rect 14642 11698 14702 11724
rect 14760 11698 14820 11724
rect 14768 11575 14834 11578
rect 14878 11575 14938 11724
rect 17844 11936 18140 11975
rect 17844 11920 17904 11936
rect 17962 11920 18022 11936
rect 18080 11920 18140 11936
rect 18780 11936 19076 11975
rect 18780 11920 18840 11936
rect 18898 11920 18958 11936
rect 19016 11920 19076 11936
rect 20988 11936 21284 11975
rect 20988 11920 21048 11936
rect 21106 11920 21166 11936
rect 21224 11920 21284 11936
rect 21912 11940 22208 11979
rect 21912 11924 21972 11940
rect 22030 11924 22090 11940
rect 22148 11924 22208 11940
rect 24120 11940 24416 11979
rect 24120 11924 24180 11940
rect 24238 11924 24298 11940
rect 24356 11924 24416 11940
rect 25056 11940 25352 11979
rect 25056 11924 25116 11940
rect 25174 11924 25234 11940
rect 25292 11924 25352 11940
rect 27264 11940 27560 11979
rect 27264 11924 27324 11940
rect 27382 11924 27442 11940
rect 27500 11924 27560 11940
rect 14768 11562 14938 11575
rect 14768 11528 14784 11562
rect 14818 11528 14938 11562
rect 14768 11515 14938 11528
rect 14768 11512 14834 11515
rect 13809 11291 14347 11308
rect 13809 11257 13828 11291
rect 13862 11257 14347 11291
rect 13809 11251 14347 11257
rect 13809 11241 13878 11251
rect 13809 11239 13874 11241
rect 13693 10901 13759 10917
rect 13693 10867 13709 10901
rect 13743 10867 13759 10901
rect 13693 10851 13759 10867
rect 13696 10791 13756 10851
rect 13814 10791 13874 11239
rect 14878 11039 14938 11515
rect 14010 10994 14938 11039
rect 15636 11434 15696 11720
rect 15754 11694 15814 11720
rect 15872 11694 15932 11720
rect 16077 11694 16137 11720
rect 15636 11417 15772 11434
rect 15636 11362 15695 11417
rect 15753 11362 15772 11417
rect 15636 11347 15772 11362
rect 15636 11035 15696 11347
rect 16195 11302 16255 11720
rect 16313 11694 16373 11720
rect 16544 11694 16604 11720
rect 16662 11694 16722 11720
rect 16780 11694 16840 11720
rect 16898 11694 16958 11720
rect 16663 11534 16722 11694
rect 16663 11533 16726 11534
rect 16660 11517 16726 11533
rect 16660 11483 16676 11517
rect 16710 11483 16726 11517
rect 16660 11467 16726 11483
rect 16763 11418 16858 11433
rect 16763 11363 16782 11418
rect 16840 11395 16858 11418
rect 17016 11395 17076 11720
rect 17134 11694 17194 11720
rect 17371 11694 17431 11720
rect 16840 11363 17076 11395
rect 16763 11346 17076 11363
rect 16195 11245 16722 11302
rect 16662 11146 16722 11245
rect 16651 11133 16732 11146
rect 16651 11078 16664 11133
rect 16722 11078 16732 11133
rect 16651 11067 16732 11078
rect 14010 10791 14070 10994
rect 15636 10990 16530 11035
rect 3848 10561 3908 10587
rect 4040 10361 4100 10387
rect 4158 10361 4218 10387
rect 4276 10361 4336 10387
rect 4394 10361 4454 10387
rect 4215 10306 4281 10314
rect 4590 10306 4650 10587
rect 6992 10561 7052 10587
rect 7184 10361 7244 10387
rect 7302 10361 7362 10387
rect 7420 10361 7480 10387
rect 7538 10361 7598 10387
rect 4215 10298 4650 10306
rect 4215 10264 4231 10298
rect 4265 10264 4650 10298
rect 4215 10255 4650 10264
rect 7359 10306 7425 10314
rect 7734 10306 7794 10587
rect 10124 10565 10184 10591
rect 10316 10365 10376 10391
rect 10434 10365 10494 10391
rect 10552 10365 10612 10391
rect 10670 10365 10730 10391
rect 7359 10298 7794 10306
rect 7359 10264 7375 10298
rect 7409 10264 7794 10298
rect 7359 10255 7794 10264
rect 10491 10310 10557 10318
rect 10866 10310 10926 10591
rect 13268 10565 13328 10591
rect 16470 10787 16530 10990
rect 16662 10787 16722 11067
rect 16780 10787 16840 11346
rect 17489 11304 17549 11720
rect 17607 11694 17667 11720
rect 17844 11694 17904 11720
rect 17962 11694 18022 11720
rect 17970 11571 18036 11574
rect 18080 11571 18140 11720
rect 17970 11558 18140 11571
rect 17970 11524 17986 11558
rect 18020 11524 18140 11558
rect 17970 11511 18140 11524
rect 17970 11508 18036 11511
rect 17011 11287 17549 11304
rect 17011 11253 17030 11287
rect 17064 11253 17549 11287
rect 17011 11247 17549 11253
rect 17011 11237 17080 11247
rect 17011 11235 17076 11237
rect 16895 10897 16961 10913
rect 16895 10863 16911 10897
rect 16945 10863 16961 10897
rect 16895 10847 16961 10863
rect 16898 10787 16958 10847
rect 17016 10787 17076 11235
rect 18080 11035 18140 11511
rect 17212 10990 18140 11035
rect 18780 11434 18840 11720
rect 18898 11694 18958 11720
rect 19016 11694 19076 11720
rect 19221 11694 19281 11720
rect 18780 11417 18916 11434
rect 18780 11362 18839 11417
rect 18897 11362 18916 11417
rect 18780 11347 18916 11362
rect 18780 11035 18840 11347
rect 19339 11302 19399 11720
rect 19457 11694 19517 11720
rect 19688 11694 19748 11720
rect 19806 11694 19866 11720
rect 19924 11694 19984 11720
rect 20042 11694 20102 11720
rect 19807 11534 19866 11694
rect 19807 11533 19870 11534
rect 19804 11517 19870 11533
rect 19804 11483 19820 11517
rect 19854 11483 19870 11517
rect 19804 11467 19870 11483
rect 19907 11418 20002 11433
rect 19907 11363 19926 11418
rect 19984 11395 20002 11418
rect 20160 11395 20220 11720
rect 20278 11694 20338 11720
rect 20515 11694 20575 11720
rect 19984 11363 20220 11395
rect 19907 11346 20220 11363
rect 19339 11245 19866 11302
rect 19806 11146 19866 11245
rect 19795 11133 19876 11146
rect 19795 11078 19808 11133
rect 19866 11078 19876 11133
rect 19795 11067 19876 11078
rect 18780 10990 19674 11035
rect 17212 10787 17272 10990
rect 19614 10787 19674 10990
rect 19806 10787 19866 11067
rect 19924 10787 19984 11346
rect 20633 11304 20693 11720
rect 20751 11694 20811 11720
rect 20988 11694 21048 11720
rect 21106 11694 21166 11720
rect 21114 11571 21180 11574
rect 21224 11571 21284 11720
rect 21114 11558 21284 11571
rect 21114 11524 21130 11558
rect 21164 11524 21284 11558
rect 21114 11511 21284 11524
rect 21114 11508 21180 11511
rect 20155 11287 20693 11304
rect 20155 11253 20174 11287
rect 20208 11253 20693 11287
rect 20155 11247 20693 11253
rect 20155 11237 20224 11247
rect 20155 11235 20220 11237
rect 20039 10897 20105 10913
rect 20039 10863 20055 10897
rect 20089 10863 20105 10897
rect 20039 10847 20105 10863
rect 20042 10787 20102 10847
rect 20160 10787 20220 11235
rect 21224 11035 21284 11511
rect 20356 10990 21284 11035
rect 21912 11438 21972 11724
rect 22030 11698 22090 11724
rect 22148 11698 22208 11724
rect 22353 11698 22413 11724
rect 21912 11421 22048 11438
rect 21912 11366 21971 11421
rect 22029 11366 22048 11421
rect 21912 11351 22048 11366
rect 21912 11039 21972 11351
rect 22471 11306 22531 11724
rect 22589 11698 22649 11724
rect 22820 11698 22880 11724
rect 22938 11698 22998 11724
rect 23056 11698 23116 11724
rect 23174 11698 23234 11724
rect 22939 11538 22998 11698
rect 22939 11537 23002 11538
rect 22936 11521 23002 11537
rect 22936 11487 22952 11521
rect 22986 11487 23002 11521
rect 22936 11471 23002 11487
rect 23039 11422 23134 11437
rect 23039 11367 23058 11422
rect 23116 11399 23134 11422
rect 23292 11399 23352 11724
rect 23410 11698 23470 11724
rect 23647 11698 23707 11724
rect 23116 11367 23352 11399
rect 23039 11350 23352 11367
rect 22471 11249 22998 11306
rect 22938 11150 22998 11249
rect 22927 11137 23008 11150
rect 22927 11082 22940 11137
rect 22998 11082 23008 11137
rect 22927 11071 23008 11082
rect 21912 10994 22806 11039
rect 20356 10787 20416 10990
rect 22746 10791 22806 10994
rect 22938 10791 22998 11071
rect 23056 10791 23116 11350
rect 23765 11308 23825 11724
rect 23883 11698 23943 11724
rect 24120 11698 24180 11724
rect 24238 11698 24298 11724
rect 24246 11575 24312 11578
rect 24356 11575 24416 11724
rect 24246 11562 24416 11575
rect 24246 11528 24262 11562
rect 24296 11528 24416 11562
rect 24246 11515 24416 11528
rect 24246 11512 24312 11515
rect 23287 11291 23825 11308
rect 23287 11257 23306 11291
rect 23340 11257 23825 11291
rect 23287 11251 23825 11257
rect 23287 11241 23356 11251
rect 23287 11239 23352 11241
rect 23171 10901 23237 10917
rect 23171 10867 23187 10901
rect 23221 10867 23237 10901
rect 23171 10851 23237 10867
rect 23174 10791 23234 10851
rect 23292 10791 23352 11239
rect 24356 11039 24416 11515
rect 23488 10994 24416 11039
rect 25056 11438 25116 11724
rect 25174 11698 25234 11724
rect 25292 11698 25352 11724
rect 25497 11698 25557 11724
rect 25056 11421 25192 11438
rect 25056 11366 25115 11421
rect 25173 11366 25192 11421
rect 25056 11351 25192 11366
rect 25056 11039 25116 11351
rect 25615 11306 25675 11724
rect 25733 11698 25793 11724
rect 25964 11698 26024 11724
rect 26082 11698 26142 11724
rect 26200 11698 26260 11724
rect 26318 11698 26378 11724
rect 26083 11538 26142 11698
rect 26083 11537 26146 11538
rect 26080 11521 26146 11537
rect 26080 11487 26096 11521
rect 26130 11487 26146 11521
rect 26080 11471 26146 11487
rect 26183 11422 26278 11437
rect 26183 11367 26202 11422
rect 26260 11399 26278 11422
rect 26436 11399 26496 11724
rect 26554 11698 26614 11724
rect 26791 11698 26851 11724
rect 26260 11367 26496 11399
rect 26183 11350 26496 11367
rect 25615 11249 26142 11306
rect 26082 11150 26142 11249
rect 26071 11137 26152 11150
rect 26071 11082 26084 11137
rect 26142 11082 26152 11137
rect 26071 11071 26152 11082
rect 25056 10994 25950 11039
rect 23488 10791 23548 10994
rect 25890 10791 25950 10994
rect 26082 10791 26142 11071
rect 26200 10791 26260 11350
rect 26909 11308 26969 11724
rect 27027 11698 27087 11724
rect 27264 11698 27324 11724
rect 27382 11698 27442 11724
rect 27390 11575 27456 11578
rect 27500 11575 27560 11724
rect 27390 11562 27560 11575
rect 27390 11528 27406 11562
rect 27440 11528 27560 11562
rect 27390 11515 27560 11528
rect 27390 11512 27456 11515
rect 26431 11291 26969 11308
rect 26431 11257 26450 11291
rect 26484 11257 26969 11291
rect 26431 11251 26969 11257
rect 26431 11241 26500 11251
rect 26431 11239 26496 11241
rect 26315 10901 26381 10917
rect 26315 10867 26331 10901
rect 26365 10867 26381 10901
rect 26315 10851 26381 10867
rect 26318 10791 26378 10851
rect 26436 10791 26496 11239
rect 27500 11039 27560 11515
rect 26632 10994 27560 11039
rect 26632 10791 26692 10994
rect 13460 10365 13520 10391
rect 13578 10365 13638 10391
rect 13696 10365 13756 10391
rect 13814 10365 13874 10391
rect 10491 10302 10926 10310
rect 10491 10268 10507 10302
rect 10541 10268 10926 10302
rect 10491 10259 10926 10268
rect 13635 10310 13701 10318
rect 14010 10310 14070 10591
rect 16470 10561 16530 10587
rect 16662 10361 16722 10387
rect 16780 10361 16840 10387
rect 16898 10361 16958 10387
rect 17016 10361 17076 10387
rect 13635 10302 14070 10310
rect 13635 10268 13651 10302
rect 13685 10268 14070 10302
rect 13635 10259 14070 10268
rect 16837 10306 16903 10314
rect 17212 10306 17272 10587
rect 19614 10561 19674 10587
rect 19806 10361 19866 10387
rect 19924 10361 19984 10387
rect 20042 10361 20102 10387
rect 20160 10361 20220 10387
rect 16837 10298 17272 10306
rect 16837 10264 16853 10298
rect 16887 10264 17272 10298
rect 4215 10248 4281 10255
rect 7359 10248 7425 10255
rect 10491 10252 10557 10259
rect 13635 10252 13701 10259
rect 16837 10255 17272 10264
rect 19981 10306 20047 10314
rect 20356 10306 20416 10587
rect 22746 10565 22806 10591
rect 22938 10365 22998 10391
rect 23056 10365 23116 10391
rect 23174 10365 23234 10391
rect 23292 10365 23352 10391
rect 19981 10298 20416 10306
rect 19981 10264 19997 10298
rect 20031 10264 20416 10298
rect 19981 10255 20416 10264
rect 23113 10310 23179 10318
rect 23488 10310 23548 10591
rect 25890 10565 25950 10591
rect 26082 10365 26142 10391
rect 26200 10365 26260 10391
rect 26318 10365 26378 10391
rect 26436 10365 26496 10391
rect 23113 10302 23548 10310
rect 23113 10268 23129 10302
rect 23163 10268 23548 10302
rect 23113 10259 23548 10268
rect 26257 10310 26323 10318
rect 26632 10310 26692 10591
rect 26257 10302 26692 10310
rect 26257 10268 26273 10302
rect 26307 10268 26692 10302
rect 26257 10259 26692 10268
rect 16837 10248 16903 10255
rect 19981 10248 20047 10255
rect 23113 10252 23179 10259
rect 26257 10252 26323 10259
rect 3445 9403 3741 9442
rect 3445 9388 3505 9403
rect 3563 9388 3623 9403
rect 3681 9388 3741 9403
rect 3912 9403 4208 9442
rect 3912 9388 3972 9403
rect 4030 9388 4090 9403
rect 4148 9388 4208 9403
rect 4266 9403 4562 9442
rect 4266 9388 4326 9403
rect 4384 9388 4444 9403
rect 4502 9388 4562 9403
rect 4739 9403 5035 9442
rect 4739 9388 4799 9403
rect 4857 9388 4917 9403
rect 4975 9388 5035 9403
rect 6589 9403 6885 9442
rect 6589 9388 6649 9403
rect 6707 9388 6767 9403
rect 6825 9388 6885 9403
rect 7056 9403 7352 9442
rect 7056 9388 7116 9403
rect 7174 9388 7234 9403
rect 7292 9388 7352 9403
rect 7410 9403 7706 9442
rect 7410 9388 7470 9403
rect 7528 9388 7588 9403
rect 7646 9388 7706 9403
rect 7883 9403 8179 9442
rect 7883 9388 7943 9403
rect 8001 9388 8061 9403
rect 8119 9388 8179 9403
rect 9721 9407 10017 9446
rect 9721 9392 9781 9407
rect 9839 9392 9899 9407
rect 9957 9392 10017 9407
rect 10188 9407 10484 9446
rect 10188 9392 10248 9407
rect 10306 9392 10366 9407
rect 10424 9392 10484 9407
rect 10542 9407 10838 9446
rect 10542 9392 10602 9407
rect 10660 9392 10720 9407
rect 10778 9392 10838 9407
rect 11015 9407 11311 9446
rect 11015 9392 11075 9407
rect 11133 9392 11193 9407
rect 11251 9392 11311 9407
rect 12865 9407 13161 9446
rect 12865 9392 12925 9407
rect 12983 9392 13043 9407
rect 13101 9392 13161 9407
rect 13332 9407 13628 9446
rect 13332 9392 13392 9407
rect 13450 9392 13510 9407
rect 13568 9392 13628 9407
rect 13686 9407 13982 9446
rect 13686 9392 13746 9407
rect 13804 9392 13864 9407
rect 13922 9392 13982 9407
rect 14159 9407 14455 9446
rect 14159 9392 14219 9407
rect 14277 9392 14337 9407
rect 14395 9392 14455 9407
rect 16067 9403 16363 9442
rect 3004 9204 3300 9243
rect 3004 9188 3064 9204
rect 3122 9188 3182 9204
rect 3240 9188 3300 9204
rect 5212 9204 5508 9243
rect 5212 9188 5272 9204
rect 5330 9188 5390 9204
rect 5448 9188 5508 9204
rect 6148 9204 6444 9243
rect 6148 9188 6208 9204
rect 6266 9188 6326 9204
rect 6384 9188 6444 9204
rect 8356 9204 8652 9243
rect 8356 9188 8416 9204
rect 8474 9188 8534 9204
rect 8592 9188 8652 9204
rect 9280 9208 9576 9247
rect 9280 9192 9340 9208
rect 9398 9192 9458 9208
rect 9516 9192 9576 9208
rect 11488 9208 11784 9247
rect 11488 9192 11548 9208
rect 11606 9192 11666 9208
rect 11724 9192 11784 9208
rect 12424 9208 12720 9247
rect 12424 9192 12484 9208
rect 12542 9192 12602 9208
rect 12660 9192 12720 9208
rect 16067 9388 16127 9403
rect 16185 9388 16245 9403
rect 16303 9388 16363 9403
rect 16534 9403 16830 9442
rect 16534 9388 16594 9403
rect 16652 9388 16712 9403
rect 16770 9388 16830 9403
rect 16888 9403 17184 9442
rect 16888 9388 16948 9403
rect 17006 9388 17066 9403
rect 17124 9388 17184 9403
rect 17361 9403 17657 9442
rect 17361 9388 17421 9403
rect 17479 9388 17539 9403
rect 17597 9388 17657 9403
rect 19211 9403 19507 9442
rect 19211 9388 19271 9403
rect 19329 9388 19389 9403
rect 19447 9388 19507 9403
rect 19678 9403 19974 9442
rect 19678 9388 19738 9403
rect 19796 9388 19856 9403
rect 19914 9388 19974 9403
rect 20032 9403 20328 9442
rect 20032 9388 20092 9403
rect 20150 9388 20210 9403
rect 20268 9388 20328 9403
rect 20505 9403 20801 9442
rect 20505 9388 20565 9403
rect 20623 9388 20683 9403
rect 20741 9388 20801 9403
rect 22343 9407 22639 9446
rect 22343 9392 22403 9407
rect 22461 9392 22521 9407
rect 22579 9392 22639 9407
rect 22810 9407 23106 9446
rect 22810 9392 22870 9407
rect 22928 9392 22988 9407
rect 23046 9392 23106 9407
rect 23164 9407 23460 9446
rect 23164 9392 23224 9407
rect 23282 9392 23342 9407
rect 23400 9392 23460 9407
rect 23637 9407 23933 9446
rect 23637 9392 23697 9407
rect 23755 9392 23815 9407
rect 23873 9392 23933 9407
rect 25487 9407 25783 9446
rect 25487 9392 25547 9407
rect 25605 9392 25665 9407
rect 25723 9392 25783 9407
rect 25954 9407 26250 9446
rect 25954 9392 26014 9407
rect 26072 9392 26132 9407
rect 26190 9392 26250 9407
rect 26308 9407 26604 9446
rect 26308 9392 26368 9407
rect 26426 9392 26486 9407
rect 26544 9392 26604 9407
rect 26781 9407 27077 9446
rect 26781 9392 26841 9407
rect 26899 9392 26959 9407
rect 27017 9392 27077 9407
rect 14632 9208 14928 9247
rect 14632 9192 14692 9208
rect 14750 9192 14810 9208
rect 14868 9192 14928 9208
rect 15626 9204 15922 9243
rect 15626 9188 15686 9204
rect 15744 9188 15804 9204
rect 15862 9188 15922 9204
rect 3004 8702 3064 8988
rect 3122 8962 3182 8988
rect 3240 8962 3300 8988
rect 3445 8962 3505 8988
rect 3004 8685 3140 8702
rect 3004 8630 3063 8685
rect 3121 8630 3140 8685
rect 3004 8615 3140 8630
rect 3004 8303 3064 8615
rect 3563 8570 3623 8988
rect 3681 8962 3741 8988
rect 3912 8962 3972 8988
rect 4030 8962 4090 8988
rect 4148 8962 4208 8988
rect 4266 8962 4326 8988
rect 4031 8802 4090 8962
rect 4031 8801 4094 8802
rect 4028 8785 4094 8801
rect 4028 8751 4044 8785
rect 4078 8751 4094 8785
rect 4028 8735 4094 8751
rect 4131 8686 4226 8701
rect 4131 8631 4150 8686
rect 4208 8663 4226 8686
rect 4384 8663 4444 8988
rect 4502 8962 4562 8988
rect 4739 8962 4799 8988
rect 4208 8631 4444 8663
rect 4131 8614 4444 8631
rect 3563 8513 4090 8570
rect 4030 8414 4090 8513
rect 4019 8401 4100 8414
rect 4019 8346 4032 8401
rect 4090 8346 4100 8401
rect 4019 8335 4100 8346
rect 3004 8258 3898 8303
rect 3838 8055 3898 8258
rect 4030 8055 4090 8335
rect 4148 8055 4208 8614
rect 4857 8572 4917 8988
rect 4975 8962 5035 8988
rect 5212 8962 5272 8988
rect 5330 8962 5390 8988
rect 5338 8839 5404 8842
rect 5448 8839 5508 8988
rect 5338 8826 5508 8839
rect 5338 8792 5354 8826
rect 5388 8792 5508 8826
rect 5338 8779 5508 8792
rect 5338 8776 5404 8779
rect 4379 8555 4917 8572
rect 4379 8521 4398 8555
rect 4432 8521 4917 8555
rect 4379 8515 4917 8521
rect 4379 8505 4448 8515
rect 4379 8503 4444 8505
rect 4263 8165 4329 8181
rect 4263 8131 4279 8165
rect 4313 8131 4329 8165
rect 4263 8115 4329 8131
rect 4266 8055 4326 8115
rect 4384 8055 4444 8503
rect 5448 8303 5508 8779
rect 4580 8258 5508 8303
rect 6148 8702 6208 8988
rect 6266 8962 6326 8988
rect 6384 8962 6444 8988
rect 6589 8962 6649 8988
rect 6148 8685 6284 8702
rect 6148 8630 6207 8685
rect 6265 8630 6284 8685
rect 6148 8615 6284 8630
rect 6148 8303 6208 8615
rect 6707 8570 6767 8988
rect 6825 8962 6885 8988
rect 7056 8962 7116 8988
rect 7174 8962 7234 8988
rect 7292 8962 7352 8988
rect 7410 8962 7470 8988
rect 7175 8802 7234 8962
rect 7175 8801 7238 8802
rect 7172 8785 7238 8801
rect 7172 8751 7188 8785
rect 7222 8751 7238 8785
rect 7172 8735 7238 8751
rect 7275 8686 7370 8701
rect 7275 8631 7294 8686
rect 7352 8663 7370 8686
rect 7528 8663 7588 8988
rect 7646 8962 7706 8988
rect 7883 8962 7943 8988
rect 7352 8631 7588 8663
rect 7275 8614 7588 8631
rect 6707 8513 7234 8570
rect 7174 8414 7234 8513
rect 7163 8401 7244 8414
rect 7163 8346 7176 8401
rect 7234 8346 7244 8401
rect 7163 8335 7244 8346
rect 6148 8258 7042 8303
rect 4580 8055 4640 8258
rect 6982 8055 7042 8258
rect 7174 8055 7234 8335
rect 7292 8055 7352 8614
rect 8001 8572 8061 8988
rect 8119 8962 8179 8988
rect 8356 8962 8416 8988
rect 8474 8962 8534 8988
rect 8482 8839 8548 8842
rect 8592 8839 8652 8988
rect 8482 8826 8652 8839
rect 8482 8792 8498 8826
rect 8532 8792 8652 8826
rect 8482 8779 8652 8792
rect 8482 8776 8548 8779
rect 7523 8555 8061 8572
rect 7523 8521 7542 8555
rect 7576 8521 8061 8555
rect 7523 8515 8061 8521
rect 7523 8505 7592 8515
rect 7523 8503 7588 8505
rect 7407 8165 7473 8181
rect 7407 8131 7423 8165
rect 7457 8131 7473 8165
rect 7407 8115 7473 8131
rect 7410 8055 7470 8115
rect 7528 8055 7588 8503
rect 8592 8303 8652 8779
rect 7724 8258 8652 8303
rect 9280 8706 9340 8992
rect 9398 8966 9458 8992
rect 9516 8966 9576 8992
rect 9721 8966 9781 8992
rect 9280 8689 9416 8706
rect 9280 8634 9339 8689
rect 9397 8634 9416 8689
rect 9280 8619 9416 8634
rect 9280 8307 9340 8619
rect 9839 8574 9899 8992
rect 9957 8966 10017 8992
rect 10188 8966 10248 8992
rect 10306 8966 10366 8992
rect 10424 8966 10484 8992
rect 10542 8966 10602 8992
rect 10307 8806 10366 8966
rect 10307 8805 10370 8806
rect 10304 8789 10370 8805
rect 10304 8755 10320 8789
rect 10354 8755 10370 8789
rect 10304 8739 10370 8755
rect 10407 8690 10502 8705
rect 10407 8635 10426 8690
rect 10484 8667 10502 8690
rect 10660 8667 10720 8992
rect 10778 8966 10838 8992
rect 11015 8966 11075 8992
rect 10484 8635 10720 8667
rect 10407 8618 10720 8635
rect 9839 8517 10366 8574
rect 10306 8418 10366 8517
rect 10295 8405 10376 8418
rect 10295 8350 10308 8405
rect 10366 8350 10376 8405
rect 10295 8339 10376 8350
rect 9280 8262 10174 8307
rect 7724 8055 7784 8258
rect 10114 8059 10174 8262
rect 10306 8059 10366 8339
rect 10424 8059 10484 8618
rect 11133 8576 11193 8992
rect 11251 8966 11311 8992
rect 11488 8966 11548 8992
rect 11606 8966 11666 8992
rect 11614 8843 11680 8846
rect 11724 8843 11784 8992
rect 11614 8830 11784 8843
rect 11614 8796 11630 8830
rect 11664 8796 11784 8830
rect 11614 8783 11784 8796
rect 11614 8780 11680 8783
rect 10655 8559 11193 8576
rect 10655 8525 10674 8559
rect 10708 8525 11193 8559
rect 10655 8519 11193 8525
rect 10655 8509 10724 8519
rect 10655 8507 10720 8509
rect 10539 8169 10605 8185
rect 10539 8135 10555 8169
rect 10589 8135 10605 8169
rect 10539 8119 10605 8135
rect 10542 8059 10602 8119
rect 10660 8059 10720 8507
rect 11724 8307 11784 8783
rect 10856 8262 11784 8307
rect 12424 8706 12484 8992
rect 12542 8966 12602 8992
rect 12660 8966 12720 8992
rect 12865 8966 12925 8992
rect 12424 8689 12560 8706
rect 12424 8634 12483 8689
rect 12541 8634 12560 8689
rect 12424 8619 12560 8634
rect 12424 8307 12484 8619
rect 12983 8574 13043 8992
rect 13101 8966 13161 8992
rect 13332 8966 13392 8992
rect 13450 8966 13510 8992
rect 13568 8966 13628 8992
rect 13686 8966 13746 8992
rect 13451 8806 13510 8966
rect 13451 8805 13514 8806
rect 13448 8789 13514 8805
rect 13448 8755 13464 8789
rect 13498 8755 13514 8789
rect 13448 8739 13514 8755
rect 13551 8690 13646 8705
rect 13551 8635 13570 8690
rect 13628 8667 13646 8690
rect 13804 8667 13864 8992
rect 13922 8966 13982 8992
rect 14159 8966 14219 8992
rect 13628 8635 13864 8667
rect 13551 8618 13864 8635
rect 12983 8517 13510 8574
rect 13450 8418 13510 8517
rect 13439 8405 13520 8418
rect 13439 8350 13452 8405
rect 13510 8350 13520 8405
rect 13439 8339 13520 8350
rect 12424 8262 13318 8307
rect 10856 8059 10916 8262
rect 13258 8059 13318 8262
rect 13450 8059 13510 8339
rect 13568 8059 13628 8618
rect 14277 8576 14337 8992
rect 14395 8966 14455 8992
rect 14632 8966 14692 8992
rect 14750 8966 14810 8992
rect 14758 8843 14824 8846
rect 14868 8843 14928 8992
rect 17834 9204 18130 9243
rect 17834 9188 17894 9204
rect 17952 9188 18012 9204
rect 18070 9188 18130 9204
rect 18770 9204 19066 9243
rect 18770 9188 18830 9204
rect 18888 9188 18948 9204
rect 19006 9188 19066 9204
rect 20978 9204 21274 9243
rect 20978 9188 21038 9204
rect 21096 9188 21156 9204
rect 21214 9188 21274 9204
rect 21902 9208 22198 9247
rect 21902 9192 21962 9208
rect 22020 9192 22080 9208
rect 22138 9192 22198 9208
rect 24110 9208 24406 9247
rect 24110 9192 24170 9208
rect 24228 9192 24288 9208
rect 24346 9192 24406 9208
rect 25046 9208 25342 9247
rect 25046 9192 25106 9208
rect 25164 9192 25224 9208
rect 25282 9192 25342 9208
rect 27254 9208 27550 9247
rect 27254 9192 27314 9208
rect 27372 9192 27432 9208
rect 27490 9192 27550 9208
rect 14758 8830 14928 8843
rect 14758 8796 14774 8830
rect 14808 8796 14928 8830
rect 14758 8783 14928 8796
rect 14758 8780 14824 8783
rect 13799 8559 14337 8576
rect 13799 8525 13818 8559
rect 13852 8525 14337 8559
rect 13799 8519 14337 8525
rect 13799 8509 13868 8519
rect 13799 8507 13864 8509
rect 13683 8169 13749 8185
rect 13683 8135 13699 8169
rect 13733 8135 13749 8169
rect 13683 8119 13749 8135
rect 13686 8059 13746 8119
rect 13804 8059 13864 8507
rect 14868 8307 14928 8783
rect 14000 8262 14928 8307
rect 15626 8702 15686 8988
rect 15744 8962 15804 8988
rect 15862 8962 15922 8988
rect 16067 8962 16127 8988
rect 15626 8685 15762 8702
rect 15626 8630 15685 8685
rect 15743 8630 15762 8685
rect 15626 8615 15762 8630
rect 15626 8303 15686 8615
rect 16185 8570 16245 8988
rect 16303 8962 16363 8988
rect 16534 8962 16594 8988
rect 16652 8962 16712 8988
rect 16770 8962 16830 8988
rect 16888 8962 16948 8988
rect 16653 8802 16712 8962
rect 16653 8801 16716 8802
rect 16650 8785 16716 8801
rect 16650 8751 16666 8785
rect 16700 8751 16716 8785
rect 16650 8735 16716 8751
rect 16753 8686 16848 8701
rect 16753 8631 16772 8686
rect 16830 8663 16848 8686
rect 17006 8663 17066 8988
rect 17124 8962 17184 8988
rect 17361 8962 17421 8988
rect 16830 8631 17066 8663
rect 16753 8614 17066 8631
rect 16185 8513 16712 8570
rect 16652 8414 16712 8513
rect 16641 8401 16722 8414
rect 16641 8346 16654 8401
rect 16712 8346 16722 8401
rect 16641 8335 16722 8346
rect 14000 8059 14060 8262
rect 15626 8258 16520 8303
rect 3838 7829 3898 7855
rect 4030 7629 4090 7655
rect 4148 7629 4208 7655
rect 4266 7629 4326 7655
rect 4384 7629 4444 7655
rect 4205 7574 4271 7582
rect 4580 7574 4640 7855
rect 6982 7829 7042 7855
rect 7174 7629 7234 7655
rect 7292 7629 7352 7655
rect 7410 7629 7470 7655
rect 7528 7629 7588 7655
rect 4205 7566 4640 7574
rect 4205 7532 4221 7566
rect 4255 7532 4640 7566
rect 4205 7523 4640 7532
rect 7349 7574 7415 7582
rect 7724 7574 7784 7855
rect 10114 7833 10174 7859
rect 10306 7633 10366 7659
rect 10424 7633 10484 7659
rect 10542 7633 10602 7659
rect 10660 7633 10720 7659
rect 7349 7566 7784 7574
rect 7349 7532 7365 7566
rect 7399 7532 7784 7566
rect 7349 7523 7784 7532
rect 10481 7578 10547 7586
rect 10856 7578 10916 7859
rect 13258 7833 13318 7859
rect 16460 8055 16520 8258
rect 16652 8055 16712 8335
rect 16770 8055 16830 8614
rect 17479 8572 17539 8988
rect 17597 8962 17657 8988
rect 17834 8962 17894 8988
rect 17952 8962 18012 8988
rect 17960 8839 18026 8842
rect 18070 8839 18130 8988
rect 17960 8826 18130 8839
rect 17960 8792 17976 8826
rect 18010 8792 18130 8826
rect 17960 8779 18130 8792
rect 17960 8776 18026 8779
rect 17001 8555 17539 8572
rect 17001 8521 17020 8555
rect 17054 8521 17539 8555
rect 17001 8515 17539 8521
rect 17001 8505 17070 8515
rect 17001 8503 17066 8505
rect 16885 8165 16951 8181
rect 16885 8131 16901 8165
rect 16935 8131 16951 8165
rect 16885 8115 16951 8131
rect 16888 8055 16948 8115
rect 17006 8055 17066 8503
rect 18070 8303 18130 8779
rect 17202 8258 18130 8303
rect 18770 8702 18830 8988
rect 18888 8962 18948 8988
rect 19006 8962 19066 8988
rect 19211 8962 19271 8988
rect 18770 8685 18906 8702
rect 18770 8630 18829 8685
rect 18887 8630 18906 8685
rect 18770 8615 18906 8630
rect 18770 8303 18830 8615
rect 19329 8570 19389 8988
rect 19447 8962 19507 8988
rect 19678 8962 19738 8988
rect 19796 8962 19856 8988
rect 19914 8962 19974 8988
rect 20032 8962 20092 8988
rect 19797 8802 19856 8962
rect 19797 8801 19860 8802
rect 19794 8785 19860 8801
rect 19794 8751 19810 8785
rect 19844 8751 19860 8785
rect 19794 8735 19860 8751
rect 19897 8686 19992 8701
rect 19897 8631 19916 8686
rect 19974 8663 19992 8686
rect 20150 8663 20210 8988
rect 20268 8962 20328 8988
rect 20505 8962 20565 8988
rect 19974 8631 20210 8663
rect 19897 8614 20210 8631
rect 19329 8513 19856 8570
rect 19796 8414 19856 8513
rect 19785 8401 19866 8414
rect 19785 8346 19798 8401
rect 19856 8346 19866 8401
rect 19785 8335 19866 8346
rect 18770 8258 19664 8303
rect 17202 8055 17262 8258
rect 19604 8055 19664 8258
rect 19796 8055 19856 8335
rect 19914 8055 19974 8614
rect 20623 8572 20683 8988
rect 20741 8962 20801 8988
rect 20978 8962 21038 8988
rect 21096 8962 21156 8988
rect 21104 8839 21170 8842
rect 21214 8839 21274 8988
rect 21104 8826 21274 8839
rect 21104 8792 21120 8826
rect 21154 8792 21274 8826
rect 21104 8779 21274 8792
rect 21104 8776 21170 8779
rect 20145 8555 20683 8572
rect 20145 8521 20164 8555
rect 20198 8521 20683 8555
rect 20145 8515 20683 8521
rect 20145 8505 20214 8515
rect 20145 8503 20210 8505
rect 20029 8165 20095 8181
rect 20029 8131 20045 8165
rect 20079 8131 20095 8165
rect 20029 8115 20095 8131
rect 20032 8055 20092 8115
rect 20150 8055 20210 8503
rect 21214 8303 21274 8779
rect 20346 8258 21274 8303
rect 21902 8706 21962 8992
rect 22020 8966 22080 8992
rect 22138 8966 22198 8992
rect 22343 8966 22403 8992
rect 21902 8689 22038 8706
rect 21902 8634 21961 8689
rect 22019 8634 22038 8689
rect 21902 8619 22038 8634
rect 21902 8307 21962 8619
rect 22461 8574 22521 8992
rect 22579 8966 22639 8992
rect 22810 8966 22870 8992
rect 22928 8966 22988 8992
rect 23046 8966 23106 8992
rect 23164 8966 23224 8992
rect 22929 8806 22988 8966
rect 22929 8805 22992 8806
rect 22926 8789 22992 8805
rect 22926 8755 22942 8789
rect 22976 8755 22992 8789
rect 22926 8739 22992 8755
rect 23029 8690 23124 8705
rect 23029 8635 23048 8690
rect 23106 8667 23124 8690
rect 23282 8667 23342 8992
rect 23400 8966 23460 8992
rect 23637 8966 23697 8992
rect 23106 8635 23342 8667
rect 23029 8618 23342 8635
rect 22461 8517 22988 8574
rect 22928 8418 22988 8517
rect 22917 8405 22998 8418
rect 22917 8350 22930 8405
rect 22988 8350 22998 8405
rect 22917 8339 22998 8350
rect 21902 8262 22796 8307
rect 20346 8055 20406 8258
rect 22736 8059 22796 8262
rect 22928 8059 22988 8339
rect 23046 8059 23106 8618
rect 23755 8576 23815 8992
rect 23873 8966 23933 8992
rect 24110 8966 24170 8992
rect 24228 8966 24288 8992
rect 24236 8843 24302 8846
rect 24346 8843 24406 8992
rect 24236 8830 24406 8843
rect 24236 8796 24252 8830
rect 24286 8796 24406 8830
rect 24236 8783 24406 8796
rect 24236 8780 24302 8783
rect 23277 8559 23815 8576
rect 23277 8525 23296 8559
rect 23330 8525 23815 8559
rect 23277 8519 23815 8525
rect 23277 8509 23346 8519
rect 23277 8507 23342 8509
rect 23161 8169 23227 8185
rect 23161 8135 23177 8169
rect 23211 8135 23227 8169
rect 23161 8119 23227 8135
rect 23164 8059 23224 8119
rect 23282 8059 23342 8507
rect 24346 8307 24406 8783
rect 23478 8262 24406 8307
rect 25046 8706 25106 8992
rect 25164 8966 25224 8992
rect 25282 8966 25342 8992
rect 25487 8966 25547 8992
rect 25046 8689 25182 8706
rect 25046 8634 25105 8689
rect 25163 8634 25182 8689
rect 25046 8619 25182 8634
rect 25046 8307 25106 8619
rect 25605 8574 25665 8992
rect 25723 8966 25783 8992
rect 25954 8966 26014 8992
rect 26072 8966 26132 8992
rect 26190 8966 26250 8992
rect 26308 8966 26368 8992
rect 26073 8806 26132 8966
rect 26073 8805 26136 8806
rect 26070 8789 26136 8805
rect 26070 8755 26086 8789
rect 26120 8755 26136 8789
rect 26070 8739 26136 8755
rect 26173 8690 26268 8705
rect 26173 8635 26192 8690
rect 26250 8667 26268 8690
rect 26426 8667 26486 8992
rect 26544 8966 26604 8992
rect 26781 8966 26841 8992
rect 26250 8635 26486 8667
rect 26173 8618 26486 8635
rect 25605 8517 26132 8574
rect 26072 8418 26132 8517
rect 26061 8405 26142 8418
rect 26061 8350 26074 8405
rect 26132 8350 26142 8405
rect 26061 8339 26142 8350
rect 25046 8262 25940 8307
rect 23478 8059 23538 8262
rect 25880 8059 25940 8262
rect 26072 8059 26132 8339
rect 26190 8059 26250 8618
rect 26899 8576 26959 8992
rect 27017 8966 27077 8992
rect 27254 8966 27314 8992
rect 27372 8966 27432 8992
rect 27380 8843 27446 8846
rect 27490 8843 27550 8992
rect 27380 8830 27550 8843
rect 27380 8796 27396 8830
rect 27430 8796 27550 8830
rect 27380 8783 27550 8796
rect 27380 8780 27446 8783
rect 26421 8559 26959 8576
rect 26421 8525 26440 8559
rect 26474 8525 26959 8559
rect 26421 8519 26959 8525
rect 26421 8509 26490 8519
rect 26421 8507 26486 8509
rect 26305 8169 26371 8185
rect 26305 8135 26321 8169
rect 26355 8135 26371 8169
rect 26305 8119 26371 8135
rect 26308 8059 26368 8119
rect 26426 8059 26486 8507
rect 27490 8307 27550 8783
rect 26622 8262 27550 8307
rect 26622 8059 26682 8262
rect 13450 7633 13510 7659
rect 13568 7633 13628 7659
rect 13686 7633 13746 7659
rect 13804 7633 13864 7659
rect 10481 7570 10916 7578
rect 10481 7536 10497 7570
rect 10531 7536 10916 7570
rect 10481 7527 10916 7536
rect 13625 7578 13691 7586
rect 14000 7578 14060 7859
rect 16460 7829 16520 7855
rect 16652 7629 16712 7655
rect 16770 7629 16830 7655
rect 16888 7629 16948 7655
rect 17006 7629 17066 7655
rect 13625 7570 14060 7578
rect 13625 7536 13641 7570
rect 13675 7536 14060 7570
rect 13625 7527 14060 7536
rect 16827 7574 16893 7582
rect 17202 7574 17262 7855
rect 19604 7829 19664 7855
rect 19796 7629 19856 7655
rect 19914 7629 19974 7655
rect 20032 7629 20092 7655
rect 20150 7629 20210 7655
rect 16827 7566 17262 7574
rect 16827 7532 16843 7566
rect 16877 7532 17262 7566
rect 4205 7516 4271 7523
rect 7349 7516 7415 7523
rect 10481 7520 10547 7527
rect 13625 7520 13691 7527
rect 16827 7523 17262 7532
rect 19971 7574 20037 7582
rect 20346 7574 20406 7855
rect 22736 7833 22796 7859
rect 22928 7633 22988 7659
rect 23046 7633 23106 7659
rect 23164 7633 23224 7659
rect 23282 7633 23342 7659
rect 19971 7566 20406 7574
rect 19971 7532 19987 7566
rect 20021 7532 20406 7566
rect 19971 7523 20406 7532
rect 23103 7578 23169 7586
rect 23478 7578 23538 7859
rect 25880 7833 25940 7859
rect 26072 7633 26132 7659
rect 26190 7633 26250 7659
rect 26308 7633 26368 7659
rect 26426 7633 26486 7659
rect 23103 7570 23538 7578
rect 23103 7536 23119 7570
rect 23153 7536 23538 7570
rect 23103 7527 23538 7536
rect 26247 7578 26313 7586
rect 26622 7578 26682 7859
rect 26247 7570 26682 7578
rect 26247 7536 26263 7570
rect 26297 7536 26682 7570
rect 26247 7527 26682 7536
rect 16827 7516 16893 7523
rect 19971 7516 20037 7523
rect 23103 7520 23169 7527
rect 26247 7520 26313 7527
rect 19473 6559 19533 6585
rect 19591 6559 19651 6585
rect 19709 6559 19769 6585
rect 20211 6563 20271 6589
rect 20329 6563 20389 6589
rect 20447 6563 20507 6589
rect 3225 6458 3521 6509
rect 3225 6443 3285 6458
rect 3343 6443 3403 6458
rect 3461 6443 3521 6458
rect 3579 6443 3639 6469
rect 3697 6443 3757 6469
rect 3815 6443 3875 6469
rect 5293 6460 5589 6511
rect 5293 6445 5353 6460
rect 5411 6445 5471 6460
rect 5529 6445 5589 6460
rect 5647 6445 5707 6471
rect 5765 6445 5825 6471
rect 5883 6445 5943 6471
rect 7362 6458 7658 6509
rect 2741 6243 2801 6269
rect 2859 6243 2919 6269
rect 2977 6243 3037 6269
rect 4062 6260 4358 6311
rect 4062 6243 4122 6260
rect 4180 6243 4240 6260
rect 4298 6243 4358 6260
rect 4809 6245 4869 6271
rect 4927 6245 4987 6271
rect 5045 6245 5105 6271
rect 7362 6443 7422 6458
rect 7480 6443 7540 6458
rect 7598 6443 7658 6458
rect 7716 6443 7776 6469
rect 7834 6443 7894 6469
rect 7952 6443 8012 6469
rect 9430 6460 9726 6511
rect 9430 6445 9490 6460
rect 9548 6445 9608 6460
rect 9666 6445 9726 6460
rect 9784 6445 9844 6471
rect 9902 6445 9962 6471
rect 10020 6445 10080 6471
rect 11499 6460 11795 6511
rect 11499 6445 11559 6460
rect 11617 6445 11677 6460
rect 11735 6445 11795 6460
rect 11853 6445 11913 6471
rect 11971 6445 12031 6471
rect 12089 6445 12149 6471
rect 13567 6462 13863 6513
rect 13567 6447 13627 6462
rect 13685 6447 13745 6462
rect 13803 6447 13863 6462
rect 13921 6447 13981 6473
rect 14039 6447 14099 6473
rect 14157 6447 14217 6473
rect 15636 6460 15932 6511
rect 6130 6262 6426 6313
rect 6130 6245 6190 6262
rect 6248 6245 6308 6262
rect 6366 6245 6426 6262
rect 6878 6243 6938 6269
rect 6996 6243 7056 6269
rect 7114 6243 7174 6269
rect 2741 6026 2801 6043
rect 2859 6026 2919 6043
rect 2977 6026 3037 6043
rect 3225 6026 3285 6043
rect 2741 5975 3285 6026
rect 3343 6017 3403 6043
rect 3461 6017 3521 6043
rect 3579 6024 3639 6043
rect 3697 6024 3757 6043
rect 3815 6024 3875 6043
rect 4062 6024 4122 6043
rect 4180 6024 4240 6043
rect 2866 5696 2926 5975
rect 3579 5973 4122 6024
rect 4164 6017 4240 6024
rect 4298 6017 4358 6043
rect 4809 6028 4869 6045
rect 4927 6028 4987 6045
rect 5045 6028 5105 6045
rect 5293 6028 5353 6045
rect 4164 5973 4239 6017
rect 4809 5977 5353 6028
rect 5411 6019 5471 6045
rect 5529 6019 5589 6045
rect 5647 6026 5707 6045
rect 5765 6026 5825 6045
rect 5883 6026 5943 6045
rect 6130 6026 6190 6045
rect 6248 6026 6308 6045
rect 4164 5886 4224 5973
rect 4096 5876 4224 5886
rect 4096 5842 4112 5876
rect 4146 5842 4224 5876
rect 3168 5773 3464 5833
rect 3168 5750 3228 5773
rect 3286 5750 3346 5773
rect 3404 5750 3464 5773
rect 3522 5774 3818 5834
rect 4096 5832 4224 5842
rect 3522 5750 3582 5774
rect 3640 5750 3700 5774
rect 3758 5750 3818 5774
rect 2702 5682 2926 5696
rect 2702 5648 2718 5682
rect 2752 5648 2926 5682
rect 2702 5636 2926 5648
rect 2866 5123 2926 5636
rect 3168 5324 3228 5350
rect 3136 5183 3203 5190
rect 3286 5183 3346 5350
rect 3404 5324 3464 5350
rect 3522 5324 3582 5350
rect 3136 5174 3346 5183
rect 3136 5140 3152 5174
rect 3186 5140 3346 5174
rect 3136 5124 3346 5140
rect 2866 5107 3017 5123
rect 2866 5073 2967 5107
rect 3001 5073 3017 5107
rect 2866 5057 3017 5073
rect 2866 5018 2926 5057
rect 3286 5018 3346 5124
rect 3640 5183 3700 5350
rect 3758 5324 3818 5350
rect 3783 5183 3850 5190
rect 3640 5174 3850 5183
rect 3640 5140 3800 5174
rect 3834 5140 3850 5174
rect 3640 5124 3850 5140
rect 3402 5090 3468 5106
rect 3402 5056 3418 5090
rect 3452 5056 3468 5090
rect 3402 5040 3468 5056
rect 3520 5091 3586 5106
rect 3520 5057 3536 5091
rect 3570 5057 3586 5091
rect 3520 5041 3586 5057
rect 3404 5018 3464 5040
rect 3522 5018 3582 5041
rect 3640 5018 3700 5124
rect 4164 5122 4224 5832
rect 4934 5698 4994 5977
rect 5647 5975 6190 6026
rect 6232 6019 6308 6026
rect 6366 6019 6426 6045
rect 8199 6260 8495 6311
rect 8199 6243 8259 6260
rect 8317 6243 8377 6260
rect 8435 6243 8495 6260
rect 8946 6245 9006 6271
rect 9064 6245 9124 6271
rect 9182 6245 9242 6271
rect 10267 6262 10563 6313
rect 10267 6245 10327 6262
rect 10385 6245 10445 6262
rect 10503 6245 10563 6262
rect 11015 6245 11075 6271
rect 11133 6245 11193 6271
rect 11251 6245 11311 6271
rect 12336 6262 12632 6313
rect 12336 6245 12396 6262
rect 12454 6245 12514 6262
rect 12572 6245 12632 6262
rect 13083 6247 13143 6273
rect 13201 6247 13261 6273
rect 13319 6247 13379 6273
rect 15636 6445 15696 6460
rect 15754 6445 15814 6460
rect 15872 6445 15932 6460
rect 15990 6445 16050 6471
rect 16108 6445 16168 6471
rect 16226 6445 16286 6471
rect 17704 6462 18000 6513
rect 17704 6447 17764 6462
rect 17822 6447 17882 6462
rect 17940 6447 18000 6462
rect 18058 6447 18118 6473
rect 18176 6447 18236 6473
rect 18294 6447 18354 6473
rect 14404 6264 14700 6315
rect 14404 6247 14464 6264
rect 14522 6247 14582 6264
rect 14640 6247 14700 6264
rect 15152 6245 15212 6271
rect 15270 6245 15330 6271
rect 15388 6245 15448 6271
rect 6878 6026 6938 6043
rect 6996 6026 7056 6043
rect 7114 6026 7174 6043
rect 7362 6026 7422 6043
rect 6232 5975 6307 6019
rect 6878 5975 7422 6026
rect 7480 6017 7540 6043
rect 7598 6017 7658 6043
rect 7716 6024 7776 6043
rect 7834 6024 7894 6043
rect 7952 6024 8012 6043
rect 8199 6024 8259 6043
rect 8317 6024 8377 6043
rect 6232 5888 6292 5975
rect 6164 5878 6292 5888
rect 6164 5844 6180 5878
rect 6214 5844 6292 5878
rect 5236 5775 5532 5835
rect 5236 5752 5296 5775
rect 5354 5752 5414 5775
rect 5472 5752 5532 5775
rect 5590 5776 5886 5836
rect 6164 5834 6292 5844
rect 5590 5752 5650 5776
rect 5708 5752 5768 5776
rect 5826 5752 5886 5776
rect 4770 5684 4994 5698
rect 4770 5650 4786 5684
rect 4820 5650 4994 5684
rect 4770 5638 4994 5650
rect 4074 5106 4224 5122
rect 4074 5072 4090 5106
rect 4124 5072 4224 5106
rect 4074 5056 4224 5072
rect 4164 5018 4224 5056
rect 4934 5125 4994 5638
rect 5236 5326 5296 5352
rect 5204 5185 5271 5192
rect 5354 5185 5414 5352
rect 5472 5326 5532 5352
rect 5590 5326 5650 5352
rect 5204 5176 5414 5185
rect 5204 5142 5220 5176
rect 5254 5142 5414 5176
rect 5204 5126 5414 5142
rect 4934 5109 5085 5125
rect 4934 5075 5035 5109
rect 5069 5075 5085 5109
rect 4934 5059 5085 5075
rect 4934 5020 4994 5059
rect 5354 5020 5414 5126
rect 5708 5185 5768 5352
rect 5826 5326 5886 5352
rect 5851 5185 5918 5192
rect 5708 5176 5918 5185
rect 5708 5142 5868 5176
rect 5902 5142 5918 5176
rect 5708 5126 5918 5142
rect 5470 5092 5536 5108
rect 5470 5058 5486 5092
rect 5520 5058 5536 5092
rect 5470 5042 5536 5058
rect 5588 5093 5654 5108
rect 5588 5059 5604 5093
rect 5638 5059 5654 5093
rect 5588 5043 5654 5059
rect 5472 5020 5532 5042
rect 5590 5020 5650 5043
rect 5708 5020 5768 5126
rect 6232 5124 6292 5834
rect 7003 5696 7063 5975
rect 7716 5973 8259 6024
rect 8301 6017 8377 6024
rect 8435 6017 8495 6043
rect 8946 6028 9006 6045
rect 9064 6028 9124 6045
rect 9182 6028 9242 6045
rect 9430 6028 9490 6045
rect 8301 5973 8376 6017
rect 8946 5977 9490 6028
rect 9548 6019 9608 6045
rect 9666 6019 9726 6045
rect 9784 6026 9844 6045
rect 9902 6026 9962 6045
rect 10020 6026 10080 6045
rect 10267 6026 10327 6045
rect 10385 6026 10445 6045
rect 8301 5886 8361 5973
rect 8233 5876 8361 5886
rect 8233 5842 8249 5876
rect 8283 5842 8361 5876
rect 7305 5773 7601 5833
rect 7305 5750 7365 5773
rect 7423 5750 7483 5773
rect 7541 5750 7601 5773
rect 7659 5774 7955 5834
rect 8233 5832 8361 5842
rect 7659 5750 7719 5774
rect 7777 5750 7837 5774
rect 7895 5750 7955 5774
rect 6839 5682 7063 5696
rect 6839 5648 6855 5682
rect 6889 5648 7063 5682
rect 6839 5636 7063 5648
rect 6142 5108 6292 5124
rect 6142 5074 6158 5108
rect 6192 5074 6292 5108
rect 6142 5058 6292 5074
rect 6232 5020 6292 5058
rect 7003 5123 7063 5636
rect 7305 5324 7365 5350
rect 7273 5183 7340 5190
rect 7423 5183 7483 5350
rect 7541 5324 7601 5350
rect 7659 5324 7719 5350
rect 7273 5174 7483 5183
rect 7273 5140 7289 5174
rect 7323 5140 7483 5174
rect 7273 5124 7483 5140
rect 7003 5107 7154 5123
rect 7003 5073 7104 5107
rect 7138 5073 7154 5107
rect 7003 5057 7154 5073
rect 2866 4792 2926 4818
rect 4164 4792 4224 4818
rect 4934 4794 4994 4820
rect 7003 5018 7063 5057
rect 7423 5018 7483 5124
rect 7777 5183 7837 5350
rect 7895 5324 7955 5350
rect 7920 5183 7987 5190
rect 7777 5174 7987 5183
rect 7777 5140 7937 5174
rect 7971 5140 7987 5174
rect 7777 5124 7987 5140
rect 7539 5090 7605 5106
rect 7539 5056 7555 5090
rect 7589 5056 7605 5090
rect 7539 5040 7605 5056
rect 7657 5091 7723 5106
rect 7657 5057 7673 5091
rect 7707 5057 7723 5091
rect 7657 5041 7723 5057
rect 7541 5018 7601 5040
rect 7659 5018 7719 5041
rect 7777 5018 7837 5124
rect 8301 5122 8361 5832
rect 9071 5698 9131 5977
rect 9784 5975 10327 6026
rect 10369 6019 10445 6026
rect 10503 6019 10563 6045
rect 11015 6028 11075 6045
rect 11133 6028 11193 6045
rect 11251 6028 11311 6045
rect 11499 6028 11559 6045
rect 10369 5975 10444 6019
rect 11015 5977 11559 6028
rect 11617 6019 11677 6045
rect 11735 6019 11795 6045
rect 11853 6026 11913 6045
rect 11971 6026 12031 6045
rect 12089 6026 12149 6045
rect 12336 6026 12396 6045
rect 12454 6026 12514 6045
rect 10369 5888 10429 5975
rect 10301 5878 10429 5888
rect 10301 5844 10317 5878
rect 10351 5844 10429 5878
rect 9373 5775 9669 5835
rect 9373 5752 9433 5775
rect 9491 5752 9551 5775
rect 9609 5752 9669 5775
rect 9727 5776 10023 5836
rect 10301 5834 10429 5844
rect 9727 5752 9787 5776
rect 9845 5752 9905 5776
rect 9963 5752 10023 5776
rect 8907 5684 9131 5698
rect 8907 5650 8923 5684
rect 8957 5650 9131 5684
rect 8907 5638 9131 5650
rect 8211 5106 8361 5122
rect 8211 5072 8227 5106
rect 8261 5072 8361 5106
rect 8211 5056 8361 5072
rect 8301 5018 8361 5056
rect 9071 5125 9131 5638
rect 9373 5326 9433 5352
rect 9341 5185 9408 5192
rect 9491 5185 9551 5352
rect 9609 5326 9669 5352
rect 9727 5326 9787 5352
rect 9341 5176 9551 5185
rect 9341 5142 9357 5176
rect 9391 5142 9551 5176
rect 9341 5126 9551 5142
rect 9071 5109 9222 5125
rect 9071 5075 9172 5109
rect 9206 5075 9222 5109
rect 9071 5059 9222 5075
rect 9071 5020 9131 5059
rect 9491 5020 9551 5126
rect 9845 5185 9905 5352
rect 9963 5326 10023 5352
rect 9988 5185 10055 5192
rect 9845 5176 10055 5185
rect 9845 5142 10005 5176
rect 10039 5142 10055 5176
rect 9845 5126 10055 5142
rect 9607 5092 9673 5108
rect 9607 5058 9623 5092
rect 9657 5058 9673 5092
rect 9607 5042 9673 5058
rect 9725 5093 9791 5108
rect 9725 5059 9741 5093
rect 9775 5059 9791 5093
rect 9725 5043 9791 5059
rect 9609 5020 9669 5042
rect 9727 5020 9787 5043
rect 9845 5020 9905 5126
rect 10369 5124 10429 5834
rect 11140 5698 11200 5977
rect 11853 5975 12396 6026
rect 12438 6019 12514 6026
rect 12572 6019 12632 6045
rect 13083 6030 13143 6047
rect 13201 6030 13261 6047
rect 13319 6030 13379 6047
rect 13567 6030 13627 6047
rect 12438 5975 12513 6019
rect 13083 5979 13627 6030
rect 13685 6021 13745 6047
rect 13803 6021 13863 6047
rect 13921 6028 13981 6047
rect 14039 6028 14099 6047
rect 14157 6028 14217 6047
rect 14404 6028 14464 6047
rect 14522 6028 14582 6047
rect 12438 5888 12498 5975
rect 12370 5878 12498 5888
rect 12370 5844 12386 5878
rect 12420 5844 12498 5878
rect 11442 5775 11738 5835
rect 11442 5752 11502 5775
rect 11560 5752 11620 5775
rect 11678 5752 11738 5775
rect 11796 5776 12092 5836
rect 12370 5834 12498 5844
rect 11796 5752 11856 5776
rect 11914 5752 11974 5776
rect 12032 5752 12092 5776
rect 10976 5684 11200 5698
rect 10976 5650 10992 5684
rect 11026 5650 11200 5684
rect 10976 5638 11200 5650
rect 10279 5108 10429 5124
rect 10279 5074 10295 5108
rect 10329 5074 10429 5108
rect 10279 5058 10429 5074
rect 10369 5020 10429 5058
rect 11140 5125 11200 5638
rect 11442 5326 11502 5352
rect 11410 5185 11477 5192
rect 11560 5185 11620 5352
rect 11678 5326 11738 5352
rect 11796 5326 11856 5352
rect 11410 5176 11620 5185
rect 11410 5142 11426 5176
rect 11460 5142 11620 5176
rect 11410 5126 11620 5142
rect 11140 5109 11291 5125
rect 11140 5075 11241 5109
rect 11275 5075 11291 5109
rect 11140 5059 11291 5075
rect 11140 5020 11200 5059
rect 11560 5020 11620 5126
rect 11914 5185 11974 5352
rect 12032 5326 12092 5352
rect 12057 5185 12124 5192
rect 11914 5176 12124 5185
rect 11914 5142 12074 5176
rect 12108 5142 12124 5176
rect 11914 5126 12124 5142
rect 11676 5092 11742 5108
rect 11676 5058 11692 5092
rect 11726 5058 11742 5092
rect 11676 5042 11742 5058
rect 11794 5093 11860 5108
rect 11794 5059 11810 5093
rect 11844 5059 11860 5093
rect 11794 5043 11860 5059
rect 11678 5020 11738 5042
rect 11796 5020 11856 5043
rect 11914 5020 11974 5126
rect 12438 5124 12498 5834
rect 13208 5700 13268 5979
rect 13921 5977 14464 6028
rect 14506 6021 14582 6028
rect 14640 6021 14700 6047
rect 16473 6262 16769 6313
rect 16473 6245 16533 6262
rect 16591 6245 16651 6262
rect 16709 6245 16769 6262
rect 17220 6247 17280 6273
rect 17338 6247 17398 6273
rect 17456 6247 17516 6273
rect 20949 6559 21009 6585
rect 21067 6559 21127 6585
rect 21185 6559 21245 6585
rect 19473 6343 19533 6359
rect 19591 6343 19651 6359
rect 19709 6343 19769 6359
rect 18541 6264 18837 6315
rect 19473 6307 19769 6343
rect 20211 6341 20271 6363
rect 20329 6341 20389 6363
rect 20447 6341 20507 6363
rect 21691 6557 21751 6583
rect 21809 6557 21869 6583
rect 21927 6557 21987 6583
rect 22431 6557 22491 6583
rect 22549 6557 22609 6583
rect 22667 6557 22727 6583
rect 23169 6557 23229 6583
rect 23287 6557 23347 6583
rect 23405 6557 23465 6583
rect 23907 6557 23967 6583
rect 24025 6557 24085 6583
rect 24143 6557 24203 6583
rect 24645 6557 24705 6583
rect 24763 6557 24823 6583
rect 24881 6557 24941 6583
rect 18541 6247 18601 6264
rect 18659 6247 18719 6264
rect 18777 6247 18837 6264
rect 19591 6265 19651 6307
rect 20211 6305 20507 6341
rect 20949 6341 21009 6359
rect 21067 6341 21127 6359
rect 21185 6341 21245 6359
rect 20949 6305 21245 6341
rect 21691 6341 21751 6357
rect 21809 6341 21869 6357
rect 21927 6341 21987 6357
rect 21691 6305 21987 6341
rect 22431 6341 22491 6357
rect 22549 6341 22609 6357
rect 22667 6341 22727 6357
rect 22431 6305 22727 6341
rect 23169 6341 23229 6357
rect 23287 6341 23347 6357
rect 23405 6341 23465 6357
rect 23169 6305 23465 6341
rect 23907 6341 23967 6357
rect 24025 6341 24085 6357
rect 24143 6341 24203 6357
rect 23907 6305 24203 6341
rect 24645 6341 24705 6357
rect 24763 6341 24823 6357
rect 24881 6341 24941 6357
rect 24645 6305 24941 6341
rect 19591 6231 19603 6265
rect 19637 6231 19651 6265
rect 19591 6173 19651 6231
rect 20329 6263 20389 6305
rect 20329 6229 20341 6263
rect 20375 6229 20389 6263
rect 20329 6175 20389 6229
rect 21067 6263 21127 6305
rect 21067 6229 21079 6263
rect 21113 6229 21127 6263
rect 15152 6028 15212 6045
rect 15270 6028 15330 6045
rect 15388 6028 15448 6045
rect 15636 6028 15696 6045
rect 14506 5977 14581 6021
rect 15152 5977 15696 6028
rect 15754 6019 15814 6045
rect 15872 6019 15932 6045
rect 15990 6026 16050 6045
rect 16108 6026 16168 6045
rect 16226 6026 16286 6045
rect 16473 6026 16533 6045
rect 16591 6026 16651 6045
rect 14506 5890 14566 5977
rect 14438 5880 14566 5890
rect 14438 5846 14454 5880
rect 14488 5846 14566 5880
rect 13510 5777 13806 5837
rect 13510 5754 13570 5777
rect 13628 5754 13688 5777
rect 13746 5754 13806 5777
rect 13864 5778 14160 5838
rect 14438 5836 14566 5846
rect 13864 5754 13924 5778
rect 13982 5754 14042 5778
rect 14100 5754 14160 5778
rect 13044 5686 13268 5700
rect 13044 5652 13060 5686
rect 13094 5652 13268 5686
rect 13044 5640 13268 5652
rect 12348 5108 12498 5124
rect 12348 5074 12364 5108
rect 12398 5074 12498 5108
rect 12348 5058 12498 5074
rect 12438 5020 12498 5058
rect 13208 5127 13268 5640
rect 13510 5328 13570 5354
rect 13478 5187 13545 5194
rect 13628 5187 13688 5354
rect 13746 5328 13806 5354
rect 13864 5328 13924 5354
rect 13478 5178 13688 5187
rect 13478 5144 13494 5178
rect 13528 5144 13688 5178
rect 13478 5128 13688 5144
rect 13208 5111 13359 5127
rect 13208 5077 13309 5111
rect 13343 5077 13359 5111
rect 13208 5061 13359 5077
rect 13208 5022 13268 5061
rect 13628 5022 13688 5128
rect 13982 5187 14042 5354
rect 14100 5328 14160 5354
rect 14125 5187 14192 5194
rect 13982 5178 14192 5187
rect 13982 5144 14142 5178
rect 14176 5144 14192 5178
rect 13982 5128 14192 5144
rect 13744 5094 13810 5110
rect 13744 5060 13760 5094
rect 13794 5060 13810 5094
rect 13744 5044 13810 5060
rect 13862 5095 13928 5110
rect 13862 5061 13878 5095
rect 13912 5061 13928 5095
rect 13862 5045 13928 5061
rect 13746 5022 13806 5044
rect 13864 5022 13924 5045
rect 13982 5022 14042 5128
rect 14506 5126 14566 5836
rect 15277 5698 15337 5977
rect 15990 5975 16533 6026
rect 16575 6019 16651 6026
rect 16709 6019 16769 6045
rect 17220 6030 17280 6047
rect 17338 6030 17398 6047
rect 17456 6030 17516 6047
rect 17704 6030 17764 6047
rect 16575 5975 16650 6019
rect 17220 5979 17764 6030
rect 17822 6021 17882 6047
rect 17940 6021 18000 6047
rect 18058 6028 18118 6047
rect 18176 6028 18236 6047
rect 18294 6028 18354 6047
rect 18541 6028 18601 6047
rect 18659 6028 18719 6047
rect 16575 5888 16635 5975
rect 16507 5878 16635 5888
rect 16507 5844 16523 5878
rect 16557 5844 16635 5878
rect 15579 5775 15875 5835
rect 15579 5752 15639 5775
rect 15697 5752 15757 5775
rect 15815 5752 15875 5775
rect 15933 5776 16229 5836
rect 16507 5834 16635 5844
rect 15933 5752 15993 5776
rect 16051 5752 16111 5776
rect 16169 5752 16229 5776
rect 15113 5684 15337 5698
rect 15113 5650 15129 5684
rect 15163 5650 15337 5684
rect 15113 5638 15337 5650
rect 14416 5110 14566 5126
rect 14416 5076 14432 5110
rect 14466 5076 14566 5110
rect 14416 5060 14566 5076
rect 14506 5022 14566 5060
rect 15277 5125 15337 5638
rect 15579 5326 15639 5352
rect 15547 5185 15614 5192
rect 15697 5185 15757 5352
rect 15815 5326 15875 5352
rect 15933 5326 15993 5352
rect 15547 5176 15757 5185
rect 15547 5142 15563 5176
rect 15597 5142 15757 5176
rect 15547 5126 15757 5142
rect 15277 5109 15428 5125
rect 15277 5075 15378 5109
rect 15412 5075 15428 5109
rect 15277 5059 15428 5075
rect 6232 4794 6292 4820
rect 7003 4792 7063 4818
rect 3286 4592 3346 4618
rect 3404 4592 3464 4618
rect 3522 4592 3582 4618
rect 3640 4592 3700 4618
rect 5354 4594 5414 4620
rect 5472 4594 5532 4620
rect 5590 4594 5650 4620
rect 5708 4594 5768 4620
rect 8301 4792 8361 4818
rect 9071 4794 9131 4820
rect 10369 4794 10429 4820
rect 11140 4794 11200 4820
rect 12438 4794 12498 4820
rect 13208 4796 13268 4822
rect 15277 5020 15337 5059
rect 15697 5020 15757 5126
rect 16051 5185 16111 5352
rect 16169 5326 16229 5352
rect 16194 5185 16261 5192
rect 16051 5176 16261 5185
rect 16051 5142 16211 5176
rect 16245 5142 16261 5176
rect 16051 5126 16261 5142
rect 15813 5092 15879 5108
rect 15813 5058 15829 5092
rect 15863 5058 15879 5092
rect 15813 5042 15879 5058
rect 15931 5093 15997 5108
rect 15931 5059 15947 5093
rect 15981 5059 15997 5093
rect 15931 5043 15997 5059
rect 15815 5020 15875 5042
rect 15933 5020 15993 5043
rect 16051 5020 16111 5126
rect 16575 5124 16635 5834
rect 17345 5700 17405 5979
rect 18058 5977 18601 6028
rect 18643 6021 18719 6028
rect 18777 6021 18837 6047
rect 18643 5977 18718 6021
rect 18643 5890 18703 5977
rect 21067 6171 21127 6229
rect 21809 6263 21869 6305
rect 21809 6229 21821 6263
rect 21855 6229 21869 6263
rect 21809 6171 21869 6229
rect 22549 6263 22609 6305
rect 22549 6229 22561 6263
rect 22595 6229 22609 6263
rect 22549 6171 22609 6229
rect 23287 6263 23347 6305
rect 23287 6229 23299 6263
rect 23333 6229 23347 6263
rect 23287 6171 23347 6229
rect 24025 6263 24085 6305
rect 24025 6229 24037 6263
rect 24071 6229 24085 6263
rect 24025 6175 24085 6229
rect 24763 6263 24823 6305
rect 24763 6229 24775 6263
rect 24809 6229 24823 6263
rect 24763 6175 24823 6229
rect 19591 5947 19651 5973
rect 20329 5949 20389 5975
rect 21067 5945 21127 5971
rect 21809 5945 21869 5971
rect 22549 5945 22609 5971
rect 23287 5945 23347 5971
rect 24025 5949 24085 5975
rect 24763 5949 24823 5975
rect 18575 5880 18703 5890
rect 18575 5846 18591 5880
rect 18625 5846 18703 5880
rect 17647 5777 17943 5837
rect 17647 5754 17707 5777
rect 17765 5754 17825 5777
rect 17883 5754 17943 5777
rect 18001 5778 18297 5838
rect 18575 5836 18703 5846
rect 18001 5754 18061 5778
rect 18119 5754 18179 5778
rect 18237 5754 18297 5778
rect 17181 5686 17405 5700
rect 17181 5652 17197 5686
rect 17231 5652 17405 5686
rect 17181 5640 17405 5652
rect 16485 5108 16635 5124
rect 16485 5074 16501 5108
rect 16535 5074 16635 5108
rect 16485 5058 16635 5074
rect 16575 5020 16635 5058
rect 17345 5127 17405 5640
rect 17647 5328 17707 5354
rect 17615 5187 17682 5194
rect 17765 5187 17825 5354
rect 17883 5328 17943 5354
rect 18001 5328 18061 5354
rect 17615 5178 17825 5187
rect 17615 5144 17631 5178
rect 17665 5144 17825 5178
rect 17615 5128 17825 5144
rect 17345 5111 17496 5127
rect 17345 5077 17446 5111
rect 17480 5077 17496 5111
rect 17345 5061 17496 5077
rect 17345 5022 17405 5061
rect 17765 5022 17825 5128
rect 18119 5187 18179 5354
rect 18237 5328 18297 5354
rect 18262 5187 18329 5194
rect 18119 5178 18329 5187
rect 18119 5144 18279 5178
rect 18313 5144 18329 5178
rect 18119 5128 18329 5144
rect 17881 5094 17947 5110
rect 17881 5060 17897 5094
rect 17931 5060 17947 5094
rect 17881 5044 17947 5060
rect 17999 5095 18065 5110
rect 17999 5061 18015 5095
rect 18049 5061 18065 5095
rect 17999 5045 18065 5061
rect 17883 5022 17943 5044
rect 18001 5022 18061 5045
rect 18119 5022 18179 5128
rect 18643 5126 18703 5836
rect 18553 5110 18703 5126
rect 18553 5076 18569 5110
rect 18603 5076 18703 5110
rect 18553 5060 18703 5076
rect 18643 5022 18703 5060
rect 14506 4796 14566 4822
rect 15277 4794 15337 4820
rect 7423 4592 7483 4618
rect 7541 4592 7601 4618
rect 7659 4592 7719 4618
rect 7777 4592 7837 4618
rect 9491 4594 9551 4620
rect 9609 4594 9669 4620
rect 9727 4594 9787 4620
rect 9845 4594 9905 4620
rect 11560 4594 11620 4620
rect 11678 4594 11738 4620
rect 11796 4594 11856 4620
rect 11914 4594 11974 4620
rect 13628 4596 13688 4622
rect 13746 4596 13806 4622
rect 13864 4596 13924 4622
rect 13982 4596 14042 4622
rect 16575 4794 16635 4820
rect 17345 4796 17405 4822
rect 18643 4796 18703 4822
rect 15697 4594 15757 4620
rect 15815 4594 15875 4620
rect 15933 4594 15993 4620
rect 16051 4594 16111 4620
rect 17765 4596 17825 4622
rect 17883 4596 17943 4622
rect 18001 4596 18061 4622
rect 18119 4596 18179 4622
rect 747 2155 1043 2194
rect 747 2140 807 2155
rect 865 2140 925 2155
rect 983 2140 1043 2155
rect 1214 2155 1510 2194
rect 1214 2140 1274 2155
rect 1332 2140 1392 2155
rect 1450 2140 1510 2155
rect 1568 2155 1864 2194
rect 1568 2140 1628 2155
rect 1686 2140 1746 2155
rect 1804 2140 1864 2155
rect 2041 2155 2337 2194
rect 2041 2140 2101 2155
rect 2159 2140 2219 2155
rect 2277 2140 2337 2155
rect 3891 2155 4187 2194
rect 3891 2140 3951 2155
rect 4009 2140 4069 2155
rect 4127 2140 4187 2155
rect 4358 2155 4654 2194
rect 4358 2140 4418 2155
rect 4476 2140 4536 2155
rect 4594 2140 4654 2155
rect 4712 2155 5008 2194
rect 4712 2140 4772 2155
rect 4830 2140 4890 2155
rect 4948 2140 5008 2155
rect 5185 2155 5481 2194
rect 5185 2140 5245 2155
rect 5303 2140 5363 2155
rect 5421 2140 5481 2155
rect 7023 2159 7319 2198
rect 7023 2144 7083 2159
rect 7141 2144 7201 2159
rect 7259 2144 7319 2159
rect 7490 2159 7786 2198
rect 7490 2144 7550 2159
rect 7608 2144 7668 2159
rect 7726 2144 7786 2159
rect 7844 2159 8140 2198
rect 7844 2144 7904 2159
rect 7962 2144 8022 2159
rect 8080 2144 8140 2159
rect 8317 2159 8613 2198
rect 8317 2144 8377 2159
rect 8435 2144 8495 2159
rect 8553 2144 8613 2159
rect 10167 2159 10463 2198
rect 10167 2144 10227 2159
rect 10285 2144 10345 2159
rect 10403 2144 10463 2159
rect 10634 2159 10930 2198
rect 10634 2144 10694 2159
rect 10752 2144 10812 2159
rect 10870 2144 10930 2159
rect 10988 2159 11284 2198
rect 10988 2144 11048 2159
rect 11106 2144 11166 2159
rect 11224 2144 11284 2159
rect 11461 2159 11757 2198
rect 11461 2144 11521 2159
rect 11579 2144 11639 2159
rect 11697 2144 11757 2159
rect 13369 2155 13665 2194
rect 306 1956 602 1995
rect 306 1940 366 1956
rect 424 1940 484 1956
rect 542 1940 602 1956
rect 2514 1956 2810 1995
rect 2514 1940 2574 1956
rect 2632 1940 2692 1956
rect 2750 1940 2810 1956
rect 3450 1956 3746 1995
rect 3450 1940 3510 1956
rect 3568 1940 3628 1956
rect 3686 1940 3746 1956
rect 5658 1956 5954 1995
rect 5658 1940 5718 1956
rect 5776 1940 5836 1956
rect 5894 1940 5954 1956
rect 6582 1960 6878 1999
rect 6582 1944 6642 1960
rect 6700 1944 6760 1960
rect 6818 1944 6878 1960
rect 8790 1960 9086 1999
rect 8790 1944 8850 1960
rect 8908 1944 8968 1960
rect 9026 1944 9086 1960
rect 9726 1960 10022 1999
rect 9726 1944 9786 1960
rect 9844 1944 9904 1960
rect 9962 1944 10022 1960
rect 13369 2140 13429 2155
rect 13487 2140 13547 2155
rect 13605 2140 13665 2155
rect 13836 2155 14132 2194
rect 13836 2140 13896 2155
rect 13954 2140 14014 2155
rect 14072 2140 14132 2155
rect 14190 2155 14486 2194
rect 14190 2140 14250 2155
rect 14308 2140 14368 2155
rect 14426 2140 14486 2155
rect 14663 2155 14959 2194
rect 14663 2140 14723 2155
rect 14781 2140 14841 2155
rect 14899 2140 14959 2155
rect 16513 2155 16809 2194
rect 16513 2140 16573 2155
rect 16631 2140 16691 2155
rect 16749 2140 16809 2155
rect 16980 2155 17276 2194
rect 16980 2140 17040 2155
rect 17098 2140 17158 2155
rect 17216 2140 17276 2155
rect 17334 2155 17630 2194
rect 17334 2140 17394 2155
rect 17452 2140 17512 2155
rect 17570 2140 17630 2155
rect 17807 2155 18103 2194
rect 17807 2140 17867 2155
rect 17925 2140 17985 2155
rect 18043 2140 18103 2155
rect 19645 2159 19941 2198
rect 19645 2144 19705 2159
rect 19763 2144 19823 2159
rect 19881 2144 19941 2159
rect 20112 2159 20408 2198
rect 20112 2144 20172 2159
rect 20230 2144 20290 2159
rect 20348 2144 20408 2159
rect 20466 2159 20762 2198
rect 20466 2144 20526 2159
rect 20584 2144 20644 2159
rect 20702 2144 20762 2159
rect 20939 2159 21235 2198
rect 20939 2144 20999 2159
rect 21057 2144 21117 2159
rect 21175 2144 21235 2159
rect 22789 2159 23085 2198
rect 22789 2144 22849 2159
rect 22907 2144 22967 2159
rect 23025 2144 23085 2159
rect 23256 2159 23552 2198
rect 23256 2144 23316 2159
rect 23374 2144 23434 2159
rect 23492 2144 23552 2159
rect 23610 2159 23906 2198
rect 23610 2144 23670 2159
rect 23728 2144 23788 2159
rect 23846 2144 23906 2159
rect 24083 2159 24379 2198
rect 24083 2144 24143 2159
rect 24201 2144 24261 2159
rect 24319 2144 24379 2159
rect 11934 1960 12230 1999
rect 11934 1944 11994 1960
rect 12052 1944 12112 1960
rect 12170 1944 12230 1960
rect 12928 1956 13224 1995
rect 12928 1940 12988 1956
rect 13046 1940 13106 1956
rect 13164 1940 13224 1956
rect 306 1454 366 1740
rect 424 1714 484 1740
rect 542 1714 602 1740
rect 747 1714 807 1740
rect 306 1437 442 1454
rect 306 1382 365 1437
rect 423 1382 442 1437
rect 306 1367 442 1382
rect 306 1055 366 1367
rect 865 1322 925 1740
rect 983 1714 1043 1740
rect 1214 1714 1274 1740
rect 1332 1714 1392 1740
rect 1450 1714 1510 1740
rect 1568 1714 1628 1740
rect 1333 1554 1392 1714
rect 1333 1553 1396 1554
rect 1330 1537 1396 1553
rect 1330 1503 1346 1537
rect 1380 1503 1396 1537
rect 1330 1487 1396 1503
rect 1433 1438 1528 1453
rect 1433 1383 1452 1438
rect 1510 1415 1528 1438
rect 1686 1415 1746 1740
rect 1804 1714 1864 1740
rect 2041 1714 2101 1740
rect 1510 1383 1746 1415
rect 1433 1366 1746 1383
rect 865 1265 1392 1322
rect 1332 1166 1392 1265
rect 1321 1153 1402 1166
rect 1321 1098 1334 1153
rect 1392 1098 1402 1153
rect 1321 1087 1402 1098
rect 306 1010 1200 1055
rect 1140 807 1200 1010
rect 1332 807 1392 1087
rect 1450 807 1510 1366
rect 2159 1324 2219 1740
rect 2277 1714 2337 1740
rect 2514 1714 2574 1740
rect 2632 1714 2692 1740
rect 2640 1591 2706 1594
rect 2750 1591 2810 1740
rect 2640 1578 2810 1591
rect 2640 1544 2656 1578
rect 2690 1544 2810 1578
rect 2640 1531 2810 1544
rect 2640 1528 2706 1531
rect 1681 1307 2219 1324
rect 1681 1273 1700 1307
rect 1734 1273 2219 1307
rect 1681 1267 2219 1273
rect 1681 1257 1750 1267
rect 1681 1255 1746 1257
rect 1565 917 1631 933
rect 1565 883 1581 917
rect 1615 883 1631 917
rect 1565 867 1631 883
rect 1568 807 1628 867
rect 1686 807 1746 1255
rect 2750 1055 2810 1531
rect 1882 1010 2810 1055
rect 3450 1454 3510 1740
rect 3568 1714 3628 1740
rect 3686 1714 3746 1740
rect 3891 1714 3951 1740
rect 3450 1437 3586 1454
rect 3450 1382 3509 1437
rect 3567 1382 3586 1437
rect 3450 1367 3586 1382
rect 3450 1055 3510 1367
rect 4009 1322 4069 1740
rect 4127 1714 4187 1740
rect 4358 1714 4418 1740
rect 4476 1714 4536 1740
rect 4594 1714 4654 1740
rect 4712 1714 4772 1740
rect 4477 1554 4536 1714
rect 4477 1553 4540 1554
rect 4474 1537 4540 1553
rect 4474 1503 4490 1537
rect 4524 1503 4540 1537
rect 4474 1487 4540 1503
rect 4577 1438 4672 1453
rect 4577 1383 4596 1438
rect 4654 1415 4672 1438
rect 4830 1415 4890 1740
rect 4948 1714 5008 1740
rect 5185 1714 5245 1740
rect 4654 1383 4890 1415
rect 4577 1366 4890 1383
rect 4009 1265 4536 1322
rect 4476 1166 4536 1265
rect 4465 1153 4546 1166
rect 4465 1098 4478 1153
rect 4536 1098 4546 1153
rect 4465 1087 4546 1098
rect 3450 1010 4344 1055
rect 1882 807 1942 1010
rect 4284 807 4344 1010
rect 4476 807 4536 1087
rect 4594 807 4654 1366
rect 5303 1324 5363 1740
rect 5421 1714 5481 1740
rect 5658 1714 5718 1740
rect 5776 1714 5836 1740
rect 5784 1591 5850 1594
rect 5894 1591 5954 1740
rect 5784 1578 5954 1591
rect 5784 1544 5800 1578
rect 5834 1544 5954 1578
rect 5784 1531 5954 1544
rect 5784 1528 5850 1531
rect 4825 1307 5363 1324
rect 4825 1273 4844 1307
rect 4878 1273 5363 1307
rect 4825 1267 5363 1273
rect 4825 1257 4894 1267
rect 4825 1255 4890 1257
rect 4709 917 4775 933
rect 4709 883 4725 917
rect 4759 883 4775 917
rect 4709 867 4775 883
rect 4712 807 4772 867
rect 4830 807 4890 1255
rect 5894 1055 5954 1531
rect 5026 1010 5954 1055
rect 6582 1458 6642 1744
rect 6700 1718 6760 1744
rect 6818 1718 6878 1744
rect 7023 1718 7083 1744
rect 6582 1441 6718 1458
rect 6582 1386 6641 1441
rect 6699 1386 6718 1441
rect 6582 1371 6718 1386
rect 6582 1059 6642 1371
rect 7141 1326 7201 1744
rect 7259 1718 7319 1744
rect 7490 1718 7550 1744
rect 7608 1718 7668 1744
rect 7726 1718 7786 1744
rect 7844 1718 7904 1744
rect 7609 1558 7668 1718
rect 7609 1557 7672 1558
rect 7606 1541 7672 1557
rect 7606 1507 7622 1541
rect 7656 1507 7672 1541
rect 7606 1491 7672 1507
rect 7709 1442 7804 1457
rect 7709 1387 7728 1442
rect 7786 1419 7804 1442
rect 7962 1419 8022 1744
rect 8080 1718 8140 1744
rect 8317 1718 8377 1744
rect 7786 1387 8022 1419
rect 7709 1370 8022 1387
rect 7141 1269 7668 1326
rect 7608 1170 7668 1269
rect 7597 1157 7678 1170
rect 7597 1102 7610 1157
rect 7668 1102 7678 1157
rect 7597 1091 7678 1102
rect 6582 1014 7476 1059
rect 5026 807 5086 1010
rect 7416 811 7476 1014
rect 7608 811 7668 1091
rect 7726 811 7786 1370
rect 8435 1328 8495 1744
rect 8553 1718 8613 1744
rect 8790 1718 8850 1744
rect 8908 1718 8968 1744
rect 8916 1595 8982 1598
rect 9026 1595 9086 1744
rect 8916 1582 9086 1595
rect 8916 1548 8932 1582
rect 8966 1548 9086 1582
rect 8916 1535 9086 1548
rect 8916 1532 8982 1535
rect 7957 1311 8495 1328
rect 7957 1277 7976 1311
rect 8010 1277 8495 1311
rect 7957 1271 8495 1277
rect 7957 1261 8026 1271
rect 7957 1259 8022 1261
rect 7841 921 7907 937
rect 7841 887 7857 921
rect 7891 887 7907 921
rect 7841 871 7907 887
rect 7844 811 7904 871
rect 7962 811 8022 1259
rect 9026 1059 9086 1535
rect 8158 1014 9086 1059
rect 9726 1458 9786 1744
rect 9844 1718 9904 1744
rect 9962 1718 10022 1744
rect 10167 1718 10227 1744
rect 9726 1441 9862 1458
rect 9726 1386 9785 1441
rect 9843 1386 9862 1441
rect 9726 1371 9862 1386
rect 9726 1059 9786 1371
rect 10285 1326 10345 1744
rect 10403 1718 10463 1744
rect 10634 1718 10694 1744
rect 10752 1718 10812 1744
rect 10870 1718 10930 1744
rect 10988 1718 11048 1744
rect 10753 1558 10812 1718
rect 10753 1557 10816 1558
rect 10750 1541 10816 1557
rect 10750 1507 10766 1541
rect 10800 1507 10816 1541
rect 10750 1491 10816 1507
rect 10853 1442 10948 1457
rect 10853 1387 10872 1442
rect 10930 1419 10948 1442
rect 11106 1419 11166 1744
rect 11224 1718 11284 1744
rect 11461 1718 11521 1744
rect 10930 1387 11166 1419
rect 10853 1370 11166 1387
rect 10285 1269 10812 1326
rect 10752 1170 10812 1269
rect 10741 1157 10822 1170
rect 10741 1102 10754 1157
rect 10812 1102 10822 1157
rect 10741 1091 10822 1102
rect 9726 1014 10620 1059
rect 8158 811 8218 1014
rect 10560 811 10620 1014
rect 10752 811 10812 1091
rect 10870 811 10930 1370
rect 11579 1328 11639 1744
rect 11697 1718 11757 1744
rect 11934 1718 11994 1744
rect 12052 1718 12112 1744
rect 12060 1595 12126 1598
rect 12170 1595 12230 1744
rect 15136 1956 15432 1995
rect 15136 1940 15196 1956
rect 15254 1940 15314 1956
rect 15372 1940 15432 1956
rect 16072 1956 16368 1995
rect 16072 1940 16132 1956
rect 16190 1940 16250 1956
rect 16308 1940 16368 1956
rect 18280 1956 18576 1995
rect 18280 1940 18340 1956
rect 18398 1940 18458 1956
rect 18516 1940 18576 1956
rect 19204 1960 19500 1999
rect 19204 1944 19264 1960
rect 19322 1944 19382 1960
rect 19440 1944 19500 1960
rect 21412 1960 21708 1999
rect 21412 1944 21472 1960
rect 21530 1944 21590 1960
rect 21648 1944 21708 1960
rect 22348 1960 22644 1999
rect 22348 1944 22408 1960
rect 22466 1944 22526 1960
rect 22584 1944 22644 1960
rect 24556 1960 24852 1999
rect 24556 1944 24616 1960
rect 24674 1944 24734 1960
rect 24792 1944 24852 1960
rect 12060 1582 12230 1595
rect 12060 1548 12076 1582
rect 12110 1548 12230 1582
rect 12060 1535 12230 1548
rect 12060 1532 12126 1535
rect 11101 1311 11639 1328
rect 11101 1277 11120 1311
rect 11154 1277 11639 1311
rect 11101 1271 11639 1277
rect 11101 1261 11170 1271
rect 11101 1259 11166 1261
rect 10985 921 11051 937
rect 10985 887 11001 921
rect 11035 887 11051 921
rect 10985 871 11051 887
rect 10988 811 11048 871
rect 11106 811 11166 1259
rect 12170 1059 12230 1535
rect 11302 1014 12230 1059
rect 12928 1454 12988 1740
rect 13046 1714 13106 1740
rect 13164 1714 13224 1740
rect 13369 1714 13429 1740
rect 12928 1437 13064 1454
rect 12928 1382 12987 1437
rect 13045 1382 13064 1437
rect 12928 1367 13064 1382
rect 12928 1055 12988 1367
rect 13487 1322 13547 1740
rect 13605 1714 13665 1740
rect 13836 1714 13896 1740
rect 13954 1714 14014 1740
rect 14072 1714 14132 1740
rect 14190 1714 14250 1740
rect 13955 1554 14014 1714
rect 13955 1553 14018 1554
rect 13952 1537 14018 1553
rect 13952 1503 13968 1537
rect 14002 1503 14018 1537
rect 13952 1487 14018 1503
rect 14055 1438 14150 1453
rect 14055 1383 14074 1438
rect 14132 1415 14150 1438
rect 14308 1415 14368 1740
rect 14426 1714 14486 1740
rect 14663 1714 14723 1740
rect 14132 1383 14368 1415
rect 14055 1366 14368 1383
rect 13487 1265 14014 1322
rect 13954 1166 14014 1265
rect 13943 1153 14024 1166
rect 13943 1098 13956 1153
rect 14014 1098 14024 1153
rect 13943 1087 14024 1098
rect 11302 811 11362 1014
rect 12928 1010 13822 1055
rect 1140 581 1200 607
rect 1332 381 1392 407
rect 1450 381 1510 407
rect 1568 381 1628 407
rect 1686 381 1746 407
rect 1507 326 1573 334
rect 1882 326 1942 607
rect 4284 581 4344 607
rect 4476 381 4536 407
rect 4594 381 4654 407
rect 4712 381 4772 407
rect 4830 381 4890 407
rect 1507 318 1942 326
rect 1507 284 1523 318
rect 1557 284 1942 318
rect 1507 275 1942 284
rect 4651 326 4717 334
rect 5026 326 5086 607
rect 7416 585 7476 611
rect 7608 385 7668 411
rect 7726 385 7786 411
rect 7844 385 7904 411
rect 7962 385 8022 411
rect 4651 318 5086 326
rect 4651 284 4667 318
rect 4701 284 5086 318
rect 4651 275 5086 284
rect 7783 330 7849 338
rect 8158 330 8218 611
rect 10560 585 10620 611
rect 13762 807 13822 1010
rect 13954 807 14014 1087
rect 14072 807 14132 1366
rect 14781 1324 14841 1740
rect 14899 1714 14959 1740
rect 15136 1714 15196 1740
rect 15254 1714 15314 1740
rect 15262 1591 15328 1594
rect 15372 1591 15432 1740
rect 15262 1578 15432 1591
rect 15262 1544 15278 1578
rect 15312 1544 15432 1578
rect 15262 1531 15432 1544
rect 15262 1528 15328 1531
rect 14303 1307 14841 1324
rect 14303 1273 14322 1307
rect 14356 1273 14841 1307
rect 14303 1267 14841 1273
rect 14303 1257 14372 1267
rect 14303 1255 14368 1257
rect 14187 917 14253 933
rect 14187 883 14203 917
rect 14237 883 14253 917
rect 14187 867 14253 883
rect 14190 807 14250 867
rect 14308 807 14368 1255
rect 15372 1055 15432 1531
rect 14504 1010 15432 1055
rect 16072 1454 16132 1740
rect 16190 1714 16250 1740
rect 16308 1714 16368 1740
rect 16513 1714 16573 1740
rect 16072 1437 16208 1454
rect 16072 1382 16131 1437
rect 16189 1382 16208 1437
rect 16072 1367 16208 1382
rect 16072 1055 16132 1367
rect 16631 1322 16691 1740
rect 16749 1714 16809 1740
rect 16980 1714 17040 1740
rect 17098 1714 17158 1740
rect 17216 1714 17276 1740
rect 17334 1714 17394 1740
rect 17099 1554 17158 1714
rect 17099 1553 17162 1554
rect 17096 1537 17162 1553
rect 17096 1503 17112 1537
rect 17146 1503 17162 1537
rect 17096 1487 17162 1503
rect 17199 1438 17294 1453
rect 17199 1383 17218 1438
rect 17276 1415 17294 1438
rect 17452 1415 17512 1740
rect 17570 1714 17630 1740
rect 17807 1714 17867 1740
rect 17276 1383 17512 1415
rect 17199 1366 17512 1383
rect 16631 1265 17158 1322
rect 17098 1166 17158 1265
rect 17087 1153 17168 1166
rect 17087 1098 17100 1153
rect 17158 1098 17168 1153
rect 17087 1087 17168 1098
rect 16072 1010 16966 1055
rect 14504 807 14564 1010
rect 16906 807 16966 1010
rect 17098 807 17158 1087
rect 17216 807 17276 1366
rect 17925 1324 17985 1740
rect 18043 1714 18103 1740
rect 18280 1714 18340 1740
rect 18398 1714 18458 1740
rect 18406 1591 18472 1594
rect 18516 1591 18576 1740
rect 18406 1578 18576 1591
rect 18406 1544 18422 1578
rect 18456 1544 18576 1578
rect 18406 1531 18576 1544
rect 18406 1528 18472 1531
rect 17447 1307 17985 1324
rect 17447 1273 17466 1307
rect 17500 1273 17985 1307
rect 17447 1267 17985 1273
rect 17447 1257 17516 1267
rect 17447 1255 17512 1257
rect 17331 917 17397 933
rect 17331 883 17347 917
rect 17381 883 17397 917
rect 17331 867 17397 883
rect 17334 807 17394 867
rect 17452 807 17512 1255
rect 18516 1055 18576 1531
rect 17648 1010 18576 1055
rect 19204 1458 19264 1744
rect 19322 1718 19382 1744
rect 19440 1718 19500 1744
rect 19645 1718 19705 1744
rect 19204 1441 19340 1458
rect 19204 1386 19263 1441
rect 19321 1386 19340 1441
rect 19204 1371 19340 1386
rect 19204 1059 19264 1371
rect 19763 1326 19823 1744
rect 19881 1718 19941 1744
rect 20112 1718 20172 1744
rect 20230 1718 20290 1744
rect 20348 1718 20408 1744
rect 20466 1718 20526 1744
rect 20231 1558 20290 1718
rect 20231 1557 20294 1558
rect 20228 1541 20294 1557
rect 20228 1507 20244 1541
rect 20278 1507 20294 1541
rect 20228 1491 20294 1507
rect 20331 1442 20426 1457
rect 20331 1387 20350 1442
rect 20408 1419 20426 1442
rect 20584 1419 20644 1744
rect 20702 1718 20762 1744
rect 20939 1718 20999 1744
rect 20408 1387 20644 1419
rect 20331 1370 20644 1387
rect 19763 1269 20290 1326
rect 20230 1170 20290 1269
rect 20219 1157 20300 1170
rect 20219 1102 20232 1157
rect 20290 1102 20300 1157
rect 20219 1091 20300 1102
rect 19204 1014 20098 1059
rect 17648 807 17708 1010
rect 20038 811 20098 1014
rect 20230 811 20290 1091
rect 20348 811 20408 1370
rect 21057 1328 21117 1744
rect 21175 1718 21235 1744
rect 21412 1718 21472 1744
rect 21530 1718 21590 1744
rect 21538 1595 21604 1598
rect 21648 1595 21708 1744
rect 21538 1582 21708 1595
rect 21538 1548 21554 1582
rect 21588 1548 21708 1582
rect 21538 1535 21708 1548
rect 21538 1532 21604 1535
rect 20579 1311 21117 1328
rect 20579 1277 20598 1311
rect 20632 1277 21117 1311
rect 20579 1271 21117 1277
rect 20579 1261 20648 1271
rect 20579 1259 20644 1261
rect 20463 921 20529 937
rect 20463 887 20479 921
rect 20513 887 20529 921
rect 20463 871 20529 887
rect 20466 811 20526 871
rect 20584 811 20644 1259
rect 21648 1059 21708 1535
rect 20780 1014 21708 1059
rect 22348 1458 22408 1744
rect 22466 1718 22526 1744
rect 22584 1718 22644 1744
rect 22789 1718 22849 1744
rect 22348 1441 22484 1458
rect 22348 1386 22407 1441
rect 22465 1386 22484 1441
rect 22348 1371 22484 1386
rect 22348 1059 22408 1371
rect 22907 1326 22967 1744
rect 23025 1718 23085 1744
rect 23256 1718 23316 1744
rect 23374 1718 23434 1744
rect 23492 1718 23552 1744
rect 23610 1718 23670 1744
rect 23375 1558 23434 1718
rect 23375 1557 23438 1558
rect 23372 1541 23438 1557
rect 23372 1507 23388 1541
rect 23422 1507 23438 1541
rect 23372 1491 23438 1507
rect 23475 1442 23570 1457
rect 23475 1387 23494 1442
rect 23552 1419 23570 1442
rect 23728 1419 23788 1744
rect 23846 1718 23906 1744
rect 24083 1718 24143 1744
rect 23552 1387 23788 1419
rect 23475 1370 23788 1387
rect 22907 1269 23434 1326
rect 23374 1170 23434 1269
rect 23363 1157 23444 1170
rect 23363 1102 23376 1157
rect 23434 1102 23444 1157
rect 23363 1091 23444 1102
rect 22348 1014 23242 1059
rect 20780 811 20840 1014
rect 23182 811 23242 1014
rect 23374 811 23434 1091
rect 23492 811 23552 1370
rect 24201 1328 24261 1744
rect 24319 1718 24379 1744
rect 24556 1718 24616 1744
rect 24674 1718 24734 1744
rect 24682 1595 24748 1598
rect 24792 1595 24852 1744
rect 24682 1582 24852 1595
rect 24682 1548 24698 1582
rect 24732 1548 24852 1582
rect 24682 1535 24852 1548
rect 24682 1532 24748 1535
rect 23723 1311 24261 1328
rect 23723 1277 23742 1311
rect 23776 1277 24261 1311
rect 23723 1271 24261 1277
rect 23723 1261 23792 1271
rect 23723 1259 23788 1261
rect 23607 921 23673 937
rect 23607 887 23623 921
rect 23657 887 23673 921
rect 23607 871 23673 887
rect 23610 811 23670 871
rect 23728 811 23788 1259
rect 24792 1059 24852 1535
rect 23924 1014 24852 1059
rect 23924 811 23984 1014
rect 10752 385 10812 411
rect 10870 385 10930 411
rect 10988 385 11048 411
rect 11106 385 11166 411
rect 7783 322 8218 330
rect 7783 288 7799 322
rect 7833 288 8218 322
rect 7783 279 8218 288
rect 10927 330 10993 338
rect 11302 330 11362 611
rect 13762 581 13822 607
rect 13954 381 14014 407
rect 14072 381 14132 407
rect 14190 381 14250 407
rect 14308 381 14368 407
rect 10927 322 11362 330
rect 10927 288 10943 322
rect 10977 288 11362 322
rect 10927 279 11362 288
rect 14129 326 14195 334
rect 14504 326 14564 607
rect 16906 581 16966 607
rect 17098 381 17158 407
rect 17216 381 17276 407
rect 17334 381 17394 407
rect 17452 381 17512 407
rect 14129 318 14564 326
rect 14129 284 14145 318
rect 14179 284 14564 318
rect 1507 268 1573 275
rect 4651 268 4717 275
rect 7783 272 7849 279
rect 10927 272 10993 279
rect 14129 275 14564 284
rect 17273 326 17339 334
rect 17648 326 17708 607
rect 20038 585 20098 611
rect 20230 385 20290 411
rect 20348 385 20408 411
rect 20466 385 20526 411
rect 20584 385 20644 411
rect 17273 318 17708 326
rect 17273 284 17289 318
rect 17323 284 17708 318
rect 17273 275 17708 284
rect 20405 330 20471 338
rect 20780 330 20840 611
rect 23182 585 23242 611
rect 23374 385 23434 411
rect 23492 385 23552 411
rect 23610 385 23670 411
rect 23728 385 23788 411
rect 20405 322 20840 330
rect 20405 288 20421 322
rect 20455 288 20840 322
rect 20405 279 20840 288
rect 23549 330 23615 338
rect 23924 330 23984 611
rect 23549 322 23984 330
rect 23549 288 23565 322
rect 23599 288 23984 322
rect 23549 279 23984 288
rect 14129 268 14195 275
rect 17273 268 17339 275
rect 20405 272 20471 279
rect 23549 272 23615 279
rect 779 -1737 1075 -1698
rect 779 -1752 839 -1737
rect 897 -1752 957 -1737
rect 1015 -1752 1075 -1737
rect 1246 -1737 1542 -1698
rect 1246 -1752 1306 -1737
rect 1364 -1752 1424 -1737
rect 1482 -1752 1542 -1737
rect 1600 -1737 1896 -1698
rect 1600 -1752 1660 -1737
rect 1718 -1752 1778 -1737
rect 1836 -1752 1896 -1737
rect 2073 -1737 2369 -1698
rect 2073 -1752 2133 -1737
rect 2191 -1752 2251 -1737
rect 2309 -1752 2369 -1737
rect 3923 -1737 4219 -1698
rect 3923 -1752 3983 -1737
rect 4041 -1752 4101 -1737
rect 4159 -1752 4219 -1737
rect 4390 -1737 4686 -1698
rect 4390 -1752 4450 -1737
rect 4508 -1752 4568 -1737
rect 4626 -1752 4686 -1737
rect 4744 -1737 5040 -1698
rect 4744 -1752 4804 -1737
rect 4862 -1752 4922 -1737
rect 4980 -1752 5040 -1737
rect 5217 -1737 5513 -1698
rect 5217 -1752 5277 -1737
rect 5335 -1752 5395 -1737
rect 5453 -1752 5513 -1737
rect 7055 -1733 7351 -1694
rect 7055 -1748 7115 -1733
rect 7173 -1748 7233 -1733
rect 7291 -1748 7351 -1733
rect 7522 -1733 7818 -1694
rect 7522 -1748 7582 -1733
rect 7640 -1748 7700 -1733
rect 7758 -1748 7818 -1733
rect 7876 -1733 8172 -1694
rect 7876 -1748 7936 -1733
rect 7994 -1748 8054 -1733
rect 8112 -1748 8172 -1733
rect 8349 -1733 8645 -1694
rect 8349 -1748 8409 -1733
rect 8467 -1748 8527 -1733
rect 8585 -1748 8645 -1733
rect 10199 -1733 10495 -1694
rect 10199 -1748 10259 -1733
rect 10317 -1748 10377 -1733
rect 10435 -1748 10495 -1733
rect 10666 -1733 10962 -1694
rect 10666 -1748 10726 -1733
rect 10784 -1748 10844 -1733
rect 10902 -1748 10962 -1733
rect 11020 -1733 11316 -1694
rect 11020 -1748 11080 -1733
rect 11138 -1748 11198 -1733
rect 11256 -1748 11316 -1733
rect 11493 -1733 11789 -1694
rect 11493 -1748 11553 -1733
rect 11611 -1748 11671 -1733
rect 11729 -1748 11789 -1733
rect 13401 -1737 13697 -1698
rect 338 -1936 634 -1897
rect 338 -1952 398 -1936
rect 456 -1952 516 -1936
rect 574 -1952 634 -1936
rect 2546 -1936 2842 -1897
rect 2546 -1952 2606 -1936
rect 2664 -1952 2724 -1936
rect 2782 -1952 2842 -1936
rect 3482 -1936 3778 -1897
rect 3482 -1952 3542 -1936
rect 3600 -1952 3660 -1936
rect 3718 -1952 3778 -1936
rect 5690 -1936 5986 -1897
rect 5690 -1952 5750 -1936
rect 5808 -1952 5868 -1936
rect 5926 -1952 5986 -1936
rect 6614 -1932 6910 -1893
rect 6614 -1948 6674 -1932
rect 6732 -1948 6792 -1932
rect 6850 -1948 6910 -1932
rect 8822 -1932 9118 -1893
rect 8822 -1948 8882 -1932
rect 8940 -1948 9000 -1932
rect 9058 -1948 9118 -1932
rect 9758 -1932 10054 -1893
rect 9758 -1948 9818 -1932
rect 9876 -1948 9936 -1932
rect 9994 -1948 10054 -1932
rect 13401 -1752 13461 -1737
rect 13519 -1752 13579 -1737
rect 13637 -1752 13697 -1737
rect 13868 -1737 14164 -1698
rect 13868 -1752 13928 -1737
rect 13986 -1752 14046 -1737
rect 14104 -1752 14164 -1737
rect 14222 -1737 14518 -1698
rect 14222 -1752 14282 -1737
rect 14340 -1752 14400 -1737
rect 14458 -1752 14518 -1737
rect 14695 -1737 14991 -1698
rect 14695 -1752 14755 -1737
rect 14813 -1752 14873 -1737
rect 14931 -1752 14991 -1737
rect 16545 -1737 16841 -1698
rect 16545 -1752 16605 -1737
rect 16663 -1752 16723 -1737
rect 16781 -1752 16841 -1737
rect 17012 -1737 17308 -1698
rect 17012 -1752 17072 -1737
rect 17130 -1752 17190 -1737
rect 17248 -1752 17308 -1737
rect 17366 -1737 17662 -1698
rect 17366 -1752 17426 -1737
rect 17484 -1752 17544 -1737
rect 17602 -1752 17662 -1737
rect 17839 -1737 18135 -1698
rect 17839 -1752 17899 -1737
rect 17957 -1752 18017 -1737
rect 18075 -1752 18135 -1737
rect 19677 -1733 19973 -1694
rect 19677 -1748 19737 -1733
rect 19795 -1748 19855 -1733
rect 19913 -1748 19973 -1733
rect 20144 -1733 20440 -1694
rect 20144 -1748 20204 -1733
rect 20262 -1748 20322 -1733
rect 20380 -1748 20440 -1733
rect 20498 -1733 20794 -1694
rect 20498 -1748 20558 -1733
rect 20616 -1748 20676 -1733
rect 20734 -1748 20794 -1733
rect 20971 -1733 21267 -1694
rect 20971 -1748 21031 -1733
rect 21089 -1748 21149 -1733
rect 21207 -1748 21267 -1733
rect 22821 -1733 23117 -1694
rect 22821 -1748 22881 -1733
rect 22939 -1748 22999 -1733
rect 23057 -1748 23117 -1733
rect 23288 -1733 23584 -1694
rect 23288 -1748 23348 -1733
rect 23406 -1748 23466 -1733
rect 23524 -1748 23584 -1733
rect 23642 -1733 23938 -1694
rect 23642 -1748 23702 -1733
rect 23760 -1748 23820 -1733
rect 23878 -1748 23938 -1733
rect 24115 -1733 24411 -1694
rect 24115 -1748 24175 -1733
rect 24233 -1748 24293 -1733
rect 24351 -1748 24411 -1733
rect 11966 -1932 12262 -1893
rect 11966 -1948 12026 -1932
rect 12084 -1948 12144 -1932
rect 12202 -1948 12262 -1932
rect 12960 -1936 13256 -1897
rect 12960 -1952 13020 -1936
rect 13078 -1952 13138 -1936
rect 13196 -1952 13256 -1936
rect 338 -2438 398 -2152
rect 456 -2178 516 -2152
rect 574 -2178 634 -2152
rect 779 -2178 839 -2152
rect 338 -2455 474 -2438
rect 338 -2510 397 -2455
rect 455 -2510 474 -2455
rect 338 -2525 474 -2510
rect 338 -2837 398 -2525
rect 897 -2570 957 -2152
rect 1015 -2178 1075 -2152
rect 1246 -2178 1306 -2152
rect 1364 -2178 1424 -2152
rect 1482 -2178 1542 -2152
rect 1600 -2178 1660 -2152
rect 1365 -2338 1424 -2178
rect 1365 -2339 1428 -2338
rect 1362 -2355 1428 -2339
rect 1362 -2389 1378 -2355
rect 1412 -2389 1428 -2355
rect 1362 -2405 1428 -2389
rect 1465 -2454 1560 -2439
rect 1465 -2509 1484 -2454
rect 1542 -2477 1560 -2454
rect 1718 -2477 1778 -2152
rect 1836 -2178 1896 -2152
rect 2073 -2178 2133 -2152
rect 1542 -2509 1778 -2477
rect 1465 -2526 1778 -2509
rect 897 -2627 1424 -2570
rect 1364 -2726 1424 -2627
rect 1353 -2739 1434 -2726
rect 1353 -2794 1366 -2739
rect 1424 -2794 1434 -2739
rect 1353 -2805 1434 -2794
rect 338 -2882 1232 -2837
rect 1172 -3085 1232 -2882
rect 1364 -3085 1424 -2805
rect 1482 -3085 1542 -2526
rect 2191 -2568 2251 -2152
rect 2309 -2178 2369 -2152
rect 2546 -2178 2606 -2152
rect 2664 -2178 2724 -2152
rect 2672 -2301 2738 -2298
rect 2782 -2301 2842 -2152
rect 2672 -2314 2842 -2301
rect 2672 -2348 2688 -2314
rect 2722 -2348 2842 -2314
rect 2672 -2361 2842 -2348
rect 2672 -2364 2738 -2361
rect 1713 -2585 2251 -2568
rect 1713 -2619 1732 -2585
rect 1766 -2619 2251 -2585
rect 1713 -2625 2251 -2619
rect 1713 -2635 1782 -2625
rect 1713 -2637 1778 -2635
rect 1597 -2975 1663 -2959
rect 1597 -3009 1613 -2975
rect 1647 -3009 1663 -2975
rect 1597 -3025 1663 -3009
rect 1600 -3085 1660 -3025
rect 1718 -3085 1778 -2637
rect 2782 -2837 2842 -2361
rect 1914 -2882 2842 -2837
rect 3482 -2438 3542 -2152
rect 3600 -2178 3660 -2152
rect 3718 -2178 3778 -2152
rect 3923 -2178 3983 -2152
rect 3482 -2455 3618 -2438
rect 3482 -2510 3541 -2455
rect 3599 -2510 3618 -2455
rect 3482 -2525 3618 -2510
rect 3482 -2837 3542 -2525
rect 4041 -2570 4101 -2152
rect 4159 -2178 4219 -2152
rect 4390 -2178 4450 -2152
rect 4508 -2178 4568 -2152
rect 4626 -2178 4686 -2152
rect 4744 -2178 4804 -2152
rect 4509 -2338 4568 -2178
rect 4509 -2339 4572 -2338
rect 4506 -2355 4572 -2339
rect 4506 -2389 4522 -2355
rect 4556 -2389 4572 -2355
rect 4506 -2405 4572 -2389
rect 4609 -2454 4704 -2439
rect 4609 -2509 4628 -2454
rect 4686 -2477 4704 -2454
rect 4862 -2477 4922 -2152
rect 4980 -2178 5040 -2152
rect 5217 -2178 5277 -2152
rect 4686 -2509 4922 -2477
rect 4609 -2526 4922 -2509
rect 4041 -2627 4568 -2570
rect 4508 -2726 4568 -2627
rect 4497 -2739 4578 -2726
rect 4497 -2794 4510 -2739
rect 4568 -2794 4578 -2739
rect 4497 -2805 4578 -2794
rect 3482 -2882 4376 -2837
rect 1914 -3085 1974 -2882
rect 4316 -3085 4376 -2882
rect 4508 -3085 4568 -2805
rect 4626 -3085 4686 -2526
rect 5335 -2568 5395 -2152
rect 5453 -2178 5513 -2152
rect 5690 -2178 5750 -2152
rect 5808 -2178 5868 -2152
rect 5816 -2301 5882 -2298
rect 5926 -2301 5986 -2152
rect 5816 -2314 5986 -2301
rect 5816 -2348 5832 -2314
rect 5866 -2348 5986 -2314
rect 5816 -2361 5986 -2348
rect 5816 -2364 5882 -2361
rect 4857 -2585 5395 -2568
rect 4857 -2619 4876 -2585
rect 4910 -2619 5395 -2585
rect 4857 -2625 5395 -2619
rect 4857 -2635 4926 -2625
rect 4857 -2637 4922 -2635
rect 4741 -2975 4807 -2959
rect 4741 -3009 4757 -2975
rect 4791 -3009 4807 -2975
rect 4741 -3025 4807 -3009
rect 4744 -3085 4804 -3025
rect 4862 -3085 4922 -2637
rect 5926 -2837 5986 -2361
rect 5058 -2882 5986 -2837
rect 6614 -2434 6674 -2148
rect 6732 -2174 6792 -2148
rect 6850 -2174 6910 -2148
rect 7055 -2174 7115 -2148
rect 6614 -2451 6750 -2434
rect 6614 -2506 6673 -2451
rect 6731 -2506 6750 -2451
rect 6614 -2521 6750 -2506
rect 6614 -2833 6674 -2521
rect 7173 -2566 7233 -2148
rect 7291 -2174 7351 -2148
rect 7522 -2174 7582 -2148
rect 7640 -2174 7700 -2148
rect 7758 -2174 7818 -2148
rect 7876 -2174 7936 -2148
rect 7641 -2334 7700 -2174
rect 7641 -2335 7704 -2334
rect 7638 -2351 7704 -2335
rect 7638 -2385 7654 -2351
rect 7688 -2385 7704 -2351
rect 7638 -2401 7704 -2385
rect 7741 -2450 7836 -2435
rect 7741 -2505 7760 -2450
rect 7818 -2473 7836 -2450
rect 7994 -2473 8054 -2148
rect 8112 -2174 8172 -2148
rect 8349 -2174 8409 -2148
rect 7818 -2505 8054 -2473
rect 7741 -2522 8054 -2505
rect 7173 -2623 7700 -2566
rect 7640 -2722 7700 -2623
rect 7629 -2735 7710 -2722
rect 7629 -2790 7642 -2735
rect 7700 -2790 7710 -2735
rect 7629 -2801 7710 -2790
rect 6614 -2878 7508 -2833
rect 5058 -3085 5118 -2882
rect 7448 -3081 7508 -2878
rect 7640 -3081 7700 -2801
rect 7758 -3081 7818 -2522
rect 8467 -2564 8527 -2148
rect 8585 -2174 8645 -2148
rect 8822 -2174 8882 -2148
rect 8940 -2174 9000 -2148
rect 8948 -2297 9014 -2294
rect 9058 -2297 9118 -2148
rect 8948 -2310 9118 -2297
rect 8948 -2344 8964 -2310
rect 8998 -2344 9118 -2310
rect 8948 -2357 9118 -2344
rect 8948 -2360 9014 -2357
rect 7989 -2581 8527 -2564
rect 7989 -2615 8008 -2581
rect 8042 -2615 8527 -2581
rect 7989 -2621 8527 -2615
rect 7989 -2631 8058 -2621
rect 7989 -2633 8054 -2631
rect 7873 -2971 7939 -2955
rect 7873 -3005 7889 -2971
rect 7923 -3005 7939 -2971
rect 7873 -3021 7939 -3005
rect 7876 -3081 7936 -3021
rect 7994 -3081 8054 -2633
rect 9058 -2833 9118 -2357
rect 8190 -2878 9118 -2833
rect 9758 -2434 9818 -2148
rect 9876 -2174 9936 -2148
rect 9994 -2174 10054 -2148
rect 10199 -2174 10259 -2148
rect 9758 -2451 9894 -2434
rect 9758 -2506 9817 -2451
rect 9875 -2506 9894 -2451
rect 9758 -2521 9894 -2506
rect 9758 -2833 9818 -2521
rect 10317 -2566 10377 -2148
rect 10435 -2174 10495 -2148
rect 10666 -2174 10726 -2148
rect 10784 -2174 10844 -2148
rect 10902 -2174 10962 -2148
rect 11020 -2174 11080 -2148
rect 10785 -2334 10844 -2174
rect 10785 -2335 10848 -2334
rect 10782 -2351 10848 -2335
rect 10782 -2385 10798 -2351
rect 10832 -2385 10848 -2351
rect 10782 -2401 10848 -2385
rect 10885 -2450 10980 -2435
rect 10885 -2505 10904 -2450
rect 10962 -2473 10980 -2450
rect 11138 -2473 11198 -2148
rect 11256 -2174 11316 -2148
rect 11493 -2174 11553 -2148
rect 10962 -2505 11198 -2473
rect 10885 -2522 11198 -2505
rect 10317 -2623 10844 -2566
rect 10784 -2722 10844 -2623
rect 10773 -2735 10854 -2722
rect 10773 -2790 10786 -2735
rect 10844 -2790 10854 -2735
rect 10773 -2801 10854 -2790
rect 9758 -2878 10652 -2833
rect 8190 -3081 8250 -2878
rect 10592 -3081 10652 -2878
rect 10784 -3081 10844 -2801
rect 10902 -3081 10962 -2522
rect 11611 -2564 11671 -2148
rect 11729 -2174 11789 -2148
rect 11966 -2174 12026 -2148
rect 12084 -2174 12144 -2148
rect 12092 -2297 12158 -2294
rect 12202 -2297 12262 -2148
rect 15168 -1936 15464 -1897
rect 15168 -1952 15228 -1936
rect 15286 -1952 15346 -1936
rect 15404 -1952 15464 -1936
rect 16104 -1936 16400 -1897
rect 16104 -1952 16164 -1936
rect 16222 -1952 16282 -1936
rect 16340 -1952 16400 -1936
rect 18312 -1936 18608 -1897
rect 18312 -1952 18372 -1936
rect 18430 -1952 18490 -1936
rect 18548 -1952 18608 -1936
rect 19236 -1932 19532 -1893
rect 19236 -1948 19296 -1932
rect 19354 -1948 19414 -1932
rect 19472 -1948 19532 -1932
rect 21444 -1932 21740 -1893
rect 21444 -1948 21504 -1932
rect 21562 -1948 21622 -1932
rect 21680 -1948 21740 -1932
rect 22380 -1932 22676 -1893
rect 22380 -1948 22440 -1932
rect 22498 -1948 22558 -1932
rect 22616 -1948 22676 -1932
rect 24588 -1932 24884 -1893
rect 24588 -1948 24648 -1932
rect 24706 -1948 24766 -1932
rect 24824 -1948 24884 -1932
rect 12092 -2310 12262 -2297
rect 12092 -2344 12108 -2310
rect 12142 -2344 12262 -2310
rect 12092 -2357 12262 -2344
rect 12092 -2360 12158 -2357
rect 11133 -2581 11671 -2564
rect 11133 -2615 11152 -2581
rect 11186 -2615 11671 -2581
rect 11133 -2621 11671 -2615
rect 11133 -2631 11202 -2621
rect 11133 -2633 11198 -2631
rect 11017 -2971 11083 -2955
rect 11017 -3005 11033 -2971
rect 11067 -3005 11083 -2971
rect 11017 -3021 11083 -3005
rect 11020 -3081 11080 -3021
rect 11138 -3081 11198 -2633
rect 12202 -2833 12262 -2357
rect 11334 -2878 12262 -2833
rect 12960 -2438 13020 -2152
rect 13078 -2178 13138 -2152
rect 13196 -2178 13256 -2152
rect 13401 -2178 13461 -2152
rect 12960 -2455 13096 -2438
rect 12960 -2510 13019 -2455
rect 13077 -2510 13096 -2455
rect 12960 -2525 13096 -2510
rect 12960 -2837 13020 -2525
rect 13519 -2570 13579 -2152
rect 13637 -2178 13697 -2152
rect 13868 -2178 13928 -2152
rect 13986 -2178 14046 -2152
rect 14104 -2178 14164 -2152
rect 14222 -2178 14282 -2152
rect 13987 -2338 14046 -2178
rect 13987 -2339 14050 -2338
rect 13984 -2355 14050 -2339
rect 13984 -2389 14000 -2355
rect 14034 -2389 14050 -2355
rect 13984 -2405 14050 -2389
rect 14087 -2454 14182 -2439
rect 14087 -2509 14106 -2454
rect 14164 -2477 14182 -2454
rect 14340 -2477 14400 -2152
rect 14458 -2178 14518 -2152
rect 14695 -2178 14755 -2152
rect 14164 -2509 14400 -2477
rect 14087 -2526 14400 -2509
rect 13519 -2627 14046 -2570
rect 13986 -2726 14046 -2627
rect 13975 -2739 14056 -2726
rect 13975 -2794 13988 -2739
rect 14046 -2794 14056 -2739
rect 13975 -2805 14056 -2794
rect 11334 -3081 11394 -2878
rect 12960 -2882 13854 -2837
rect 1172 -3311 1232 -3285
rect 1364 -3511 1424 -3485
rect 1482 -3511 1542 -3485
rect 1600 -3511 1660 -3485
rect 1718 -3511 1778 -3485
rect 1539 -3566 1605 -3558
rect 1914 -3566 1974 -3285
rect 4316 -3311 4376 -3285
rect 4508 -3511 4568 -3485
rect 4626 -3511 4686 -3485
rect 4744 -3511 4804 -3485
rect 4862 -3511 4922 -3485
rect 1539 -3574 1974 -3566
rect 1539 -3608 1555 -3574
rect 1589 -3608 1974 -3574
rect 1539 -3617 1974 -3608
rect 4683 -3566 4749 -3558
rect 5058 -3566 5118 -3285
rect 7448 -3307 7508 -3281
rect 7640 -3507 7700 -3481
rect 7758 -3507 7818 -3481
rect 7876 -3507 7936 -3481
rect 7994 -3507 8054 -3481
rect 4683 -3574 5118 -3566
rect 4683 -3608 4699 -3574
rect 4733 -3608 5118 -3574
rect 4683 -3617 5118 -3608
rect 7815 -3562 7881 -3554
rect 8190 -3562 8250 -3281
rect 10592 -3307 10652 -3281
rect 13794 -3085 13854 -2882
rect 13986 -3085 14046 -2805
rect 14104 -3085 14164 -2526
rect 14813 -2568 14873 -2152
rect 14931 -2178 14991 -2152
rect 15168 -2178 15228 -2152
rect 15286 -2178 15346 -2152
rect 15294 -2301 15360 -2298
rect 15404 -2301 15464 -2152
rect 15294 -2314 15464 -2301
rect 15294 -2348 15310 -2314
rect 15344 -2348 15464 -2314
rect 15294 -2361 15464 -2348
rect 15294 -2364 15360 -2361
rect 14335 -2585 14873 -2568
rect 14335 -2619 14354 -2585
rect 14388 -2619 14873 -2585
rect 14335 -2625 14873 -2619
rect 14335 -2635 14404 -2625
rect 14335 -2637 14400 -2635
rect 14219 -2975 14285 -2959
rect 14219 -3009 14235 -2975
rect 14269 -3009 14285 -2975
rect 14219 -3025 14285 -3009
rect 14222 -3085 14282 -3025
rect 14340 -3085 14400 -2637
rect 15404 -2837 15464 -2361
rect 14536 -2882 15464 -2837
rect 16104 -2438 16164 -2152
rect 16222 -2178 16282 -2152
rect 16340 -2178 16400 -2152
rect 16545 -2178 16605 -2152
rect 16104 -2455 16240 -2438
rect 16104 -2510 16163 -2455
rect 16221 -2510 16240 -2455
rect 16104 -2525 16240 -2510
rect 16104 -2837 16164 -2525
rect 16663 -2570 16723 -2152
rect 16781 -2178 16841 -2152
rect 17012 -2178 17072 -2152
rect 17130 -2178 17190 -2152
rect 17248 -2178 17308 -2152
rect 17366 -2178 17426 -2152
rect 17131 -2338 17190 -2178
rect 17131 -2339 17194 -2338
rect 17128 -2355 17194 -2339
rect 17128 -2389 17144 -2355
rect 17178 -2389 17194 -2355
rect 17128 -2405 17194 -2389
rect 17231 -2454 17326 -2439
rect 17231 -2509 17250 -2454
rect 17308 -2477 17326 -2454
rect 17484 -2477 17544 -2152
rect 17602 -2178 17662 -2152
rect 17839 -2178 17899 -2152
rect 17308 -2509 17544 -2477
rect 17231 -2526 17544 -2509
rect 16663 -2627 17190 -2570
rect 17130 -2726 17190 -2627
rect 17119 -2739 17200 -2726
rect 17119 -2794 17132 -2739
rect 17190 -2794 17200 -2739
rect 17119 -2805 17200 -2794
rect 16104 -2882 16998 -2837
rect 14536 -3085 14596 -2882
rect 16938 -3085 16998 -2882
rect 17130 -3085 17190 -2805
rect 17248 -3085 17308 -2526
rect 17957 -2568 18017 -2152
rect 18075 -2178 18135 -2152
rect 18312 -2178 18372 -2152
rect 18430 -2178 18490 -2152
rect 18438 -2301 18504 -2298
rect 18548 -2301 18608 -2152
rect 18438 -2314 18608 -2301
rect 18438 -2348 18454 -2314
rect 18488 -2348 18608 -2314
rect 18438 -2361 18608 -2348
rect 18438 -2364 18504 -2361
rect 17479 -2585 18017 -2568
rect 17479 -2619 17498 -2585
rect 17532 -2619 18017 -2585
rect 17479 -2625 18017 -2619
rect 17479 -2635 17548 -2625
rect 17479 -2637 17544 -2635
rect 17363 -2975 17429 -2959
rect 17363 -3009 17379 -2975
rect 17413 -3009 17429 -2975
rect 17363 -3025 17429 -3009
rect 17366 -3085 17426 -3025
rect 17484 -3085 17544 -2637
rect 18548 -2837 18608 -2361
rect 17680 -2882 18608 -2837
rect 19236 -2434 19296 -2148
rect 19354 -2174 19414 -2148
rect 19472 -2174 19532 -2148
rect 19677 -2174 19737 -2148
rect 19236 -2451 19372 -2434
rect 19236 -2506 19295 -2451
rect 19353 -2506 19372 -2451
rect 19236 -2521 19372 -2506
rect 19236 -2833 19296 -2521
rect 19795 -2566 19855 -2148
rect 19913 -2174 19973 -2148
rect 20144 -2174 20204 -2148
rect 20262 -2174 20322 -2148
rect 20380 -2174 20440 -2148
rect 20498 -2174 20558 -2148
rect 20263 -2334 20322 -2174
rect 20263 -2335 20326 -2334
rect 20260 -2351 20326 -2335
rect 20260 -2385 20276 -2351
rect 20310 -2385 20326 -2351
rect 20260 -2401 20326 -2385
rect 20363 -2450 20458 -2435
rect 20363 -2505 20382 -2450
rect 20440 -2473 20458 -2450
rect 20616 -2473 20676 -2148
rect 20734 -2174 20794 -2148
rect 20971 -2174 21031 -2148
rect 20440 -2505 20676 -2473
rect 20363 -2522 20676 -2505
rect 19795 -2623 20322 -2566
rect 20262 -2722 20322 -2623
rect 20251 -2735 20332 -2722
rect 20251 -2790 20264 -2735
rect 20322 -2790 20332 -2735
rect 20251 -2801 20332 -2790
rect 19236 -2878 20130 -2833
rect 17680 -3085 17740 -2882
rect 20070 -3081 20130 -2878
rect 20262 -3081 20322 -2801
rect 20380 -3081 20440 -2522
rect 21089 -2564 21149 -2148
rect 21207 -2174 21267 -2148
rect 21444 -2174 21504 -2148
rect 21562 -2174 21622 -2148
rect 21570 -2297 21636 -2294
rect 21680 -2297 21740 -2148
rect 21570 -2310 21740 -2297
rect 21570 -2344 21586 -2310
rect 21620 -2344 21740 -2310
rect 21570 -2357 21740 -2344
rect 21570 -2360 21636 -2357
rect 20611 -2581 21149 -2564
rect 20611 -2615 20630 -2581
rect 20664 -2615 21149 -2581
rect 20611 -2621 21149 -2615
rect 20611 -2631 20680 -2621
rect 20611 -2633 20676 -2631
rect 20495 -2971 20561 -2955
rect 20495 -3005 20511 -2971
rect 20545 -3005 20561 -2971
rect 20495 -3021 20561 -3005
rect 20498 -3081 20558 -3021
rect 20616 -3081 20676 -2633
rect 21680 -2833 21740 -2357
rect 20812 -2878 21740 -2833
rect 22380 -2434 22440 -2148
rect 22498 -2174 22558 -2148
rect 22616 -2174 22676 -2148
rect 22821 -2174 22881 -2148
rect 22380 -2451 22516 -2434
rect 22380 -2506 22439 -2451
rect 22497 -2506 22516 -2451
rect 22380 -2521 22516 -2506
rect 22380 -2833 22440 -2521
rect 22939 -2566 22999 -2148
rect 23057 -2174 23117 -2148
rect 23288 -2174 23348 -2148
rect 23406 -2174 23466 -2148
rect 23524 -2174 23584 -2148
rect 23642 -2174 23702 -2148
rect 23407 -2334 23466 -2174
rect 23407 -2335 23470 -2334
rect 23404 -2351 23470 -2335
rect 23404 -2385 23420 -2351
rect 23454 -2385 23470 -2351
rect 23404 -2401 23470 -2385
rect 23507 -2450 23602 -2435
rect 23507 -2505 23526 -2450
rect 23584 -2473 23602 -2450
rect 23760 -2473 23820 -2148
rect 23878 -2174 23938 -2148
rect 24115 -2174 24175 -2148
rect 23584 -2505 23820 -2473
rect 23507 -2522 23820 -2505
rect 22939 -2623 23466 -2566
rect 23406 -2722 23466 -2623
rect 23395 -2735 23476 -2722
rect 23395 -2790 23408 -2735
rect 23466 -2790 23476 -2735
rect 23395 -2801 23476 -2790
rect 22380 -2878 23274 -2833
rect 20812 -3081 20872 -2878
rect 23214 -3081 23274 -2878
rect 23406 -3081 23466 -2801
rect 23524 -3081 23584 -2522
rect 24233 -2564 24293 -2148
rect 24351 -2174 24411 -2148
rect 24588 -2174 24648 -2148
rect 24706 -2174 24766 -2148
rect 24714 -2297 24780 -2294
rect 24824 -2297 24884 -2148
rect 24714 -2310 24884 -2297
rect 24714 -2344 24730 -2310
rect 24764 -2344 24884 -2310
rect 24714 -2357 24884 -2344
rect 24714 -2360 24780 -2357
rect 23755 -2581 24293 -2564
rect 23755 -2615 23774 -2581
rect 23808 -2615 24293 -2581
rect 23755 -2621 24293 -2615
rect 23755 -2631 23824 -2621
rect 23755 -2633 23820 -2631
rect 23639 -2971 23705 -2955
rect 23639 -3005 23655 -2971
rect 23689 -3005 23705 -2971
rect 23639 -3021 23705 -3005
rect 23642 -3081 23702 -3021
rect 23760 -3081 23820 -2633
rect 24824 -2833 24884 -2357
rect 23956 -2878 24884 -2833
rect 23956 -3081 24016 -2878
rect 10784 -3507 10844 -3481
rect 10902 -3507 10962 -3481
rect 11020 -3507 11080 -3481
rect 11138 -3507 11198 -3481
rect 7815 -3570 8250 -3562
rect 7815 -3604 7831 -3570
rect 7865 -3604 8250 -3570
rect 7815 -3613 8250 -3604
rect 10959 -3562 11025 -3554
rect 11334 -3562 11394 -3281
rect 13794 -3311 13854 -3285
rect 13986 -3511 14046 -3485
rect 14104 -3511 14164 -3485
rect 14222 -3511 14282 -3485
rect 14340 -3511 14400 -3485
rect 10959 -3570 11394 -3562
rect 10959 -3604 10975 -3570
rect 11009 -3604 11394 -3570
rect 10959 -3613 11394 -3604
rect 14161 -3566 14227 -3558
rect 14536 -3566 14596 -3285
rect 16938 -3311 16998 -3285
rect 17130 -3511 17190 -3485
rect 17248 -3511 17308 -3485
rect 17366 -3511 17426 -3485
rect 17484 -3511 17544 -3485
rect 14161 -3574 14596 -3566
rect 14161 -3608 14177 -3574
rect 14211 -3608 14596 -3574
rect 1539 -3624 1605 -3617
rect 4683 -3624 4749 -3617
rect 7815 -3620 7881 -3613
rect 10959 -3620 11025 -3613
rect 14161 -3617 14596 -3608
rect 17305 -3566 17371 -3558
rect 17680 -3566 17740 -3285
rect 20070 -3307 20130 -3281
rect 20262 -3507 20322 -3481
rect 20380 -3507 20440 -3481
rect 20498 -3507 20558 -3481
rect 20616 -3507 20676 -3481
rect 17305 -3574 17740 -3566
rect 17305 -3608 17321 -3574
rect 17355 -3608 17740 -3574
rect 17305 -3617 17740 -3608
rect 20437 -3562 20503 -3554
rect 20812 -3562 20872 -3281
rect 23214 -3307 23274 -3281
rect 23406 -3507 23466 -3481
rect 23524 -3507 23584 -3481
rect 23642 -3507 23702 -3481
rect 23760 -3507 23820 -3481
rect 20437 -3570 20872 -3562
rect 20437 -3604 20453 -3570
rect 20487 -3604 20872 -3570
rect 20437 -3613 20872 -3604
rect 23581 -3562 23647 -3554
rect 23956 -3562 24016 -3281
rect 23581 -3570 24016 -3562
rect 23581 -3604 23597 -3570
rect 23631 -3604 24016 -3570
rect 23581 -3613 24016 -3604
rect 14161 -3624 14227 -3617
rect 17305 -3624 17371 -3617
rect 20437 -3620 20503 -3613
rect 23581 -3620 23647 -3613
<< polycont >>
rect 571 21234 629 21289
rect 1552 21355 1586 21389
rect 1658 21235 1716 21290
rect 1540 20950 1598 21005
rect 2862 21396 2896 21430
rect 1906 21125 1940 21159
rect 1787 20735 1821 20769
rect 3715 21234 3773 21289
rect 4696 21355 4730 21389
rect 4802 21235 4860 21290
rect 4684 20950 4742 21005
rect 6006 21396 6040 21430
rect 5050 21125 5084 21159
rect 4931 20735 4965 20769
rect 6847 21238 6905 21293
rect 7828 21359 7862 21393
rect 7934 21239 7992 21294
rect 7816 20954 7874 21009
rect 9138 21400 9172 21434
rect 8182 21129 8216 21163
rect 8063 20739 8097 20773
rect 9991 21238 10049 21293
rect 10972 21359 11006 21393
rect 11078 21239 11136 21294
rect 10960 20954 11018 21009
rect 12282 21400 12316 21434
rect 11326 21129 11360 21163
rect 11207 20739 11241 20773
rect 13193 21234 13251 21289
rect 14174 21355 14208 21389
rect 14280 21235 14338 21290
rect 14162 20950 14220 21005
rect 1729 20136 1763 20170
rect 4873 20136 4907 20170
rect 15484 21396 15518 21430
rect 14528 21125 14562 21159
rect 14409 20735 14443 20769
rect 16337 21234 16395 21289
rect 17318 21355 17352 21389
rect 17424 21235 17482 21290
rect 17306 20950 17364 21005
rect 18628 21396 18662 21430
rect 17672 21125 17706 21159
rect 17553 20735 17587 20769
rect 19469 21238 19527 21293
rect 20450 21359 20484 21393
rect 20556 21239 20614 21294
rect 20438 20954 20496 21009
rect 21760 21400 21794 21434
rect 20804 21129 20838 21163
rect 20685 20739 20719 20773
rect 22613 21238 22671 21293
rect 23594 21359 23628 21393
rect 23700 21239 23758 21294
rect 23582 20954 23640 21009
rect 24904 21400 24938 21434
rect 23948 21129 23982 21163
rect 23829 20739 23863 20773
rect 8005 20140 8039 20174
rect 11149 20140 11183 20174
rect 14351 20136 14385 20170
rect 17495 20136 17529 20170
rect 20627 20140 20661 20174
rect 23771 20140 23805 20174
rect 14582 16934 14616 16968
rect 15750 16934 15784 16968
rect 16918 16934 16952 16968
rect 18086 16934 18120 16968
rect 19260 16936 19294 16970
rect 20428 16936 20462 16970
rect 21596 16936 21630 16970
rect 22764 16936 22798 16970
rect 14582 16826 14616 16860
rect 15750 16826 15784 16860
rect 16918 16826 16952 16860
rect 3676 16329 3710 16363
rect 3558 16212 3592 16246
rect 5124 16329 5158 16363
rect 5006 16212 5040 16246
rect 6622 16331 6656 16365
rect 6504 16214 6538 16248
rect 8070 16331 8104 16365
rect 7952 16214 7986 16248
rect 9590 16329 9624 16363
rect 9472 16212 9506 16246
rect 11038 16329 11072 16363
rect 10920 16212 10954 16246
rect 12536 16331 12570 16365
rect 12418 16214 12452 16248
rect 18086 16826 18120 16860
rect 19260 16828 19294 16862
rect 20428 16828 20462 16862
rect 13984 16331 14018 16365
rect 13866 16214 13900 16248
rect 14877 16063 14911 16097
rect 21596 16828 21630 16862
rect 22764 16828 22798 16862
rect 16045 16063 16079 16097
rect 17213 16063 17247 16097
rect 18381 16063 18415 16097
rect 19555 16065 19589 16099
rect 20723 16065 20757 16099
rect 3205 15702 3239 15736
rect 3323 15702 3357 15736
rect 4653 15702 4687 15736
rect 4771 15702 4805 15736
rect 6151 15704 6185 15738
rect 6269 15704 6303 15738
rect 7599 15704 7633 15738
rect 7717 15704 7751 15738
rect 9119 15702 9153 15736
rect 9237 15702 9271 15736
rect 10567 15702 10601 15736
rect 10685 15702 10719 15736
rect 12065 15704 12099 15738
rect 12183 15704 12217 15738
rect 13513 15704 13547 15738
rect 21891 16065 21925 16099
rect 23059 16065 23093 16099
rect 13631 15704 13665 15738
rect 3073 14096 3131 14151
rect 4054 14217 4088 14251
rect 4160 14097 4218 14152
rect 4042 13812 4100 13867
rect 5364 14258 5398 14292
rect 4408 13987 4442 14021
rect 4289 13597 4323 13631
rect 6217 14096 6275 14151
rect 7198 14217 7232 14251
rect 7304 14097 7362 14152
rect 7186 13812 7244 13867
rect 8508 14258 8542 14292
rect 7552 13987 7586 14021
rect 7433 13597 7467 13631
rect 9349 14100 9407 14155
rect 10330 14221 10364 14255
rect 10436 14101 10494 14156
rect 10318 13816 10376 13871
rect 11640 14262 11674 14296
rect 10684 13991 10718 14025
rect 10565 13601 10599 13635
rect 12493 14100 12551 14155
rect 13474 14221 13508 14255
rect 13580 14101 13638 14156
rect 13462 13816 13520 13871
rect 14784 14262 14818 14296
rect 13828 13991 13862 14025
rect 13709 13601 13743 13635
rect 15695 14096 15753 14151
rect 16676 14217 16710 14251
rect 16782 14097 16840 14152
rect 16664 13812 16722 13867
rect 4231 12998 4265 13032
rect 7375 12998 7409 13032
rect 17986 14258 18020 14292
rect 17030 13987 17064 14021
rect 16911 13597 16945 13631
rect 18839 14096 18897 14151
rect 19820 14217 19854 14251
rect 19926 14097 19984 14152
rect 19808 13812 19866 13867
rect 21130 14258 21164 14292
rect 20174 13987 20208 14021
rect 20055 13597 20089 13631
rect 21971 14100 22029 14155
rect 22952 14221 22986 14255
rect 23058 14101 23116 14156
rect 22940 13816 22998 13871
rect 24262 14262 24296 14296
rect 23306 13991 23340 14025
rect 23187 13601 23221 13635
rect 25115 14100 25173 14155
rect 26096 14221 26130 14255
rect 26202 14101 26260 14156
rect 26084 13816 26142 13871
rect 27406 14262 27440 14296
rect 26450 13991 26484 14025
rect 26331 13601 26365 13635
rect 10507 13002 10541 13036
rect 13651 13002 13685 13036
rect 16853 12998 16887 13032
rect 19997 12998 20031 13032
rect 23129 13002 23163 13036
rect 26273 13002 26307 13036
rect 3073 11362 3131 11417
rect 4054 11483 4088 11517
rect 4160 11363 4218 11418
rect 4042 11078 4100 11133
rect 5364 11524 5398 11558
rect 4408 11253 4442 11287
rect 4289 10863 4323 10897
rect 6217 11362 6275 11417
rect 7198 11483 7232 11517
rect 7304 11363 7362 11418
rect 7186 11078 7244 11133
rect 8508 11524 8542 11558
rect 7552 11253 7586 11287
rect 7433 10863 7467 10897
rect 9349 11366 9407 11421
rect 10330 11487 10364 11521
rect 10436 11367 10494 11422
rect 10318 11082 10376 11137
rect 11640 11528 11674 11562
rect 10684 11257 10718 11291
rect 10565 10867 10599 10901
rect 12493 11366 12551 11421
rect 13474 11487 13508 11521
rect 13580 11367 13638 11422
rect 13462 11082 13520 11137
rect 14784 11528 14818 11562
rect 13828 11257 13862 11291
rect 13709 10867 13743 10901
rect 15695 11362 15753 11417
rect 16676 11483 16710 11517
rect 16782 11363 16840 11418
rect 16664 11078 16722 11133
rect 4231 10264 4265 10298
rect 7375 10264 7409 10298
rect 17986 11524 18020 11558
rect 17030 11253 17064 11287
rect 16911 10863 16945 10897
rect 18839 11362 18897 11417
rect 19820 11483 19854 11517
rect 19926 11363 19984 11418
rect 19808 11078 19866 11133
rect 21130 11524 21164 11558
rect 20174 11253 20208 11287
rect 20055 10863 20089 10897
rect 21971 11366 22029 11421
rect 22952 11487 22986 11521
rect 23058 11367 23116 11422
rect 22940 11082 22998 11137
rect 24262 11528 24296 11562
rect 23306 11257 23340 11291
rect 23187 10867 23221 10901
rect 25115 11366 25173 11421
rect 26096 11487 26130 11521
rect 26202 11367 26260 11422
rect 26084 11082 26142 11137
rect 27406 11528 27440 11562
rect 26450 11257 26484 11291
rect 26331 10867 26365 10901
rect 10507 10268 10541 10302
rect 13651 10268 13685 10302
rect 16853 10264 16887 10298
rect 19997 10264 20031 10298
rect 23129 10268 23163 10302
rect 26273 10268 26307 10302
rect 3063 8630 3121 8685
rect 4044 8751 4078 8785
rect 4150 8631 4208 8686
rect 4032 8346 4090 8401
rect 5354 8792 5388 8826
rect 4398 8521 4432 8555
rect 4279 8131 4313 8165
rect 6207 8630 6265 8685
rect 7188 8751 7222 8785
rect 7294 8631 7352 8686
rect 7176 8346 7234 8401
rect 8498 8792 8532 8826
rect 7542 8521 7576 8555
rect 7423 8131 7457 8165
rect 9339 8634 9397 8689
rect 10320 8755 10354 8789
rect 10426 8635 10484 8690
rect 10308 8350 10366 8405
rect 11630 8796 11664 8830
rect 10674 8525 10708 8559
rect 10555 8135 10589 8169
rect 12483 8634 12541 8689
rect 13464 8755 13498 8789
rect 13570 8635 13628 8690
rect 13452 8350 13510 8405
rect 14774 8796 14808 8830
rect 13818 8525 13852 8559
rect 13699 8135 13733 8169
rect 15685 8630 15743 8685
rect 16666 8751 16700 8785
rect 16772 8631 16830 8686
rect 16654 8346 16712 8401
rect 4221 7532 4255 7566
rect 7365 7532 7399 7566
rect 17976 8792 18010 8826
rect 17020 8521 17054 8555
rect 16901 8131 16935 8165
rect 18829 8630 18887 8685
rect 19810 8751 19844 8785
rect 19916 8631 19974 8686
rect 19798 8346 19856 8401
rect 21120 8792 21154 8826
rect 20164 8521 20198 8555
rect 20045 8131 20079 8165
rect 21961 8634 22019 8689
rect 22942 8755 22976 8789
rect 23048 8635 23106 8690
rect 22930 8350 22988 8405
rect 24252 8796 24286 8830
rect 23296 8525 23330 8559
rect 23177 8135 23211 8169
rect 25105 8634 25163 8689
rect 26086 8755 26120 8789
rect 26192 8635 26250 8690
rect 26074 8350 26132 8405
rect 27396 8796 27430 8830
rect 26440 8525 26474 8559
rect 26321 8135 26355 8169
rect 10497 7536 10531 7570
rect 13641 7536 13675 7570
rect 16843 7532 16877 7566
rect 19987 7532 20021 7566
rect 23119 7536 23153 7570
rect 26263 7536 26297 7570
rect 4112 5842 4146 5876
rect 2718 5648 2752 5682
rect 3152 5140 3186 5174
rect 2967 5073 3001 5107
rect 3800 5140 3834 5174
rect 3418 5056 3452 5090
rect 3536 5057 3570 5091
rect 6180 5844 6214 5878
rect 4786 5650 4820 5684
rect 4090 5072 4124 5106
rect 5220 5142 5254 5176
rect 5035 5075 5069 5109
rect 5868 5142 5902 5176
rect 5486 5058 5520 5092
rect 5604 5059 5638 5093
rect 8249 5842 8283 5876
rect 6855 5648 6889 5682
rect 6158 5074 6192 5108
rect 7289 5140 7323 5174
rect 7104 5073 7138 5107
rect 7937 5140 7971 5174
rect 7555 5056 7589 5090
rect 7673 5057 7707 5091
rect 10317 5844 10351 5878
rect 8923 5650 8957 5684
rect 8227 5072 8261 5106
rect 9357 5142 9391 5176
rect 9172 5075 9206 5109
rect 10005 5142 10039 5176
rect 9623 5058 9657 5092
rect 9741 5059 9775 5093
rect 12386 5844 12420 5878
rect 10992 5650 11026 5684
rect 10295 5074 10329 5108
rect 11426 5142 11460 5176
rect 11241 5075 11275 5109
rect 12074 5142 12108 5176
rect 11692 5058 11726 5092
rect 11810 5059 11844 5093
rect 19603 6231 19637 6265
rect 20341 6229 20375 6263
rect 21079 6229 21113 6263
rect 14454 5846 14488 5880
rect 13060 5652 13094 5686
rect 12364 5074 12398 5108
rect 13494 5144 13528 5178
rect 13309 5077 13343 5111
rect 14142 5144 14176 5178
rect 13760 5060 13794 5094
rect 13878 5061 13912 5095
rect 16523 5844 16557 5878
rect 15129 5650 15163 5684
rect 14432 5076 14466 5110
rect 15563 5142 15597 5176
rect 15378 5075 15412 5109
rect 16211 5142 16245 5176
rect 15829 5058 15863 5092
rect 15947 5059 15981 5093
rect 21821 6229 21855 6263
rect 22561 6229 22595 6263
rect 23299 6229 23333 6263
rect 24037 6229 24071 6263
rect 24775 6229 24809 6263
rect 18591 5846 18625 5880
rect 17197 5652 17231 5686
rect 16501 5074 16535 5108
rect 17631 5144 17665 5178
rect 17446 5077 17480 5111
rect 18279 5144 18313 5178
rect 17897 5060 17931 5094
rect 18015 5061 18049 5095
rect 18569 5076 18603 5110
rect 365 1382 423 1437
rect 1346 1503 1380 1537
rect 1452 1383 1510 1438
rect 1334 1098 1392 1153
rect 2656 1544 2690 1578
rect 1700 1273 1734 1307
rect 1581 883 1615 917
rect 3509 1382 3567 1437
rect 4490 1503 4524 1537
rect 4596 1383 4654 1438
rect 4478 1098 4536 1153
rect 5800 1544 5834 1578
rect 4844 1273 4878 1307
rect 4725 883 4759 917
rect 6641 1386 6699 1441
rect 7622 1507 7656 1541
rect 7728 1387 7786 1442
rect 7610 1102 7668 1157
rect 8932 1548 8966 1582
rect 7976 1277 8010 1311
rect 7857 887 7891 921
rect 9785 1386 9843 1441
rect 10766 1507 10800 1541
rect 10872 1387 10930 1442
rect 10754 1102 10812 1157
rect 12076 1548 12110 1582
rect 11120 1277 11154 1311
rect 11001 887 11035 921
rect 12987 1382 13045 1437
rect 13968 1503 14002 1537
rect 14074 1383 14132 1438
rect 13956 1098 14014 1153
rect 1523 284 1557 318
rect 4667 284 4701 318
rect 15278 1544 15312 1578
rect 14322 1273 14356 1307
rect 14203 883 14237 917
rect 16131 1382 16189 1437
rect 17112 1503 17146 1537
rect 17218 1383 17276 1438
rect 17100 1098 17158 1153
rect 18422 1544 18456 1578
rect 17466 1273 17500 1307
rect 17347 883 17381 917
rect 19263 1386 19321 1441
rect 20244 1507 20278 1541
rect 20350 1387 20408 1442
rect 20232 1102 20290 1157
rect 21554 1548 21588 1582
rect 20598 1277 20632 1311
rect 20479 887 20513 921
rect 22407 1386 22465 1441
rect 23388 1507 23422 1541
rect 23494 1387 23552 1442
rect 23376 1102 23434 1157
rect 24698 1548 24732 1582
rect 23742 1277 23776 1311
rect 23623 887 23657 921
rect 7799 288 7833 322
rect 10943 288 10977 322
rect 14145 284 14179 318
rect 17289 284 17323 318
rect 20421 288 20455 322
rect 23565 288 23599 322
rect 397 -2510 455 -2455
rect 1378 -2389 1412 -2355
rect 1484 -2509 1542 -2454
rect 1366 -2794 1424 -2739
rect 2688 -2348 2722 -2314
rect 1732 -2619 1766 -2585
rect 1613 -3009 1647 -2975
rect 3541 -2510 3599 -2455
rect 4522 -2389 4556 -2355
rect 4628 -2509 4686 -2454
rect 4510 -2794 4568 -2739
rect 5832 -2348 5866 -2314
rect 4876 -2619 4910 -2585
rect 4757 -3009 4791 -2975
rect 6673 -2506 6731 -2451
rect 7654 -2385 7688 -2351
rect 7760 -2505 7818 -2450
rect 7642 -2790 7700 -2735
rect 8964 -2344 8998 -2310
rect 8008 -2615 8042 -2581
rect 7889 -3005 7923 -2971
rect 9817 -2506 9875 -2451
rect 10798 -2385 10832 -2351
rect 10904 -2505 10962 -2450
rect 10786 -2790 10844 -2735
rect 12108 -2344 12142 -2310
rect 11152 -2615 11186 -2581
rect 11033 -3005 11067 -2971
rect 13019 -2510 13077 -2455
rect 14000 -2389 14034 -2355
rect 14106 -2509 14164 -2454
rect 13988 -2794 14046 -2739
rect 1555 -3608 1589 -3574
rect 4699 -3608 4733 -3574
rect 15310 -2348 15344 -2314
rect 14354 -2619 14388 -2585
rect 14235 -3009 14269 -2975
rect 16163 -2510 16221 -2455
rect 17144 -2389 17178 -2355
rect 17250 -2509 17308 -2454
rect 17132 -2794 17190 -2739
rect 18454 -2348 18488 -2314
rect 17498 -2619 17532 -2585
rect 17379 -3009 17413 -2975
rect 19295 -2506 19353 -2451
rect 20276 -2385 20310 -2351
rect 20382 -2505 20440 -2450
rect 20264 -2790 20322 -2735
rect 21586 -2344 21620 -2310
rect 20630 -2615 20664 -2581
rect 20511 -3005 20545 -2971
rect 22439 -2506 22497 -2451
rect 23420 -2385 23454 -2351
rect 23526 -2505 23584 -2450
rect 23408 -2790 23466 -2735
rect 24730 -2344 24764 -2310
rect 23774 -2615 23808 -2581
rect 23655 -3005 23689 -2971
rect 7831 -3604 7865 -3570
rect 10975 -3604 11009 -3570
rect 14177 -3608 14211 -3574
rect 17321 -3608 17355 -3574
rect 20453 -3604 20487 -3570
rect 23597 -3604 23631 -3570
<< locali >>
rect 1636 22250 1864 22268
rect 1636 22174 1652 22250
rect 1848 22174 1864 22250
rect 1636 22158 1864 22174
rect 4780 22250 5008 22268
rect 4780 22174 4796 22250
rect 4992 22174 5008 22250
rect 4780 22158 5008 22174
rect 7912 22254 8140 22272
rect 7912 22178 7928 22254
rect 8124 22178 8140 22254
rect 7912 22162 8140 22178
rect 11056 22254 11284 22272
rect 11056 22178 11072 22254
rect 11268 22178 11284 22254
rect 11056 22162 11284 22178
rect 14258 22250 14486 22268
rect 14258 22174 14274 22250
rect 14470 22174 14486 22250
rect 14258 22158 14486 22174
rect 17402 22250 17630 22268
rect 17402 22174 17418 22250
rect 17614 22174 17630 22250
rect 17402 22158 17630 22174
rect 20534 22254 20762 22272
rect 20534 22178 20550 22254
rect 20746 22178 20762 22254
rect 20534 22162 20762 22178
rect 23678 22254 23906 22272
rect 23678 22178 23694 22254
rect 23890 22178 23906 22254
rect 23678 22162 23906 22178
rect 907 22033 1177 22072
rect 907 21980 941 22033
rect 466 21831 736 21870
rect 466 21780 500 21831
rect 466 21588 500 21604
rect 584 21780 618 21796
rect 584 21553 618 21604
rect 702 21780 736 21831
rect 702 21588 736 21604
rect 820 21780 854 21796
rect 820 21553 854 21604
rect 907 21588 941 21604
rect 1025 21980 1059 21996
rect 584 21514 854 21553
rect 1025 21553 1059 21604
rect 1143 21980 1177 22033
rect 1374 22032 1644 22071
rect 1143 21588 1177 21604
rect 1261 21980 1295 21996
rect 1261 21553 1295 21604
rect 1374 21980 1408 22032
rect 1374 21588 1408 21604
rect 1492 21980 1526 21996
rect 1492 21553 1526 21604
rect 1610 21980 1644 22032
rect 1846 22032 2116 22071
rect 1610 21588 1644 21604
rect 1728 21980 1762 21996
rect 1728 21553 1762 21604
rect 1846 21980 1880 22032
rect 1846 21588 1880 21604
rect 1964 21980 1998 21996
rect 1964 21553 1998 21604
rect 2082 21980 2116 22032
rect 2319 22032 2589 22071
rect 2082 21588 2116 21604
rect 2201 21980 2235 21996
rect 2201 21553 2235 21604
rect 2319 21980 2353 22032
rect 2319 21588 2353 21604
rect 2437 21980 2471 21996
rect 2437 21553 2471 21604
rect 2555 21980 2589 22032
rect 4051 22033 4321 22072
rect 4051 21980 4085 22033
rect 2792 21830 3062 21867
rect 2555 21588 2589 21604
rect 2674 21780 2708 21796
rect 1025 21514 2471 21553
rect 2674 21550 2708 21604
rect 2792 21780 2826 21830
rect 2792 21588 2826 21604
rect 2910 21780 2944 21796
rect 2910 21550 2944 21604
rect 3028 21780 3062 21830
rect 3028 21588 3062 21604
rect 3610 21831 3880 21870
rect 3610 21780 3644 21831
rect 3610 21588 3644 21604
rect 3728 21780 3762 21796
rect 2674 21511 2944 21550
rect 3728 21553 3762 21604
rect 3846 21780 3880 21831
rect 3846 21588 3880 21604
rect 3964 21780 3998 21796
rect 3964 21553 3998 21604
rect 4051 21588 4085 21604
rect 4169 21980 4203 21996
rect 3728 21514 3998 21553
rect 4169 21553 4203 21604
rect 4287 21980 4321 22033
rect 4518 22032 4788 22071
rect 4287 21588 4321 21604
rect 4405 21980 4439 21996
rect 4405 21553 4439 21604
rect 4518 21980 4552 22032
rect 4518 21588 4552 21604
rect 4636 21980 4670 21996
rect 4636 21553 4670 21604
rect 4754 21980 4788 22032
rect 4990 22032 5260 22071
rect 4754 21588 4788 21604
rect 4872 21980 4906 21996
rect 4872 21553 4906 21604
rect 4990 21980 5024 22032
rect 4990 21588 5024 21604
rect 5108 21980 5142 21996
rect 5108 21553 5142 21604
rect 5226 21980 5260 22032
rect 5463 22032 5733 22071
rect 5226 21588 5260 21604
rect 5345 21980 5379 21996
rect 5345 21553 5379 21604
rect 5463 21980 5497 22032
rect 5463 21588 5497 21604
rect 5581 21980 5615 21996
rect 5581 21553 5615 21604
rect 5699 21980 5733 22032
rect 7183 22037 7453 22076
rect 7183 21984 7217 22037
rect 5936 21830 6206 21867
rect 5699 21588 5733 21604
rect 5818 21780 5852 21796
rect 4169 21514 5615 21553
rect 5818 21550 5852 21604
rect 5936 21780 5970 21830
rect 5936 21588 5970 21604
rect 6054 21780 6088 21796
rect 6054 21550 6088 21604
rect 6172 21780 6206 21830
rect 6172 21588 6206 21604
rect 6742 21835 7012 21874
rect 6742 21784 6776 21835
rect 6742 21592 6776 21608
rect 6860 21784 6894 21800
rect 5818 21511 6088 21550
rect 6860 21557 6894 21608
rect 6978 21784 7012 21835
rect 6978 21592 7012 21608
rect 7096 21784 7130 21800
rect 7096 21557 7130 21608
rect 7183 21592 7217 21608
rect 7301 21984 7335 22000
rect 6860 21518 7130 21557
rect 7301 21557 7335 21608
rect 7419 21984 7453 22037
rect 7650 22036 7920 22075
rect 7419 21592 7453 21608
rect 7537 21984 7571 22000
rect 7537 21557 7571 21608
rect 7650 21984 7684 22036
rect 7650 21592 7684 21608
rect 7768 21984 7802 22000
rect 7768 21557 7802 21608
rect 7886 21984 7920 22036
rect 8122 22036 8392 22075
rect 7886 21592 7920 21608
rect 8004 21984 8038 22000
rect 8004 21557 8038 21608
rect 8122 21984 8156 22036
rect 8122 21592 8156 21608
rect 8240 21984 8274 22000
rect 8240 21557 8274 21608
rect 8358 21984 8392 22036
rect 8595 22036 8865 22075
rect 8358 21592 8392 21608
rect 8477 21984 8511 22000
rect 8477 21557 8511 21608
rect 8595 21984 8629 22036
rect 8595 21592 8629 21608
rect 8713 21984 8747 22000
rect 8713 21557 8747 21608
rect 8831 21984 8865 22036
rect 10327 22037 10597 22076
rect 10327 21984 10361 22037
rect 9068 21834 9338 21871
rect 8831 21592 8865 21608
rect 8950 21784 8984 21800
rect 7301 21518 8747 21557
rect 8950 21554 8984 21608
rect 9068 21784 9102 21834
rect 9068 21592 9102 21608
rect 9186 21784 9220 21800
rect 9186 21554 9220 21608
rect 9304 21784 9338 21834
rect 9304 21592 9338 21608
rect 9886 21835 10156 21874
rect 9886 21784 9920 21835
rect 9886 21592 9920 21608
rect 10004 21784 10038 21800
rect 8950 21515 9220 21554
rect 10004 21557 10038 21608
rect 10122 21784 10156 21835
rect 10122 21592 10156 21608
rect 10240 21784 10274 21800
rect 10240 21557 10274 21608
rect 10327 21592 10361 21608
rect 10445 21984 10479 22000
rect 10004 21518 10274 21557
rect 10445 21557 10479 21608
rect 10563 21984 10597 22037
rect 10794 22036 11064 22075
rect 10563 21592 10597 21608
rect 10681 21984 10715 22000
rect 10681 21557 10715 21608
rect 10794 21984 10828 22036
rect 10794 21592 10828 21608
rect 10912 21984 10946 22000
rect 10912 21557 10946 21608
rect 11030 21984 11064 22036
rect 11266 22036 11536 22075
rect 11030 21592 11064 21608
rect 11148 21984 11182 22000
rect 11148 21557 11182 21608
rect 11266 21984 11300 22036
rect 11266 21592 11300 21608
rect 11384 21984 11418 22000
rect 11384 21557 11418 21608
rect 11502 21984 11536 22036
rect 11739 22036 12009 22075
rect 11502 21592 11536 21608
rect 11621 21984 11655 22000
rect 11621 21557 11655 21608
rect 11739 21984 11773 22036
rect 11739 21592 11773 21608
rect 11857 21984 11891 22000
rect 11857 21557 11891 21608
rect 11975 21984 12009 22036
rect 13529 22033 13799 22072
rect 13529 21980 13563 22033
rect 12212 21834 12482 21871
rect 11975 21592 12009 21608
rect 12094 21784 12128 21800
rect 10445 21518 11891 21557
rect 12094 21554 12128 21608
rect 12212 21784 12246 21834
rect 12212 21592 12246 21608
rect 12330 21784 12364 21800
rect 12330 21554 12364 21608
rect 12448 21784 12482 21834
rect 12448 21592 12482 21608
rect 13088 21831 13358 21870
rect 13088 21780 13122 21831
rect 13088 21588 13122 21604
rect 13206 21780 13240 21796
rect 12094 21515 12364 21554
rect 13206 21553 13240 21604
rect 13324 21780 13358 21831
rect 13324 21588 13358 21604
rect 13442 21780 13476 21796
rect 13442 21553 13476 21604
rect 13529 21588 13563 21604
rect 13647 21980 13681 21996
rect 13206 21514 13476 21553
rect 13647 21553 13681 21604
rect 13765 21980 13799 22033
rect 13996 22032 14266 22071
rect 13765 21588 13799 21604
rect 13883 21980 13917 21996
rect 13883 21553 13917 21604
rect 13996 21980 14030 22032
rect 13996 21588 14030 21604
rect 14114 21980 14148 21996
rect 14114 21553 14148 21604
rect 14232 21980 14266 22032
rect 14468 22032 14738 22071
rect 14232 21588 14266 21604
rect 14350 21980 14384 21996
rect 14350 21553 14384 21604
rect 14468 21980 14502 22032
rect 14468 21588 14502 21604
rect 14586 21980 14620 21996
rect 14586 21553 14620 21604
rect 14704 21980 14738 22032
rect 14941 22032 15211 22071
rect 14704 21588 14738 21604
rect 14823 21980 14857 21996
rect 14823 21553 14857 21604
rect 14941 21980 14975 22032
rect 14941 21588 14975 21604
rect 15059 21980 15093 21996
rect 15059 21553 15093 21604
rect 15177 21980 15211 22032
rect 16673 22033 16943 22072
rect 16673 21980 16707 22033
rect 15414 21830 15684 21867
rect 15177 21588 15211 21604
rect 15296 21780 15330 21796
rect 13647 21514 15093 21553
rect 15296 21550 15330 21604
rect 15414 21780 15448 21830
rect 15414 21588 15448 21604
rect 15532 21780 15566 21796
rect 15532 21550 15566 21604
rect 15650 21780 15684 21830
rect 15650 21588 15684 21604
rect 16232 21831 16502 21870
rect 16232 21780 16266 21831
rect 16232 21588 16266 21604
rect 16350 21780 16384 21796
rect 15296 21511 15566 21550
rect 16350 21553 16384 21604
rect 16468 21780 16502 21831
rect 16468 21588 16502 21604
rect 16586 21780 16620 21796
rect 16586 21553 16620 21604
rect 16673 21588 16707 21604
rect 16791 21980 16825 21996
rect 16350 21514 16620 21553
rect 16791 21553 16825 21604
rect 16909 21980 16943 22033
rect 17140 22032 17410 22071
rect 16909 21588 16943 21604
rect 17027 21980 17061 21996
rect 17027 21553 17061 21604
rect 17140 21980 17174 22032
rect 17140 21588 17174 21604
rect 17258 21980 17292 21996
rect 17258 21553 17292 21604
rect 17376 21980 17410 22032
rect 17612 22032 17882 22071
rect 17376 21588 17410 21604
rect 17494 21980 17528 21996
rect 17494 21553 17528 21604
rect 17612 21980 17646 22032
rect 17612 21588 17646 21604
rect 17730 21980 17764 21996
rect 17730 21553 17764 21604
rect 17848 21980 17882 22032
rect 18085 22032 18355 22071
rect 17848 21588 17882 21604
rect 17967 21980 18001 21996
rect 17967 21553 18001 21604
rect 18085 21980 18119 22032
rect 18085 21588 18119 21604
rect 18203 21980 18237 21996
rect 18203 21553 18237 21604
rect 18321 21980 18355 22032
rect 19805 22037 20075 22076
rect 19805 21984 19839 22037
rect 18558 21830 18828 21867
rect 18321 21588 18355 21604
rect 18440 21780 18474 21796
rect 16791 21514 18237 21553
rect 18440 21550 18474 21604
rect 18558 21780 18592 21830
rect 18558 21588 18592 21604
rect 18676 21780 18710 21796
rect 18676 21550 18710 21604
rect 18794 21780 18828 21830
rect 18794 21588 18828 21604
rect 19364 21835 19634 21874
rect 19364 21784 19398 21835
rect 19364 21592 19398 21608
rect 19482 21784 19516 21800
rect 18440 21511 18710 21550
rect 19482 21557 19516 21608
rect 19600 21784 19634 21835
rect 19600 21592 19634 21608
rect 19718 21784 19752 21800
rect 19718 21557 19752 21608
rect 19805 21592 19839 21608
rect 19923 21984 19957 22000
rect 19482 21518 19752 21557
rect 19923 21557 19957 21608
rect 20041 21984 20075 22037
rect 20272 22036 20542 22075
rect 20041 21592 20075 21608
rect 20159 21984 20193 22000
rect 20159 21557 20193 21608
rect 20272 21984 20306 22036
rect 20272 21592 20306 21608
rect 20390 21984 20424 22000
rect 20390 21557 20424 21608
rect 20508 21984 20542 22036
rect 20744 22036 21014 22075
rect 20508 21592 20542 21608
rect 20626 21984 20660 22000
rect 20626 21557 20660 21608
rect 20744 21984 20778 22036
rect 20744 21592 20778 21608
rect 20862 21984 20896 22000
rect 20862 21557 20896 21608
rect 20980 21984 21014 22036
rect 21217 22036 21487 22075
rect 20980 21592 21014 21608
rect 21099 21984 21133 22000
rect 21099 21557 21133 21608
rect 21217 21984 21251 22036
rect 21217 21592 21251 21608
rect 21335 21984 21369 22000
rect 21335 21557 21369 21608
rect 21453 21984 21487 22036
rect 22949 22037 23219 22076
rect 22949 21984 22983 22037
rect 21690 21834 21960 21871
rect 21453 21592 21487 21608
rect 21572 21784 21606 21800
rect 19923 21518 21369 21557
rect 21572 21554 21606 21608
rect 21690 21784 21724 21834
rect 21690 21592 21724 21608
rect 21808 21784 21842 21800
rect 21808 21554 21842 21608
rect 21926 21784 21960 21834
rect 21926 21592 21960 21608
rect 22508 21835 22778 21874
rect 22508 21784 22542 21835
rect 22508 21592 22542 21608
rect 22626 21784 22660 21800
rect 21572 21515 21842 21554
rect 22626 21557 22660 21608
rect 22744 21784 22778 21835
rect 22744 21592 22778 21608
rect 22862 21784 22896 21800
rect 22862 21557 22896 21608
rect 22949 21592 22983 21608
rect 23067 21984 23101 22000
rect 22626 21518 22896 21557
rect 23067 21557 23101 21608
rect 23185 21984 23219 22037
rect 23416 22036 23686 22075
rect 23185 21592 23219 21608
rect 23303 21984 23337 22000
rect 23303 21557 23337 21608
rect 23416 21984 23450 22036
rect 23416 21592 23450 21608
rect 23534 21984 23568 22000
rect 23534 21557 23568 21608
rect 23652 21984 23686 22036
rect 23888 22036 24158 22075
rect 23652 21592 23686 21608
rect 23770 21984 23804 22000
rect 23770 21557 23804 21608
rect 23888 21984 23922 22036
rect 23888 21592 23922 21608
rect 24006 21984 24040 22000
rect 24006 21557 24040 21608
rect 24124 21984 24158 22036
rect 24361 22036 24631 22075
rect 24124 21592 24158 21608
rect 24243 21984 24277 22000
rect 24243 21557 24277 21608
rect 24361 21984 24395 22036
rect 24361 21592 24395 21608
rect 24479 21984 24513 22000
rect 24479 21557 24513 21608
rect 24597 21984 24631 22036
rect 24834 21834 25104 21871
rect 24597 21592 24631 21608
rect 24716 21784 24750 21800
rect 23067 21518 24513 21557
rect 24716 21554 24750 21608
rect 24834 21784 24868 21834
rect 24834 21592 24868 21608
rect 24952 21784 24986 21800
rect 24952 21554 24986 21608
rect 25070 21784 25104 21834
rect 25070 21592 25104 21608
rect 24716 21515 24986 21554
rect 1552 21389 1586 21405
rect 2846 21396 2862 21430
rect 2896 21396 2912 21430
rect 1552 21339 1586 21355
rect 4696 21389 4730 21405
rect 5990 21396 6006 21430
rect 6040 21396 6056 21430
rect 4696 21339 4730 21355
rect 7828 21393 7862 21409
rect 9122 21400 9138 21434
rect 9172 21400 9188 21434
rect 7828 21343 7862 21359
rect 10972 21393 11006 21409
rect 12266 21400 12282 21434
rect 12316 21400 12332 21434
rect 10972 21343 11006 21359
rect 14174 21389 14208 21405
rect 15468 21396 15484 21430
rect 15518 21396 15534 21430
rect 14174 21339 14208 21355
rect 17318 21389 17352 21405
rect 18612 21396 18628 21430
rect 18662 21396 18678 21430
rect 17318 21339 17352 21355
rect 20450 21393 20484 21409
rect 21744 21400 21760 21434
rect 21794 21400 21810 21434
rect 20450 21343 20484 21359
rect 23594 21393 23628 21409
rect 24888 21400 24904 21434
rect 24938 21400 24954 21434
rect 23594 21343 23628 21359
rect 323 21290 380 21294
rect 323 21230 327 21290
rect 376 21230 380 21290
rect 323 21226 380 21230
rect 555 21289 647 21306
rect 555 21234 571 21289
rect 631 21234 647 21289
rect 555 21221 647 21234
rect 1640 21290 1732 21303
rect 1640 21235 1656 21290
rect 1716 21235 1732 21290
rect 1640 21218 1732 21235
rect 3699 21289 3791 21306
rect 3699 21234 3715 21289
rect 3775 21234 3791 21289
rect 3699 21221 3791 21234
rect 4784 21290 4876 21303
rect 4784 21235 4800 21290
rect 4860 21235 4876 21290
rect 4784 21218 4876 21235
rect 6831 21293 6923 21310
rect 6831 21238 6847 21293
rect 6907 21238 6923 21293
rect 6831 21225 6923 21238
rect 7916 21294 8008 21307
rect 7916 21239 7932 21294
rect 7992 21239 8008 21294
rect 7916 21222 8008 21239
rect 9975 21293 10067 21310
rect 9975 21238 9991 21293
rect 10051 21238 10067 21293
rect 9975 21225 10067 21238
rect 11060 21294 11152 21307
rect 11060 21239 11076 21294
rect 11136 21239 11152 21294
rect 11060 21222 11152 21239
rect 13177 21289 13269 21306
rect 13177 21234 13193 21289
rect 13253 21234 13269 21289
rect 13177 21221 13269 21234
rect 14262 21290 14354 21303
rect 14262 21235 14278 21290
rect 14338 21235 14354 21290
rect 14262 21218 14354 21235
rect 16321 21289 16413 21306
rect 16321 21234 16337 21289
rect 16397 21234 16413 21289
rect 16321 21221 16413 21234
rect 17406 21290 17498 21303
rect 17406 21235 17422 21290
rect 17482 21235 17498 21290
rect 17406 21218 17498 21235
rect 19453 21293 19545 21310
rect 19453 21238 19469 21293
rect 19529 21238 19545 21293
rect 19453 21225 19545 21238
rect 20538 21294 20630 21307
rect 20538 21239 20554 21294
rect 20614 21239 20630 21294
rect 20538 21222 20630 21239
rect 22597 21293 22689 21310
rect 22597 21238 22613 21293
rect 22673 21238 22689 21293
rect 22597 21225 22689 21238
rect 23682 21294 23774 21307
rect 23682 21239 23698 21294
rect 23758 21239 23774 21294
rect 23682 21222 23774 21239
rect 1906 21159 1940 21175
rect 1906 21109 1940 21125
rect 3467 21174 3524 21178
rect 3467 21114 3471 21174
rect 3520 21114 3524 21174
rect 3467 21110 3524 21114
rect 5050 21159 5084 21175
rect 5050 21109 5084 21125
rect 8182 21163 8216 21179
rect 8182 21113 8216 21129
rect 9617 21178 9812 21182
rect 9617 21118 9747 21178
rect 9796 21118 9812 21178
rect 9617 21110 9812 21118
rect 11326 21163 11360 21179
rect 15868 21178 16122 21179
rect 19221 21178 19278 21182
rect 11326 21113 11360 21129
rect 14528 21159 14562 21175
rect 9617 21107 9675 21110
rect 14528 21109 14562 21125
rect 15868 21174 16146 21178
rect 15868 21114 16093 21174
rect 16142 21114 16146 21174
rect 15868 21110 16146 21114
rect 17672 21159 17706 21175
rect 9444 21050 9675 21107
rect 323 21006 380 21010
rect 323 20946 327 21006
rect 376 20946 380 21006
rect 323 20942 380 20946
rect 1522 21005 1614 21018
rect 1522 20950 1538 21005
rect 1598 20950 1614 21005
rect 1522 20933 1614 20950
rect 3467 21006 3524 21010
rect 3467 20946 3471 21006
rect 3520 20946 3524 21006
rect 3467 20942 3524 20946
rect 4666 21005 6073 21018
rect 4666 20950 4682 21005
rect 4742 20950 6073 21005
rect 4666 20933 6073 20950
rect 6599 21010 6656 21014
rect 6599 20950 6603 21010
rect 6652 20950 6656 21010
rect 6599 20946 6656 20950
rect 7798 21009 7890 21022
rect 7798 20954 7814 21009
rect 7874 20954 7890 21009
rect 7798 20937 7890 20954
rect 5993 20876 6073 20933
rect 9444 20876 9521 21050
rect 9743 21010 9800 21014
rect 9743 20950 9747 21010
rect 9796 20950 9800 21010
rect 9743 20946 9800 20950
rect 10942 21009 11814 21022
rect 10942 20954 10958 21009
rect 11018 20954 11814 21009
rect 10942 20937 11814 20954
rect 12945 21006 13002 21010
rect 12945 20946 12949 21006
rect 12998 20946 13002 21006
rect 12945 20942 13002 20946
rect 14144 21005 14236 21018
rect 14144 20950 14160 21005
rect 14220 20950 14236 21005
rect 5993 20823 9521 20876
rect 11737 20882 11814 20937
rect 14144 20933 14236 20950
rect 15868 20882 15936 21110
rect 17672 21109 17706 21125
rect 19221 21118 19225 21178
rect 19274 21118 19278 21178
rect 19221 21114 19278 21118
rect 20804 21163 20838 21179
rect 20804 21113 20838 21129
rect 22171 21178 22422 21182
rect 22171 21118 22369 21178
rect 22418 21118 22422 21178
rect 22171 21114 22422 21118
rect 23948 21163 23982 21179
rect 16089 21006 16146 21010
rect 16089 20946 16093 21006
rect 16142 20946 16146 21006
rect 16089 20942 16146 20946
rect 17288 21005 18225 21018
rect 17288 20950 17304 21005
rect 17364 20950 18225 21005
rect 17288 20933 18225 20950
rect 19221 21010 19278 21014
rect 19221 20950 19225 21010
rect 19274 20950 19278 21010
rect 19221 20946 19278 20950
rect 20420 21009 20512 21022
rect 20420 20954 20436 21009
rect 20496 20954 20512 21009
rect 20420 20937 20512 20954
rect 11737 20820 15936 20882
rect 18150 20888 18225 20933
rect 22171 20888 22228 21114
rect 23948 21113 23982 21129
rect 23564 21009 23656 21022
rect 23564 20954 23580 21009
rect 23640 20954 23656 21009
rect 23564 20937 23656 20954
rect 18150 20823 22228 20888
rect 1787 20769 1821 20785
rect 1787 20719 1821 20735
rect 4931 20769 4965 20785
rect 4931 20719 4965 20735
rect 8063 20773 8097 20789
rect 8063 20723 8097 20739
rect 11207 20773 11241 20789
rect 11207 20723 11241 20739
rect 14409 20769 14443 20785
rect 14409 20719 14443 20735
rect 17553 20769 17587 20785
rect 17553 20719 17587 20735
rect 20685 20773 20719 20789
rect 20685 20723 20719 20739
rect 23829 20773 23863 20789
rect 23829 20723 23863 20739
rect 1300 20647 1334 20663
rect 1300 20455 1334 20471
rect 1418 20659 1452 20663
rect 1492 20659 1526 20663
rect 1418 20647 1526 20659
rect 1452 20471 1492 20647
rect 1418 20459 1492 20471
rect 1418 20455 1452 20459
rect 1492 20255 1526 20271
rect 1610 20647 1644 20663
rect 1610 20255 1644 20271
rect 1728 20647 1762 20663
rect 1728 20255 1762 20271
rect 1846 20647 1880 20663
rect 1846 20255 1880 20271
rect 1964 20659 1998 20663
rect 2042 20659 2076 20663
rect 1964 20647 2076 20659
rect 1998 20471 2042 20647
rect 1998 20459 2076 20471
rect 2042 20455 2076 20459
rect 2160 20647 2194 20663
rect 2160 20455 2194 20471
rect 4444 20647 4478 20663
rect 4444 20455 4478 20471
rect 4562 20659 4596 20663
rect 4636 20659 4670 20663
rect 4562 20647 4670 20659
rect 4596 20471 4636 20647
rect 4562 20459 4636 20471
rect 4562 20455 4596 20459
rect 1964 20255 1998 20271
rect 4636 20255 4670 20271
rect 4754 20647 4788 20663
rect 4754 20255 4788 20271
rect 4872 20647 4906 20663
rect 4872 20255 4906 20271
rect 4990 20647 5024 20663
rect 4990 20255 5024 20271
rect 5108 20659 5142 20663
rect 5186 20659 5220 20663
rect 5108 20647 5220 20659
rect 5142 20471 5186 20647
rect 5142 20459 5220 20471
rect 5186 20455 5220 20459
rect 5304 20647 5338 20663
rect 5304 20455 5338 20471
rect 7576 20651 7610 20667
rect 7576 20459 7610 20475
rect 7694 20663 7728 20667
rect 7768 20663 7802 20667
rect 7694 20651 7802 20663
rect 7728 20475 7768 20651
rect 7694 20463 7768 20475
rect 7694 20459 7728 20463
rect 5108 20255 5142 20271
rect 7768 20259 7802 20275
rect 7886 20651 7920 20667
rect 7886 20259 7920 20275
rect 8004 20651 8038 20667
rect 8004 20259 8038 20275
rect 8122 20651 8156 20667
rect 8122 20259 8156 20275
rect 8240 20663 8274 20667
rect 8318 20663 8352 20667
rect 8240 20651 8352 20663
rect 8274 20475 8318 20651
rect 8274 20463 8352 20475
rect 8318 20459 8352 20463
rect 8436 20651 8470 20667
rect 8436 20459 8470 20475
rect 10720 20651 10754 20667
rect 10720 20459 10754 20475
rect 10838 20663 10872 20667
rect 10912 20663 10946 20667
rect 10838 20651 10946 20663
rect 10872 20475 10912 20651
rect 10838 20463 10912 20475
rect 10838 20459 10872 20463
rect 8240 20259 8274 20275
rect 10912 20259 10946 20275
rect 11030 20651 11064 20667
rect 11030 20259 11064 20275
rect 11148 20651 11182 20667
rect 11148 20259 11182 20275
rect 11266 20651 11300 20667
rect 11266 20259 11300 20275
rect 11384 20663 11418 20667
rect 11462 20663 11496 20667
rect 11384 20651 11496 20663
rect 11418 20475 11462 20651
rect 11418 20463 11496 20475
rect 11462 20459 11496 20463
rect 11580 20651 11614 20667
rect 11580 20459 11614 20475
rect 13922 20647 13956 20663
rect 13922 20455 13956 20471
rect 14040 20659 14074 20663
rect 14114 20659 14148 20663
rect 14040 20647 14148 20659
rect 14074 20471 14114 20647
rect 14040 20459 14114 20471
rect 14040 20455 14074 20459
rect 11384 20259 11418 20275
rect 14114 20255 14148 20271
rect 14232 20647 14266 20663
rect 14232 20255 14266 20271
rect 14350 20647 14384 20663
rect 14350 20255 14384 20271
rect 14468 20647 14502 20663
rect 14468 20255 14502 20271
rect 14586 20659 14620 20663
rect 14664 20659 14698 20663
rect 14586 20647 14698 20659
rect 14620 20471 14664 20647
rect 14620 20459 14698 20471
rect 14664 20455 14698 20459
rect 14782 20647 14816 20663
rect 14782 20455 14816 20471
rect 17066 20647 17100 20663
rect 17066 20455 17100 20471
rect 17184 20659 17218 20663
rect 17258 20659 17292 20663
rect 17184 20647 17292 20659
rect 17218 20471 17258 20647
rect 17184 20459 17258 20471
rect 17184 20455 17218 20459
rect 14586 20255 14620 20271
rect 17258 20255 17292 20271
rect 17376 20647 17410 20663
rect 17376 20255 17410 20271
rect 17494 20647 17528 20663
rect 17494 20255 17528 20271
rect 17612 20647 17646 20663
rect 17612 20255 17646 20271
rect 17730 20659 17764 20663
rect 17808 20659 17842 20663
rect 17730 20647 17842 20659
rect 17764 20471 17808 20647
rect 17764 20459 17842 20471
rect 17808 20455 17842 20459
rect 17926 20647 17960 20663
rect 17926 20455 17960 20471
rect 20198 20651 20232 20667
rect 20198 20459 20232 20475
rect 20316 20663 20350 20667
rect 20390 20663 20424 20667
rect 20316 20651 20424 20663
rect 20350 20475 20390 20651
rect 20316 20463 20390 20475
rect 20316 20459 20350 20463
rect 17730 20255 17764 20271
rect 20390 20259 20424 20275
rect 20508 20651 20542 20667
rect 20508 20259 20542 20275
rect 20626 20651 20660 20667
rect 20626 20259 20660 20275
rect 20744 20651 20778 20667
rect 20744 20259 20778 20275
rect 20862 20663 20896 20667
rect 20940 20663 20974 20667
rect 20862 20651 20974 20663
rect 20896 20475 20940 20651
rect 20896 20463 20974 20475
rect 20940 20459 20974 20463
rect 21058 20651 21092 20667
rect 21058 20459 21092 20475
rect 23342 20651 23376 20667
rect 23342 20459 23376 20475
rect 23460 20663 23494 20667
rect 23534 20663 23568 20667
rect 23460 20651 23568 20663
rect 23494 20475 23534 20651
rect 23460 20463 23534 20475
rect 23460 20459 23494 20463
rect 20862 20259 20896 20275
rect 23534 20259 23568 20275
rect 23652 20651 23686 20667
rect 23652 20259 23686 20275
rect 23770 20651 23804 20667
rect 23770 20259 23804 20275
rect 23888 20651 23922 20667
rect 23888 20259 23922 20275
rect 24006 20663 24040 20667
rect 24084 20663 24118 20667
rect 24006 20651 24118 20663
rect 24040 20475 24084 20651
rect 24040 20463 24118 20475
rect 24084 20459 24118 20463
rect 24202 20651 24236 20667
rect 24202 20459 24236 20475
rect 24006 20259 24040 20275
rect 1713 20136 1729 20170
rect 1763 20136 1779 20170
rect 4857 20136 4873 20170
rect 4907 20136 4923 20170
rect 7989 20140 8005 20174
rect 8039 20140 8055 20174
rect 11133 20140 11149 20174
rect 11183 20140 11199 20174
rect 14335 20136 14351 20170
rect 14385 20136 14401 20170
rect 17479 20136 17495 20170
rect 17529 20136 17545 20170
rect 20611 20140 20627 20174
rect 20661 20140 20677 20174
rect 23755 20140 23771 20174
rect 23805 20140 23821 20174
rect 7970 20022 8106 20026
rect 1694 20018 1830 20022
rect 1694 20004 1732 20018
rect 1790 20004 1830 20018
rect 1694 19958 1710 20004
rect 1814 19958 1830 20004
rect 1694 19936 1830 19958
rect 4838 20018 4974 20022
rect 4838 20004 4876 20018
rect 4934 20004 4974 20018
rect 4838 19958 4854 20004
rect 4958 19958 4974 20004
rect 4838 19936 4974 19958
rect 7970 20008 8008 20022
rect 8066 20008 8106 20022
rect 7970 19962 7986 20008
rect 8090 19962 8106 20008
rect 7970 19940 8106 19962
rect 11114 20022 11250 20026
rect 20592 20022 20728 20026
rect 11114 20008 11152 20022
rect 11210 20008 11250 20022
rect 11114 19962 11130 20008
rect 11234 19962 11250 20008
rect 11114 19940 11250 19962
rect 14316 20018 14452 20022
rect 14316 20004 14354 20018
rect 14412 20004 14452 20018
rect 14316 19958 14332 20004
rect 14436 19958 14452 20004
rect 14316 19936 14452 19958
rect 17460 20018 17596 20022
rect 17460 20004 17498 20018
rect 17556 20004 17596 20018
rect 17460 19958 17476 20004
rect 17580 19958 17596 20004
rect 17460 19936 17596 19958
rect 20592 20008 20630 20022
rect 20688 20008 20728 20022
rect 20592 19962 20608 20008
rect 20712 19962 20728 20008
rect 20592 19940 20728 19962
rect 23736 20022 23872 20026
rect 23736 20008 23774 20022
rect 23832 20008 23872 20022
rect 23736 19962 23752 20008
rect 23856 19962 23872 20008
rect 23736 19940 23872 19962
rect 15168 17046 15372 17058
rect 15168 16974 15200 17046
rect 15344 16974 15372 17046
rect 15168 16972 15230 16974
rect 15310 16972 15372 16974
rect 14566 16934 14582 16968
rect 14616 16934 14632 16968
rect 15168 16956 15372 16972
rect 16336 17046 16540 17058
rect 16336 16974 16368 17046
rect 16512 16974 16540 17046
rect 16336 16972 16398 16974
rect 16478 16972 16540 16974
rect 15734 16934 15750 16968
rect 15784 16934 15800 16968
rect 16336 16956 16540 16972
rect 17504 17046 17708 17058
rect 17504 16974 17536 17046
rect 17680 16974 17708 17046
rect 17504 16972 17566 16974
rect 17646 16972 17708 16974
rect 16902 16934 16918 16968
rect 16952 16934 16968 16968
rect 17504 16956 17708 16972
rect 18672 17046 18876 17058
rect 18672 16974 18704 17046
rect 18848 16974 18876 17046
rect 18672 16972 18734 16974
rect 18814 16972 18876 16974
rect 18070 16934 18086 16968
rect 18120 16934 18136 16968
rect 18672 16956 18876 16972
rect 19846 17048 20050 17060
rect 19846 16976 19878 17048
rect 20022 16976 20050 17048
rect 19846 16974 19908 16976
rect 19988 16974 20050 16976
rect 19244 16936 19260 16970
rect 19294 16936 19310 16970
rect 19846 16958 20050 16974
rect 21014 17048 21218 17060
rect 21014 16976 21046 17048
rect 21190 16976 21218 17048
rect 21014 16974 21076 16976
rect 21156 16974 21218 16976
rect 20412 16936 20428 16970
rect 20462 16936 20478 16970
rect 21014 16958 21218 16974
rect 22182 17048 22386 17060
rect 22182 16976 22214 17048
rect 22358 16976 22386 17048
rect 22182 16974 22244 16976
rect 22324 16974 22386 16976
rect 21580 16936 21596 16970
rect 21630 16936 21646 16970
rect 22182 16958 22386 16974
rect 23350 17048 23554 17060
rect 23350 16976 23382 17048
rect 23526 16976 23554 17048
rect 23350 16974 23412 16976
rect 23492 16974 23554 16976
rect 22748 16936 22764 16970
rect 22798 16936 22814 16970
rect 23350 16958 23554 16974
rect 3198 16839 3366 16855
rect 3198 16769 3214 16839
rect 3350 16769 3366 16839
rect 3198 16753 3366 16769
rect 4646 16839 4814 16855
rect 4646 16769 4662 16839
rect 4798 16769 4814 16839
rect 4646 16753 4814 16769
rect 6144 16841 6312 16857
rect 6144 16771 6160 16841
rect 6296 16771 6312 16841
rect 6144 16755 6312 16771
rect 7592 16841 7760 16857
rect 7592 16771 7608 16841
rect 7744 16771 7760 16841
rect 7592 16755 7760 16771
rect 9112 16839 9280 16855
rect 9112 16769 9128 16839
rect 9264 16769 9280 16839
rect 9112 16753 9280 16769
rect 10560 16839 10728 16855
rect 10560 16769 10576 16839
rect 10712 16769 10728 16839
rect 10560 16753 10728 16769
rect 12058 16841 12226 16857
rect 12058 16771 12074 16841
rect 12210 16771 12226 16841
rect 12058 16755 12226 16771
rect 13506 16841 13674 16857
rect 13506 16771 13522 16841
rect 13658 16771 13674 16841
rect 14566 16826 14582 16860
rect 14616 16826 14632 16860
rect 15734 16826 15750 16860
rect 15784 16826 15800 16860
rect 16902 16826 16918 16860
rect 16952 16826 16968 16860
rect 18070 16826 18086 16860
rect 18120 16826 18136 16860
rect 19244 16828 19260 16862
rect 19294 16828 19310 16862
rect 20412 16828 20428 16862
rect 20462 16828 20478 16862
rect 21580 16828 21596 16862
rect 21630 16828 21646 16862
rect 22748 16828 22764 16862
rect 22798 16828 22814 16862
rect 13506 16755 13674 16771
rect 14672 16796 14706 16812
rect 3735 16649 4005 16683
rect 2909 16599 2943 16615
rect 2909 16407 2943 16423
rect 3027 16599 3061 16615
rect 3027 16407 3061 16423
rect 3145 16599 3179 16615
rect 3145 16407 3179 16423
rect 3263 16599 3297 16615
rect 3263 16407 3297 16423
rect 3381 16599 3415 16615
rect 3381 16407 3415 16423
rect 3499 16599 3533 16615
rect 3499 16407 3533 16423
rect 3617 16599 3651 16615
rect 3617 16407 3651 16423
rect 3735 16599 3769 16649
rect 3735 16407 3769 16423
rect 3853 16599 3887 16615
rect 3853 16407 3887 16423
rect 3971 16599 4005 16649
rect 5183 16649 5453 16683
rect 3971 16407 4005 16423
rect 4357 16599 4391 16615
rect 4357 16407 4391 16423
rect 4475 16599 4509 16615
rect 4475 16407 4509 16423
rect 4593 16599 4627 16615
rect 4593 16407 4627 16423
rect 4711 16599 4745 16615
rect 4711 16407 4745 16423
rect 4829 16599 4863 16615
rect 4829 16407 4863 16423
rect 4947 16599 4981 16615
rect 4947 16407 4981 16423
rect 5065 16599 5099 16615
rect 5065 16407 5099 16423
rect 5183 16599 5217 16649
rect 5183 16407 5217 16423
rect 5301 16599 5335 16615
rect 5301 16407 5335 16423
rect 5419 16599 5453 16649
rect 6681 16651 6951 16685
rect 5419 16407 5453 16423
rect 5855 16601 5889 16617
rect 5855 16409 5889 16425
rect 5973 16601 6007 16617
rect 5973 16409 6007 16425
rect 6091 16601 6125 16617
rect 6091 16409 6125 16425
rect 6209 16601 6243 16617
rect 6209 16409 6243 16425
rect 6327 16601 6361 16617
rect 6327 16409 6361 16425
rect 6445 16601 6479 16617
rect 6445 16409 6479 16425
rect 6563 16601 6597 16617
rect 6563 16409 6597 16425
rect 6681 16601 6715 16651
rect 6681 16409 6715 16425
rect 6799 16601 6833 16617
rect 6799 16409 6833 16425
rect 6917 16601 6951 16651
rect 8129 16651 8399 16685
rect 6917 16409 6951 16425
rect 7303 16601 7337 16617
rect 7303 16409 7337 16425
rect 7421 16601 7455 16617
rect 7421 16409 7455 16425
rect 7539 16601 7573 16617
rect 7539 16409 7573 16425
rect 7657 16601 7691 16617
rect 7657 16409 7691 16425
rect 7775 16601 7809 16617
rect 7775 16409 7809 16425
rect 7893 16601 7927 16617
rect 7893 16409 7927 16425
rect 8011 16601 8045 16617
rect 8011 16409 8045 16425
rect 8129 16601 8163 16651
rect 8129 16409 8163 16425
rect 8247 16601 8281 16617
rect 8247 16409 8281 16425
rect 8365 16601 8399 16651
rect 9649 16649 9919 16683
rect 8365 16409 8399 16425
rect 8823 16599 8857 16615
rect 8823 16407 8857 16423
rect 8941 16599 8975 16615
rect 8941 16407 8975 16423
rect 9059 16599 9093 16615
rect 9059 16407 9093 16423
rect 9177 16599 9211 16615
rect 9177 16407 9211 16423
rect 9295 16599 9329 16615
rect 9295 16407 9329 16423
rect 9413 16599 9447 16615
rect 9413 16407 9447 16423
rect 9531 16599 9565 16615
rect 9531 16407 9565 16423
rect 9649 16599 9683 16649
rect 9649 16407 9683 16423
rect 9767 16599 9801 16615
rect 9767 16407 9801 16423
rect 9885 16599 9919 16649
rect 11097 16649 11367 16683
rect 9885 16407 9919 16423
rect 10271 16599 10305 16615
rect 10271 16407 10305 16423
rect 10389 16599 10423 16615
rect 10389 16407 10423 16423
rect 10507 16599 10541 16615
rect 10507 16407 10541 16423
rect 10625 16599 10659 16615
rect 10625 16407 10659 16423
rect 10743 16599 10777 16615
rect 10743 16407 10777 16423
rect 10861 16599 10895 16615
rect 10861 16407 10895 16423
rect 10979 16599 11013 16615
rect 10979 16407 11013 16423
rect 11097 16599 11131 16649
rect 11097 16407 11131 16423
rect 11215 16599 11249 16615
rect 11215 16407 11249 16423
rect 11333 16599 11367 16649
rect 12595 16651 12865 16685
rect 11333 16407 11367 16423
rect 11769 16601 11803 16617
rect 11769 16409 11803 16425
rect 11887 16601 11921 16617
rect 11887 16409 11921 16425
rect 12005 16601 12039 16617
rect 12005 16409 12039 16425
rect 12123 16601 12157 16617
rect 12123 16409 12157 16425
rect 12241 16601 12275 16617
rect 12241 16409 12275 16425
rect 12359 16601 12393 16617
rect 12359 16409 12393 16425
rect 12477 16601 12511 16617
rect 12477 16409 12511 16425
rect 12595 16601 12629 16651
rect 12595 16409 12629 16425
rect 12713 16601 12747 16617
rect 12713 16409 12747 16425
rect 12831 16601 12865 16651
rect 14043 16651 14313 16685
rect 12831 16409 12865 16425
rect 13217 16601 13251 16617
rect 13217 16409 13251 16425
rect 13335 16601 13369 16617
rect 13335 16409 13369 16425
rect 13453 16601 13487 16617
rect 13453 16409 13487 16425
rect 13571 16601 13605 16617
rect 13571 16409 13605 16425
rect 13689 16601 13723 16617
rect 13689 16409 13723 16425
rect 13807 16601 13841 16617
rect 13807 16409 13841 16425
rect 13925 16601 13959 16617
rect 13925 16409 13959 16425
rect 14043 16601 14077 16651
rect 14043 16409 14077 16425
rect 14161 16601 14195 16617
rect 14161 16409 14195 16425
rect 14279 16601 14313 16651
rect 14279 16409 14313 16425
rect 14672 16404 14706 16420
rect 14790 16796 14824 16812
rect 14790 16404 14824 16420
rect 14908 16796 14942 16812
rect 14908 16404 14942 16420
rect 15026 16796 15060 16812
rect 15026 16404 15060 16420
rect 15144 16796 15178 16812
rect 15144 16404 15178 16420
rect 15262 16796 15296 16812
rect 15262 16404 15296 16420
rect 15380 16796 15414 16812
rect 15380 16404 15414 16420
rect 15840 16796 15874 16812
rect 15840 16404 15874 16420
rect 15958 16796 15992 16812
rect 15958 16404 15992 16420
rect 16076 16796 16110 16812
rect 16076 16404 16110 16420
rect 16194 16796 16228 16812
rect 16194 16404 16228 16420
rect 16312 16796 16346 16812
rect 16312 16404 16346 16420
rect 16430 16796 16464 16812
rect 16430 16404 16464 16420
rect 16548 16796 16582 16812
rect 16548 16404 16582 16420
rect 17008 16794 17042 16810
rect 17008 16402 17042 16418
rect 17126 16794 17160 16810
rect 17126 16402 17160 16418
rect 17244 16794 17278 16810
rect 17244 16402 17278 16418
rect 17362 16794 17396 16810
rect 17362 16402 17396 16418
rect 17480 16794 17514 16810
rect 17480 16402 17514 16418
rect 17598 16794 17632 16810
rect 17598 16402 17632 16418
rect 17716 16794 17750 16810
rect 17716 16402 17750 16418
rect 18176 16796 18210 16812
rect 18176 16404 18210 16420
rect 18294 16796 18328 16812
rect 18294 16404 18328 16420
rect 18412 16796 18446 16812
rect 18412 16404 18446 16420
rect 18530 16796 18564 16812
rect 18530 16404 18564 16420
rect 18648 16796 18682 16812
rect 18648 16404 18682 16420
rect 18766 16796 18800 16812
rect 18766 16404 18800 16420
rect 18884 16796 18918 16812
rect 18884 16404 18918 16420
rect 19350 16798 19384 16814
rect 19350 16406 19384 16422
rect 19468 16798 19502 16814
rect 19468 16406 19502 16422
rect 19586 16798 19620 16814
rect 19586 16406 19620 16422
rect 19704 16798 19738 16814
rect 19704 16406 19738 16422
rect 19822 16798 19856 16814
rect 19822 16406 19856 16422
rect 19940 16798 19974 16814
rect 19940 16406 19974 16422
rect 20058 16798 20092 16814
rect 20058 16406 20092 16422
rect 20518 16796 20552 16812
rect 20518 16404 20552 16420
rect 20636 16796 20670 16812
rect 20636 16404 20670 16420
rect 20754 16796 20788 16812
rect 20754 16404 20788 16420
rect 20872 16796 20906 16812
rect 20872 16404 20906 16420
rect 20990 16796 21024 16812
rect 20990 16404 21024 16420
rect 21108 16796 21142 16812
rect 21108 16404 21142 16420
rect 21226 16796 21260 16812
rect 21226 16404 21260 16420
rect 21686 16798 21720 16814
rect 21686 16406 21720 16422
rect 21804 16798 21838 16814
rect 21804 16406 21838 16422
rect 21922 16798 21956 16814
rect 21922 16406 21956 16422
rect 22040 16798 22074 16814
rect 22040 16406 22074 16422
rect 22158 16798 22192 16814
rect 22158 16406 22192 16422
rect 22276 16798 22310 16814
rect 22276 16406 22310 16422
rect 22394 16798 22428 16814
rect 22394 16406 22428 16422
rect 22854 16796 22888 16812
rect 22854 16404 22888 16420
rect 22972 16796 23006 16812
rect 22972 16404 23006 16420
rect 23090 16796 23124 16812
rect 23090 16404 23124 16420
rect 23208 16796 23242 16812
rect 23208 16404 23242 16420
rect 23326 16796 23360 16812
rect 23326 16404 23360 16420
rect 23444 16796 23478 16812
rect 23444 16404 23478 16420
rect 23562 16796 23596 16812
rect 23562 16404 23596 16420
rect 3660 16329 3676 16363
rect 3710 16329 3726 16363
rect 5108 16329 5124 16363
rect 5158 16329 5174 16363
rect 6606 16331 6622 16365
rect 6656 16331 6672 16365
rect 8054 16331 8070 16365
rect 8104 16331 8120 16365
rect 9574 16329 9590 16363
rect 9624 16329 9640 16363
rect 11022 16329 11038 16363
rect 11072 16329 11088 16363
rect 12520 16331 12536 16365
rect 12570 16331 12586 16365
rect 13968 16331 13984 16365
rect 14018 16331 14034 16365
rect 3542 16212 3558 16246
rect 3592 16212 3608 16246
rect 4990 16212 5006 16246
rect 5040 16212 5056 16246
rect 6488 16214 6504 16248
rect 6538 16214 6554 16248
rect 7936 16214 7952 16248
rect 7986 16214 8002 16248
rect 9456 16212 9472 16246
rect 9506 16212 9522 16246
rect 10904 16212 10920 16246
rect 10954 16212 10970 16246
rect 12402 16214 12418 16248
rect 12452 16214 12468 16248
rect 13850 16214 13866 16248
rect 13900 16214 13916 16248
rect 3146 16162 3180 16178
rect 3146 15770 3180 15786
rect 3264 16162 3298 16178
rect 3264 15770 3298 15786
rect 3382 16162 3416 16178
rect 3499 16162 3533 16178
rect 3499 15970 3533 15986
rect 3617 16162 3651 16178
rect 3617 15970 3651 15986
rect 4594 16162 4628 16178
rect 3382 15770 3416 15786
rect 4594 15770 4628 15786
rect 4712 16162 4746 16178
rect 4712 15770 4746 15786
rect 4830 16162 4864 16178
rect 4947 16162 4981 16178
rect 4947 15970 4981 15986
rect 5065 16162 5099 16178
rect 5065 15970 5099 15986
rect 6092 16164 6126 16180
rect 4830 15770 4864 15786
rect 6092 15772 6126 15788
rect 6210 16164 6244 16180
rect 6210 15772 6244 15788
rect 6328 16164 6362 16180
rect 6445 16164 6479 16180
rect 6445 15972 6479 15988
rect 6563 16164 6597 16180
rect 6563 15972 6597 15988
rect 7540 16164 7574 16180
rect 6328 15772 6362 15788
rect 7540 15772 7574 15788
rect 7658 16164 7692 16180
rect 7658 15772 7692 15788
rect 7776 16164 7810 16180
rect 7893 16164 7927 16180
rect 7893 15972 7927 15988
rect 8011 16164 8045 16180
rect 8011 15972 8045 15988
rect 9060 16162 9094 16178
rect 7776 15772 7810 15788
rect 9060 15770 9094 15786
rect 9178 16162 9212 16178
rect 9178 15770 9212 15786
rect 9296 16162 9330 16178
rect 9413 16162 9447 16178
rect 9413 15970 9447 15986
rect 9531 16162 9565 16178
rect 9531 15970 9565 15986
rect 10508 16162 10542 16178
rect 9296 15770 9330 15786
rect 10508 15770 10542 15786
rect 10626 16162 10660 16178
rect 10626 15770 10660 15786
rect 10744 16162 10778 16178
rect 10861 16162 10895 16178
rect 10861 15970 10895 15986
rect 10979 16162 11013 16178
rect 10979 15970 11013 15986
rect 12006 16164 12040 16180
rect 10744 15770 10778 15786
rect 12006 15772 12040 15788
rect 12124 16164 12158 16180
rect 12124 15772 12158 15788
rect 12242 16164 12276 16180
rect 12359 16164 12393 16180
rect 12359 15972 12393 15988
rect 12477 16164 12511 16180
rect 12477 15972 12511 15988
rect 13454 16164 13488 16180
rect 12242 15772 12276 15788
rect 13454 15772 13488 15788
rect 13572 16164 13606 16180
rect 13572 15772 13606 15788
rect 13690 16164 13724 16180
rect 13807 16164 13841 16180
rect 13807 15972 13841 15988
rect 13925 16164 13959 16180
rect 17956 16134 18756 16168
rect 14861 16063 14877 16097
rect 14911 16063 14927 16097
rect 16029 16063 16045 16097
rect 16079 16063 16095 16097
rect 17197 16063 17213 16097
rect 17247 16063 17263 16097
rect 13925 15972 13959 15988
rect 14582 16010 14616 16026
rect 14582 15818 14616 15834
rect 14700 16010 14734 16026
rect 14700 15818 14734 15834
rect 14818 16010 14852 16026
rect 14818 15818 14852 15834
rect 14936 16010 14970 16026
rect 14936 15818 14970 15834
rect 15102 16006 15136 16022
rect 13690 15772 13724 15788
rect 3189 15702 3205 15736
rect 3239 15702 3255 15736
rect 3307 15702 3323 15736
rect 3357 15702 3373 15736
rect 4637 15702 4653 15736
rect 4687 15702 4703 15736
rect 4755 15702 4771 15736
rect 4805 15702 4821 15736
rect 6135 15704 6151 15738
rect 6185 15704 6201 15738
rect 6253 15704 6269 15738
rect 6303 15704 6319 15738
rect 7583 15704 7599 15738
rect 7633 15704 7649 15738
rect 7701 15704 7717 15738
rect 7751 15704 7767 15738
rect 9103 15702 9119 15736
rect 9153 15702 9169 15736
rect 9221 15702 9237 15736
rect 9271 15702 9287 15736
rect 10551 15702 10567 15736
rect 10601 15702 10617 15736
rect 10669 15702 10685 15736
rect 10719 15702 10735 15736
rect 12049 15704 12065 15738
rect 12099 15704 12115 15738
rect 12167 15704 12183 15738
rect 12217 15704 12233 15738
rect 13497 15704 13513 15738
rect 13547 15704 13563 15738
rect 13615 15704 13631 15738
rect 13665 15704 13681 15738
rect 15102 15730 15136 15830
rect 15220 16006 15254 16022
rect 15220 15814 15254 15830
rect 15338 16006 15372 16022
rect 15338 15730 15372 15830
rect 15456 16006 15490 16022
rect 15456 15814 15490 15830
rect 15750 16012 15784 16028
rect 15750 15820 15784 15836
rect 15868 16012 15902 16028
rect 15868 15820 15902 15836
rect 15986 16012 16020 16028
rect 15986 15820 16020 15836
rect 16104 16012 16138 16028
rect 16104 15820 16138 15836
rect 16269 16012 16303 16028
rect 14726 15706 14868 15718
rect 14726 15702 14766 15706
rect 14832 15702 14868 15706
rect 3422 15631 3590 15649
rect 3422 15575 3438 15631
rect 3572 15575 3590 15631
rect 3422 15559 3590 15575
rect 4870 15631 5038 15649
rect 4870 15575 4886 15631
rect 5020 15575 5038 15631
rect 4870 15559 5038 15575
rect 6368 15633 6536 15651
rect 6368 15577 6384 15633
rect 6518 15577 6536 15633
rect 6368 15561 6536 15577
rect 7816 15633 7984 15651
rect 7816 15577 7832 15633
rect 7966 15577 7984 15633
rect 7816 15561 7984 15577
rect 9336 15631 9504 15649
rect 9336 15575 9352 15631
rect 9486 15575 9504 15631
rect 9336 15559 9504 15575
rect 10784 15631 10952 15649
rect 10784 15575 10800 15631
rect 10934 15575 10952 15631
rect 10784 15559 10952 15575
rect 12282 15633 12450 15651
rect 12282 15577 12298 15633
rect 12432 15577 12450 15633
rect 12282 15561 12450 15577
rect 13730 15633 13898 15651
rect 13730 15577 13746 15633
rect 13880 15577 13898 15633
rect 14726 15636 14744 15702
rect 14862 15636 14868 15702
rect 15102 15696 15372 15730
rect 16269 15742 16303 15836
rect 16387 16012 16421 16028
rect 16387 15820 16421 15836
rect 16505 16012 16539 16028
rect 16505 15742 16539 15836
rect 16623 16012 16657 16028
rect 16623 15820 16657 15836
rect 16918 16012 16952 16028
rect 16918 15820 16952 15836
rect 17036 16012 17070 16028
rect 17036 15820 17070 15836
rect 17154 16012 17188 16028
rect 17154 15820 17188 15836
rect 17272 16012 17306 16028
rect 17272 15820 17306 15836
rect 17437 16012 17471 16028
rect 15894 15706 16036 15718
rect 16269 15708 16539 15742
rect 17437 15725 17471 15836
rect 17555 16012 17589 16028
rect 17555 15820 17589 15836
rect 17673 16012 17707 16028
rect 17673 15725 17707 15836
rect 17791 16012 17825 16028
rect 17791 15820 17825 15836
rect 15894 15702 15934 15706
rect 16000 15702 16036 15706
rect 14726 15610 14868 15636
rect 13730 15561 13898 15577
rect 15194 15523 15239 15696
rect 15894 15636 15912 15702
rect 16030 15636 16036 15702
rect 15894 15610 16036 15636
rect 2574 15469 15239 15523
rect 2574 14322 2666 15469
rect 16387 15435 16421 15708
rect 17062 15706 17204 15718
rect 17062 15702 17102 15706
rect 17168 15702 17204 15706
rect 17062 15636 17080 15702
rect 17198 15636 17204 15702
rect 17437 15689 17707 15725
rect 17062 15610 17204 15636
rect 5797 15381 16421 15435
rect 4138 15112 4366 15130
rect 4138 15036 4154 15112
rect 4350 15036 4366 15112
rect 4138 15020 4366 15036
rect 3409 14895 3679 14934
rect 3409 14842 3443 14895
rect 2968 14693 3238 14732
rect 2968 14642 3002 14693
rect 2968 14450 3002 14466
rect 3086 14642 3120 14658
rect 3086 14415 3120 14466
rect 3204 14642 3238 14693
rect 3204 14450 3238 14466
rect 3322 14642 3356 14658
rect 3322 14415 3356 14466
rect 3409 14450 3443 14466
rect 3527 14842 3561 14858
rect 3086 14376 3356 14415
rect 3527 14415 3561 14466
rect 3645 14842 3679 14895
rect 3876 14894 4146 14933
rect 3645 14450 3679 14466
rect 3763 14842 3797 14858
rect 3763 14415 3797 14466
rect 3876 14842 3910 14894
rect 3876 14450 3910 14466
rect 3994 14842 4028 14858
rect 3994 14415 4028 14466
rect 4112 14842 4146 14894
rect 4348 14894 4618 14933
rect 4112 14450 4146 14466
rect 4230 14842 4264 14858
rect 4230 14415 4264 14466
rect 4348 14842 4382 14894
rect 4348 14450 4382 14466
rect 4466 14842 4500 14858
rect 4466 14415 4500 14466
rect 4584 14842 4618 14894
rect 4821 14894 5091 14933
rect 4584 14450 4618 14466
rect 4703 14842 4737 14858
rect 4703 14415 4737 14466
rect 4821 14842 4855 14894
rect 4821 14450 4855 14466
rect 4939 14842 4973 14858
rect 4939 14415 4973 14466
rect 5057 14842 5091 14894
rect 5294 14692 5564 14729
rect 5057 14450 5091 14466
rect 5176 14642 5210 14658
rect 3527 14376 4973 14415
rect 5176 14412 5210 14466
rect 5294 14642 5328 14692
rect 5294 14450 5328 14466
rect 5412 14642 5446 14658
rect 5412 14412 5446 14466
rect 5530 14642 5564 14692
rect 5530 14450 5564 14466
rect 5176 14373 5446 14412
rect 2574 13881 2667 14322
rect 4054 14251 4088 14267
rect 5348 14258 5364 14292
rect 5398 14258 5414 14292
rect 4054 14201 4088 14217
rect 3057 14151 3149 14168
rect 3057 14096 3073 14151
rect 3133 14096 3149 14151
rect 3057 14083 3149 14096
rect 4142 14152 4234 14165
rect 4142 14097 4158 14152
rect 4218 14097 4234 14152
rect 4142 14080 4234 14097
rect 2825 14036 2882 14040
rect 2825 13976 2829 14036
rect 2878 13976 2882 14036
rect 2825 13972 2882 13976
rect 4408 14021 4442 14037
rect 4408 13971 4442 13987
rect 2574 13868 2885 13881
rect 2574 13808 2829 13868
rect 2878 13808 2885 13868
rect 2574 13795 2885 13808
rect 4024 13867 4116 13880
rect 4024 13812 4040 13867
rect 4100 13812 4116 13867
rect 4024 13795 4116 13812
rect 5797 13872 5875 15381
rect 17523 15347 17572 15689
rect 8921 15299 17572 15347
rect 7282 15112 7510 15130
rect 7282 15036 7298 15112
rect 7494 15036 7510 15112
rect 7282 15020 7510 15036
rect 6553 14895 6823 14934
rect 6553 14842 6587 14895
rect 6112 14693 6382 14732
rect 6112 14642 6146 14693
rect 6112 14450 6146 14466
rect 6230 14642 6264 14658
rect 6230 14415 6264 14466
rect 6348 14642 6382 14693
rect 6348 14450 6382 14466
rect 6466 14642 6500 14658
rect 6466 14415 6500 14466
rect 6553 14450 6587 14466
rect 6671 14842 6705 14858
rect 6230 14376 6500 14415
rect 6671 14415 6705 14466
rect 6789 14842 6823 14895
rect 7020 14894 7290 14933
rect 6789 14450 6823 14466
rect 6907 14842 6941 14858
rect 6907 14415 6941 14466
rect 7020 14842 7054 14894
rect 7020 14450 7054 14466
rect 7138 14842 7172 14858
rect 7138 14415 7172 14466
rect 7256 14842 7290 14894
rect 7492 14894 7762 14933
rect 7256 14450 7290 14466
rect 7374 14842 7408 14858
rect 7374 14415 7408 14466
rect 7492 14842 7526 14894
rect 7492 14450 7526 14466
rect 7610 14842 7644 14858
rect 7610 14415 7644 14466
rect 7728 14842 7762 14894
rect 7965 14894 8235 14933
rect 7728 14450 7762 14466
rect 7847 14842 7881 14858
rect 7847 14415 7881 14466
rect 7965 14842 7999 14894
rect 7965 14450 7999 14466
rect 8083 14842 8117 14858
rect 8083 14415 8117 14466
rect 8201 14842 8235 14894
rect 8438 14692 8708 14729
rect 8201 14450 8235 14466
rect 8320 14642 8354 14658
rect 6671 14376 8117 14415
rect 8320 14412 8354 14466
rect 8438 14642 8472 14692
rect 8438 14450 8472 14466
rect 8556 14642 8590 14658
rect 8556 14412 8590 14466
rect 8674 14642 8708 14692
rect 8674 14450 8708 14466
rect 8320 14373 8590 14412
rect 7198 14251 7232 14267
rect 8492 14258 8508 14292
rect 8542 14258 8558 14292
rect 7198 14201 7232 14217
rect 6201 14151 6293 14168
rect 6201 14096 6217 14151
rect 6277 14096 6293 14151
rect 6201 14083 6293 14096
rect 7286 14152 7378 14165
rect 7286 14097 7302 14152
rect 7362 14097 7378 14152
rect 7286 14080 7378 14097
rect 5969 14036 6026 14040
rect 5969 13976 5973 14036
rect 6022 13976 6026 14036
rect 5969 13972 6026 13976
rect 7552 14021 7586 14037
rect 7552 13971 7586 13987
rect 5797 13868 6026 13872
rect 5797 13808 5973 13868
rect 6022 13808 6026 13868
rect 5797 13804 6026 13808
rect 7168 13867 7260 13880
rect 7168 13812 7184 13867
rect 7244 13812 7260 13867
rect 7168 13795 7260 13812
rect 8921 13876 8989 15299
rect 17956 15265 18029 16134
rect 18365 16063 18381 16097
rect 18415 16063 18431 16097
rect 18722 16096 18756 16134
rect 18606 16062 18876 16096
rect 19539 16065 19555 16099
rect 19589 16065 19605 16099
rect 20707 16065 20723 16099
rect 20757 16065 20773 16099
rect 21875 16065 21891 16099
rect 21925 16065 21941 16099
rect 23043 16065 23059 16099
rect 23093 16065 23109 16099
rect 18086 16012 18120 16028
rect 18086 15820 18120 15836
rect 18204 16012 18238 16028
rect 18204 15820 18238 15836
rect 18322 16012 18356 16028
rect 18322 15820 18356 15836
rect 18440 16012 18474 16028
rect 18440 15820 18474 15836
rect 18606 16012 18640 16062
rect 18606 15820 18640 15836
rect 18724 16012 18758 16028
rect 18724 15820 18758 15836
rect 18842 16012 18876 16062
rect 18842 15820 18876 15836
rect 18960 16012 18994 16028
rect 18960 15820 18994 15836
rect 19260 16012 19294 16028
rect 19260 15820 19294 15836
rect 19378 16012 19412 16028
rect 19378 15820 19412 15836
rect 19496 16012 19530 16028
rect 19496 15820 19530 15836
rect 19614 16012 19648 16028
rect 19614 15820 19648 15836
rect 19778 16008 19812 16024
rect 19778 15732 19812 15832
rect 19896 16008 19930 16024
rect 19896 15816 19930 15832
rect 20014 16008 20048 16024
rect 20014 15732 20048 15832
rect 20132 16008 20166 16024
rect 20132 15816 20166 15832
rect 20428 16012 20462 16028
rect 20428 15820 20462 15836
rect 20546 16012 20580 16028
rect 20546 15820 20580 15836
rect 20664 16012 20698 16028
rect 20664 15820 20698 15836
rect 20782 16012 20816 16028
rect 20782 15820 20816 15836
rect 20947 16007 20981 16023
rect 18230 15706 18372 15718
rect 18230 15702 18270 15706
rect 18336 15702 18372 15706
rect 18230 15636 18248 15702
rect 18366 15636 18372 15702
rect 18230 15610 18372 15636
rect 19404 15708 19546 15720
rect 19404 15704 19444 15708
rect 19510 15704 19546 15708
rect 19404 15638 19422 15704
rect 19540 15638 19546 15704
rect 19778 15697 20048 15732
rect 20947 15746 20981 15831
rect 21065 16007 21099 16023
rect 21065 15815 21099 15831
rect 21183 16007 21217 16023
rect 21183 15746 21217 15831
rect 21301 16007 21335 16023
rect 21301 15815 21335 15831
rect 21596 16014 21630 16030
rect 21596 15822 21630 15838
rect 21714 16014 21748 16030
rect 21714 15822 21748 15838
rect 21832 16014 21866 16030
rect 21832 15822 21866 15838
rect 21950 16014 21984 16030
rect 21950 15822 21984 15838
rect 22115 16007 22149 16023
rect 20572 15708 20714 15720
rect 20947 15711 21217 15746
rect 22115 15746 22149 15831
rect 22233 16007 22267 16023
rect 22233 15815 22267 15831
rect 22351 16007 22385 16023
rect 22351 15746 22385 15831
rect 22469 16007 22503 16023
rect 22469 15815 22503 15831
rect 22764 16014 22798 16030
rect 22764 15822 22798 15838
rect 22882 16014 22916 16030
rect 22882 15822 22916 15838
rect 23000 16014 23034 16030
rect 23000 15822 23034 15838
rect 23118 16014 23152 16030
rect 23118 15822 23152 15838
rect 23283 16008 23317 16024
rect 20572 15704 20612 15708
rect 20678 15704 20714 15708
rect 19404 15612 19546 15638
rect 19900 15464 19958 15697
rect 20572 15638 20590 15704
rect 20708 15638 20714 15704
rect 20572 15612 20714 15638
rect 15037 15211 18029 15265
rect 18249 15405 19958 15464
rect 10414 15116 10642 15134
rect 10414 15040 10430 15116
rect 10626 15040 10642 15116
rect 10414 15024 10642 15040
rect 13558 15116 13786 15134
rect 13558 15040 13574 15116
rect 13770 15040 13786 15116
rect 13558 15024 13786 15040
rect 9685 14899 9955 14938
rect 9685 14846 9719 14899
rect 9244 14697 9514 14736
rect 9244 14646 9278 14697
rect 9244 14454 9278 14470
rect 9362 14646 9396 14662
rect 9362 14419 9396 14470
rect 9480 14646 9514 14697
rect 9480 14454 9514 14470
rect 9598 14646 9632 14662
rect 9598 14419 9632 14470
rect 9685 14454 9719 14470
rect 9803 14846 9837 14862
rect 9362 14380 9632 14419
rect 9803 14419 9837 14470
rect 9921 14846 9955 14899
rect 10152 14898 10422 14937
rect 9921 14454 9955 14470
rect 10039 14846 10073 14862
rect 10039 14419 10073 14470
rect 10152 14846 10186 14898
rect 10152 14454 10186 14470
rect 10270 14846 10304 14862
rect 10270 14419 10304 14470
rect 10388 14846 10422 14898
rect 10624 14898 10894 14937
rect 10388 14454 10422 14470
rect 10506 14846 10540 14862
rect 10506 14419 10540 14470
rect 10624 14846 10658 14898
rect 10624 14454 10658 14470
rect 10742 14846 10776 14862
rect 10742 14419 10776 14470
rect 10860 14846 10894 14898
rect 11097 14898 11367 14937
rect 10860 14454 10894 14470
rect 10979 14846 11013 14862
rect 10979 14419 11013 14470
rect 11097 14846 11131 14898
rect 11097 14454 11131 14470
rect 11215 14846 11249 14862
rect 11215 14419 11249 14470
rect 11333 14846 11367 14898
rect 12829 14899 13099 14938
rect 12829 14846 12863 14899
rect 11570 14696 11840 14733
rect 11333 14454 11367 14470
rect 11452 14646 11486 14662
rect 9803 14380 11249 14419
rect 11452 14416 11486 14470
rect 11570 14646 11604 14696
rect 11570 14454 11604 14470
rect 11688 14646 11722 14662
rect 11688 14416 11722 14470
rect 11806 14646 11840 14696
rect 11806 14454 11840 14470
rect 12388 14697 12658 14736
rect 12388 14646 12422 14697
rect 12388 14454 12422 14470
rect 12506 14646 12540 14662
rect 11452 14377 11722 14416
rect 12506 14419 12540 14470
rect 12624 14646 12658 14697
rect 12624 14454 12658 14470
rect 12742 14646 12776 14662
rect 12742 14419 12776 14470
rect 12829 14454 12863 14470
rect 12947 14846 12981 14862
rect 12506 14380 12776 14419
rect 12947 14419 12981 14470
rect 13065 14846 13099 14899
rect 13296 14898 13566 14937
rect 13065 14454 13099 14470
rect 13183 14846 13217 14862
rect 13183 14419 13217 14470
rect 13296 14846 13330 14898
rect 13296 14454 13330 14470
rect 13414 14846 13448 14862
rect 13414 14419 13448 14470
rect 13532 14846 13566 14898
rect 13768 14898 14038 14937
rect 13532 14454 13566 14470
rect 13650 14846 13684 14862
rect 13650 14419 13684 14470
rect 13768 14846 13802 14898
rect 13768 14454 13802 14470
rect 13886 14846 13920 14862
rect 13886 14419 13920 14470
rect 14004 14846 14038 14898
rect 14241 14898 14511 14937
rect 14004 14454 14038 14470
rect 14123 14846 14157 14862
rect 14123 14419 14157 14470
rect 14241 14846 14275 14898
rect 14241 14454 14275 14470
rect 14359 14846 14393 14862
rect 14359 14419 14393 14470
rect 14477 14846 14511 14898
rect 14714 14696 14984 14733
rect 14477 14454 14511 14470
rect 14596 14646 14630 14662
rect 12947 14380 14393 14419
rect 14596 14416 14630 14470
rect 14714 14646 14748 14696
rect 14714 14454 14748 14470
rect 14832 14646 14866 14662
rect 14832 14416 14866 14470
rect 14950 14646 14984 14696
rect 14950 14454 14984 14470
rect 14596 14377 14866 14416
rect 10330 14255 10364 14271
rect 11624 14262 11640 14296
rect 11674 14262 11690 14296
rect 10330 14205 10364 14221
rect 13474 14255 13508 14271
rect 14768 14262 14784 14296
rect 14818 14262 14834 14296
rect 13474 14205 13508 14221
rect 9333 14155 9425 14172
rect 9333 14100 9349 14155
rect 9409 14100 9425 14155
rect 9333 14087 9425 14100
rect 10418 14156 10510 14169
rect 10418 14101 10434 14156
rect 10494 14101 10510 14156
rect 10418 14084 10510 14101
rect 12477 14155 12569 14172
rect 12477 14100 12493 14155
rect 12553 14100 12569 14155
rect 12477 14087 12569 14100
rect 13562 14156 13654 14169
rect 13562 14101 13578 14156
rect 13638 14101 13654 14156
rect 13562 14084 13654 14101
rect 9101 14040 9158 14044
rect 9101 13980 9105 14040
rect 9154 13980 9158 14040
rect 9101 13976 9158 13980
rect 10684 14025 10718 14041
rect 10684 13975 10718 13991
rect 12245 14040 12302 14044
rect 12245 13980 12249 14040
rect 12298 13980 12302 14040
rect 12245 13976 12302 13980
rect 13828 14025 13862 14041
rect 13828 13975 13862 13991
rect 8921 13872 9159 13876
rect 8921 13812 9105 13872
rect 9154 13812 9159 13872
rect 8921 13807 9159 13812
rect 10300 13871 10392 13884
rect 10300 13816 10316 13871
rect 10376 13816 10392 13871
rect 10300 13799 10392 13816
rect 13444 13877 13536 13884
rect 15037 13877 15109 15211
rect 16760 15112 16988 15130
rect 16760 15036 16776 15112
rect 16972 15036 16988 15112
rect 16760 15020 16988 15036
rect 16031 14895 16301 14934
rect 16031 14842 16065 14895
rect 15590 14693 15860 14732
rect 15590 14642 15624 14693
rect 15590 14450 15624 14466
rect 15708 14642 15742 14658
rect 15708 14415 15742 14466
rect 15826 14642 15860 14693
rect 15826 14450 15860 14466
rect 15944 14642 15978 14658
rect 15944 14415 15978 14466
rect 16031 14450 16065 14466
rect 16149 14842 16183 14858
rect 15708 14376 15978 14415
rect 16149 14415 16183 14466
rect 16267 14842 16301 14895
rect 16498 14894 16768 14933
rect 16267 14450 16301 14466
rect 16385 14842 16419 14858
rect 16385 14415 16419 14466
rect 16498 14842 16532 14894
rect 16498 14450 16532 14466
rect 16616 14842 16650 14858
rect 16616 14415 16650 14466
rect 16734 14842 16768 14894
rect 16970 14894 17240 14933
rect 16734 14450 16768 14466
rect 16852 14842 16886 14858
rect 16852 14415 16886 14466
rect 16970 14842 17004 14894
rect 16970 14450 17004 14466
rect 17088 14842 17122 14858
rect 17088 14415 17122 14466
rect 17206 14842 17240 14894
rect 17443 14894 17713 14933
rect 17206 14450 17240 14466
rect 17325 14842 17359 14858
rect 17325 14415 17359 14466
rect 17443 14842 17477 14894
rect 17443 14450 17477 14466
rect 17561 14842 17595 14858
rect 17561 14415 17595 14466
rect 17679 14842 17713 14894
rect 17916 14692 18186 14729
rect 17679 14450 17713 14466
rect 17798 14642 17832 14658
rect 16149 14376 17595 14415
rect 17798 14412 17832 14466
rect 17916 14642 17950 14692
rect 17916 14450 17950 14466
rect 18034 14642 18068 14658
rect 18034 14412 18068 14466
rect 18152 14642 18186 14692
rect 18152 14450 18186 14466
rect 17798 14373 18068 14412
rect 16676 14251 16710 14267
rect 17970 14258 17986 14292
rect 18020 14258 18036 14292
rect 16676 14201 16710 14217
rect 15679 14151 15771 14168
rect 15679 14096 15695 14151
rect 15755 14096 15771 14151
rect 15679 14083 15771 14096
rect 16764 14152 16856 14165
rect 16764 14097 16780 14152
rect 16840 14097 16856 14152
rect 16764 14080 16856 14097
rect 15447 14036 15504 14040
rect 15447 13976 15451 14036
rect 15500 13976 15504 14036
rect 15447 13972 15504 13976
rect 17030 14021 17064 14037
rect 17030 13971 17064 13987
rect 13444 13871 15109 13877
rect 13444 13816 13462 13871
rect 13520 13816 15109 13871
rect 13444 13806 15109 13816
rect 16646 13872 16738 13880
rect 18249 13872 18328 15405
rect 21052 15369 21119 15711
rect 21740 15708 21882 15720
rect 22115 15711 22385 15746
rect 23283 15741 23317 15832
rect 23401 16008 23435 16024
rect 23401 15816 23435 15832
rect 23519 16008 23553 16024
rect 23519 15741 23553 15832
rect 23637 16008 23671 16024
rect 23637 15816 23671 15832
rect 21740 15704 21780 15708
rect 21846 15704 21882 15708
rect 21740 15638 21758 15704
rect 21876 15638 21882 15704
rect 21740 15612 21882 15638
rect 16646 13867 18328 13872
rect 16646 13812 16664 13867
rect 16722 13812 18328 13867
rect 13444 13799 13536 13806
rect 16646 13801 18328 13812
rect 18402 15305 21119 15369
rect 22229 15346 22272 15711
rect 22908 15708 23050 15720
rect 22908 15704 22948 15708
rect 23014 15704 23050 15708
rect 23283 15704 24717 15741
rect 22908 15638 22926 15704
rect 23044 15638 23050 15704
rect 22908 15612 23050 15638
rect 18402 13872 18470 15305
rect 21531 15287 22272 15346
rect 19904 15112 20132 15130
rect 19904 15036 19920 15112
rect 20116 15036 20132 15112
rect 19904 15020 20132 15036
rect 19175 14895 19445 14934
rect 19175 14842 19209 14895
rect 18734 14693 19004 14732
rect 18734 14642 18768 14693
rect 18734 14450 18768 14466
rect 18852 14642 18886 14658
rect 18852 14415 18886 14466
rect 18970 14642 19004 14693
rect 18970 14450 19004 14466
rect 19088 14642 19122 14658
rect 19088 14415 19122 14466
rect 19175 14450 19209 14466
rect 19293 14842 19327 14858
rect 18852 14376 19122 14415
rect 19293 14415 19327 14466
rect 19411 14842 19445 14895
rect 19642 14894 19912 14933
rect 19411 14450 19445 14466
rect 19529 14842 19563 14858
rect 19529 14415 19563 14466
rect 19642 14842 19676 14894
rect 19642 14450 19676 14466
rect 19760 14842 19794 14858
rect 19760 14415 19794 14466
rect 19878 14842 19912 14894
rect 20114 14894 20384 14933
rect 19878 14450 19912 14466
rect 19996 14842 20030 14858
rect 19996 14415 20030 14466
rect 20114 14842 20148 14894
rect 20114 14450 20148 14466
rect 20232 14842 20266 14858
rect 20232 14415 20266 14466
rect 20350 14842 20384 14894
rect 20587 14894 20857 14933
rect 20350 14450 20384 14466
rect 20469 14842 20503 14858
rect 20469 14415 20503 14466
rect 20587 14842 20621 14894
rect 20587 14450 20621 14466
rect 20705 14842 20739 14858
rect 20705 14415 20739 14466
rect 20823 14842 20857 14894
rect 21060 14692 21330 14729
rect 20823 14450 20857 14466
rect 20942 14642 20976 14658
rect 19293 14376 20739 14415
rect 20942 14412 20976 14466
rect 21060 14642 21094 14692
rect 21060 14450 21094 14466
rect 21178 14642 21212 14658
rect 21178 14412 21212 14466
rect 21296 14642 21330 14692
rect 21296 14450 21330 14466
rect 20942 14373 21212 14412
rect 19820 14251 19854 14267
rect 21114 14258 21130 14292
rect 21164 14258 21180 14292
rect 19820 14201 19854 14217
rect 21531 14234 21598 15287
rect 23036 15116 23264 15134
rect 23036 15040 23052 15116
rect 23248 15040 23264 15116
rect 23036 15024 23264 15040
rect 22307 14899 22577 14938
rect 22307 14846 22341 14899
rect 21866 14697 22136 14736
rect 21866 14646 21900 14697
rect 21866 14454 21900 14470
rect 21984 14646 22018 14662
rect 21984 14419 22018 14470
rect 22102 14646 22136 14697
rect 22102 14454 22136 14470
rect 22220 14646 22254 14662
rect 22220 14419 22254 14470
rect 22307 14454 22341 14470
rect 22425 14846 22459 14862
rect 21984 14380 22254 14419
rect 22425 14419 22459 14470
rect 22543 14846 22577 14899
rect 22774 14898 23044 14937
rect 22543 14454 22577 14470
rect 22661 14846 22695 14862
rect 22661 14419 22695 14470
rect 22774 14846 22808 14898
rect 22774 14454 22808 14470
rect 22892 14846 22926 14862
rect 22892 14419 22926 14470
rect 23010 14846 23044 14898
rect 23246 14898 23516 14937
rect 23010 14454 23044 14470
rect 23128 14846 23162 14862
rect 23128 14419 23162 14470
rect 23246 14846 23280 14898
rect 23246 14454 23280 14470
rect 23364 14846 23398 14862
rect 23364 14419 23398 14470
rect 23482 14846 23516 14898
rect 23719 14898 23989 14937
rect 23482 14454 23516 14470
rect 23601 14846 23635 14862
rect 23601 14419 23635 14470
rect 23719 14846 23753 14898
rect 23719 14454 23753 14470
rect 23837 14846 23871 14862
rect 23837 14419 23871 14470
rect 23955 14846 23989 14898
rect 24192 14696 24462 14733
rect 23955 14454 23989 14470
rect 24074 14646 24108 14662
rect 22425 14380 23871 14419
rect 24074 14416 24108 14470
rect 24192 14646 24226 14696
rect 24192 14454 24226 14470
rect 24310 14646 24344 14662
rect 24310 14416 24344 14470
rect 24428 14646 24462 14696
rect 24428 14454 24462 14470
rect 24074 14377 24344 14416
rect 22952 14255 22986 14271
rect 24246 14262 24262 14296
rect 24296 14262 24312 14296
rect 18823 14151 18915 14168
rect 18823 14096 18839 14151
rect 18899 14096 18915 14151
rect 18823 14083 18915 14096
rect 19908 14152 20000 14165
rect 19908 14097 19924 14152
rect 19984 14097 20000 14152
rect 19908 14080 20000 14097
rect 18591 14036 18648 14040
rect 18591 13976 18595 14036
rect 18644 13976 18648 14036
rect 18591 13972 18648 13976
rect 20174 14021 20208 14037
rect 20174 13971 20208 13987
rect 18402 13868 18648 13872
rect 18402 13808 18595 13868
rect 18644 13808 18648 13868
rect 18402 13804 18648 13808
rect 19790 13867 19882 13880
rect 19790 13812 19806 13867
rect 19866 13812 19882 13867
rect 16646 13795 16738 13801
rect 19790 13795 19882 13812
rect 21531 13875 21599 14234
rect 22952 14205 22986 14221
rect 21955 14155 22047 14172
rect 21955 14100 21971 14155
rect 22031 14100 22047 14155
rect 21955 14087 22047 14100
rect 23040 14156 23132 14169
rect 23040 14101 23056 14156
rect 23116 14101 23132 14156
rect 23040 14084 23132 14101
rect 21723 14040 21780 14044
rect 21723 13980 21727 14040
rect 21776 13980 21780 14040
rect 21723 13976 21780 13980
rect 23306 14025 23340 14041
rect 23306 13975 23340 13991
rect 21723 13875 21780 13876
rect 21531 13872 21780 13875
rect 21531 13812 21727 13872
rect 21776 13812 21780 13872
rect 21531 13808 21780 13812
rect 22922 13871 23014 13884
rect 22922 13816 22938 13871
rect 22998 13816 23014 13871
rect 21531 13807 21777 13808
rect 22922 13799 23014 13816
rect 24679 13876 24717 15704
rect 26180 15116 26408 15134
rect 26180 15040 26196 15116
rect 26392 15040 26408 15116
rect 26180 15024 26408 15040
rect 25451 14899 25721 14938
rect 25451 14846 25485 14899
rect 25010 14697 25280 14736
rect 25010 14646 25044 14697
rect 25010 14454 25044 14470
rect 25128 14646 25162 14662
rect 25128 14419 25162 14470
rect 25246 14646 25280 14697
rect 25246 14454 25280 14470
rect 25364 14646 25398 14662
rect 25364 14419 25398 14470
rect 25451 14454 25485 14470
rect 25569 14846 25603 14862
rect 25128 14380 25398 14419
rect 25569 14419 25603 14470
rect 25687 14846 25721 14899
rect 25918 14898 26188 14937
rect 25687 14454 25721 14470
rect 25805 14846 25839 14862
rect 25805 14419 25839 14470
rect 25918 14846 25952 14898
rect 25918 14454 25952 14470
rect 26036 14846 26070 14862
rect 26036 14419 26070 14470
rect 26154 14846 26188 14898
rect 26390 14898 26660 14937
rect 26154 14454 26188 14470
rect 26272 14846 26306 14862
rect 26272 14419 26306 14470
rect 26390 14846 26424 14898
rect 26390 14454 26424 14470
rect 26508 14846 26542 14862
rect 26508 14419 26542 14470
rect 26626 14846 26660 14898
rect 26863 14898 27133 14937
rect 26626 14454 26660 14470
rect 26745 14846 26779 14862
rect 26745 14419 26779 14470
rect 26863 14846 26897 14898
rect 26863 14454 26897 14470
rect 26981 14846 27015 14862
rect 26981 14419 27015 14470
rect 27099 14846 27133 14898
rect 27336 14696 27606 14733
rect 27099 14454 27133 14470
rect 27218 14646 27252 14662
rect 25569 14380 27015 14419
rect 27218 14416 27252 14470
rect 27336 14646 27370 14696
rect 27336 14454 27370 14470
rect 27454 14646 27488 14662
rect 27454 14416 27488 14470
rect 27572 14646 27606 14696
rect 27572 14454 27606 14470
rect 27218 14377 27488 14416
rect 26096 14255 26130 14271
rect 27390 14262 27406 14296
rect 27440 14262 27456 14296
rect 26096 14205 26130 14221
rect 25099 14155 25191 14172
rect 25099 14100 25115 14155
rect 25175 14100 25191 14155
rect 25099 14087 25191 14100
rect 26184 14156 26276 14169
rect 26184 14101 26200 14156
rect 26260 14101 26276 14156
rect 26184 14084 26276 14101
rect 24867 14040 24924 14044
rect 24867 13980 24871 14040
rect 24920 13980 24924 14040
rect 24867 13976 24924 13980
rect 26450 14025 26484 14041
rect 26450 13975 26484 13991
rect 24679 13872 24933 13876
rect 24679 13812 24871 13872
rect 24920 13812 24933 13872
rect 24679 13808 24933 13812
rect 26066 13871 26158 13884
rect 26066 13816 26082 13871
rect 26142 13816 26158 13871
rect 26066 13799 26158 13816
rect 4289 13631 4323 13647
rect 4289 13581 4323 13597
rect 7433 13631 7467 13647
rect 7433 13581 7467 13597
rect 10565 13635 10599 13651
rect 10565 13585 10599 13601
rect 13709 13635 13743 13651
rect 13709 13585 13743 13601
rect 16911 13631 16945 13647
rect 16911 13581 16945 13597
rect 20055 13631 20089 13647
rect 20055 13581 20089 13597
rect 23187 13635 23221 13651
rect 23187 13585 23221 13601
rect 26331 13635 26365 13651
rect 26331 13585 26365 13601
rect 3802 13509 3836 13525
rect 3802 13317 3836 13333
rect 3920 13521 3954 13525
rect 3994 13521 4028 13525
rect 3920 13509 4028 13521
rect 3954 13333 3994 13509
rect 3920 13321 3994 13333
rect 3920 13317 3954 13321
rect 3994 13117 4028 13133
rect 4112 13509 4146 13525
rect 4112 13117 4146 13133
rect 4230 13509 4264 13525
rect 4230 13117 4264 13133
rect 4348 13509 4382 13525
rect 4348 13117 4382 13133
rect 4466 13521 4500 13525
rect 4544 13521 4578 13525
rect 4466 13509 4578 13521
rect 4500 13333 4544 13509
rect 4500 13321 4578 13333
rect 4544 13317 4578 13321
rect 4662 13509 4696 13525
rect 4662 13317 4696 13333
rect 6946 13509 6980 13525
rect 6946 13317 6980 13333
rect 7064 13521 7098 13525
rect 7138 13521 7172 13525
rect 7064 13509 7172 13521
rect 7098 13333 7138 13509
rect 7064 13321 7138 13333
rect 7064 13317 7098 13321
rect 4466 13117 4500 13133
rect 7138 13117 7172 13133
rect 7256 13509 7290 13525
rect 7256 13117 7290 13133
rect 7374 13509 7408 13525
rect 7374 13117 7408 13133
rect 7492 13509 7526 13525
rect 7492 13117 7526 13133
rect 7610 13521 7644 13525
rect 7688 13521 7722 13525
rect 7610 13509 7722 13521
rect 7644 13333 7688 13509
rect 7644 13321 7722 13333
rect 7688 13317 7722 13321
rect 7806 13509 7840 13525
rect 7806 13317 7840 13333
rect 10078 13513 10112 13529
rect 10078 13321 10112 13337
rect 10196 13525 10230 13529
rect 10270 13525 10304 13529
rect 10196 13513 10304 13525
rect 10230 13337 10270 13513
rect 10196 13325 10270 13337
rect 10196 13321 10230 13325
rect 7610 13117 7644 13133
rect 10270 13121 10304 13137
rect 10388 13513 10422 13529
rect 10388 13121 10422 13137
rect 10506 13513 10540 13529
rect 10506 13121 10540 13137
rect 10624 13513 10658 13529
rect 10624 13121 10658 13137
rect 10742 13525 10776 13529
rect 10820 13525 10854 13529
rect 10742 13513 10854 13525
rect 10776 13337 10820 13513
rect 10776 13325 10854 13337
rect 10820 13321 10854 13325
rect 10938 13513 10972 13529
rect 10938 13321 10972 13337
rect 13222 13513 13256 13529
rect 13222 13321 13256 13337
rect 13340 13525 13374 13529
rect 13414 13525 13448 13529
rect 13340 13513 13448 13525
rect 13374 13337 13414 13513
rect 13340 13325 13414 13337
rect 13340 13321 13374 13325
rect 10742 13121 10776 13137
rect 13414 13121 13448 13137
rect 13532 13513 13566 13529
rect 13532 13121 13566 13137
rect 13650 13513 13684 13529
rect 13650 13121 13684 13137
rect 13768 13513 13802 13529
rect 13768 13121 13802 13137
rect 13886 13525 13920 13529
rect 13964 13525 13998 13529
rect 13886 13513 13998 13525
rect 13920 13337 13964 13513
rect 13920 13325 13998 13337
rect 13964 13321 13998 13325
rect 14082 13513 14116 13529
rect 14082 13321 14116 13337
rect 16424 13509 16458 13525
rect 16424 13317 16458 13333
rect 16542 13521 16576 13525
rect 16616 13521 16650 13525
rect 16542 13509 16650 13521
rect 16576 13333 16616 13509
rect 16542 13321 16616 13333
rect 16542 13317 16576 13321
rect 13886 13121 13920 13137
rect 16616 13117 16650 13133
rect 16734 13509 16768 13525
rect 16734 13117 16768 13133
rect 16852 13509 16886 13525
rect 16852 13117 16886 13133
rect 16970 13509 17004 13525
rect 16970 13117 17004 13133
rect 17088 13521 17122 13525
rect 17166 13521 17200 13525
rect 17088 13509 17200 13521
rect 17122 13333 17166 13509
rect 17122 13321 17200 13333
rect 17166 13317 17200 13321
rect 17284 13509 17318 13525
rect 17284 13317 17318 13333
rect 19568 13509 19602 13525
rect 19568 13317 19602 13333
rect 19686 13521 19720 13525
rect 19760 13521 19794 13525
rect 19686 13509 19794 13521
rect 19720 13333 19760 13509
rect 19686 13321 19760 13333
rect 19686 13317 19720 13321
rect 17088 13117 17122 13133
rect 19760 13117 19794 13133
rect 19878 13509 19912 13525
rect 19878 13117 19912 13133
rect 19996 13509 20030 13525
rect 19996 13117 20030 13133
rect 20114 13509 20148 13525
rect 20114 13117 20148 13133
rect 20232 13521 20266 13525
rect 20310 13521 20344 13525
rect 20232 13509 20344 13521
rect 20266 13333 20310 13509
rect 20266 13321 20344 13333
rect 20310 13317 20344 13321
rect 20428 13509 20462 13525
rect 20428 13317 20462 13333
rect 22700 13513 22734 13529
rect 22700 13321 22734 13337
rect 22818 13525 22852 13529
rect 22892 13525 22926 13529
rect 22818 13513 22926 13525
rect 22852 13337 22892 13513
rect 22818 13325 22892 13337
rect 22818 13321 22852 13325
rect 20232 13117 20266 13133
rect 22892 13121 22926 13137
rect 23010 13513 23044 13529
rect 23010 13121 23044 13137
rect 23128 13513 23162 13529
rect 23128 13121 23162 13137
rect 23246 13513 23280 13529
rect 23246 13121 23280 13137
rect 23364 13525 23398 13529
rect 23442 13525 23476 13529
rect 23364 13513 23476 13525
rect 23398 13337 23442 13513
rect 23398 13325 23476 13337
rect 23442 13321 23476 13325
rect 23560 13513 23594 13529
rect 23560 13321 23594 13337
rect 25844 13513 25878 13529
rect 25844 13321 25878 13337
rect 25962 13525 25996 13529
rect 26036 13525 26070 13529
rect 25962 13513 26070 13525
rect 25996 13337 26036 13513
rect 25962 13325 26036 13337
rect 25962 13321 25996 13325
rect 23364 13121 23398 13137
rect 26036 13121 26070 13137
rect 26154 13513 26188 13529
rect 26154 13121 26188 13137
rect 26272 13513 26306 13529
rect 26272 13121 26306 13137
rect 26390 13513 26424 13529
rect 26390 13121 26424 13137
rect 26508 13525 26542 13529
rect 26586 13525 26620 13529
rect 26508 13513 26620 13525
rect 26542 13337 26586 13513
rect 26542 13325 26620 13337
rect 26586 13321 26620 13325
rect 26704 13513 26738 13529
rect 26704 13321 26738 13337
rect 26508 13121 26542 13137
rect 4215 12998 4231 13032
rect 4265 12998 4281 13032
rect 7359 12998 7375 13032
rect 7409 12998 7425 13032
rect 10491 13002 10507 13036
rect 10541 13002 10557 13036
rect 13635 13002 13651 13036
rect 13685 13002 13701 13036
rect 16837 12998 16853 13032
rect 16887 12998 16903 13032
rect 19981 12998 19997 13032
rect 20031 12998 20047 13032
rect 23113 13002 23129 13036
rect 23163 13002 23179 13036
rect 26257 13002 26273 13036
rect 26307 13002 26323 13036
rect 10472 12884 10608 12888
rect 4196 12880 4332 12884
rect 4196 12866 4234 12880
rect 4292 12866 4332 12880
rect 4196 12820 4212 12866
rect 4316 12820 4332 12866
rect 4196 12798 4332 12820
rect 7340 12880 7476 12884
rect 7340 12866 7378 12880
rect 7436 12866 7476 12880
rect 7340 12820 7356 12866
rect 7460 12820 7476 12866
rect 7340 12798 7476 12820
rect 10472 12870 10510 12884
rect 10568 12870 10608 12884
rect 10472 12824 10488 12870
rect 10592 12824 10608 12870
rect 10472 12802 10608 12824
rect 13616 12884 13752 12888
rect 23094 12884 23230 12888
rect 13616 12870 13654 12884
rect 13712 12870 13752 12884
rect 13616 12824 13632 12870
rect 13736 12824 13752 12870
rect 13616 12802 13752 12824
rect 16818 12880 16954 12884
rect 16818 12866 16856 12880
rect 16914 12866 16954 12880
rect 16818 12820 16834 12866
rect 16938 12820 16954 12866
rect 16818 12798 16954 12820
rect 19962 12880 20098 12884
rect 19962 12866 20000 12880
rect 20058 12866 20098 12880
rect 19962 12820 19978 12866
rect 20082 12820 20098 12866
rect 19962 12798 20098 12820
rect 23094 12870 23132 12884
rect 23190 12870 23230 12884
rect 23094 12824 23110 12870
rect 23214 12824 23230 12870
rect 23094 12802 23230 12824
rect 26238 12884 26374 12888
rect 26238 12870 26276 12884
rect 26334 12870 26374 12884
rect 26238 12824 26254 12870
rect 26358 12824 26374 12870
rect 26238 12802 26374 12824
rect 4138 12378 4366 12396
rect 4138 12302 4154 12378
rect 4350 12302 4366 12378
rect 4138 12286 4366 12302
rect 7282 12378 7510 12396
rect 7282 12302 7298 12378
rect 7494 12302 7510 12378
rect 7282 12286 7510 12302
rect 10414 12382 10642 12400
rect 10414 12306 10430 12382
rect 10626 12306 10642 12382
rect 10414 12290 10642 12306
rect 13558 12382 13786 12400
rect 13558 12306 13574 12382
rect 13770 12306 13786 12382
rect 13558 12290 13786 12306
rect 16760 12378 16988 12396
rect 16760 12302 16776 12378
rect 16972 12302 16988 12378
rect 16760 12286 16988 12302
rect 19904 12378 20132 12396
rect 19904 12302 19920 12378
rect 20116 12302 20132 12378
rect 19904 12286 20132 12302
rect 23036 12382 23264 12400
rect 23036 12306 23052 12382
rect 23248 12306 23264 12382
rect 23036 12290 23264 12306
rect 26180 12382 26408 12400
rect 26180 12306 26196 12382
rect 26392 12306 26408 12382
rect 26180 12290 26408 12306
rect 3409 12161 3679 12200
rect 3409 12108 3443 12161
rect 2968 11959 3238 11998
rect 2968 11908 3002 11959
rect 2968 11716 3002 11732
rect 3086 11908 3120 11924
rect 3086 11681 3120 11732
rect 3204 11908 3238 11959
rect 3204 11716 3238 11732
rect 3322 11908 3356 11924
rect 3322 11681 3356 11732
rect 3409 11716 3443 11732
rect 3527 12108 3561 12124
rect 3086 11642 3356 11681
rect 3527 11681 3561 11732
rect 3645 12108 3679 12161
rect 3876 12160 4146 12199
rect 3645 11716 3679 11732
rect 3763 12108 3797 12124
rect 3763 11681 3797 11732
rect 3876 12108 3910 12160
rect 3876 11716 3910 11732
rect 3994 12108 4028 12124
rect 3994 11681 4028 11732
rect 4112 12108 4146 12160
rect 4348 12160 4618 12199
rect 4112 11716 4146 11732
rect 4230 12108 4264 12124
rect 4230 11681 4264 11732
rect 4348 12108 4382 12160
rect 4348 11716 4382 11732
rect 4466 12108 4500 12124
rect 4466 11681 4500 11732
rect 4584 12108 4618 12160
rect 4821 12160 5091 12199
rect 4584 11716 4618 11732
rect 4703 12108 4737 12124
rect 4703 11681 4737 11732
rect 4821 12108 4855 12160
rect 4821 11716 4855 11732
rect 4939 12108 4973 12124
rect 4939 11681 4973 11732
rect 5057 12108 5091 12160
rect 6553 12161 6823 12200
rect 6553 12108 6587 12161
rect 5294 11958 5564 11995
rect 5057 11716 5091 11732
rect 5176 11908 5210 11924
rect 3527 11642 4973 11681
rect 5176 11678 5210 11732
rect 5294 11908 5328 11958
rect 5294 11716 5328 11732
rect 5412 11908 5446 11924
rect 5412 11678 5446 11732
rect 5530 11908 5564 11958
rect 5530 11716 5564 11732
rect 6112 11959 6382 11998
rect 6112 11908 6146 11959
rect 6112 11716 6146 11732
rect 6230 11908 6264 11924
rect 5176 11639 5446 11678
rect 6230 11681 6264 11732
rect 6348 11908 6382 11959
rect 6348 11716 6382 11732
rect 6466 11908 6500 11924
rect 6466 11681 6500 11732
rect 6553 11716 6587 11732
rect 6671 12108 6705 12124
rect 6230 11642 6500 11681
rect 6671 11681 6705 11732
rect 6789 12108 6823 12161
rect 7020 12160 7290 12199
rect 6789 11716 6823 11732
rect 6907 12108 6941 12124
rect 6907 11681 6941 11732
rect 7020 12108 7054 12160
rect 7020 11716 7054 11732
rect 7138 12108 7172 12124
rect 7138 11681 7172 11732
rect 7256 12108 7290 12160
rect 7492 12160 7762 12199
rect 7256 11716 7290 11732
rect 7374 12108 7408 12124
rect 7374 11681 7408 11732
rect 7492 12108 7526 12160
rect 7492 11716 7526 11732
rect 7610 12108 7644 12124
rect 7610 11681 7644 11732
rect 7728 12108 7762 12160
rect 7965 12160 8235 12199
rect 7728 11716 7762 11732
rect 7847 12108 7881 12124
rect 7847 11681 7881 11732
rect 7965 12108 7999 12160
rect 7965 11716 7999 11732
rect 8083 12108 8117 12124
rect 8083 11681 8117 11732
rect 8201 12108 8235 12160
rect 9685 12165 9955 12204
rect 9685 12112 9719 12165
rect 8438 11958 8708 11995
rect 8201 11716 8235 11732
rect 8320 11908 8354 11924
rect 6671 11642 8117 11681
rect 8320 11678 8354 11732
rect 8438 11908 8472 11958
rect 8438 11716 8472 11732
rect 8556 11908 8590 11924
rect 8556 11678 8590 11732
rect 8674 11908 8708 11958
rect 8674 11716 8708 11732
rect 9244 11963 9514 12002
rect 9244 11912 9278 11963
rect 9244 11720 9278 11736
rect 9362 11912 9396 11928
rect 8320 11639 8590 11678
rect 9362 11685 9396 11736
rect 9480 11912 9514 11963
rect 9480 11720 9514 11736
rect 9598 11912 9632 11928
rect 9598 11685 9632 11736
rect 9685 11720 9719 11736
rect 9803 12112 9837 12128
rect 9362 11646 9632 11685
rect 9803 11685 9837 11736
rect 9921 12112 9955 12165
rect 10152 12164 10422 12203
rect 9921 11720 9955 11736
rect 10039 12112 10073 12128
rect 10039 11685 10073 11736
rect 10152 12112 10186 12164
rect 10152 11720 10186 11736
rect 10270 12112 10304 12128
rect 10270 11685 10304 11736
rect 10388 12112 10422 12164
rect 10624 12164 10894 12203
rect 10388 11720 10422 11736
rect 10506 12112 10540 12128
rect 10506 11685 10540 11736
rect 10624 12112 10658 12164
rect 10624 11720 10658 11736
rect 10742 12112 10776 12128
rect 10742 11685 10776 11736
rect 10860 12112 10894 12164
rect 11097 12164 11367 12203
rect 10860 11720 10894 11736
rect 10979 12112 11013 12128
rect 10979 11685 11013 11736
rect 11097 12112 11131 12164
rect 11097 11720 11131 11736
rect 11215 12112 11249 12128
rect 11215 11685 11249 11736
rect 11333 12112 11367 12164
rect 12829 12165 13099 12204
rect 12829 12112 12863 12165
rect 11570 11962 11840 11999
rect 11333 11720 11367 11736
rect 11452 11912 11486 11928
rect 9803 11646 11249 11685
rect 11452 11682 11486 11736
rect 11570 11912 11604 11962
rect 11570 11720 11604 11736
rect 11688 11912 11722 11928
rect 11688 11682 11722 11736
rect 11806 11912 11840 11962
rect 11806 11720 11840 11736
rect 12388 11963 12658 12002
rect 12388 11912 12422 11963
rect 12388 11720 12422 11736
rect 12506 11912 12540 11928
rect 11452 11643 11722 11682
rect 12506 11685 12540 11736
rect 12624 11912 12658 11963
rect 12624 11720 12658 11736
rect 12742 11912 12776 11928
rect 12742 11685 12776 11736
rect 12829 11720 12863 11736
rect 12947 12112 12981 12128
rect 12506 11646 12776 11685
rect 12947 11685 12981 11736
rect 13065 12112 13099 12165
rect 13296 12164 13566 12203
rect 13065 11720 13099 11736
rect 13183 12112 13217 12128
rect 13183 11685 13217 11736
rect 13296 12112 13330 12164
rect 13296 11720 13330 11736
rect 13414 12112 13448 12128
rect 13414 11685 13448 11736
rect 13532 12112 13566 12164
rect 13768 12164 14038 12203
rect 13532 11720 13566 11736
rect 13650 12112 13684 12128
rect 13650 11685 13684 11736
rect 13768 12112 13802 12164
rect 13768 11720 13802 11736
rect 13886 12112 13920 12128
rect 13886 11685 13920 11736
rect 14004 12112 14038 12164
rect 14241 12164 14511 12203
rect 14004 11720 14038 11736
rect 14123 12112 14157 12128
rect 14123 11685 14157 11736
rect 14241 12112 14275 12164
rect 14241 11720 14275 11736
rect 14359 12112 14393 12128
rect 14359 11685 14393 11736
rect 14477 12112 14511 12164
rect 16031 12161 16301 12200
rect 16031 12108 16065 12161
rect 14714 11962 14984 11999
rect 14477 11720 14511 11736
rect 14596 11912 14630 11928
rect 12947 11646 14393 11685
rect 14596 11682 14630 11736
rect 14714 11912 14748 11962
rect 14714 11720 14748 11736
rect 14832 11912 14866 11928
rect 14832 11682 14866 11736
rect 14950 11912 14984 11962
rect 14950 11720 14984 11736
rect 15590 11959 15860 11998
rect 15590 11908 15624 11959
rect 15590 11716 15624 11732
rect 15708 11908 15742 11924
rect 14596 11643 14866 11682
rect 15708 11681 15742 11732
rect 15826 11908 15860 11959
rect 15826 11716 15860 11732
rect 15944 11908 15978 11924
rect 15944 11681 15978 11732
rect 16031 11716 16065 11732
rect 16149 12108 16183 12124
rect 15708 11642 15978 11681
rect 16149 11681 16183 11732
rect 16267 12108 16301 12161
rect 16498 12160 16768 12199
rect 16267 11716 16301 11732
rect 16385 12108 16419 12124
rect 16385 11681 16419 11732
rect 16498 12108 16532 12160
rect 16498 11716 16532 11732
rect 16616 12108 16650 12124
rect 16616 11681 16650 11732
rect 16734 12108 16768 12160
rect 16970 12160 17240 12199
rect 16734 11716 16768 11732
rect 16852 12108 16886 12124
rect 16852 11681 16886 11732
rect 16970 12108 17004 12160
rect 16970 11716 17004 11732
rect 17088 12108 17122 12124
rect 17088 11681 17122 11732
rect 17206 12108 17240 12160
rect 17443 12160 17713 12199
rect 17206 11716 17240 11732
rect 17325 12108 17359 12124
rect 17325 11681 17359 11732
rect 17443 12108 17477 12160
rect 17443 11716 17477 11732
rect 17561 12108 17595 12124
rect 17561 11681 17595 11732
rect 17679 12108 17713 12160
rect 19175 12161 19445 12200
rect 19175 12108 19209 12161
rect 17916 11958 18186 11995
rect 17679 11716 17713 11732
rect 17798 11908 17832 11924
rect 16149 11642 17595 11681
rect 17798 11678 17832 11732
rect 17916 11908 17950 11958
rect 17916 11716 17950 11732
rect 18034 11908 18068 11924
rect 18034 11678 18068 11732
rect 18152 11908 18186 11958
rect 18152 11716 18186 11732
rect 18734 11959 19004 11998
rect 18734 11908 18768 11959
rect 18734 11716 18768 11732
rect 18852 11908 18886 11924
rect 17798 11639 18068 11678
rect 18852 11681 18886 11732
rect 18970 11908 19004 11959
rect 18970 11716 19004 11732
rect 19088 11908 19122 11924
rect 19088 11681 19122 11732
rect 19175 11716 19209 11732
rect 19293 12108 19327 12124
rect 18852 11642 19122 11681
rect 19293 11681 19327 11732
rect 19411 12108 19445 12161
rect 19642 12160 19912 12199
rect 19411 11716 19445 11732
rect 19529 12108 19563 12124
rect 19529 11681 19563 11732
rect 19642 12108 19676 12160
rect 19642 11716 19676 11732
rect 19760 12108 19794 12124
rect 19760 11681 19794 11732
rect 19878 12108 19912 12160
rect 20114 12160 20384 12199
rect 19878 11716 19912 11732
rect 19996 12108 20030 12124
rect 19996 11681 20030 11732
rect 20114 12108 20148 12160
rect 20114 11716 20148 11732
rect 20232 12108 20266 12124
rect 20232 11681 20266 11732
rect 20350 12108 20384 12160
rect 20587 12160 20857 12199
rect 20350 11716 20384 11732
rect 20469 12108 20503 12124
rect 20469 11681 20503 11732
rect 20587 12108 20621 12160
rect 20587 11716 20621 11732
rect 20705 12108 20739 12124
rect 20705 11681 20739 11732
rect 20823 12108 20857 12160
rect 22307 12165 22577 12204
rect 22307 12112 22341 12165
rect 21060 11958 21330 11995
rect 20823 11716 20857 11732
rect 20942 11908 20976 11924
rect 19293 11642 20739 11681
rect 20942 11678 20976 11732
rect 21060 11908 21094 11958
rect 21060 11716 21094 11732
rect 21178 11908 21212 11924
rect 21178 11678 21212 11732
rect 21296 11908 21330 11958
rect 21296 11716 21330 11732
rect 21866 11963 22136 12002
rect 21866 11912 21900 11963
rect 21866 11720 21900 11736
rect 21984 11912 22018 11928
rect 20942 11639 21212 11678
rect 21984 11685 22018 11736
rect 22102 11912 22136 11963
rect 22102 11720 22136 11736
rect 22220 11912 22254 11928
rect 22220 11685 22254 11736
rect 22307 11720 22341 11736
rect 22425 12112 22459 12128
rect 21984 11646 22254 11685
rect 22425 11685 22459 11736
rect 22543 12112 22577 12165
rect 22774 12164 23044 12203
rect 22543 11720 22577 11736
rect 22661 12112 22695 12128
rect 22661 11685 22695 11736
rect 22774 12112 22808 12164
rect 22774 11720 22808 11736
rect 22892 12112 22926 12128
rect 22892 11685 22926 11736
rect 23010 12112 23044 12164
rect 23246 12164 23516 12203
rect 23010 11720 23044 11736
rect 23128 12112 23162 12128
rect 23128 11685 23162 11736
rect 23246 12112 23280 12164
rect 23246 11720 23280 11736
rect 23364 12112 23398 12128
rect 23364 11685 23398 11736
rect 23482 12112 23516 12164
rect 23719 12164 23989 12203
rect 23482 11720 23516 11736
rect 23601 12112 23635 12128
rect 23601 11685 23635 11736
rect 23719 12112 23753 12164
rect 23719 11720 23753 11736
rect 23837 12112 23871 12128
rect 23837 11685 23871 11736
rect 23955 12112 23989 12164
rect 25451 12165 25721 12204
rect 25451 12112 25485 12165
rect 24192 11962 24462 11999
rect 23955 11720 23989 11736
rect 24074 11912 24108 11928
rect 22425 11646 23871 11685
rect 24074 11682 24108 11736
rect 24192 11912 24226 11962
rect 24192 11720 24226 11736
rect 24310 11912 24344 11928
rect 24310 11682 24344 11736
rect 24428 11912 24462 11962
rect 24428 11720 24462 11736
rect 25010 11963 25280 12002
rect 25010 11912 25044 11963
rect 25010 11720 25044 11736
rect 25128 11912 25162 11928
rect 24074 11643 24344 11682
rect 25128 11685 25162 11736
rect 25246 11912 25280 11963
rect 25246 11720 25280 11736
rect 25364 11912 25398 11928
rect 25364 11685 25398 11736
rect 25451 11720 25485 11736
rect 25569 12112 25603 12128
rect 25128 11646 25398 11685
rect 25569 11685 25603 11736
rect 25687 12112 25721 12165
rect 25918 12164 26188 12203
rect 25687 11720 25721 11736
rect 25805 12112 25839 12128
rect 25805 11685 25839 11736
rect 25918 12112 25952 12164
rect 25918 11720 25952 11736
rect 26036 12112 26070 12128
rect 26036 11685 26070 11736
rect 26154 12112 26188 12164
rect 26390 12164 26660 12203
rect 26154 11720 26188 11736
rect 26272 12112 26306 12128
rect 26272 11685 26306 11736
rect 26390 12112 26424 12164
rect 26390 11720 26424 11736
rect 26508 12112 26542 12128
rect 26508 11685 26542 11736
rect 26626 12112 26660 12164
rect 26863 12164 27133 12203
rect 26626 11720 26660 11736
rect 26745 12112 26779 12128
rect 26745 11685 26779 11736
rect 26863 12112 26897 12164
rect 26863 11720 26897 11736
rect 26981 12112 27015 12128
rect 26981 11685 27015 11736
rect 27099 12112 27133 12164
rect 27336 11962 27606 11999
rect 27099 11720 27133 11736
rect 27218 11912 27252 11928
rect 25569 11646 27015 11685
rect 27218 11682 27252 11736
rect 27336 11912 27370 11962
rect 27336 11720 27370 11736
rect 27454 11912 27488 11928
rect 27454 11682 27488 11736
rect 27572 11912 27606 11962
rect 27572 11720 27606 11736
rect 27218 11643 27488 11682
rect 4054 11517 4088 11533
rect 5348 11524 5364 11558
rect 5398 11524 5414 11558
rect 4054 11467 4088 11483
rect 7198 11517 7232 11533
rect 8492 11524 8508 11558
rect 8542 11524 8558 11558
rect 7198 11467 7232 11483
rect 10330 11521 10364 11537
rect 11624 11528 11640 11562
rect 11674 11528 11690 11562
rect 10330 11471 10364 11487
rect 13474 11521 13508 11537
rect 14768 11528 14784 11562
rect 14818 11528 14834 11562
rect 13474 11471 13508 11487
rect 16676 11517 16710 11533
rect 17970 11524 17986 11558
rect 18020 11524 18036 11558
rect 16676 11467 16710 11483
rect 19820 11517 19854 11533
rect 21114 11524 21130 11558
rect 21164 11524 21180 11558
rect 19820 11467 19854 11483
rect 22952 11521 22986 11537
rect 24246 11528 24262 11562
rect 24296 11528 24312 11562
rect 22952 11471 22986 11487
rect 26096 11521 26130 11537
rect 27390 11528 27406 11562
rect 27440 11528 27456 11562
rect 26096 11471 26130 11487
rect 3057 11417 3149 11434
rect 3057 11362 3073 11417
rect 3133 11362 3149 11417
rect 3057 11349 3149 11362
rect 4142 11418 4234 11431
rect 4142 11363 4158 11418
rect 4218 11363 4234 11418
rect 4142 11346 4234 11363
rect 6201 11417 6293 11434
rect 6201 11362 6217 11417
rect 6277 11362 6293 11417
rect 6201 11349 6293 11362
rect 7286 11418 7378 11431
rect 7286 11363 7302 11418
rect 7362 11363 7378 11418
rect 7286 11346 7378 11363
rect 9333 11421 9425 11438
rect 9333 11366 9349 11421
rect 9409 11366 9425 11421
rect 9333 11353 9425 11366
rect 10418 11422 10510 11435
rect 10418 11367 10434 11422
rect 10494 11367 10510 11422
rect 10418 11350 10510 11367
rect 12477 11421 12569 11438
rect 12477 11366 12493 11421
rect 12553 11366 12569 11421
rect 12477 11353 12569 11366
rect 13562 11422 13654 11435
rect 13562 11367 13578 11422
rect 13638 11367 13654 11422
rect 13562 11350 13654 11367
rect 15679 11417 15771 11434
rect 15679 11362 15695 11417
rect 15755 11362 15771 11417
rect 15679 11349 15771 11362
rect 16764 11418 16856 11431
rect 16764 11363 16780 11418
rect 16840 11363 16856 11418
rect 16764 11346 16856 11363
rect 18591 11418 18648 11422
rect 18591 11358 18595 11418
rect 18644 11358 18648 11418
rect 18591 11354 18648 11358
rect 18823 11417 18915 11434
rect 18823 11362 18839 11417
rect 18899 11362 18915 11417
rect 18823 11349 18915 11362
rect 19908 11418 20000 11431
rect 19908 11363 19924 11418
rect 19984 11363 20000 11418
rect 19908 11346 20000 11363
rect 21955 11421 22047 11438
rect 21955 11366 21971 11421
rect 22031 11366 22047 11421
rect 21955 11353 22047 11366
rect 23040 11422 23132 11435
rect 23040 11367 23056 11422
rect 23116 11367 23132 11422
rect 23040 11350 23132 11367
rect 25099 11421 25191 11438
rect 25099 11366 25115 11421
rect 25175 11366 25191 11421
rect 25099 11353 25191 11366
rect 26184 11422 26276 11435
rect 26184 11367 26200 11422
rect 26260 11367 26276 11422
rect 26184 11350 26276 11367
rect 9101 11306 9158 11310
rect 2825 11302 2882 11306
rect 2825 11242 2829 11302
rect 2878 11242 2882 11302
rect 2825 11238 2882 11242
rect 4408 11287 4442 11303
rect 4408 11237 4442 11253
rect 5969 11302 6026 11306
rect 5969 11242 5973 11302
rect 6022 11242 6026 11302
rect 5969 11238 6026 11242
rect 7552 11287 7586 11303
rect 7552 11237 7586 11253
rect 9101 11246 9105 11306
rect 9154 11246 9158 11306
rect 9101 11242 9158 11246
rect 10684 11291 10718 11307
rect 10684 11241 10718 11257
rect 12245 11306 12302 11310
rect 12245 11246 12249 11306
rect 12298 11246 12302 11306
rect 12245 11242 12302 11246
rect 13828 11291 13862 11307
rect 21723 11306 21780 11310
rect 13828 11241 13862 11257
rect 15447 11302 15504 11306
rect 15447 11242 15451 11302
rect 15500 11242 15504 11302
rect 15447 11238 15504 11242
rect 17030 11287 17064 11303
rect 17030 11237 17064 11253
rect 18591 11302 18648 11306
rect 18591 11242 18595 11302
rect 18644 11242 18648 11302
rect 18591 11238 18648 11242
rect 20174 11287 20208 11303
rect 20174 11237 20208 11253
rect 21723 11246 21727 11306
rect 21776 11246 21780 11306
rect 21723 11242 21780 11246
rect 23306 11291 23340 11307
rect 23306 11241 23340 11257
rect 24867 11306 24924 11310
rect 24867 11246 24871 11306
rect 24920 11246 24924 11306
rect 24867 11242 24924 11246
rect 26450 11291 26484 11307
rect 26450 11241 26484 11257
rect 2825 11134 2882 11138
rect 2825 11074 2829 11134
rect 2878 11074 2882 11134
rect 2825 11070 2882 11074
rect 4024 11133 4116 11146
rect 4024 11078 4040 11133
rect 4100 11078 4116 11133
rect 4024 11061 4116 11078
rect 5969 11134 6026 11138
rect 5969 11074 5973 11134
rect 6022 11074 6026 11134
rect 5969 11070 6026 11074
rect 7168 11133 7260 11146
rect 7168 11078 7184 11133
rect 7244 11078 7260 11133
rect 7168 11061 7260 11078
rect 9101 11138 9158 11142
rect 9101 11078 9105 11138
rect 9154 11078 9158 11138
rect 9101 11074 9158 11078
rect 10300 11137 10392 11150
rect 10300 11082 10316 11137
rect 10376 11082 10392 11137
rect 10300 11065 10392 11082
rect 12245 11138 12302 11142
rect 12245 11078 12249 11138
rect 12298 11078 12302 11138
rect 12245 11074 12302 11078
rect 13444 11137 13536 11150
rect 13444 11082 13460 11137
rect 13520 11082 13536 11137
rect 13444 11065 13536 11082
rect 15447 11134 15504 11138
rect 15447 11074 15451 11134
rect 15500 11074 15504 11134
rect 15447 11070 15504 11074
rect 16646 11133 16738 11146
rect 16646 11078 16662 11133
rect 16722 11078 16738 11133
rect 16646 11061 16738 11078
rect 18591 11134 18648 11138
rect 18591 11074 18595 11134
rect 18644 11074 18648 11134
rect 18591 11070 18648 11074
rect 19790 11133 19882 11146
rect 19790 11078 19806 11133
rect 19866 11078 19882 11133
rect 19790 11061 19882 11078
rect 21723 11138 21780 11142
rect 21723 11078 21727 11138
rect 21776 11078 21780 11138
rect 21723 11074 21780 11078
rect 22922 11137 23014 11150
rect 22922 11082 22938 11137
rect 22998 11082 23014 11137
rect 22922 11065 23014 11082
rect 24867 11138 24924 11142
rect 24867 11078 24871 11138
rect 24920 11078 24924 11138
rect 24867 11074 24924 11078
rect 26066 11137 26158 11150
rect 26066 11082 26082 11137
rect 26142 11082 26158 11137
rect 26066 11065 26158 11082
rect 4289 10897 4323 10913
rect 4289 10847 4323 10863
rect 7433 10897 7467 10913
rect 7433 10847 7467 10863
rect 10565 10901 10599 10917
rect 10565 10851 10599 10867
rect 13709 10901 13743 10917
rect 13709 10851 13743 10867
rect 16911 10897 16945 10913
rect 16911 10847 16945 10863
rect 20055 10897 20089 10913
rect 20055 10847 20089 10863
rect 23187 10901 23221 10917
rect 23187 10851 23221 10867
rect 26331 10901 26365 10917
rect 26331 10851 26365 10867
rect 3802 10775 3836 10791
rect 3802 10583 3836 10599
rect 3920 10787 3954 10791
rect 3994 10787 4028 10791
rect 3920 10775 4028 10787
rect 3954 10599 3994 10775
rect 3920 10587 3994 10599
rect 3920 10583 3954 10587
rect 3994 10383 4028 10399
rect 4112 10775 4146 10791
rect 4112 10383 4146 10399
rect 4230 10775 4264 10791
rect 4230 10383 4264 10399
rect 4348 10775 4382 10791
rect 4348 10383 4382 10399
rect 4466 10787 4500 10791
rect 4544 10787 4578 10791
rect 4466 10775 4578 10787
rect 4500 10599 4544 10775
rect 4500 10587 4578 10599
rect 4544 10583 4578 10587
rect 4662 10775 4696 10791
rect 4662 10583 4696 10599
rect 6946 10775 6980 10791
rect 6946 10583 6980 10599
rect 7064 10787 7098 10791
rect 7138 10787 7172 10791
rect 7064 10775 7172 10787
rect 7098 10599 7138 10775
rect 7064 10587 7138 10599
rect 7064 10583 7098 10587
rect 4466 10383 4500 10399
rect 7138 10383 7172 10399
rect 7256 10775 7290 10791
rect 7256 10383 7290 10399
rect 7374 10775 7408 10791
rect 7374 10383 7408 10399
rect 7492 10775 7526 10791
rect 7492 10383 7526 10399
rect 7610 10787 7644 10791
rect 7688 10787 7722 10791
rect 7610 10775 7722 10787
rect 7644 10599 7688 10775
rect 7644 10587 7722 10599
rect 7688 10583 7722 10587
rect 7806 10775 7840 10791
rect 7806 10583 7840 10599
rect 10078 10779 10112 10795
rect 10078 10587 10112 10603
rect 10196 10791 10230 10795
rect 10270 10791 10304 10795
rect 10196 10779 10304 10791
rect 10230 10603 10270 10779
rect 10196 10591 10270 10603
rect 10196 10587 10230 10591
rect 7610 10383 7644 10399
rect 10270 10387 10304 10403
rect 10388 10779 10422 10795
rect 10388 10387 10422 10403
rect 10506 10779 10540 10795
rect 10506 10387 10540 10403
rect 10624 10779 10658 10795
rect 10624 10387 10658 10403
rect 10742 10791 10776 10795
rect 10820 10791 10854 10795
rect 10742 10779 10854 10791
rect 10776 10603 10820 10779
rect 10776 10591 10854 10603
rect 10820 10587 10854 10591
rect 10938 10779 10972 10795
rect 10938 10587 10972 10603
rect 13222 10779 13256 10795
rect 13222 10587 13256 10603
rect 13340 10791 13374 10795
rect 13414 10791 13448 10795
rect 13340 10779 13448 10791
rect 13374 10603 13414 10779
rect 13340 10591 13414 10603
rect 13340 10587 13374 10591
rect 10742 10387 10776 10403
rect 13414 10387 13448 10403
rect 13532 10779 13566 10795
rect 13532 10387 13566 10403
rect 13650 10779 13684 10795
rect 13650 10387 13684 10403
rect 13768 10779 13802 10795
rect 13768 10387 13802 10403
rect 13886 10791 13920 10795
rect 13964 10791 13998 10795
rect 13886 10779 13998 10791
rect 13920 10603 13964 10779
rect 13920 10591 13998 10603
rect 13964 10587 13998 10591
rect 14082 10779 14116 10795
rect 14082 10587 14116 10603
rect 16424 10775 16458 10791
rect 16424 10583 16458 10599
rect 16542 10787 16576 10791
rect 16616 10787 16650 10791
rect 16542 10775 16650 10787
rect 16576 10599 16616 10775
rect 16542 10587 16616 10599
rect 16542 10583 16576 10587
rect 13886 10387 13920 10403
rect 16616 10383 16650 10399
rect 16734 10775 16768 10791
rect 16734 10383 16768 10399
rect 16852 10775 16886 10791
rect 16852 10383 16886 10399
rect 16970 10775 17004 10791
rect 16970 10383 17004 10399
rect 17088 10787 17122 10791
rect 17166 10787 17200 10791
rect 17088 10775 17200 10787
rect 17122 10599 17166 10775
rect 17122 10587 17200 10599
rect 17166 10583 17200 10587
rect 17284 10775 17318 10791
rect 17284 10583 17318 10599
rect 19568 10775 19602 10791
rect 19568 10583 19602 10599
rect 19686 10787 19720 10791
rect 19760 10787 19794 10791
rect 19686 10775 19794 10787
rect 19720 10599 19760 10775
rect 19686 10587 19760 10599
rect 19686 10583 19720 10587
rect 17088 10383 17122 10399
rect 19760 10383 19794 10399
rect 19878 10775 19912 10791
rect 19878 10383 19912 10399
rect 19996 10775 20030 10791
rect 19996 10383 20030 10399
rect 20114 10775 20148 10791
rect 20114 10383 20148 10399
rect 20232 10787 20266 10791
rect 20310 10787 20344 10791
rect 20232 10775 20344 10787
rect 20266 10599 20310 10775
rect 20266 10587 20344 10599
rect 20310 10583 20344 10587
rect 20428 10775 20462 10791
rect 20428 10583 20462 10599
rect 22700 10779 22734 10795
rect 22700 10587 22734 10603
rect 22818 10791 22852 10795
rect 22892 10791 22926 10795
rect 22818 10779 22926 10791
rect 22852 10603 22892 10779
rect 22818 10591 22892 10603
rect 22818 10587 22852 10591
rect 20232 10383 20266 10399
rect 22892 10387 22926 10403
rect 23010 10779 23044 10795
rect 23010 10387 23044 10403
rect 23128 10779 23162 10795
rect 23128 10387 23162 10403
rect 23246 10779 23280 10795
rect 23246 10387 23280 10403
rect 23364 10791 23398 10795
rect 23442 10791 23476 10795
rect 23364 10779 23476 10791
rect 23398 10603 23442 10779
rect 23398 10591 23476 10603
rect 23442 10587 23476 10591
rect 23560 10779 23594 10795
rect 23560 10587 23594 10603
rect 25844 10779 25878 10795
rect 25844 10587 25878 10603
rect 25962 10791 25996 10795
rect 26036 10791 26070 10795
rect 25962 10779 26070 10791
rect 25996 10603 26036 10779
rect 25962 10591 26036 10603
rect 25962 10587 25996 10591
rect 23364 10387 23398 10403
rect 26036 10387 26070 10403
rect 26154 10779 26188 10795
rect 26154 10387 26188 10403
rect 26272 10779 26306 10795
rect 26272 10387 26306 10403
rect 26390 10779 26424 10795
rect 26390 10387 26424 10403
rect 26508 10791 26542 10795
rect 26586 10791 26620 10795
rect 26508 10779 26620 10791
rect 26542 10603 26586 10779
rect 26542 10591 26620 10603
rect 26586 10587 26620 10591
rect 26704 10779 26738 10795
rect 26704 10587 26738 10603
rect 26508 10387 26542 10403
rect 4215 10264 4231 10298
rect 4265 10264 4281 10298
rect 7359 10264 7375 10298
rect 7409 10264 7425 10298
rect 10491 10268 10507 10302
rect 10541 10268 10557 10302
rect 13635 10268 13651 10302
rect 13685 10268 13701 10302
rect 16837 10264 16853 10298
rect 16887 10264 16903 10298
rect 19981 10264 19997 10298
rect 20031 10264 20047 10298
rect 23113 10268 23129 10302
rect 23163 10268 23179 10302
rect 26257 10268 26273 10302
rect 26307 10268 26323 10302
rect 10472 10150 10608 10154
rect 4196 10146 4332 10150
rect 4196 10132 4234 10146
rect 4292 10132 4332 10146
rect 4196 10086 4212 10132
rect 4316 10086 4332 10132
rect 4196 10064 4332 10086
rect 7340 10146 7476 10150
rect 7340 10132 7378 10146
rect 7436 10132 7476 10146
rect 7340 10086 7356 10132
rect 7460 10086 7476 10132
rect 7340 10064 7476 10086
rect 10472 10136 10510 10150
rect 10568 10136 10608 10150
rect 10472 10090 10488 10136
rect 10592 10090 10608 10136
rect 10472 10068 10608 10090
rect 13616 10150 13752 10154
rect 23094 10150 23230 10154
rect 13616 10136 13654 10150
rect 13712 10136 13752 10150
rect 13616 10090 13632 10136
rect 13736 10090 13752 10136
rect 13616 10068 13752 10090
rect 16818 10146 16954 10150
rect 16818 10132 16856 10146
rect 16914 10132 16954 10146
rect 16818 10086 16834 10132
rect 16938 10086 16954 10132
rect 16818 10064 16954 10086
rect 19962 10146 20098 10150
rect 19962 10132 20000 10146
rect 20058 10132 20098 10146
rect 19962 10086 19978 10132
rect 20082 10086 20098 10132
rect 19962 10064 20098 10086
rect 23094 10136 23132 10150
rect 23190 10136 23230 10150
rect 23094 10090 23110 10136
rect 23214 10090 23230 10136
rect 23094 10068 23230 10090
rect 26238 10150 26374 10154
rect 26238 10136 26276 10150
rect 26334 10136 26374 10150
rect 26238 10090 26254 10136
rect 26358 10090 26374 10136
rect 26238 10068 26374 10090
rect 4128 9646 4356 9664
rect 4128 9570 4144 9646
rect 4340 9570 4356 9646
rect 4128 9554 4356 9570
rect 7272 9646 7500 9664
rect 7272 9570 7288 9646
rect 7484 9570 7500 9646
rect 7272 9554 7500 9570
rect 10404 9650 10632 9668
rect 10404 9574 10420 9650
rect 10616 9574 10632 9650
rect 10404 9558 10632 9574
rect 13548 9650 13776 9668
rect 13548 9574 13564 9650
rect 13760 9574 13776 9650
rect 13548 9558 13776 9574
rect 16750 9646 16978 9664
rect 16750 9570 16766 9646
rect 16962 9570 16978 9646
rect 16750 9554 16978 9570
rect 19894 9646 20122 9664
rect 19894 9570 19910 9646
rect 20106 9570 20122 9646
rect 19894 9554 20122 9570
rect 23026 9650 23254 9668
rect 23026 9574 23042 9650
rect 23238 9574 23254 9650
rect 23026 9558 23254 9574
rect 26170 9650 26398 9668
rect 26170 9574 26186 9650
rect 26382 9574 26398 9650
rect 26170 9558 26398 9574
rect 3399 9429 3669 9468
rect 3399 9376 3433 9429
rect 2958 9227 3228 9266
rect 2958 9176 2992 9227
rect 2958 8984 2992 9000
rect 3076 9176 3110 9192
rect 3076 8949 3110 9000
rect 3194 9176 3228 9227
rect 3194 8984 3228 9000
rect 3312 9176 3346 9192
rect 3312 8949 3346 9000
rect 3399 8984 3433 9000
rect 3517 9376 3551 9392
rect 3076 8910 3346 8949
rect 3517 8949 3551 9000
rect 3635 9376 3669 9429
rect 3866 9428 4136 9467
rect 3635 8984 3669 9000
rect 3753 9376 3787 9392
rect 3753 8949 3787 9000
rect 3866 9376 3900 9428
rect 3866 8984 3900 9000
rect 3984 9376 4018 9392
rect 3984 8949 4018 9000
rect 4102 9376 4136 9428
rect 4338 9428 4608 9467
rect 4102 8984 4136 9000
rect 4220 9376 4254 9392
rect 4220 8949 4254 9000
rect 4338 9376 4372 9428
rect 4338 8984 4372 9000
rect 4456 9376 4490 9392
rect 4456 8949 4490 9000
rect 4574 9376 4608 9428
rect 4811 9428 5081 9467
rect 4574 8984 4608 9000
rect 4693 9376 4727 9392
rect 4693 8949 4727 9000
rect 4811 9376 4845 9428
rect 4811 8984 4845 9000
rect 4929 9376 4963 9392
rect 4929 8949 4963 9000
rect 5047 9376 5081 9428
rect 6543 9429 6813 9468
rect 6543 9376 6577 9429
rect 5284 9226 5554 9263
rect 5047 8984 5081 9000
rect 5166 9176 5200 9192
rect 3517 8910 4963 8949
rect 5166 8946 5200 9000
rect 5284 9176 5318 9226
rect 5284 8984 5318 9000
rect 5402 9176 5436 9192
rect 5402 8946 5436 9000
rect 5520 9176 5554 9226
rect 5520 8984 5554 9000
rect 6102 9227 6372 9266
rect 6102 9176 6136 9227
rect 6102 8984 6136 9000
rect 6220 9176 6254 9192
rect 5166 8907 5436 8946
rect 6220 8949 6254 9000
rect 6338 9176 6372 9227
rect 6338 8984 6372 9000
rect 6456 9176 6490 9192
rect 6456 8949 6490 9000
rect 6543 8984 6577 9000
rect 6661 9376 6695 9392
rect 6220 8910 6490 8949
rect 6661 8949 6695 9000
rect 6779 9376 6813 9429
rect 7010 9428 7280 9467
rect 6779 8984 6813 9000
rect 6897 9376 6931 9392
rect 6897 8949 6931 9000
rect 7010 9376 7044 9428
rect 7010 8984 7044 9000
rect 7128 9376 7162 9392
rect 7128 8949 7162 9000
rect 7246 9376 7280 9428
rect 7482 9428 7752 9467
rect 7246 8984 7280 9000
rect 7364 9376 7398 9392
rect 7364 8949 7398 9000
rect 7482 9376 7516 9428
rect 7482 8984 7516 9000
rect 7600 9376 7634 9392
rect 7600 8949 7634 9000
rect 7718 9376 7752 9428
rect 7955 9428 8225 9467
rect 7718 8984 7752 9000
rect 7837 9376 7871 9392
rect 7837 8949 7871 9000
rect 7955 9376 7989 9428
rect 7955 8984 7989 9000
rect 8073 9376 8107 9392
rect 8073 8949 8107 9000
rect 8191 9376 8225 9428
rect 9675 9433 9945 9472
rect 9675 9380 9709 9433
rect 8428 9226 8698 9263
rect 8191 8984 8225 9000
rect 8310 9176 8344 9192
rect 6661 8910 8107 8949
rect 8310 8946 8344 9000
rect 8428 9176 8462 9226
rect 8428 8984 8462 9000
rect 8546 9176 8580 9192
rect 8546 8946 8580 9000
rect 8664 9176 8698 9226
rect 8664 8984 8698 9000
rect 9234 9231 9504 9270
rect 9234 9180 9268 9231
rect 9234 8988 9268 9004
rect 9352 9180 9386 9196
rect 8310 8907 8580 8946
rect 9352 8953 9386 9004
rect 9470 9180 9504 9231
rect 9470 8988 9504 9004
rect 9588 9180 9622 9196
rect 9588 8953 9622 9004
rect 9675 8988 9709 9004
rect 9793 9380 9827 9396
rect 9352 8914 9622 8953
rect 9793 8953 9827 9004
rect 9911 9380 9945 9433
rect 10142 9432 10412 9471
rect 9911 8988 9945 9004
rect 10029 9380 10063 9396
rect 10029 8953 10063 9004
rect 10142 9380 10176 9432
rect 10142 8988 10176 9004
rect 10260 9380 10294 9396
rect 10260 8953 10294 9004
rect 10378 9380 10412 9432
rect 10614 9432 10884 9471
rect 10378 8988 10412 9004
rect 10496 9380 10530 9396
rect 10496 8953 10530 9004
rect 10614 9380 10648 9432
rect 10614 8988 10648 9004
rect 10732 9380 10766 9396
rect 10732 8953 10766 9004
rect 10850 9380 10884 9432
rect 11087 9432 11357 9471
rect 10850 8988 10884 9004
rect 10969 9380 11003 9396
rect 10969 8953 11003 9004
rect 11087 9380 11121 9432
rect 11087 8988 11121 9004
rect 11205 9380 11239 9396
rect 11205 8953 11239 9004
rect 11323 9380 11357 9432
rect 12819 9433 13089 9472
rect 12819 9380 12853 9433
rect 11560 9230 11830 9267
rect 11323 8988 11357 9004
rect 11442 9180 11476 9196
rect 9793 8914 11239 8953
rect 11442 8950 11476 9004
rect 11560 9180 11594 9230
rect 11560 8988 11594 9004
rect 11678 9180 11712 9196
rect 11678 8950 11712 9004
rect 11796 9180 11830 9230
rect 11796 8988 11830 9004
rect 12378 9231 12648 9270
rect 12378 9180 12412 9231
rect 12378 8988 12412 9004
rect 12496 9180 12530 9196
rect 11442 8911 11712 8950
rect 12496 8953 12530 9004
rect 12614 9180 12648 9231
rect 12614 8988 12648 9004
rect 12732 9180 12766 9196
rect 12732 8953 12766 9004
rect 12819 8988 12853 9004
rect 12937 9380 12971 9396
rect 12496 8914 12766 8953
rect 12937 8953 12971 9004
rect 13055 9380 13089 9433
rect 13286 9432 13556 9471
rect 13055 8988 13089 9004
rect 13173 9380 13207 9396
rect 13173 8953 13207 9004
rect 13286 9380 13320 9432
rect 13286 8988 13320 9004
rect 13404 9380 13438 9396
rect 13404 8953 13438 9004
rect 13522 9380 13556 9432
rect 13758 9432 14028 9471
rect 13522 8988 13556 9004
rect 13640 9380 13674 9396
rect 13640 8953 13674 9004
rect 13758 9380 13792 9432
rect 13758 8988 13792 9004
rect 13876 9380 13910 9396
rect 13876 8953 13910 9004
rect 13994 9380 14028 9432
rect 14231 9432 14501 9471
rect 13994 8988 14028 9004
rect 14113 9380 14147 9396
rect 14113 8953 14147 9004
rect 14231 9380 14265 9432
rect 14231 8988 14265 9004
rect 14349 9380 14383 9396
rect 14349 8953 14383 9004
rect 14467 9380 14501 9432
rect 16021 9429 16291 9468
rect 16021 9376 16055 9429
rect 14704 9230 14974 9267
rect 14467 8988 14501 9004
rect 14586 9180 14620 9196
rect 12937 8914 14383 8953
rect 14586 8950 14620 9004
rect 14704 9180 14738 9230
rect 14704 8988 14738 9004
rect 14822 9180 14856 9196
rect 14822 8950 14856 9004
rect 14940 9180 14974 9230
rect 14940 8988 14974 9004
rect 15580 9227 15850 9266
rect 15580 9176 15614 9227
rect 15580 8984 15614 9000
rect 15698 9176 15732 9192
rect 14586 8911 14856 8950
rect 15698 8949 15732 9000
rect 15816 9176 15850 9227
rect 15816 8984 15850 9000
rect 15934 9176 15968 9192
rect 15934 8949 15968 9000
rect 16021 8984 16055 9000
rect 16139 9376 16173 9392
rect 15698 8910 15968 8949
rect 16139 8949 16173 9000
rect 16257 9376 16291 9429
rect 16488 9428 16758 9467
rect 16257 8984 16291 9000
rect 16375 9376 16409 9392
rect 16375 8949 16409 9000
rect 16488 9376 16522 9428
rect 16488 8984 16522 9000
rect 16606 9376 16640 9392
rect 16606 8949 16640 9000
rect 16724 9376 16758 9428
rect 16960 9428 17230 9467
rect 16724 8984 16758 9000
rect 16842 9376 16876 9392
rect 16842 8949 16876 9000
rect 16960 9376 16994 9428
rect 16960 8984 16994 9000
rect 17078 9376 17112 9392
rect 17078 8949 17112 9000
rect 17196 9376 17230 9428
rect 17433 9428 17703 9467
rect 17196 8984 17230 9000
rect 17315 9376 17349 9392
rect 17315 8949 17349 9000
rect 17433 9376 17467 9428
rect 17433 8984 17467 9000
rect 17551 9376 17585 9392
rect 17551 8949 17585 9000
rect 17669 9376 17703 9428
rect 19165 9429 19435 9468
rect 19165 9376 19199 9429
rect 17906 9226 18176 9263
rect 17669 8984 17703 9000
rect 17788 9176 17822 9192
rect 16139 8910 17585 8949
rect 17788 8946 17822 9000
rect 17906 9176 17940 9226
rect 17906 8984 17940 9000
rect 18024 9176 18058 9192
rect 18024 8946 18058 9000
rect 18142 9176 18176 9226
rect 18142 8984 18176 9000
rect 18724 9227 18994 9266
rect 18724 9176 18758 9227
rect 18724 8984 18758 9000
rect 18842 9176 18876 9192
rect 17788 8907 18058 8946
rect 18842 8949 18876 9000
rect 18960 9176 18994 9227
rect 18960 8984 18994 9000
rect 19078 9176 19112 9192
rect 19078 8949 19112 9000
rect 19165 8984 19199 9000
rect 19283 9376 19317 9392
rect 18842 8910 19112 8949
rect 19283 8949 19317 9000
rect 19401 9376 19435 9429
rect 19632 9428 19902 9467
rect 19401 8984 19435 9000
rect 19519 9376 19553 9392
rect 19519 8949 19553 9000
rect 19632 9376 19666 9428
rect 19632 8984 19666 9000
rect 19750 9376 19784 9392
rect 19750 8949 19784 9000
rect 19868 9376 19902 9428
rect 20104 9428 20374 9467
rect 19868 8984 19902 9000
rect 19986 9376 20020 9392
rect 19986 8949 20020 9000
rect 20104 9376 20138 9428
rect 20104 8984 20138 9000
rect 20222 9376 20256 9392
rect 20222 8949 20256 9000
rect 20340 9376 20374 9428
rect 20577 9428 20847 9467
rect 20340 8984 20374 9000
rect 20459 9376 20493 9392
rect 20459 8949 20493 9000
rect 20577 9376 20611 9428
rect 20577 8984 20611 9000
rect 20695 9376 20729 9392
rect 20695 8949 20729 9000
rect 20813 9376 20847 9428
rect 22297 9433 22567 9472
rect 22297 9380 22331 9433
rect 21050 9226 21320 9263
rect 20813 8984 20847 9000
rect 20932 9176 20966 9192
rect 19283 8910 20729 8949
rect 20932 8946 20966 9000
rect 21050 9176 21084 9226
rect 21050 8984 21084 9000
rect 21168 9176 21202 9192
rect 21168 8946 21202 9000
rect 21286 9176 21320 9226
rect 21286 8984 21320 9000
rect 21856 9231 22126 9270
rect 21856 9180 21890 9231
rect 21856 8988 21890 9004
rect 21974 9180 22008 9196
rect 20932 8907 21202 8946
rect 21974 8953 22008 9004
rect 22092 9180 22126 9231
rect 22092 8988 22126 9004
rect 22210 9180 22244 9196
rect 22210 8953 22244 9004
rect 22297 8988 22331 9004
rect 22415 9380 22449 9396
rect 21974 8914 22244 8953
rect 22415 8953 22449 9004
rect 22533 9380 22567 9433
rect 22764 9432 23034 9471
rect 22533 8988 22567 9004
rect 22651 9380 22685 9396
rect 22651 8953 22685 9004
rect 22764 9380 22798 9432
rect 22764 8988 22798 9004
rect 22882 9380 22916 9396
rect 22882 8953 22916 9004
rect 23000 9380 23034 9432
rect 23236 9432 23506 9471
rect 23000 8988 23034 9004
rect 23118 9380 23152 9396
rect 23118 8953 23152 9004
rect 23236 9380 23270 9432
rect 23236 8988 23270 9004
rect 23354 9380 23388 9396
rect 23354 8953 23388 9004
rect 23472 9380 23506 9432
rect 23709 9432 23979 9471
rect 23472 8988 23506 9004
rect 23591 9380 23625 9396
rect 23591 8953 23625 9004
rect 23709 9380 23743 9432
rect 23709 8988 23743 9004
rect 23827 9380 23861 9396
rect 23827 8953 23861 9004
rect 23945 9380 23979 9432
rect 25441 9433 25711 9472
rect 25441 9380 25475 9433
rect 24182 9230 24452 9267
rect 23945 8988 23979 9004
rect 24064 9180 24098 9196
rect 22415 8914 23861 8953
rect 24064 8950 24098 9004
rect 24182 9180 24216 9230
rect 24182 8988 24216 9004
rect 24300 9180 24334 9196
rect 24300 8950 24334 9004
rect 24418 9180 24452 9230
rect 24418 8988 24452 9004
rect 25000 9231 25270 9270
rect 25000 9180 25034 9231
rect 25000 8988 25034 9004
rect 25118 9180 25152 9196
rect 24064 8911 24334 8950
rect 25118 8953 25152 9004
rect 25236 9180 25270 9231
rect 25236 8988 25270 9004
rect 25354 9180 25388 9196
rect 25354 8953 25388 9004
rect 25441 8988 25475 9004
rect 25559 9380 25593 9396
rect 25118 8914 25388 8953
rect 25559 8953 25593 9004
rect 25677 9380 25711 9433
rect 25908 9432 26178 9471
rect 25677 8988 25711 9004
rect 25795 9380 25829 9396
rect 25795 8953 25829 9004
rect 25908 9380 25942 9432
rect 25908 8988 25942 9004
rect 26026 9380 26060 9396
rect 26026 8953 26060 9004
rect 26144 9380 26178 9432
rect 26380 9432 26650 9471
rect 26144 8988 26178 9004
rect 26262 9380 26296 9396
rect 26262 8953 26296 9004
rect 26380 9380 26414 9432
rect 26380 8988 26414 9004
rect 26498 9380 26532 9396
rect 26498 8953 26532 9004
rect 26616 9380 26650 9432
rect 26853 9432 27123 9471
rect 26616 8988 26650 9004
rect 26735 9380 26769 9396
rect 26735 8953 26769 9004
rect 26853 9380 26887 9432
rect 26853 8988 26887 9004
rect 26971 9380 27005 9396
rect 26971 8953 27005 9004
rect 27089 9380 27123 9432
rect 27326 9230 27596 9267
rect 27089 8988 27123 9004
rect 27208 9180 27242 9196
rect 25559 8914 27005 8953
rect 27208 8950 27242 9004
rect 27326 9180 27360 9230
rect 27326 8988 27360 9004
rect 27444 9180 27478 9196
rect 27444 8950 27478 9004
rect 27562 9180 27596 9230
rect 27562 8988 27596 9004
rect 27208 8911 27478 8950
rect 4044 8785 4078 8801
rect 5338 8792 5354 8826
rect 5388 8792 5404 8826
rect 4044 8735 4078 8751
rect 7188 8785 7222 8801
rect 8482 8792 8498 8826
rect 8532 8792 8548 8826
rect 7188 8735 7222 8751
rect 10320 8789 10354 8805
rect 11614 8796 11630 8830
rect 11664 8796 11680 8830
rect 10320 8739 10354 8755
rect 13464 8789 13498 8805
rect 14758 8796 14774 8830
rect 14808 8796 14824 8830
rect 13464 8739 13498 8755
rect 16666 8785 16700 8801
rect 17960 8792 17976 8826
rect 18010 8792 18026 8826
rect 16666 8735 16700 8751
rect 19810 8785 19844 8801
rect 21104 8792 21120 8826
rect 21154 8792 21170 8826
rect 19810 8735 19844 8751
rect 22942 8789 22976 8805
rect 24236 8796 24252 8830
rect 24286 8796 24302 8830
rect 22942 8739 22976 8755
rect 26086 8789 26120 8805
rect 27380 8796 27396 8830
rect 27430 8796 27446 8830
rect 26086 8739 26120 8755
rect 2815 8686 2872 8690
rect 2815 8626 2819 8686
rect 2868 8626 2872 8686
rect 2815 8622 2872 8626
rect 3047 8685 3139 8702
rect 3047 8630 3063 8685
rect 3123 8630 3139 8685
rect 3047 8617 3139 8630
rect 4132 8686 4224 8699
rect 4132 8631 4148 8686
rect 4208 8631 4224 8686
rect 4132 8614 4224 8631
rect 5959 8686 6016 8690
rect 5959 8626 5963 8686
rect 6012 8626 6016 8686
rect 5959 8622 6016 8626
rect 6191 8685 6283 8702
rect 6191 8630 6207 8685
rect 6267 8630 6283 8685
rect 6191 8617 6283 8630
rect 7276 8686 7368 8699
rect 7276 8631 7292 8686
rect 7352 8631 7368 8686
rect 7276 8614 7368 8631
rect 9091 8690 9148 8694
rect 9091 8630 9095 8690
rect 9144 8630 9148 8690
rect 9091 8626 9148 8630
rect 9323 8689 9415 8706
rect 9323 8634 9339 8689
rect 9399 8634 9415 8689
rect 9323 8621 9415 8634
rect 10408 8690 10500 8703
rect 10408 8635 10424 8690
rect 10484 8635 10500 8690
rect 10408 8618 10500 8635
rect 12235 8690 12292 8694
rect 12235 8630 12239 8690
rect 12288 8630 12292 8690
rect 12235 8626 12292 8630
rect 12467 8689 12559 8706
rect 12467 8634 12483 8689
rect 12543 8634 12559 8689
rect 12467 8621 12559 8634
rect 13552 8690 13644 8703
rect 13552 8635 13568 8690
rect 13628 8635 13644 8690
rect 13552 8618 13644 8635
rect 15437 8686 15494 8690
rect 15437 8626 15441 8686
rect 15490 8626 15494 8686
rect 15437 8622 15494 8626
rect 15669 8685 15761 8702
rect 15669 8630 15685 8685
rect 15745 8630 15761 8685
rect 15669 8617 15761 8630
rect 16754 8686 16846 8699
rect 16754 8631 16770 8686
rect 16830 8631 16846 8686
rect 16754 8614 16846 8631
rect 18581 8686 18638 8690
rect 18581 8626 18585 8686
rect 18634 8626 18638 8686
rect 18581 8622 18638 8626
rect 18813 8685 18905 8702
rect 18813 8630 18829 8685
rect 18889 8630 18905 8685
rect 18813 8617 18905 8630
rect 19898 8686 19990 8699
rect 19898 8631 19914 8686
rect 19974 8631 19990 8686
rect 19898 8614 19990 8631
rect 21713 8690 21770 8694
rect 21713 8630 21717 8690
rect 21766 8630 21770 8690
rect 21713 8626 21770 8630
rect 21945 8689 22037 8706
rect 21945 8634 21961 8689
rect 22021 8634 22037 8689
rect 21945 8621 22037 8634
rect 23030 8690 23122 8703
rect 23030 8635 23046 8690
rect 23106 8635 23122 8690
rect 23030 8618 23122 8635
rect 24857 8690 24914 8694
rect 24857 8630 24861 8690
rect 24910 8630 24914 8690
rect 24857 8626 24914 8630
rect 25089 8689 25181 8706
rect 25089 8634 25105 8689
rect 25165 8634 25181 8689
rect 25089 8621 25181 8634
rect 26174 8690 26266 8703
rect 26174 8635 26190 8690
rect 26250 8635 26266 8690
rect 26174 8618 26266 8635
rect 9091 8576 9148 8578
rect 8893 8574 9148 8576
rect 12235 8575 12292 8578
rect 21713 8576 21770 8578
rect 2535 8570 2651 8571
rect 2815 8570 2872 8574
rect 5959 8572 6016 8574
rect 2535 8510 2819 8570
rect 2868 8510 2872 8570
rect 2535 8506 2872 8510
rect 4398 8555 4432 8571
rect 2536 6944 2600 8506
rect 4398 8505 4432 8521
rect 5763 8570 6016 8572
rect 5763 8510 5963 8570
rect 6012 8510 6016 8570
rect 5763 8508 6016 8510
rect 2815 8402 2872 8406
rect 2815 8342 2819 8402
rect 2868 8342 2872 8402
rect 2815 8338 2872 8342
rect 4014 8401 4106 8414
rect 4014 8346 4030 8401
rect 4090 8346 4106 8401
rect 4014 8329 4106 8346
rect 4279 8165 4313 8181
rect 4279 8115 4313 8131
rect 3792 8043 3826 8059
rect 3792 7851 3826 7867
rect 3910 8055 3944 8059
rect 3984 8055 4018 8059
rect 3910 8043 4018 8055
rect 3944 7867 3984 8043
rect 3910 7855 3984 7867
rect 3910 7851 3944 7855
rect 3984 7651 4018 7667
rect 4102 8043 4136 8059
rect 4102 7651 4136 7667
rect 4220 8043 4254 8059
rect 4220 7651 4254 7667
rect 4338 8043 4372 8059
rect 4338 7651 4372 7667
rect 4456 8055 4490 8059
rect 4534 8055 4568 8059
rect 4456 8043 4568 8055
rect 4490 7867 4534 8043
rect 4490 7855 4568 7867
rect 4534 7851 4568 7855
rect 4652 8043 4686 8059
rect 4652 7851 4686 7867
rect 4456 7651 4490 7667
rect 4205 7532 4221 7566
rect 4255 7532 4271 7566
rect 4186 7414 4322 7418
rect 4186 7400 4224 7414
rect 4282 7400 4322 7414
rect 4186 7354 4202 7400
rect 4306 7354 4322 7400
rect 4186 7332 4322 7354
rect 2536 6880 4535 6944
rect 3446 6702 3648 6722
rect 3446 6658 3480 6702
rect 3602 6658 3648 6702
rect 3446 6648 3532 6658
rect 3570 6648 3648 6658
rect 3446 6630 3648 6648
rect 3533 6484 3803 6519
rect 3179 6431 3213 6447
rect 2695 6285 2965 6320
rect 2695 6231 2729 6285
rect 2695 6039 2729 6055
rect 2813 6231 2847 6247
rect 2813 6039 2847 6055
rect 2931 6231 2965 6285
rect 2931 6039 2965 6055
rect 3049 6231 3083 6247
rect 3049 6039 3083 6055
rect 3179 6039 3213 6055
rect 3297 6431 3331 6447
rect 3297 6039 3331 6055
rect 3415 6431 3449 6447
rect 3415 6039 3449 6055
rect 3533 6431 3567 6484
rect 3533 6039 3567 6055
rect 3651 6431 3685 6447
rect 3651 6039 3685 6055
rect 3769 6431 3803 6484
rect 3769 6039 3803 6055
rect 3887 6431 3921 6447
rect 3887 6039 3921 6055
rect 4016 6231 4050 6247
rect 4016 6039 4050 6055
rect 4134 6231 4168 6247
rect 4134 6039 4168 6055
rect 4252 6231 4286 6247
rect 4252 6039 4286 6055
rect 4370 6231 4404 6247
rect 4370 6039 4404 6055
rect 4096 5842 4102 5876
rect 4156 5842 4162 5876
rect 3122 5738 3156 5754
rect 2665 5636 2702 5696
rect 2665 5580 2730 5636
rect 2665 4154 2729 5580
rect 3240 5738 3274 5754
rect 3122 5346 3156 5362
rect 3239 5362 3240 5409
rect 3358 5738 3392 5754
rect 3274 5362 3275 5409
rect 3239 5304 3275 5362
rect 3476 5738 3510 5754
rect 3358 5346 3392 5362
rect 3474 5362 3476 5409
rect 3474 5304 3510 5362
rect 3594 5738 3628 5754
rect 3594 5346 3628 5362
rect 3712 5738 3746 5754
rect 3830 5738 3864 5754
rect 3746 5362 3748 5408
rect 3712 5304 3748 5362
rect 3830 5346 3864 5362
rect 3239 5264 4334 5304
rect 3258 5263 4334 5264
rect 3136 5174 3203 5190
rect 3136 5140 3152 5174
rect 3186 5140 3203 5174
rect 3136 5124 3203 5140
rect 2967 5107 3001 5123
rect 2967 5057 3001 5073
rect 3313 5022 3347 5263
rect 4471 5317 4535 6880
rect 5763 6928 5827 8508
rect 5959 8506 6016 8508
rect 7542 8555 7576 8571
rect 7542 8505 7576 8521
rect 8893 8514 9095 8574
rect 9144 8514 9148 8574
rect 8893 8512 9148 8514
rect 5959 8402 6016 8406
rect 5959 8342 5963 8402
rect 6012 8342 6016 8402
rect 5959 8338 6016 8342
rect 7158 8401 7250 8414
rect 7158 8346 7174 8401
rect 7234 8346 7250 8401
rect 7158 8329 7250 8346
rect 7423 8165 7457 8181
rect 7423 8115 7457 8131
rect 8893 8072 8957 8512
rect 9091 8510 9148 8512
rect 10674 8559 10708 8575
rect 10674 8509 10708 8525
rect 12019 8574 12292 8575
rect 12019 8514 12239 8574
rect 12288 8514 12292 8574
rect 12019 8511 12292 8514
rect 9091 8406 9148 8410
rect 9091 8346 9095 8406
rect 9144 8346 9148 8406
rect 9091 8342 9148 8346
rect 10290 8405 10382 8418
rect 10290 8350 10306 8405
rect 10366 8350 10382 8405
rect 10290 8333 10382 8350
rect 10555 8169 10589 8185
rect 10555 8119 10589 8135
rect 6936 8043 6970 8059
rect 6936 7851 6970 7867
rect 7054 8055 7088 8059
rect 7128 8055 7162 8059
rect 7054 8043 7162 8055
rect 7088 7867 7128 8043
rect 7054 7855 7128 7867
rect 7054 7851 7088 7855
rect 7128 7651 7162 7667
rect 7246 8043 7280 8059
rect 7246 7651 7280 7667
rect 7364 8043 7398 8059
rect 7364 7651 7398 7667
rect 7482 8043 7516 8059
rect 7482 7651 7516 7667
rect 7600 8055 7634 8059
rect 7678 8055 7712 8059
rect 7600 8043 7712 8055
rect 7634 7867 7678 8043
rect 7634 7855 7712 7867
rect 7678 7851 7712 7855
rect 7796 8043 7830 8059
rect 7796 7851 7830 7867
rect 8632 8008 8957 8072
rect 10068 8047 10102 8063
rect 7600 7651 7634 7667
rect 7349 7532 7365 7566
rect 7399 7532 7415 7566
rect 7330 7414 7466 7418
rect 7330 7400 7368 7414
rect 7426 7400 7466 7414
rect 7330 7354 7346 7400
rect 7450 7354 7466 7400
rect 7330 7332 7466 7354
rect 5763 6864 6601 6928
rect 5514 6704 5716 6724
rect 5514 6660 5548 6704
rect 5670 6660 5716 6704
rect 5514 6650 5600 6660
rect 5638 6650 5716 6660
rect 5514 6632 5716 6650
rect 5601 6486 5871 6521
rect 5247 6433 5281 6449
rect 4763 6287 5033 6322
rect 4763 6233 4797 6287
rect 4763 6041 4797 6057
rect 4881 6233 4915 6249
rect 4881 6041 4915 6057
rect 4999 6233 5033 6287
rect 4999 6041 5033 6057
rect 5117 6233 5151 6249
rect 5117 6041 5151 6057
rect 5247 6041 5281 6057
rect 5365 6433 5399 6449
rect 5365 6041 5399 6057
rect 5483 6433 5517 6449
rect 5483 6041 5517 6057
rect 5601 6433 5635 6486
rect 5601 6041 5635 6057
rect 5719 6433 5753 6449
rect 5719 6041 5753 6057
rect 5837 6433 5871 6486
rect 5837 6041 5871 6057
rect 5955 6433 5989 6449
rect 5955 6041 5989 6057
rect 6084 6233 6118 6249
rect 6084 6041 6118 6057
rect 6202 6233 6236 6249
rect 6202 6041 6236 6057
rect 6320 6233 6354 6249
rect 6320 6041 6354 6057
rect 6438 6233 6472 6249
rect 6438 6041 6472 6057
rect 6164 5844 6170 5878
rect 6224 5844 6230 5878
rect 5190 5740 5224 5756
rect 5308 5740 5342 5756
rect 5190 5348 5224 5364
rect 5307 5364 5308 5411
rect 5426 5740 5460 5756
rect 5342 5364 5343 5411
rect 4436 5253 4535 5317
rect 5307 5306 5343 5364
rect 5544 5740 5578 5756
rect 5426 5348 5460 5364
rect 5542 5364 5544 5411
rect 5542 5306 5578 5364
rect 5662 5740 5696 5756
rect 5662 5348 5696 5364
rect 5780 5740 5814 5756
rect 5898 5740 5932 5756
rect 5814 5364 5816 5410
rect 5780 5306 5816 5364
rect 5898 5348 5932 5364
rect 5307 5266 6402 5306
rect 5326 5265 6402 5266
rect 3783 5174 3850 5190
rect 3783 5140 3800 5174
rect 3834 5140 3850 5174
rect 3783 5124 3850 5140
rect 5204 5176 5271 5192
rect 5204 5142 5220 5176
rect 5254 5142 5271 5176
rect 5204 5126 5271 5142
rect 4090 5106 4124 5122
rect 3402 5056 3418 5090
rect 3452 5056 3468 5090
rect 3520 5057 3536 5091
rect 3570 5057 3586 5091
rect 4090 5056 4124 5072
rect 5035 5109 5069 5125
rect 5035 5059 5069 5075
rect 5381 5024 5415 5265
rect 6544 5306 6600 6864
rect 7583 6702 7785 6722
rect 7583 6658 7617 6702
rect 7739 6658 7785 6702
rect 7583 6648 7669 6658
rect 7707 6648 7785 6658
rect 7583 6630 7785 6648
rect 7670 6484 7940 6519
rect 7316 6431 7350 6447
rect 6832 6285 7102 6320
rect 6832 6231 6866 6285
rect 6832 6039 6866 6055
rect 6950 6231 6984 6247
rect 6950 6039 6984 6055
rect 7068 6231 7102 6285
rect 7068 6039 7102 6055
rect 7186 6231 7220 6247
rect 7186 6039 7220 6055
rect 7316 6039 7350 6055
rect 7434 6431 7468 6447
rect 7434 6039 7468 6055
rect 7552 6431 7586 6447
rect 7552 6039 7586 6055
rect 7670 6431 7704 6484
rect 7670 6039 7704 6055
rect 7788 6431 7822 6447
rect 7788 6039 7822 6055
rect 7906 6431 7940 6484
rect 7906 6039 7940 6055
rect 8024 6431 8058 6447
rect 8024 6039 8058 6055
rect 8153 6231 8187 6247
rect 8153 6039 8187 6055
rect 8271 6231 8305 6247
rect 8271 6039 8305 6055
rect 8389 6231 8423 6247
rect 8389 6039 8423 6055
rect 8507 6231 8541 6247
rect 8507 6039 8541 6055
rect 8233 5842 8239 5876
rect 8293 5842 8299 5876
rect 7259 5738 7293 5754
rect 7377 5738 7411 5754
rect 7259 5346 7293 5362
rect 7376 5362 7377 5409
rect 7495 5738 7529 5754
rect 7411 5362 7412 5409
rect 6504 5265 6600 5306
rect 7376 5304 7412 5362
rect 7613 5738 7647 5754
rect 7495 5346 7529 5362
rect 7611 5362 7613 5409
rect 7611 5304 7647 5362
rect 7731 5738 7765 5754
rect 7731 5346 7765 5362
rect 7849 5738 7883 5754
rect 7967 5738 8001 5754
rect 7883 5362 7885 5408
rect 7849 5304 7885 5362
rect 7967 5346 8001 5362
rect 7376 5264 8471 5304
rect 7395 5263 8471 5264
rect 5851 5176 5918 5192
rect 5851 5142 5868 5176
rect 5902 5142 5918 5176
rect 5851 5126 5918 5142
rect 7273 5174 7340 5190
rect 7273 5140 7289 5174
rect 7323 5140 7340 5174
rect 7273 5124 7340 5140
rect 6158 5108 6192 5124
rect 5470 5058 5486 5092
rect 5520 5058 5536 5092
rect 5588 5059 5604 5093
rect 5638 5059 5654 5093
rect 6158 5058 6192 5074
rect 7104 5107 7138 5123
rect 7104 5057 7138 5073
rect 2820 5006 2854 5022
rect 2820 4814 2854 4830
rect 2938 5006 2972 5022
rect 2938 4814 2972 4830
rect 3240 5006 3274 5022
rect 3313 5006 3392 5022
rect 3313 4976 3358 5006
rect 3240 4563 3275 4630
rect 3358 4614 3392 4630
rect 3476 5006 3510 5022
rect 3476 4614 3510 4630
rect 3594 5006 3628 5022
rect 3712 5006 3746 5022
rect 4118 5006 4152 5022
rect 4118 4814 4152 4830
rect 4236 5006 4270 5022
rect 4236 4814 4270 4830
rect 4888 5008 4922 5024
rect 4888 4816 4922 4832
rect 5006 5008 5040 5024
rect 5006 4816 5040 4832
rect 5308 5008 5342 5024
rect 3594 4614 3628 4630
rect 3711 4563 3746 4630
rect 3240 4528 3746 4563
rect 5381 5008 5460 5024
rect 5381 4978 5426 5008
rect 5308 4565 5343 4632
rect 5426 4616 5460 4632
rect 5544 5008 5578 5024
rect 5544 4616 5578 4632
rect 5662 5008 5696 5024
rect 5780 5008 5814 5024
rect 6186 5008 6220 5024
rect 6186 4816 6220 4832
rect 6304 5008 6338 5024
rect 7450 5022 7484 5263
rect 8632 5315 8696 8008
rect 10068 7855 10102 7871
rect 10186 8059 10220 8063
rect 10260 8059 10294 8063
rect 10186 8047 10294 8059
rect 10220 7871 10260 8047
rect 10186 7859 10260 7871
rect 10186 7855 10220 7859
rect 10260 7655 10294 7671
rect 10378 8047 10412 8063
rect 10378 7655 10412 7671
rect 10496 8047 10530 8063
rect 10496 7655 10530 7671
rect 10614 8047 10648 8063
rect 10614 7655 10648 7671
rect 10732 8059 10766 8063
rect 10810 8059 10844 8063
rect 10732 8047 10844 8059
rect 10766 7871 10810 8047
rect 10766 7859 10844 7871
rect 10810 7855 10844 7859
rect 10928 8047 10962 8063
rect 10928 7855 10962 7871
rect 10732 7655 10766 7671
rect 10481 7536 10497 7570
rect 10531 7536 10547 7570
rect 10462 7418 10598 7422
rect 10462 7404 10500 7418
rect 10558 7404 10598 7418
rect 10462 7358 10478 7404
rect 10582 7358 10598 7404
rect 10462 7336 10598 7358
rect 12019 7246 12083 8511
rect 12235 8510 12292 8511
rect 13818 8559 13852 8575
rect 21497 8574 21770 8576
rect 15437 8572 15494 8574
rect 18581 8573 18638 8574
rect 13818 8509 13852 8525
rect 15193 8570 15495 8572
rect 15193 8510 15441 8570
rect 15490 8510 15495 8570
rect 15193 8508 15495 8510
rect 17020 8555 17054 8571
rect 12235 8406 12292 8410
rect 12235 8346 12239 8406
rect 12288 8346 12292 8406
rect 12235 8342 12292 8346
rect 13434 8405 13526 8418
rect 13434 8350 13450 8405
rect 13510 8350 13526 8405
rect 13434 8333 13526 8350
rect 13699 8169 13733 8185
rect 13699 8119 13733 8135
rect 13212 8047 13246 8063
rect 13212 7855 13246 7871
rect 13330 8059 13364 8063
rect 13404 8059 13438 8063
rect 13330 8047 13438 8059
rect 13364 7871 13404 8047
rect 13330 7859 13404 7871
rect 13330 7855 13364 7859
rect 13404 7655 13438 7671
rect 13522 8047 13556 8063
rect 13522 7655 13556 7671
rect 13640 8047 13674 8063
rect 13640 7655 13674 7671
rect 13758 8047 13792 8063
rect 13758 7655 13792 7671
rect 13876 8059 13910 8063
rect 13954 8059 13988 8063
rect 13876 8047 13988 8059
rect 13910 7871 13954 8047
rect 13910 7859 13988 7871
rect 13954 7855 13988 7859
rect 14072 8047 14106 8063
rect 14072 7855 14106 7871
rect 13876 7655 13910 7671
rect 13625 7536 13641 7570
rect 13675 7536 13691 7570
rect 13606 7418 13742 7422
rect 13606 7404 13644 7418
rect 13702 7404 13742 7418
rect 13606 7358 13622 7404
rect 13726 7358 13742 7404
rect 13606 7336 13742 7358
rect 15193 7273 15257 8508
rect 15437 8506 15494 8508
rect 17020 8505 17054 8521
rect 18355 8570 18638 8573
rect 18355 8510 18585 8570
rect 18634 8510 18638 8570
rect 18355 8509 18638 8510
rect 15437 8402 15494 8406
rect 15437 8342 15441 8402
rect 15490 8342 15494 8402
rect 15437 8338 15494 8342
rect 16636 8401 16728 8414
rect 16636 8346 16652 8401
rect 16712 8346 16728 8401
rect 16636 8329 16728 8346
rect 16901 8165 16935 8181
rect 16901 8115 16935 8131
rect 16414 8043 16448 8059
rect 16414 7851 16448 7867
rect 16532 8055 16566 8059
rect 16606 8055 16640 8059
rect 16532 8043 16640 8055
rect 16566 7867 16606 8043
rect 16532 7855 16606 7867
rect 16532 7851 16566 7855
rect 16606 7651 16640 7667
rect 16724 8043 16758 8059
rect 16724 7651 16758 7667
rect 16842 8043 16876 8059
rect 16842 7651 16876 7667
rect 16960 8043 16994 8059
rect 16960 7651 16994 7667
rect 17078 8055 17112 8059
rect 17156 8055 17190 8059
rect 17078 8043 17190 8055
rect 17112 7867 17156 8043
rect 17112 7855 17190 7867
rect 17156 7851 17190 7855
rect 17274 8043 17308 8059
rect 17274 7851 17308 7867
rect 17078 7651 17112 7667
rect 16827 7532 16843 7566
rect 16877 7532 16893 7566
rect 16808 7414 16944 7418
rect 16808 7400 16846 7414
rect 16904 7400 16944 7414
rect 16808 7354 16824 7400
rect 16928 7354 16944 7400
rect 16808 7332 16944 7354
rect 10713 7182 12083 7246
rect 12779 7209 15257 7273
rect 9651 6704 9853 6724
rect 9651 6660 9685 6704
rect 9807 6660 9853 6704
rect 9651 6650 9737 6660
rect 9775 6650 9853 6660
rect 9651 6632 9853 6650
rect 9738 6486 10008 6521
rect 9384 6433 9418 6449
rect 8900 6287 9170 6322
rect 8900 6233 8934 6287
rect 8900 6041 8934 6057
rect 9018 6233 9052 6249
rect 9018 6041 9052 6057
rect 9136 6233 9170 6287
rect 9136 6041 9170 6057
rect 9254 6233 9288 6249
rect 9254 6041 9288 6057
rect 9384 6041 9418 6057
rect 9502 6433 9536 6449
rect 9502 6041 9536 6057
rect 9620 6433 9654 6449
rect 9620 6041 9654 6057
rect 9738 6433 9772 6486
rect 9738 6041 9772 6057
rect 9856 6433 9890 6449
rect 9856 6041 9890 6057
rect 9974 6433 10008 6486
rect 9974 6041 10008 6057
rect 10092 6433 10126 6449
rect 10092 6041 10126 6057
rect 10221 6233 10255 6249
rect 10221 6041 10255 6057
rect 10339 6233 10373 6249
rect 10339 6041 10373 6057
rect 10457 6233 10491 6249
rect 10457 6041 10491 6057
rect 10575 6233 10609 6249
rect 10575 6041 10609 6057
rect 10301 5844 10307 5878
rect 10361 5844 10367 5878
rect 9327 5740 9361 5756
rect 9445 5740 9479 5756
rect 9327 5348 9361 5364
rect 9444 5364 9445 5411
rect 9563 5740 9597 5756
rect 9479 5364 9480 5411
rect 8573 5251 8696 5315
rect 9444 5306 9480 5364
rect 9681 5740 9715 5756
rect 9563 5348 9597 5364
rect 9679 5364 9681 5411
rect 9679 5306 9715 5364
rect 9799 5740 9833 5756
rect 9799 5348 9833 5364
rect 9917 5740 9951 5756
rect 10035 5740 10069 5756
rect 9951 5364 9953 5410
rect 9917 5306 9953 5364
rect 10035 5348 10069 5364
rect 9444 5266 10539 5306
rect 9463 5265 10539 5266
rect 7920 5174 7987 5190
rect 7920 5140 7937 5174
rect 7971 5140 7987 5174
rect 7920 5124 7987 5140
rect 9341 5176 9408 5192
rect 9341 5142 9357 5176
rect 9391 5142 9408 5176
rect 9341 5126 9408 5142
rect 8227 5106 8261 5122
rect 7539 5056 7555 5090
rect 7589 5056 7605 5090
rect 7657 5057 7673 5091
rect 7707 5057 7723 5091
rect 8227 5056 8261 5072
rect 9172 5109 9206 5125
rect 9172 5059 9206 5075
rect 9518 5024 9552 5265
rect 10713 5319 10778 7182
rect 11720 6704 11922 6724
rect 11720 6660 11754 6704
rect 11876 6660 11922 6704
rect 11720 6650 11806 6660
rect 11844 6650 11922 6660
rect 11720 6632 11922 6650
rect 11807 6486 12077 6521
rect 11453 6433 11487 6449
rect 10969 6287 11239 6322
rect 10969 6233 11003 6287
rect 10969 6041 11003 6057
rect 11087 6233 11121 6249
rect 11087 6041 11121 6057
rect 11205 6233 11239 6287
rect 11205 6041 11239 6057
rect 11323 6233 11357 6249
rect 11323 6041 11357 6057
rect 11453 6041 11487 6057
rect 11571 6433 11605 6449
rect 11571 6041 11605 6057
rect 11689 6433 11723 6449
rect 11689 6041 11723 6057
rect 11807 6433 11841 6486
rect 11807 6041 11841 6057
rect 11925 6433 11959 6449
rect 11925 6041 11959 6057
rect 12043 6433 12077 6486
rect 12043 6041 12077 6057
rect 12161 6433 12195 6449
rect 12161 6041 12195 6057
rect 12290 6233 12324 6249
rect 12290 6041 12324 6057
rect 12408 6233 12442 6249
rect 12408 6041 12442 6057
rect 12526 6233 12560 6249
rect 12526 6041 12560 6057
rect 12644 6233 12678 6249
rect 12644 6041 12678 6057
rect 12370 5844 12376 5878
rect 12430 5844 12436 5878
rect 11396 5740 11430 5756
rect 11514 5740 11548 5756
rect 11396 5348 11430 5364
rect 11513 5364 11514 5411
rect 11632 5740 11666 5756
rect 11548 5364 11549 5411
rect 10641 5255 10778 5319
rect 11513 5306 11549 5364
rect 11750 5740 11784 5756
rect 11632 5348 11666 5364
rect 11748 5364 11750 5411
rect 11748 5306 11784 5364
rect 11868 5740 11902 5756
rect 11868 5348 11902 5364
rect 11986 5740 12020 5756
rect 12104 5740 12138 5756
rect 12020 5364 12022 5410
rect 11986 5306 12022 5364
rect 12104 5348 12138 5364
rect 11513 5266 12608 5306
rect 11532 5265 12608 5266
rect 9988 5176 10055 5192
rect 9988 5142 10005 5176
rect 10039 5142 10055 5176
rect 9988 5126 10055 5142
rect 11410 5176 11477 5192
rect 11410 5142 11426 5176
rect 11460 5142 11477 5176
rect 11410 5126 11477 5142
rect 10295 5108 10329 5124
rect 9607 5058 9623 5092
rect 9657 5058 9673 5092
rect 9725 5059 9741 5093
rect 9775 5059 9791 5093
rect 10295 5058 10329 5074
rect 11241 5109 11275 5125
rect 11241 5059 11275 5075
rect 11587 5024 11621 5265
rect 12779 5306 12843 7209
rect 18355 7175 18419 8509
rect 18581 8506 18638 8509
rect 20164 8555 20198 8571
rect 20164 8505 20198 8521
rect 21497 8514 21717 8574
rect 21766 8514 21770 8574
rect 21497 8512 21770 8514
rect 18581 8402 18638 8406
rect 18581 8342 18585 8402
rect 18634 8342 18638 8402
rect 18581 8338 18638 8342
rect 19780 8401 19872 8414
rect 19780 8346 19796 8401
rect 19856 8346 19872 8401
rect 19780 8329 19872 8346
rect 20045 8165 20079 8181
rect 20045 8115 20079 8131
rect 19558 8043 19592 8059
rect 19558 7851 19592 7867
rect 19676 8055 19710 8059
rect 19750 8055 19784 8059
rect 19676 8043 19784 8055
rect 19710 7867 19750 8043
rect 19676 7855 19750 7867
rect 19676 7851 19710 7855
rect 19750 7651 19784 7667
rect 19868 8043 19902 8059
rect 19868 7651 19902 7667
rect 19986 8043 20020 8059
rect 19986 7651 20020 7667
rect 20104 8043 20138 8059
rect 20104 7651 20138 7667
rect 20222 8055 20256 8059
rect 20300 8055 20334 8059
rect 20222 8043 20334 8055
rect 20256 7867 20300 8043
rect 20256 7855 20334 7867
rect 20300 7851 20334 7855
rect 20418 8043 20452 8059
rect 20418 7851 20452 7867
rect 20222 7651 20256 7667
rect 19971 7532 19987 7566
rect 20021 7532 20037 7566
rect 19952 7414 20088 7418
rect 19952 7400 19990 7414
rect 20048 7400 20088 7414
rect 19952 7354 19968 7400
rect 20072 7354 20088 7400
rect 19952 7332 20088 7354
rect 14856 7111 18419 7175
rect 13788 6706 13990 6726
rect 13788 6662 13822 6706
rect 13944 6662 13990 6706
rect 13788 6652 13874 6662
rect 13912 6652 13990 6662
rect 13788 6634 13990 6652
rect 13875 6488 14145 6523
rect 13521 6435 13555 6451
rect 13037 6289 13307 6324
rect 13037 6235 13071 6289
rect 13037 6043 13071 6059
rect 13155 6235 13189 6251
rect 13155 6043 13189 6059
rect 13273 6235 13307 6289
rect 13273 6043 13307 6059
rect 13391 6235 13425 6251
rect 13391 6043 13425 6059
rect 13521 6043 13555 6059
rect 13639 6435 13673 6451
rect 13639 6043 13673 6059
rect 13757 6435 13791 6451
rect 13757 6043 13791 6059
rect 13875 6435 13909 6488
rect 13875 6043 13909 6059
rect 13993 6435 14027 6451
rect 13993 6043 14027 6059
rect 14111 6435 14145 6488
rect 14111 6043 14145 6059
rect 14229 6435 14263 6451
rect 14229 6043 14263 6059
rect 14358 6235 14392 6251
rect 14358 6043 14392 6059
rect 14476 6235 14510 6251
rect 14476 6043 14510 6059
rect 14594 6235 14628 6251
rect 14594 6043 14628 6059
rect 14712 6235 14746 6251
rect 14712 6043 14746 6059
rect 14438 5846 14444 5880
rect 14498 5846 14504 5880
rect 13464 5742 13498 5758
rect 13582 5742 13616 5758
rect 13464 5350 13498 5366
rect 13581 5366 13582 5413
rect 13700 5742 13734 5758
rect 13616 5366 13617 5413
rect 12710 5265 12843 5306
rect 13581 5308 13617 5366
rect 13818 5742 13852 5758
rect 13700 5350 13734 5366
rect 13816 5366 13818 5413
rect 13816 5308 13852 5366
rect 13936 5742 13970 5758
rect 13936 5350 13970 5366
rect 14054 5742 14088 5758
rect 14172 5742 14206 5758
rect 14088 5366 14090 5412
rect 14054 5308 14090 5366
rect 14172 5350 14206 5366
rect 13581 5268 14676 5308
rect 13600 5267 14676 5268
rect 12057 5176 12124 5192
rect 12057 5142 12074 5176
rect 12108 5142 12124 5176
rect 12057 5126 12124 5142
rect 13478 5178 13545 5194
rect 13478 5144 13494 5178
rect 13528 5144 13545 5178
rect 13478 5128 13545 5144
rect 12364 5108 12398 5124
rect 11676 5058 11692 5092
rect 11726 5058 11742 5092
rect 11794 5059 11810 5093
rect 11844 5059 11860 5093
rect 12364 5058 12398 5074
rect 13309 5111 13343 5127
rect 13309 5061 13343 5077
rect 13655 5026 13689 5267
rect 14856 5308 14920 7111
rect 21497 7052 21561 8512
rect 21713 8510 21770 8512
rect 23296 8559 23330 8575
rect 24857 8574 24914 8578
rect 23296 8509 23330 8525
rect 24637 8514 24861 8574
rect 24910 8514 24914 8574
rect 24637 8510 24914 8514
rect 26440 8559 26474 8575
rect 21713 8406 21770 8410
rect 21713 8346 21717 8406
rect 21766 8346 21770 8406
rect 21713 8342 21770 8346
rect 22912 8405 23004 8418
rect 22912 8350 22928 8405
rect 22988 8350 23004 8405
rect 22912 8333 23004 8350
rect 23177 8169 23211 8185
rect 23177 8119 23211 8135
rect 22690 8047 22724 8063
rect 22690 7855 22724 7871
rect 22808 8059 22842 8063
rect 22882 8059 22916 8063
rect 22808 8047 22916 8059
rect 22842 7871 22882 8047
rect 22808 7859 22882 7871
rect 22808 7855 22842 7859
rect 22882 7655 22916 7671
rect 23000 8047 23034 8063
rect 23000 7655 23034 7671
rect 23118 8047 23152 8063
rect 23118 7655 23152 7671
rect 23236 8047 23270 8063
rect 23236 7655 23270 7671
rect 23354 8059 23388 8063
rect 23432 8059 23466 8063
rect 23354 8047 23466 8059
rect 23388 7871 23432 8047
rect 23388 7859 23466 7871
rect 23432 7855 23466 7859
rect 23550 8047 23584 8063
rect 23550 7855 23584 7871
rect 23354 7655 23388 7671
rect 23103 7536 23119 7570
rect 23153 7536 23169 7570
rect 23084 7418 23220 7422
rect 23084 7404 23122 7418
rect 23180 7404 23220 7418
rect 23084 7358 23100 7404
rect 23204 7358 23220 7404
rect 23084 7336 23220 7358
rect 16934 6988 21561 7052
rect 15857 6704 16059 6724
rect 15857 6660 15891 6704
rect 16013 6660 16059 6704
rect 15857 6650 15943 6660
rect 15981 6650 16059 6660
rect 15857 6632 16059 6650
rect 15944 6486 16214 6521
rect 15590 6433 15624 6449
rect 15106 6287 15376 6322
rect 15106 6233 15140 6287
rect 15106 6041 15140 6057
rect 15224 6233 15258 6249
rect 15224 6041 15258 6057
rect 15342 6233 15376 6287
rect 15342 6041 15376 6057
rect 15460 6233 15494 6249
rect 15460 6041 15494 6057
rect 15590 6041 15624 6057
rect 15708 6433 15742 6449
rect 15708 6041 15742 6057
rect 15826 6433 15860 6449
rect 15826 6041 15860 6057
rect 15944 6433 15978 6486
rect 15944 6041 15978 6057
rect 16062 6433 16096 6449
rect 16062 6041 16096 6057
rect 16180 6433 16214 6486
rect 16180 6041 16214 6057
rect 16298 6433 16332 6449
rect 16298 6041 16332 6057
rect 16427 6233 16461 6249
rect 16427 6041 16461 6057
rect 16545 6233 16579 6249
rect 16545 6041 16579 6057
rect 16663 6233 16697 6249
rect 16663 6041 16697 6057
rect 16781 6233 16815 6249
rect 16781 6041 16815 6057
rect 16507 5844 16513 5878
rect 16567 5844 16573 5878
rect 15533 5740 15567 5756
rect 15651 5740 15685 5756
rect 15533 5348 15567 5364
rect 15650 5364 15651 5411
rect 15769 5740 15803 5756
rect 15685 5364 15686 5411
rect 14778 5267 14920 5308
rect 15650 5306 15686 5364
rect 15887 5740 15921 5756
rect 15769 5348 15803 5364
rect 15885 5364 15887 5411
rect 15885 5306 15921 5364
rect 16005 5740 16039 5756
rect 16005 5348 16039 5364
rect 16123 5740 16157 5756
rect 16241 5740 16275 5756
rect 16157 5364 16159 5410
rect 16123 5306 16159 5364
rect 16241 5348 16275 5364
rect 15650 5266 16745 5306
rect 15669 5265 16745 5266
rect 14125 5178 14192 5194
rect 14125 5144 14142 5178
rect 14176 5144 14192 5178
rect 14125 5128 14192 5144
rect 15547 5176 15614 5192
rect 15547 5142 15563 5176
rect 15597 5142 15614 5176
rect 15547 5126 15614 5142
rect 14432 5110 14466 5126
rect 13744 5060 13760 5094
rect 13794 5060 13810 5094
rect 13862 5061 13878 5095
rect 13912 5061 13928 5095
rect 14432 5060 14466 5076
rect 15378 5109 15412 5125
rect 15378 5059 15412 5075
rect 6304 4816 6338 4832
rect 6957 5006 6991 5022
rect 6957 4814 6991 4830
rect 7075 5006 7109 5022
rect 7075 4814 7109 4830
rect 7377 5006 7411 5022
rect 5662 4616 5696 4632
rect 5779 4565 5814 4632
rect 5308 4530 5814 4565
rect 7450 5006 7529 5022
rect 7450 4976 7495 5006
rect 7377 4563 7412 4630
rect 7495 4614 7529 4630
rect 7613 5006 7647 5022
rect 7613 4614 7647 4630
rect 7731 5006 7765 5022
rect 7849 5006 7883 5022
rect 8255 5006 8289 5022
rect 8255 4814 8289 4830
rect 8373 5006 8407 5022
rect 8373 4814 8407 4830
rect 9025 5008 9059 5024
rect 9025 4816 9059 4832
rect 9143 5008 9177 5024
rect 9143 4816 9177 4832
rect 9445 5008 9479 5024
rect 7731 4614 7765 4630
rect 7848 4563 7883 4630
rect 7377 4528 7883 4563
rect 9518 5008 9597 5024
rect 9518 4978 9563 5008
rect 9445 4565 9480 4632
rect 9563 4616 9597 4632
rect 9681 5008 9715 5024
rect 9681 4616 9715 4632
rect 9799 5008 9833 5024
rect 9917 5008 9951 5024
rect 10323 5008 10357 5024
rect 10323 4816 10357 4832
rect 10441 5008 10475 5024
rect 10441 4816 10475 4832
rect 11094 5008 11128 5024
rect 11094 4816 11128 4832
rect 11212 5008 11246 5024
rect 11212 4816 11246 4832
rect 11514 5008 11548 5024
rect 9799 4616 9833 4632
rect 9916 4565 9951 4632
rect 9445 4530 9951 4565
rect 11587 5008 11666 5024
rect 11587 4978 11632 5008
rect 11514 4565 11549 4632
rect 11632 4616 11666 4632
rect 11750 5008 11784 5024
rect 11750 4616 11784 4632
rect 11868 5008 11902 5024
rect 11986 5008 12020 5024
rect 12392 5008 12426 5024
rect 12392 4816 12426 4832
rect 12510 5008 12544 5024
rect 12510 4816 12544 4832
rect 13162 5010 13196 5026
rect 13162 4818 13196 4834
rect 13280 5010 13314 5026
rect 13280 4818 13314 4834
rect 13582 5010 13616 5026
rect 11868 4616 11902 4632
rect 11985 4565 12020 4632
rect 11514 4530 12020 4565
rect 13655 5010 13734 5026
rect 13655 4980 13700 5010
rect 13582 4567 13617 4634
rect 13700 4618 13734 4634
rect 13818 5010 13852 5026
rect 13818 4618 13852 4634
rect 13936 5010 13970 5026
rect 14054 5010 14088 5026
rect 14460 5010 14494 5026
rect 14460 4818 14494 4834
rect 14578 5010 14612 5026
rect 15724 5024 15758 5265
rect 16934 5306 16998 6988
rect 24637 6954 24701 8510
rect 26440 8509 26474 8525
rect 24857 8406 24914 8410
rect 24857 8346 24861 8406
rect 24910 8346 24914 8406
rect 24857 8342 24914 8346
rect 26056 8405 26148 8418
rect 26056 8350 26072 8405
rect 26132 8350 26148 8405
rect 26056 8333 26148 8350
rect 26321 8169 26355 8185
rect 26321 8119 26355 8135
rect 25834 8047 25868 8063
rect 25834 7855 25868 7871
rect 25952 8059 25986 8063
rect 26026 8059 26060 8063
rect 25952 8047 26060 8059
rect 25986 7871 26026 8047
rect 25952 7859 26026 7871
rect 25952 7855 25986 7859
rect 26026 7655 26060 7671
rect 26144 8047 26178 8063
rect 26144 7655 26178 7671
rect 26262 8047 26296 8063
rect 26262 7655 26296 7671
rect 26380 8047 26414 8063
rect 26380 7655 26414 7671
rect 26498 8059 26532 8063
rect 26576 8059 26610 8063
rect 26498 8047 26610 8059
rect 26532 7871 26576 8047
rect 26532 7859 26610 7871
rect 26576 7855 26610 7859
rect 26694 8047 26728 8063
rect 26694 7855 26728 7871
rect 26498 7655 26532 7671
rect 26247 7536 26263 7570
rect 26297 7536 26313 7570
rect 26228 7418 26364 7422
rect 26228 7404 26266 7418
rect 26324 7404 26364 7418
rect 26228 7358 26244 7404
rect 26348 7358 26364 7404
rect 26228 7336 26364 7358
rect 18985 6890 24701 6954
rect 17925 6706 18127 6726
rect 17925 6662 17959 6706
rect 18081 6662 18127 6706
rect 17925 6652 18011 6662
rect 18049 6652 18127 6662
rect 17925 6634 18127 6652
rect 18012 6488 18282 6523
rect 17658 6435 17692 6451
rect 17174 6289 17444 6324
rect 17174 6235 17208 6289
rect 17174 6043 17208 6059
rect 17292 6235 17326 6251
rect 17292 6043 17326 6059
rect 17410 6235 17444 6289
rect 17410 6043 17444 6059
rect 17528 6235 17562 6251
rect 17528 6043 17562 6059
rect 17658 6043 17692 6059
rect 17776 6435 17810 6451
rect 17776 6043 17810 6059
rect 17894 6435 17928 6451
rect 17894 6043 17928 6059
rect 18012 6435 18046 6488
rect 18012 6043 18046 6059
rect 18130 6435 18164 6451
rect 18130 6043 18164 6059
rect 18248 6435 18282 6488
rect 18248 6043 18282 6059
rect 18366 6435 18400 6451
rect 18366 6043 18400 6059
rect 18495 6235 18529 6251
rect 18495 6043 18529 6059
rect 18613 6235 18647 6251
rect 18613 6043 18647 6059
rect 18731 6235 18765 6251
rect 18731 6043 18765 6059
rect 18849 6235 18883 6251
rect 18849 6043 18883 6059
rect 18575 5846 18581 5880
rect 18635 5846 18641 5880
rect 17601 5742 17635 5758
rect 17181 5631 17247 5640
rect 17719 5742 17753 5758
rect 17601 5350 17635 5366
rect 17718 5366 17719 5413
rect 17837 5742 17871 5758
rect 17753 5366 17754 5413
rect 16847 5265 16998 5306
rect 17718 5308 17754 5366
rect 17955 5742 17989 5758
rect 17837 5350 17871 5366
rect 17953 5366 17955 5413
rect 17953 5308 17989 5366
rect 18073 5742 18107 5758
rect 18073 5350 18107 5366
rect 18191 5742 18225 5758
rect 18309 5742 18343 5758
rect 18225 5366 18227 5412
rect 18191 5308 18227 5366
rect 18309 5350 18343 5366
rect 17718 5268 18813 5308
rect 17737 5267 18813 5268
rect 16194 5176 16261 5192
rect 16194 5142 16211 5176
rect 16245 5142 16261 5176
rect 16194 5126 16261 5142
rect 17615 5178 17682 5194
rect 17615 5144 17631 5178
rect 17665 5144 17682 5178
rect 17615 5128 17682 5144
rect 16501 5108 16535 5124
rect 15813 5058 15829 5092
rect 15863 5058 15879 5092
rect 15931 5059 15947 5093
rect 15981 5059 15997 5093
rect 16501 5058 16535 5074
rect 17446 5111 17480 5127
rect 17446 5061 17480 5077
rect 17792 5026 17826 5267
rect 18985 5308 19049 6890
rect 19517 6753 19731 6757
rect 19517 6691 19551 6753
rect 19691 6691 19731 6753
rect 19517 6673 19731 6691
rect 20255 6751 20469 6755
rect 20255 6689 20289 6751
rect 20429 6689 20469 6751
rect 20255 6671 20469 6689
rect 20993 6751 21207 6755
rect 20993 6689 21027 6751
rect 21167 6689 21207 6751
rect 20993 6671 21207 6689
rect 21735 6751 21949 6755
rect 21735 6689 21769 6751
rect 21909 6689 21949 6751
rect 21735 6671 21949 6689
rect 22475 6751 22689 6755
rect 22475 6689 22509 6751
rect 22649 6689 22689 6751
rect 22475 6671 22689 6689
rect 23213 6751 23427 6755
rect 23213 6689 23247 6751
rect 23387 6689 23427 6751
rect 23213 6671 23427 6689
rect 23951 6751 24165 6755
rect 23951 6689 23985 6751
rect 24125 6689 24165 6751
rect 23951 6671 24165 6689
rect 24689 6751 24903 6755
rect 24689 6689 24723 6751
rect 24863 6689 24903 6751
rect 24689 6671 24903 6689
rect 19545 6603 19815 6637
rect 19427 6547 19461 6563
rect 19427 6355 19461 6371
rect 19545 6547 19579 6603
rect 19545 6355 19579 6371
rect 19663 6547 19697 6563
rect 19663 6355 19697 6371
rect 19781 6547 19815 6603
rect 20283 6601 20553 6635
rect 19781 6355 19815 6371
rect 20165 6551 20199 6567
rect 20165 6359 20199 6375
rect 20283 6551 20317 6601
rect 20283 6359 20317 6375
rect 20401 6551 20435 6567
rect 20401 6359 20435 6375
rect 20519 6551 20553 6601
rect 21021 6601 21291 6635
rect 20519 6359 20553 6375
rect 20903 6547 20937 6563
rect 20903 6355 20937 6371
rect 21021 6547 21055 6601
rect 21021 6355 21055 6371
rect 21139 6547 21173 6563
rect 21139 6355 21173 6371
rect 21257 6547 21291 6601
rect 21763 6601 22033 6635
rect 21257 6355 21291 6371
rect 21645 6545 21679 6561
rect 21645 6353 21679 6369
rect 21763 6545 21797 6601
rect 21763 6353 21797 6369
rect 21881 6545 21915 6561
rect 21881 6353 21915 6369
rect 21999 6545 22033 6601
rect 22503 6601 22773 6635
rect 21999 6353 22033 6369
rect 22385 6545 22419 6561
rect 22385 6353 22419 6369
rect 22503 6545 22537 6601
rect 22503 6353 22537 6369
rect 22621 6545 22655 6561
rect 22621 6353 22655 6369
rect 22739 6545 22773 6601
rect 23241 6601 23511 6635
rect 22739 6353 22773 6369
rect 23123 6545 23157 6561
rect 23123 6353 23157 6369
rect 23241 6545 23275 6601
rect 23241 6353 23275 6369
rect 23359 6545 23393 6561
rect 23359 6353 23393 6369
rect 23477 6545 23511 6601
rect 23979 6601 24249 6635
rect 23477 6353 23511 6369
rect 23861 6545 23895 6561
rect 23861 6353 23895 6369
rect 23979 6545 24013 6601
rect 23979 6353 24013 6369
rect 24097 6545 24131 6561
rect 24097 6353 24131 6369
rect 24215 6545 24249 6601
rect 24717 6601 24987 6635
rect 24215 6353 24249 6369
rect 24599 6545 24633 6561
rect 24599 6353 24633 6369
rect 24717 6545 24751 6601
rect 24717 6353 24751 6369
rect 24835 6545 24869 6561
rect 24835 6353 24869 6369
rect 24953 6545 24987 6601
rect 24953 6353 24987 6369
rect 18915 5267 19049 5308
rect 19357 6231 19603 6265
rect 19637 6231 19653 6265
rect 18262 5178 18329 5194
rect 18262 5144 18279 5178
rect 18313 5144 18329 5178
rect 18262 5128 18329 5144
rect 18569 5110 18603 5126
rect 17881 5060 17897 5094
rect 17931 5060 17947 5094
rect 17999 5061 18015 5095
rect 18049 5061 18065 5095
rect 18569 5060 18603 5076
rect 14578 4818 14612 4834
rect 15231 5008 15265 5024
rect 15231 4816 15265 4832
rect 15349 5008 15383 5024
rect 15349 4816 15383 4832
rect 15651 5008 15685 5024
rect 13936 4618 13970 4634
rect 14053 4567 14088 4634
rect 13582 4532 14088 4567
rect 15724 5008 15803 5024
rect 15724 4978 15769 5008
rect 15651 4565 15686 4632
rect 15769 4616 15803 4632
rect 15887 5008 15921 5024
rect 15887 4616 15921 4632
rect 16005 5008 16039 5024
rect 16123 5008 16157 5024
rect 16529 5008 16563 5024
rect 16529 4816 16563 4832
rect 16647 5008 16681 5024
rect 16647 4816 16681 4832
rect 17299 5010 17333 5026
rect 17299 4818 17333 4834
rect 17417 5010 17451 5026
rect 17417 4818 17451 4834
rect 17719 5010 17753 5026
rect 16005 4616 16039 4632
rect 16122 4565 16157 4632
rect 15651 4530 16157 4565
rect 17792 5010 17871 5026
rect 17792 4980 17837 5010
rect 17719 4567 17754 4634
rect 17837 4618 17871 4634
rect 17955 5010 17989 5026
rect 17955 4618 17989 4634
rect 18073 5010 18107 5026
rect 18191 5010 18225 5026
rect 18597 5010 18631 5026
rect 18597 4818 18631 4834
rect 18715 5010 18749 5026
rect 18715 4818 18749 4834
rect 18073 4618 18107 4634
rect 18190 4567 18225 4634
rect 17719 4532 18225 4567
rect 3414 4442 3470 4458
rect 3520 4442 3578 4458
rect 3414 4386 3430 4442
rect 3562 4386 3578 4442
rect 3414 4370 3578 4386
rect 5482 4444 5538 4460
rect 5588 4444 5646 4460
rect 5482 4388 5498 4444
rect 5630 4388 5646 4444
rect 5482 4372 5646 4388
rect 7551 4442 7607 4458
rect 7657 4442 7715 4458
rect 7551 4386 7567 4442
rect 7699 4386 7715 4442
rect 7551 4370 7715 4386
rect 9619 4444 9675 4460
rect 9725 4444 9783 4460
rect 9619 4388 9635 4444
rect 9767 4388 9783 4444
rect 9619 4372 9783 4388
rect 11688 4444 11744 4460
rect 11794 4444 11852 4460
rect 11688 4388 11704 4444
rect 11836 4388 11852 4444
rect 11688 4372 11852 4388
rect 13756 4446 13812 4462
rect 13862 4446 13920 4462
rect 13756 4390 13772 4446
rect 13904 4390 13920 4446
rect 13756 4374 13920 4390
rect 15825 4444 15881 4460
rect 15931 4444 15989 4460
rect 15825 4388 15841 4444
rect 15973 4388 15989 4444
rect 15825 4372 15989 4388
rect 17893 4446 17949 4462
rect 17999 4446 18057 4462
rect 17893 4390 17909 4446
rect 18041 4390 18057 4446
rect 17893 4374 18057 4390
rect 19357 4154 19421 6231
rect 19957 6229 20341 6263
rect 20375 6229 20391 6263
rect 20677 6229 21079 6263
rect 21113 6229 21129 6263
rect 21406 6229 21821 6263
rect 21855 6229 21871 6263
rect 22229 6229 22561 6263
rect 22595 6229 22611 6263
rect 22927 6229 23299 6263
rect 23333 6229 23349 6263
rect 19545 6161 19579 6177
rect 19545 5969 19579 5985
rect 19663 6161 19697 6177
rect 19663 5969 19697 5985
rect 19465 5873 19649 5893
rect 19465 5803 19485 5873
rect 19629 5803 19649 5873
rect 19465 5797 19649 5803
rect 2665 4090 19421 4154
rect 19957 4056 20021 6229
rect 20283 6163 20317 6179
rect 20283 5971 20317 5987
rect 20401 6163 20435 6179
rect 20401 5971 20435 5987
rect 20203 5871 20387 5891
rect 20203 5801 20223 5871
rect 20367 5801 20387 5871
rect 20203 5795 20387 5801
rect 4715 4055 20021 4056
rect 4766 4004 20021 4055
rect 4715 3992 20021 4004
rect 20677 3947 20741 6229
rect 21021 6159 21055 6175
rect 21021 5967 21055 5983
rect 21139 6159 21173 6175
rect 21139 5967 21173 5983
rect 20941 5871 21125 5891
rect 20941 5801 20961 5871
rect 21105 5801 21125 5871
rect 20941 5795 21125 5801
rect 6797 3896 20741 3947
rect 6750 3883 20741 3896
rect 6750 3882 6813 3883
rect 21406 3849 21470 6229
rect 21763 6159 21797 6175
rect 21763 5967 21797 5983
rect 21881 6159 21915 6175
rect 21881 5967 21915 5983
rect 21683 5871 21867 5891
rect 21683 5801 21703 5871
rect 21847 5801 21867 5871
rect 21683 5795 21867 5801
rect 8788 3847 21470 3849
rect 8788 3793 8797 3847
rect 8844 3793 21470 3847
rect 8788 3785 21470 3793
rect 22229 3741 22293 6229
rect 22927 6228 23306 6229
rect 22503 6159 22537 6175
rect 22503 5967 22537 5983
rect 22621 6159 22655 6175
rect 22621 5967 22655 5983
rect 22423 5871 22607 5891
rect 22423 5801 22443 5871
rect 22587 5801 22607 5871
rect 22423 5795 22607 5801
rect 10887 3737 22293 3741
rect 10937 3686 22293 3737
rect 10887 3677 22293 3686
rect 22927 3643 22991 6228
rect 23717 6223 23854 6269
rect 24021 6229 24037 6263
rect 24071 6229 24087 6263
rect 24475 6223 24591 6269
rect 24759 6229 24775 6263
rect 24809 6229 24825 6263
rect 23241 6159 23275 6175
rect 23241 5967 23275 5983
rect 23359 6159 23393 6175
rect 23359 5967 23393 5983
rect 23161 5871 23345 5891
rect 23161 5801 23181 5871
rect 23325 5801 23345 5871
rect 23161 5795 23345 5801
rect 12958 3642 22991 3643
rect 13009 3589 22991 3642
rect 12958 3579 22991 3589
rect 23718 3502 23782 6223
rect 23979 6163 24013 6179
rect 23979 5971 24013 5987
rect 24097 6163 24131 6179
rect 24097 5971 24131 5987
rect 23899 5871 24083 5891
rect 23899 5801 23919 5871
rect 24063 5801 24083 5871
rect 23899 5795 24083 5801
rect 24475 4004 24539 6223
rect 24717 6163 24751 6179
rect 24717 5971 24751 5987
rect 24835 6163 24869 6179
rect 24835 5971 24869 5987
rect 24637 5871 24821 5891
rect 24637 5801 24657 5871
rect 24801 5801 24821 5871
rect 24637 5795 24821 5801
rect 15051 3498 23782 3502
rect 15051 3447 15061 3498
rect 15105 3447 23782 3498
rect 15051 3438 23782 3447
rect 24474 3404 24539 4004
rect 17129 3403 24539 3404
rect 17182 3349 24539 3403
rect 17129 3340 24539 3349
rect 17129 3339 17210 3340
rect 1430 2398 1658 2416
rect 1430 2322 1446 2398
rect 1642 2322 1658 2398
rect 1430 2306 1658 2322
rect 4574 2398 4802 2416
rect 4574 2322 4590 2398
rect 4786 2322 4802 2398
rect 4574 2306 4802 2322
rect 7706 2402 7934 2420
rect 7706 2326 7722 2402
rect 7918 2326 7934 2402
rect 7706 2310 7934 2326
rect 10850 2402 11078 2420
rect 10850 2326 10866 2402
rect 11062 2326 11078 2402
rect 10850 2310 11078 2326
rect 14052 2398 14280 2416
rect 14052 2322 14068 2398
rect 14264 2322 14280 2398
rect 14052 2306 14280 2322
rect 17196 2398 17424 2416
rect 17196 2322 17212 2398
rect 17408 2322 17424 2398
rect 17196 2306 17424 2322
rect 20328 2402 20556 2420
rect 20328 2326 20344 2402
rect 20540 2326 20556 2402
rect 20328 2310 20556 2326
rect 23472 2402 23700 2420
rect 23472 2326 23488 2402
rect 23684 2326 23700 2402
rect 23472 2310 23700 2326
rect 701 2181 971 2220
rect 701 2128 735 2181
rect 260 1979 530 2018
rect 260 1928 294 1979
rect 260 1736 294 1752
rect 378 1928 412 1944
rect 378 1701 412 1752
rect 496 1928 530 1979
rect 496 1736 530 1752
rect 614 1928 648 1944
rect 614 1701 648 1752
rect 701 1736 735 1752
rect 819 2128 853 2144
rect 378 1662 648 1701
rect 819 1701 853 1752
rect 937 2128 971 2181
rect 1168 2180 1438 2219
rect 937 1736 971 1752
rect 1055 2128 1089 2144
rect 1055 1701 1089 1752
rect 1168 2128 1202 2180
rect 1168 1736 1202 1752
rect 1286 2128 1320 2144
rect 1286 1701 1320 1752
rect 1404 2128 1438 2180
rect 1640 2180 1910 2219
rect 1404 1736 1438 1752
rect 1522 2128 1556 2144
rect 1522 1701 1556 1752
rect 1640 2128 1674 2180
rect 1640 1736 1674 1752
rect 1758 2128 1792 2144
rect 1758 1701 1792 1752
rect 1876 2128 1910 2180
rect 2113 2180 2383 2219
rect 1876 1736 1910 1752
rect 1995 2128 2029 2144
rect 1995 1701 2029 1752
rect 2113 2128 2147 2180
rect 2113 1736 2147 1752
rect 2231 2128 2265 2144
rect 2231 1701 2265 1752
rect 2349 2128 2383 2180
rect 3845 2181 4115 2220
rect 3845 2128 3879 2181
rect 2586 1978 2856 2015
rect 2349 1736 2383 1752
rect 2468 1928 2502 1944
rect 819 1662 2265 1701
rect 2468 1698 2502 1752
rect 2586 1928 2620 1978
rect 2586 1736 2620 1752
rect 2704 1928 2738 1944
rect 2704 1698 2738 1752
rect 2822 1928 2856 1978
rect 2822 1736 2856 1752
rect 3404 1979 3674 2018
rect 3404 1928 3438 1979
rect 3404 1736 3438 1752
rect 3522 1928 3556 1944
rect 2468 1659 2738 1698
rect 3522 1701 3556 1752
rect 3640 1928 3674 1979
rect 3640 1736 3674 1752
rect 3758 1928 3792 1944
rect 3758 1701 3792 1752
rect 3845 1736 3879 1752
rect 3963 2128 3997 2144
rect 3522 1662 3792 1701
rect 3963 1701 3997 1752
rect 4081 2128 4115 2181
rect 4312 2180 4582 2219
rect 4081 1736 4115 1752
rect 4199 2128 4233 2144
rect 4199 1701 4233 1752
rect 4312 2128 4346 2180
rect 4312 1736 4346 1752
rect 4430 2128 4464 2144
rect 4430 1701 4464 1752
rect 4548 2128 4582 2180
rect 4784 2180 5054 2219
rect 4548 1736 4582 1752
rect 4666 2128 4700 2144
rect 4666 1701 4700 1752
rect 4784 2128 4818 2180
rect 4784 1736 4818 1752
rect 4902 2128 4936 2144
rect 4902 1701 4936 1752
rect 5020 2128 5054 2180
rect 5257 2180 5527 2219
rect 5020 1736 5054 1752
rect 5139 2128 5173 2144
rect 5139 1701 5173 1752
rect 5257 2128 5291 2180
rect 5257 1736 5291 1752
rect 5375 2128 5409 2144
rect 5375 1701 5409 1752
rect 5493 2128 5527 2180
rect 6977 2185 7247 2224
rect 6977 2132 7011 2185
rect 5730 1978 6000 2015
rect 5493 1736 5527 1752
rect 5612 1928 5646 1944
rect 3963 1662 5409 1701
rect 5612 1698 5646 1752
rect 5730 1928 5764 1978
rect 5730 1736 5764 1752
rect 5848 1928 5882 1944
rect 5848 1698 5882 1752
rect 5966 1928 6000 1978
rect 5966 1736 6000 1752
rect 6536 1983 6806 2022
rect 6536 1932 6570 1983
rect 6536 1740 6570 1756
rect 6654 1932 6688 1948
rect 5612 1659 5882 1698
rect 6654 1705 6688 1756
rect 6772 1932 6806 1983
rect 6772 1740 6806 1756
rect 6890 1932 6924 1948
rect 6890 1705 6924 1756
rect 6977 1740 7011 1756
rect 7095 2132 7129 2148
rect 6654 1666 6924 1705
rect 7095 1705 7129 1756
rect 7213 2132 7247 2185
rect 7444 2184 7714 2223
rect 7213 1740 7247 1756
rect 7331 2132 7365 2148
rect 7331 1705 7365 1756
rect 7444 2132 7478 2184
rect 7444 1740 7478 1756
rect 7562 2132 7596 2148
rect 7562 1705 7596 1756
rect 7680 2132 7714 2184
rect 7916 2184 8186 2223
rect 7680 1740 7714 1756
rect 7798 2132 7832 2148
rect 7798 1705 7832 1756
rect 7916 2132 7950 2184
rect 7916 1740 7950 1756
rect 8034 2132 8068 2148
rect 8034 1705 8068 1756
rect 8152 2132 8186 2184
rect 8389 2184 8659 2223
rect 8152 1740 8186 1756
rect 8271 2132 8305 2148
rect 8271 1705 8305 1756
rect 8389 2132 8423 2184
rect 8389 1740 8423 1756
rect 8507 2132 8541 2148
rect 8507 1705 8541 1756
rect 8625 2132 8659 2184
rect 10121 2185 10391 2224
rect 10121 2132 10155 2185
rect 8862 1982 9132 2019
rect 8625 1740 8659 1756
rect 8744 1932 8778 1948
rect 7095 1666 8541 1705
rect 8744 1702 8778 1756
rect 8862 1932 8896 1982
rect 8862 1740 8896 1756
rect 8980 1932 9014 1948
rect 8980 1702 9014 1756
rect 9098 1932 9132 1982
rect 9098 1740 9132 1756
rect 9680 1983 9950 2022
rect 9680 1932 9714 1983
rect 9680 1740 9714 1756
rect 9798 1932 9832 1948
rect 8744 1663 9014 1702
rect 9798 1705 9832 1756
rect 9916 1932 9950 1983
rect 9916 1740 9950 1756
rect 10034 1932 10068 1948
rect 10034 1705 10068 1756
rect 10121 1740 10155 1756
rect 10239 2132 10273 2148
rect 9798 1666 10068 1705
rect 10239 1705 10273 1756
rect 10357 2132 10391 2185
rect 10588 2184 10858 2223
rect 10357 1740 10391 1756
rect 10475 2132 10509 2148
rect 10475 1705 10509 1756
rect 10588 2132 10622 2184
rect 10588 1740 10622 1756
rect 10706 2132 10740 2148
rect 10706 1705 10740 1756
rect 10824 2132 10858 2184
rect 11060 2184 11330 2223
rect 10824 1740 10858 1756
rect 10942 2132 10976 2148
rect 10942 1705 10976 1756
rect 11060 2132 11094 2184
rect 11060 1740 11094 1756
rect 11178 2132 11212 2148
rect 11178 1705 11212 1756
rect 11296 2132 11330 2184
rect 11533 2184 11803 2223
rect 11296 1740 11330 1756
rect 11415 2132 11449 2148
rect 11415 1705 11449 1756
rect 11533 2132 11567 2184
rect 11533 1740 11567 1756
rect 11651 2132 11685 2148
rect 11651 1705 11685 1756
rect 11769 2132 11803 2184
rect 13323 2181 13593 2220
rect 13323 2128 13357 2181
rect 12006 1982 12276 2019
rect 11769 1740 11803 1756
rect 11888 1932 11922 1948
rect 10239 1666 11685 1705
rect 11888 1702 11922 1756
rect 12006 1932 12040 1982
rect 12006 1740 12040 1756
rect 12124 1932 12158 1948
rect 12124 1702 12158 1756
rect 12242 1932 12276 1982
rect 12242 1740 12276 1756
rect 12882 1979 13152 2018
rect 12882 1928 12916 1979
rect 12882 1736 12916 1752
rect 13000 1928 13034 1944
rect 11888 1663 12158 1702
rect 13000 1701 13034 1752
rect 13118 1928 13152 1979
rect 13118 1736 13152 1752
rect 13236 1928 13270 1944
rect 13236 1701 13270 1752
rect 13323 1736 13357 1752
rect 13441 2128 13475 2144
rect 13000 1662 13270 1701
rect 13441 1701 13475 1752
rect 13559 2128 13593 2181
rect 13790 2180 14060 2219
rect 13559 1736 13593 1752
rect 13677 2128 13711 2144
rect 13677 1701 13711 1752
rect 13790 2128 13824 2180
rect 13790 1736 13824 1752
rect 13908 2128 13942 2144
rect 13908 1701 13942 1752
rect 14026 2128 14060 2180
rect 14262 2180 14532 2219
rect 14026 1736 14060 1752
rect 14144 2128 14178 2144
rect 14144 1701 14178 1752
rect 14262 2128 14296 2180
rect 14262 1736 14296 1752
rect 14380 2128 14414 2144
rect 14380 1701 14414 1752
rect 14498 2128 14532 2180
rect 14735 2180 15005 2219
rect 14498 1736 14532 1752
rect 14617 2128 14651 2144
rect 14617 1701 14651 1752
rect 14735 2128 14769 2180
rect 14735 1736 14769 1752
rect 14853 2128 14887 2144
rect 14853 1701 14887 1752
rect 14971 2128 15005 2180
rect 16467 2181 16737 2220
rect 16467 2128 16501 2181
rect 15208 1978 15478 2015
rect 14971 1736 15005 1752
rect 15090 1928 15124 1944
rect 13441 1662 14887 1701
rect 15090 1698 15124 1752
rect 15208 1928 15242 1978
rect 15208 1736 15242 1752
rect 15326 1928 15360 1944
rect 15326 1698 15360 1752
rect 15444 1928 15478 1978
rect 15444 1736 15478 1752
rect 16026 1979 16296 2018
rect 16026 1928 16060 1979
rect 16026 1736 16060 1752
rect 16144 1928 16178 1944
rect 15090 1659 15360 1698
rect 16144 1701 16178 1752
rect 16262 1928 16296 1979
rect 16262 1736 16296 1752
rect 16380 1928 16414 1944
rect 16380 1701 16414 1752
rect 16467 1736 16501 1752
rect 16585 2128 16619 2144
rect 16144 1662 16414 1701
rect 16585 1701 16619 1752
rect 16703 2128 16737 2181
rect 16934 2180 17204 2219
rect 16703 1736 16737 1752
rect 16821 2128 16855 2144
rect 16821 1701 16855 1752
rect 16934 2128 16968 2180
rect 16934 1736 16968 1752
rect 17052 2128 17086 2144
rect 17052 1701 17086 1752
rect 17170 2128 17204 2180
rect 17406 2180 17676 2219
rect 17170 1736 17204 1752
rect 17288 2128 17322 2144
rect 17288 1701 17322 1752
rect 17406 2128 17440 2180
rect 17406 1736 17440 1752
rect 17524 2128 17558 2144
rect 17524 1701 17558 1752
rect 17642 2128 17676 2180
rect 17879 2180 18149 2219
rect 17642 1736 17676 1752
rect 17761 2128 17795 2144
rect 17761 1701 17795 1752
rect 17879 2128 17913 2180
rect 17879 1736 17913 1752
rect 17997 2128 18031 2144
rect 17997 1701 18031 1752
rect 18115 2128 18149 2180
rect 19599 2185 19869 2224
rect 19599 2132 19633 2185
rect 18352 1978 18622 2015
rect 18115 1736 18149 1752
rect 18234 1928 18268 1944
rect 16585 1662 18031 1701
rect 18234 1698 18268 1752
rect 18352 1928 18386 1978
rect 18352 1736 18386 1752
rect 18470 1928 18504 1944
rect 18470 1698 18504 1752
rect 18588 1928 18622 1978
rect 18588 1736 18622 1752
rect 19158 1983 19428 2022
rect 19158 1932 19192 1983
rect 19158 1740 19192 1756
rect 19276 1932 19310 1948
rect 18234 1659 18504 1698
rect 19276 1705 19310 1756
rect 19394 1932 19428 1983
rect 19394 1740 19428 1756
rect 19512 1932 19546 1948
rect 19512 1705 19546 1756
rect 19599 1740 19633 1756
rect 19717 2132 19751 2148
rect 19276 1666 19546 1705
rect 19717 1705 19751 1756
rect 19835 2132 19869 2185
rect 20066 2184 20336 2223
rect 19835 1740 19869 1756
rect 19953 2132 19987 2148
rect 19953 1705 19987 1756
rect 20066 2132 20100 2184
rect 20066 1740 20100 1756
rect 20184 2132 20218 2148
rect 20184 1705 20218 1756
rect 20302 2132 20336 2184
rect 20538 2184 20808 2223
rect 20302 1740 20336 1756
rect 20420 2132 20454 2148
rect 20420 1705 20454 1756
rect 20538 2132 20572 2184
rect 20538 1740 20572 1756
rect 20656 2132 20690 2148
rect 20656 1705 20690 1756
rect 20774 2132 20808 2184
rect 21011 2184 21281 2223
rect 20774 1740 20808 1756
rect 20893 2132 20927 2148
rect 20893 1705 20927 1756
rect 21011 2132 21045 2184
rect 21011 1740 21045 1756
rect 21129 2132 21163 2148
rect 21129 1705 21163 1756
rect 21247 2132 21281 2184
rect 22743 2185 23013 2224
rect 22743 2132 22777 2185
rect 21484 1982 21754 2019
rect 21247 1740 21281 1756
rect 21366 1932 21400 1948
rect 19717 1666 21163 1705
rect 21366 1702 21400 1756
rect 21484 1932 21518 1982
rect 21484 1740 21518 1756
rect 21602 1932 21636 1948
rect 21602 1702 21636 1756
rect 21720 1932 21754 1982
rect 21720 1740 21754 1756
rect 22302 1983 22572 2022
rect 22302 1932 22336 1983
rect 22302 1740 22336 1756
rect 22420 1932 22454 1948
rect 21366 1663 21636 1702
rect 22420 1705 22454 1756
rect 22538 1932 22572 1983
rect 22538 1740 22572 1756
rect 22656 1932 22690 1948
rect 22656 1705 22690 1756
rect 22743 1740 22777 1756
rect 22861 2132 22895 2148
rect 22420 1666 22690 1705
rect 22861 1705 22895 1756
rect 22979 2132 23013 2185
rect 23210 2184 23480 2223
rect 22979 1740 23013 1756
rect 23097 2132 23131 2148
rect 23097 1705 23131 1756
rect 23210 2132 23244 2184
rect 23210 1740 23244 1756
rect 23328 2132 23362 2148
rect 23328 1705 23362 1756
rect 23446 2132 23480 2184
rect 23682 2184 23952 2223
rect 23446 1740 23480 1756
rect 23564 2132 23598 2148
rect 23564 1705 23598 1756
rect 23682 2132 23716 2184
rect 23682 1740 23716 1756
rect 23800 2132 23834 2148
rect 23800 1705 23834 1756
rect 23918 2132 23952 2184
rect 24155 2184 24425 2223
rect 23918 1740 23952 1756
rect 24037 2132 24071 2148
rect 24037 1705 24071 1756
rect 24155 2132 24189 2184
rect 24155 1740 24189 1756
rect 24273 2132 24307 2148
rect 24273 1705 24307 1756
rect 24391 2132 24425 2184
rect 24628 1982 24898 2019
rect 24391 1740 24425 1756
rect 24510 1932 24544 1948
rect 22861 1666 24307 1705
rect 24510 1702 24544 1756
rect 24628 1932 24662 1982
rect 24628 1740 24662 1756
rect 24746 1932 24780 1948
rect 24746 1702 24780 1756
rect 24864 1932 24898 1982
rect 24864 1740 24898 1756
rect 24510 1663 24780 1702
rect 1346 1537 1380 1553
rect 2640 1544 2656 1578
rect 2690 1544 2706 1578
rect 1346 1487 1380 1503
rect 4490 1537 4524 1553
rect 5784 1544 5800 1578
rect 5834 1544 5850 1578
rect 4490 1487 4524 1503
rect 7622 1541 7656 1557
rect 8916 1548 8932 1582
rect 8966 1548 8982 1582
rect 7622 1491 7656 1507
rect 10766 1541 10800 1557
rect 12060 1548 12076 1582
rect 12110 1548 12126 1582
rect 10766 1491 10800 1507
rect 13968 1537 14002 1553
rect 15262 1544 15278 1578
rect 15312 1544 15328 1578
rect 13968 1487 14002 1503
rect 17112 1537 17146 1553
rect 18406 1544 18422 1578
rect 18456 1544 18472 1578
rect 17112 1487 17146 1503
rect 20244 1541 20278 1557
rect 21538 1548 21554 1582
rect 21588 1548 21604 1582
rect 20244 1491 20278 1507
rect 23388 1541 23422 1557
rect 24682 1548 24698 1582
rect 24732 1548 24748 1582
rect 23388 1491 23422 1507
rect 117 1438 174 1442
rect 117 1378 121 1438
rect 170 1378 174 1438
rect 117 1374 174 1378
rect 349 1437 441 1454
rect 349 1382 365 1437
rect 425 1382 441 1437
rect 349 1369 441 1382
rect 1434 1438 1526 1451
rect 1434 1383 1450 1438
rect 1510 1383 1526 1438
rect 1434 1366 1526 1383
rect 3261 1438 3318 1442
rect 3261 1378 3265 1438
rect 3314 1378 3318 1438
rect 3261 1374 3318 1378
rect 3493 1437 3585 1454
rect 3493 1382 3509 1437
rect 3569 1382 3585 1437
rect 3493 1369 3585 1382
rect 4578 1438 4670 1451
rect 4578 1383 4594 1438
rect 4654 1383 4670 1438
rect 4578 1366 4670 1383
rect 6393 1442 6450 1446
rect 6393 1382 6397 1442
rect 6446 1382 6450 1442
rect 6393 1378 6450 1382
rect 6625 1441 6717 1458
rect 6625 1386 6641 1441
rect 6701 1386 6717 1441
rect 6625 1373 6717 1386
rect 7710 1442 7802 1455
rect 7710 1387 7726 1442
rect 7786 1387 7802 1442
rect 7710 1370 7802 1387
rect 9537 1442 9594 1446
rect 9537 1382 9541 1442
rect 9590 1382 9594 1442
rect 9537 1378 9594 1382
rect 9769 1441 9861 1458
rect 9769 1386 9785 1441
rect 9845 1386 9861 1441
rect 9769 1373 9861 1386
rect 10854 1442 10946 1455
rect 10854 1387 10870 1442
rect 10930 1387 10946 1442
rect 10854 1370 10946 1387
rect 12739 1438 12796 1442
rect 12739 1378 12743 1438
rect 12792 1378 12796 1438
rect 12739 1374 12796 1378
rect 12971 1437 13063 1454
rect 12971 1382 12987 1437
rect 13047 1382 13063 1437
rect 12971 1369 13063 1382
rect 14056 1438 14148 1451
rect 14056 1383 14072 1438
rect 14132 1383 14148 1438
rect 14056 1366 14148 1383
rect 15883 1438 15940 1442
rect 15883 1378 15887 1438
rect 15936 1378 15940 1438
rect 15883 1374 15940 1378
rect 16115 1437 16207 1454
rect 16115 1382 16131 1437
rect 16191 1382 16207 1437
rect 16115 1369 16207 1382
rect 17200 1438 17292 1451
rect 17200 1383 17216 1438
rect 17276 1383 17292 1438
rect 17200 1366 17292 1383
rect 19015 1442 19072 1446
rect 19015 1382 19019 1442
rect 19068 1382 19072 1442
rect 19015 1378 19072 1382
rect 19247 1441 19339 1458
rect 19247 1386 19263 1441
rect 19323 1386 19339 1441
rect 19247 1373 19339 1386
rect 20332 1442 20424 1455
rect 20332 1387 20348 1442
rect 20408 1387 20424 1442
rect 20332 1370 20424 1387
rect 22159 1442 22216 1446
rect 22159 1382 22163 1442
rect 22212 1382 22216 1442
rect 22159 1378 22216 1382
rect 22391 1441 22483 1458
rect 22391 1386 22407 1441
rect 22467 1386 22483 1441
rect 22391 1373 22483 1386
rect 23476 1442 23568 1455
rect 23476 1387 23492 1442
rect 23552 1387 23568 1442
rect 23476 1370 23568 1387
rect 6393 1326 6450 1330
rect 117 1322 174 1326
rect 117 1262 121 1322
rect 170 1262 174 1322
rect 117 1258 174 1262
rect 1700 1307 1734 1323
rect 1700 1257 1734 1273
rect 3261 1322 3318 1326
rect 3261 1262 3265 1322
rect 3314 1262 3318 1322
rect 3261 1258 3318 1262
rect 4844 1307 4878 1323
rect 4844 1257 4878 1273
rect 6393 1266 6397 1326
rect 6446 1266 6450 1326
rect 6393 1262 6450 1266
rect 7976 1311 8010 1327
rect 7976 1261 8010 1277
rect 9537 1326 9594 1330
rect 9537 1266 9541 1326
rect 9590 1266 9594 1326
rect 9537 1262 9594 1266
rect 11120 1311 11154 1327
rect 19015 1326 19072 1330
rect 11120 1261 11154 1277
rect 12739 1322 12796 1326
rect 12739 1262 12743 1322
rect 12792 1262 12796 1322
rect 12739 1258 12796 1262
rect 14322 1307 14356 1323
rect 14322 1257 14356 1273
rect 15883 1322 15940 1326
rect 15883 1262 15887 1322
rect 15936 1262 15940 1322
rect 15883 1258 15940 1262
rect 17466 1307 17500 1323
rect 17466 1257 17500 1273
rect 19015 1266 19019 1326
rect 19068 1266 19072 1326
rect 19015 1262 19072 1266
rect 20598 1311 20632 1327
rect 20598 1261 20632 1277
rect 22159 1326 22216 1330
rect 22159 1266 22163 1326
rect 22212 1266 22216 1326
rect 22159 1262 22216 1266
rect 23742 1311 23776 1327
rect 23742 1261 23776 1277
rect 117 1154 174 1158
rect 117 1094 121 1154
rect 170 1094 174 1154
rect 117 1090 174 1094
rect 1316 1153 1408 1166
rect 1316 1098 1332 1153
rect 1392 1098 1408 1153
rect 1316 1081 1408 1098
rect 3261 1154 3318 1158
rect 3261 1094 3265 1154
rect 3314 1094 3318 1154
rect 3261 1090 3318 1094
rect 4460 1153 4552 1166
rect 4460 1098 4476 1153
rect 4536 1098 4552 1153
rect 4460 1081 4552 1098
rect 6393 1158 6450 1162
rect 6393 1098 6397 1158
rect 6446 1098 6450 1158
rect 6393 1094 6450 1098
rect 7592 1157 7684 1170
rect 7592 1102 7608 1157
rect 7668 1102 7684 1157
rect 7592 1085 7684 1102
rect 9537 1158 9594 1162
rect 9537 1098 9541 1158
rect 9590 1098 9594 1158
rect 9537 1094 9594 1098
rect 10736 1157 10828 1170
rect 10736 1102 10752 1157
rect 10812 1102 10828 1157
rect 10736 1085 10828 1102
rect 12739 1154 12796 1158
rect 12739 1094 12743 1154
rect 12792 1094 12796 1154
rect 12739 1090 12796 1094
rect 13938 1153 14030 1166
rect 13938 1098 13954 1153
rect 14014 1098 14030 1153
rect 13938 1081 14030 1098
rect 15883 1154 15940 1158
rect 15883 1094 15887 1154
rect 15936 1094 15940 1154
rect 15883 1090 15940 1094
rect 17082 1153 17174 1166
rect 17082 1098 17098 1153
rect 17158 1098 17174 1153
rect 17082 1081 17174 1098
rect 19015 1158 19072 1162
rect 19015 1098 19019 1158
rect 19068 1098 19072 1158
rect 19015 1094 19072 1098
rect 20214 1157 20306 1170
rect 20214 1102 20230 1157
rect 20290 1102 20306 1157
rect 20214 1085 20306 1102
rect 22159 1158 22216 1162
rect 22159 1098 22163 1158
rect 22212 1098 22216 1158
rect 22159 1094 22216 1098
rect 23358 1157 23450 1170
rect 23358 1102 23374 1157
rect 23434 1102 23450 1157
rect 23358 1085 23450 1102
rect 1581 917 1615 933
rect 1581 867 1615 883
rect 4725 917 4759 933
rect 4725 867 4759 883
rect 7857 921 7891 937
rect 7857 871 7891 887
rect 11001 921 11035 937
rect 11001 871 11035 887
rect 14203 917 14237 933
rect 14203 867 14237 883
rect 17347 917 17381 933
rect 17347 867 17381 883
rect 20479 921 20513 937
rect 20479 871 20513 887
rect 23623 921 23657 937
rect 23623 871 23657 887
rect 1094 795 1128 811
rect 1094 603 1128 619
rect 1212 807 1246 811
rect 1286 807 1320 811
rect 1212 795 1320 807
rect 1246 619 1286 795
rect 1212 607 1286 619
rect 1212 603 1246 607
rect 1286 403 1320 419
rect 1404 795 1438 811
rect 1404 403 1438 419
rect 1522 795 1556 811
rect 1522 403 1556 419
rect 1640 795 1674 811
rect 1640 403 1674 419
rect 1758 807 1792 811
rect 1836 807 1870 811
rect 1758 795 1870 807
rect 1792 619 1836 795
rect 1792 607 1870 619
rect 1836 603 1870 607
rect 1954 795 1988 811
rect 1954 603 1988 619
rect 4238 795 4272 811
rect 4238 603 4272 619
rect 4356 807 4390 811
rect 4430 807 4464 811
rect 4356 795 4464 807
rect 4390 619 4430 795
rect 4356 607 4430 619
rect 4356 603 4390 607
rect 1758 403 1792 419
rect 4430 403 4464 419
rect 4548 795 4582 811
rect 4548 403 4582 419
rect 4666 795 4700 811
rect 4666 403 4700 419
rect 4784 795 4818 811
rect 4784 403 4818 419
rect 4902 807 4936 811
rect 4980 807 5014 811
rect 4902 795 5014 807
rect 4936 619 4980 795
rect 4936 607 5014 619
rect 4980 603 5014 607
rect 5098 795 5132 811
rect 5098 603 5132 619
rect 7370 799 7404 815
rect 7370 607 7404 623
rect 7488 811 7522 815
rect 7562 811 7596 815
rect 7488 799 7596 811
rect 7522 623 7562 799
rect 7488 611 7562 623
rect 7488 607 7522 611
rect 4902 403 4936 419
rect 7562 407 7596 423
rect 7680 799 7714 815
rect 7680 407 7714 423
rect 7798 799 7832 815
rect 7798 407 7832 423
rect 7916 799 7950 815
rect 7916 407 7950 423
rect 8034 811 8068 815
rect 8112 811 8146 815
rect 8034 799 8146 811
rect 8068 623 8112 799
rect 8068 611 8146 623
rect 8112 607 8146 611
rect 8230 799 8264 815
rect 8230 607 8264 623
rect 10514 799 10548 815
rect 10514 607 10548 623
rect 10632 811 10666 815
rect 10706 811 10740 815
rect 10632 799 10740 811
rect 10666 623 10706 799
rect 10632 611 10706 623
rect 10632 607 10666 611
rect 8034 407 8068 423
rect 10706 407 10740 423
rect 10824 799 10858 815
rect 10824 407 10858 423
rect 10942 799 10976 815
rect 10942 407 10976 423
rect 11060 799 11094 815
rect 11060 407 11094 423
rect 11178 811 11212 815
rect 11256 811 11290 815
rect 11178 799 11290 811
rect 11212 623 11256 799
rect 11212 611 11290 623
rect 11256 607 11290 611
rect 11374 799 11408 815
rect 11374 607 11408 623
rect 13716 795 13750 811
rect 13716 603 13750 619
rect 13834 807 13868 811
rect 13908 807 13942 811
rect 13834 795 13942 807
rect 13868 619 13908 795
rect 13834 607 13908 619
rect 13834 603 13868 607
rect 11178 407 11212 423
rect 13908 403 13942 419
rect 14026 795 14060 811
rect 14026 403 14060 419
rect 14144 795 14178 811
rect 14144 403 14178 419
rect 14262 795 14296 811
rect 14262 403 14296 419
rect 14380 807 14414 811
rect 14458 807 14492 811
rect 14380 795 14492 807
rect 14414 619 14458 795
rect 14414 607 14492 619
rect 14458 603 14492 607
rect 14576 795 14610 811
rect 14576 603 14610 619
rect 16860 795 16894 811
rect 16860 603 16894 619
rect 16978 807 17012 811
rect 17052 807 17086 811
rect 16978 795 17086 807
rect 17012 619 17052 795
rect 16978 607 17052 619
rect 16978 603 17012 607
rect 14380 403 14414 419
rect 17052 403 17086 419
rect 17170 795 17204 811
rect 17170 403 17204 419
rect 17288 795 17322 811
rect 17288 403 17322 419
rect 17406 795 17440 811
rect 17406 403 17440 419
rect 17524 807 17558 811
rect 17602 807 17636 811
rect 17524 795 17636 807
rect 17558 619 17602 795
rect 17558 607 17636 619
rect 17602 603 17636 607
rect 17720 795 17754 811
rect 17720 603 17754 619
rect 19992 799 20026 815
rect 19992 607 20026 623
rect 20110 811 20144 815
rect 20184 811 20218 815
rect 20110 799 20218 811
rect 20144 623 20184 799
rect 20110 611 20184 623
rect 20110 607 20144 611
rect 17524 403 17558 419
rect 20184 407 20218 423
rect 20302 799 20336 815
rect 20302 407 20336 423
rect 20420 799 20454 815
rect 20420 407 20454 423
rect 20538 799 20572 815
rect 20538 407 20572 423
rect 20656 811 20690 815
rect 20734 811 20768 815
rect 20656 799 20768 811
rect 20690 623 20734 799
rect 20690 611 20768 623
rect 20734 607 20768 611
rect 20852 799 20886 815
rect 20852 607 20886 623
rect 23136 799 23170 815
rect 23136 607 23170 623
rect 23254 811 23288 815
rect 23328 811 23362 815
rect 23254 799 23362 811
rect 23288 623 23328 799
rect 23254 611 23328 623
rect 23254 607 23288 611
rect 20656 407 20690 423
rect 23328 407 23362 423
rect 23446 799 23480 815
rect 23446 407 23480 423
rect 23564 799 23598 815
rect 23564 407 23598 423
rect 23682 799 23716 815
rect 23682 407 23716 423
rect 23800 811 23834 815
rect 23878 811 23912 815
rect 23800 799 23912 811
rect 23834 623 23878 799
rect 23834 611 23912 623
rect 23878 607 23912 611
rect 23996 799 24030 815
rect 23996 607 24030 623
rect 23800 407 23834 423
rect 1507 284 1523 318
rect 1557 284 1573 318
rect 4651 284 4667 318
rect 4701 284 4717 318
rect 7783 288 7799 322
rect 7833 288 7849 322
rect 10927 288 10943 322
rect 10977 288 10993 322
rect 14129 284 14145 318
rect 14179 284 14195 318
rect 17273 284 17289 318
rect 17323 284 17339 318
rect 20405 288 20421 322
rect 20455 288 20471 322
rect 23549 288 23565 322
rect 23599 288 23615 322
rect 7764 170 7900 174
rect 1488 166 1624 170
rect 1488 152 1526 166
rect 1584 152 1624 166
rect 1488 106 1504 152
rect 1608 106 1624 152
rect 1488 84 1624 106
rect 4632 166 4768 170
rect 4632 152 4670 166
rect 4728 152 4768 166
rect 4632 106 4648 152
rect 4752 106 4768 152
rect 4632 84 4768 106
rect 7764 156 7802 170
rect 7860 156 7900 170
rect 7764 110 7780 156
rect 7884 110 7900 156
rect 7764 88 7900 110
rect 10908 170 11044 174
rect 20386 170 20522 174
rect 10908 156 10946 170
rect 11004 156 11044 170
rect 10908 110 10924 156
rect 11028 110 11044 156
rect 10908 88 11044 110
rect 14110 166 14246 170
rect 14110 152 14148 166
rect 14206 152 14246 166
rect 14110 106 14126 152
rect 14230 106 14246 152
rect 14110 84 14246 106
rect 17254 166 17390 170
rect 17254 152 17292 166
rect 17350 152 17390 166
rect 17254 106 17270 152
rect 17374 106 17390 152
rect 17254 84 17390 106
rect 20386 156 20424 170
rect 20482 156 20522 170
rect 20386 110 20402 156
rect 20506 110 20522 156
rect 20386 88 20522 110
rect 23530 170 23666 174
rect 23530 156 23568 170
rect 23626 156 23666 170
rect 23530 110 23546 156
rect 23650 110 23666 156
rect 23530 88 23666 110
rect 1462 -1494 1690 -1476
rect 1462 -1570 1478 -1494
rect 1674 -1570 1690 -1494
rect 1462 -1586 1690 -1570
rect 4606 -1494 4834 -1476
rect 4606 -1570 4622 -1494
rect 4818 -1570 4834 -1494
rect 4606 -1586 4834 -1570
rect 7738 -1490 7966 -1472
rect 7738 -1566 7754 -1490
rect 7950 -1566 7966 -1490
rect 7738 -1582 7966 -1566
rect 10882 -1490 11110 -1472
rect 10882 -1566 10898 -1490
rect 11094 -1566 11110 -1490
rect 10882 -1582 11110 -1566
rect 14084 -1494 14312 -1476
rect 14084 -1570 14100 -1494
rect 14296 -1570 14312 -1494
rect 14084 -1586 14312 -1570
rect 17228 -1494 17456 -1476
rect 17228 -1570 17244 -1494
rect 17440 -1570 17456 -1494
rect 17228 -1586 17456 -1570
rect 20360 -1490 20588 -1472
rect 20360 -1566 20376 -1490
rect 20572 -1566 20588 -1490
rect 20360 -1582 20588 -1566
rect 23504 -1490 23732 -1472
rect 23504 -1566 23520 -1490
rect 23716 -1566 23732 -1490
rect 23504 -1582 23732 -1566
rect 733 -1711 1003 -1672
rect 733 -1764 767 -1711
rect 292 -1913 562 -1874
rect 292 -1964 326 -1913
rect 292 -2156 326 -2140
rect 410 -1964 444 -1948
rect 410 -2191 444 -2140
rect 528 -1964 562 -1913
rect 528 -2156 562 -2140
rect 646 -1964 680 -1948
rect 646 -2191 680 -2140
rect 733 -2156 767 -2140
rect 851 -1764 885 -1748
rect 410 -2230 680 -2191
rect 851 -2191 885 -2140
rect 969 -1764 1003 -1711
rect 1200 -1712 1470 -1673
rect 969 -2156 1003 -2140
rect 1087 -1764 1121 -1748
rect 1087 -2191 1121 -2140
rect 1200 -1764 1234 -1712
rect 1200 -2156 1234 -2140
rect 1318 -1764 1352 -1748
rect 1318 -2191 1352 -2140
rect 1436 -1764 1470 -1712
rect 1672 -1712 1942 -1673
rect 1436 -2156 1470 -2140
rect 1554 -1764 1588 -1748
rect 1554 -2191 1588 -2140
rect 1672 -1764 1706 -1712
rect 1672 -2156 1706 -2140
rect 1790 -1764 1824 -1748
rect 1790 -2191 1824 -2140
rect 1908 -1764 1942 -1712
rect 2145 -1712 2415 -1673
rect 1908 -2156 1942 -2140
rect 2027 -1764 2061 -1748
rect 2027 -2191 2061 -2140
rect 2145 -1764 2179 -1712
rect 2145 -2156 2179 -2140
rect 2263 -1764 2297 -1748
rect 2263 -2191 2297 -2140
rect 2381 -1764 2415 -1712
rect 3877 -1711 4147 -1672
rect 3877 -1764 3911 -1711
rect 2618 -1914 2888 -1877
rect 2381 -2156 2415 -2140
rect 2500 -1964 2534 -1948
rect 851 -2230 2297 -2191
rect 2500 -2194 2534 -2140
rect 2618 -1964 2652 -1914
rect 2618 -2156 2652 -2140
rect 2736 -1964 2770 -1948
rect 2736 -2194 2770 -2140
rect 2854 -1964 2888 -1914
rect 2854 -2156 2888 -2140
rect 3436 -1913 3706 -1874
rect 3436 -1964 3470 -1913
rect 3436 -2156 3470 -2140
rect 3554 -1964 3588 -1948
rect 2500 -2233 2770 -2194
rect 3554 -2191 3588 -2140
rect 3672 -1964 3706 -1913
rect 3672 -2156 3706 -2140
rect 3790 -1964 3824 -1948
rect 3790 -2191 3824 -2140
rect 3877 -2156 3911 -2140
rect 3995 -1764 4029 -1748
rect 3554 -2230 3824 -2191
rect 3995 -2191 4029 -2140
rect 4113 -1764 4147 -1711
rect 4344 -1712 4614 -1673
rect 4113 -2156 4147 -2140
rect 4231 -1764 4265 -1748
rect 4231 -2191 4265 -2140
rect 4344 -1764 4378 -1712
rect 4344 -2156 4378 -2140
rect 4462 -1764 4496 -1748
rect 4462 -2191 4496 -2140
rect 4580 -1764 4614 -1712
rect 4816 -1712 5086 -1673
rect 4580 -2156 4614 -2140
rect 4698 -1764 4732 -1748
rect 4698 -2191 4732 -2140
rect 4816 -1764 4850 -1712
rect 4816 -2156 4850 -2140
rect 4934 -1764 4968 -1748
rect 4934 -2191 4968 -2140
rect 5052 -1764 5086 -1712
rect 5289 -1712 5559 -1673
rect 5052 -2156 5086 -2140
rect 5171 -1764 5205 -1748
rect 5171 -2191 5205 -2140
rect 5289 -1764 5323 -1712
rect 5289 -2156 5323 -2140
rect 5407 -1764 5441 -1748
rect 5407 -2191 5441 -2140
rect 5525 -1764 5559 -1712
rect 7009 -1707 7279 -1668
rect 7009 -1760 7043 -1707
rect 5762 -1914 6032 -1877
rect 5525 -2156 5559 -2140
rect 5644 -1964 5678 -1948
rect 3995 -2230 5441 -2191
rect 5644 -2194 5678 -2140
rect 5762 -1964 5796 -1914
rect 5762 -2156 5796 -2140
rect 5880 -1964 5914 -1948
rect 5880 -2194 5914 -2140
rect 5998 -1964 6032 -1914
rect 5998 -2156 6032 -2140
rect 6568 -1909 6838 -1870
rect 6568 -1960 6602 -1909
rect 6568 -2152 6602 -2136
rect 6686 -1960 6720 -1944
rect 5644 -2233 5914 -2194
rect 6686 -2187 6720 -2136
rect 6804 -1960 6838 -1909
rect 6804 -2152 6838 -2136
rect 6922 -1960 6956 -1944
rect 6922 -2187 6956 -2136
rect 7009 -2152 7043 -2136
rect 7127 -1760 7161 -1744
rect 6686 -2226 6956 -2187
rect 7127 -2187 7161 -2136
rect 7245 -1760 7279 -1707
rect 7476 -1708 7746 -1669
rect 7245 -2152 7279 -2136
rect 7363 -1760 7397 -1744
rect 7363 -2187 7397 -2136
rect 7476 -1760 7510 -1708
rect 7476 -2152 7510 -2136
rect 7594 -1760 7628 -1744
rect 7594 -2187 7628 -2136
rect 7712 -1760 7746 -1708
rect 7948 -1708 8218 -1669
rect 7712 -2152 7746 -2136
rect 7830 -1760 7864 -1744
rect 7830 -2187 7864 -2136
rect 7948 -1760 7982 -1708
rect 7948 -2152 7982 -2136
rect 8066 -1760 8100 -1744
rect 8066 -2187 8100 -2136
rect 8184 -1760 8218 -1708
rect 8421 -1708 8691 -1669
rect 8184 -2152 8218 -2136
rect 8303 -1760 8337 -1744
rect 8303 -2187 8337 -2136
rect 8421 -1760 8455 -1708
rect 8421 -2152 8455 -2136
rect 8539 -1760 8573 -1744
rect 8539 -2187 8573 -2136
rect 8657 -1760 8691 -1708
rect 10153 -1707 10423 -1668
rect 10153 -1760 10187 -1707
rect 8894 -1910 9164 -1873
rect 8657 -2152 8691 -2136
rect 8776 -1960 8810 -1944
rect 7127 -2226 8573 -2187
rect 8776 -2190 8810 -2136
rect 8894 -1960 8928 -1910
rect 8894 -2152 8928 -2136
rect 9012 -1960 9046 -1944
rect 9012 -2190 9046 -2136
rect 9130 -1960 9164 -1910
rect 9130 -2152 9164 -2136
rect 9712 -1909 9982 -1870
rect 9712 -1960 9746 -1909
rect 9712 -2152 9746 -2136
rect 9830 -1960 9864 -1944
rect 8776 -2229 9046 -2190
rect 9830 -2187 9864 -2136
rect 9948 -1960 9982 -1909
rect 9948 -2152 9982 -2136
rect 10066 -1960 10100 -1944
rect 10066 -2187 10100 -2136
rect 10153 -2152 10187 -2136
rect 10271 -1760 10305 -1744
rect 9830 -2226 10100 -2187
rect 10271 -2187 10305 -2136
rect 10389 -1760 10423 -1707
rect 10620 -1708 10890 -1669
rect 10389 -2152 10423 -2136
rect 10507 -1760 10541 -1744
rect 10507 -2187 10541 -2136
rect 10620 -1760 10654 -1708
rect 10620 -2152 10654 -2136
rect 10738 -1760 10772 -1744
rect 10738 -2187 10772 -2136
rect 10856 -1760 10890 -1708
rect 11092 -1708 11362 -1669
rect 10856 -2152 10890 -2136
rect 10974 -1760 11008 -1744
rect 10974 -2187 11008 -2136
rect 11092 -1760 11126 -1708
rect 11092 -2152 11126 -2136
rect 11210 -1760 11244 -1744
rect 11210 -2187 11244 -2136
rect 11328 -1760 11362 -1708
rect 11565 -1708 11835 -1669
rect 11328 -2152 11362 -2136
rect 11447 -1760 11481 -1744
rect 11447 -2187 11481 -2136
rect 11565 -1760 11599 -1708
rect 11565 -2152 11599 -2136
rect 11683 -1760 11717 -1744
rect 11683 -2187 11717 -2136
rect 11801 -1760 11835 -1708
rect 13355 -1711 13625 -1672
rect 13355 -1764 13389 -1711
rect 12038 -1910 12308 -1873
rect 11801 -2152 11835 -2136
rect 11920 -1960 11954 -1944
rect 10271 -2226 11717 -2187
rect 11920 -2190 11954 -2136
rect 12038 -1960 12072 -1910
rect 12038 -2152 12072 -2136
rect 12156 -1960 12190 -1944
rect 12156 -2190 12190 -2136
rect 12274 -1960 12308 -1910
rect 12274 -2152 12308 -2136
rect 12914 -1913 13184 -1874
rect 12914 -1964 12948 -1913
rect 12914 -2156 12948 -2140
rect 13032 -1964 13066 -1948
rect 11920 -2229 12190 -2190
rect 13032 -2191 13066 -2140
rect 13150 -1964 13184 -1913
rect 13150 -2156 13184 -2140
rect 13268 -1964 13302 -1948
rect 13268 -2191 13302 -2140
rect 13355 -2156 13389 -2140
rect 13473 -1764 13507 -1748
rect 13032 -2230 13302 -2191
rect 13473 -2191 13507 -2140
rect 13591 -1764 13625 -1711
rect 13822 -1712 14092 -1673
rect 13591 -2156 13625 -2140
rect 13709 -1764 13743 -1748
rect 13709 -2191 13743 -2140
rect 13822 -1764 13856 -1712
rect 13822 -2156 13856 -2140
rect 13940 -1764 13974 -1748
rect 13940 -2191 13974 -2140
rect 14058 -1764 14092 -1712
rect 14294 -1712 14564 -1673
rect 14058 -2156 14092 -2140
rect 14176 -1764 14210 -1748
rect 14176 -2191 14210 -2140
rect 14294 -1764 14328 -1712
rect 14294 -2156 14328 -2140
rect 14412 -1764 14446 -1748
rect 14412 -2191 14446 -2140
rect 14530 -1764 14564 -1712
rect 14767 -1712 15037 -1673
rect 14530 -2156 14564 -2140
rect 14649 -1764 14683 -1748
rect 14649 -2191 14683 -2140
rect 14767 -1764 14801 -1712
rect 14767 -2156 14801 -2140
rect 14885 -1764 14919 -1748
rect 14885 -2191 14919 -2140
rect 15003 -1764 15037 -1712
rect 16499 -1711 16769 -1672
rect 16499 -1764 16533 -1711
rect 15240 -1914 15510 -1877
rect 15003 -2156 15037 -2140
rect 15122 -1964 15156 -1948
rect 13473 -2230 14919 -2191
rect 15122 -2194 15156 -2140
rect 15240 -1964 15274 -1914
rect 15240 -2156 15274 -2140
rect 15358 -1964 15392 -1948
rect 15358 -2194 15392 -2140
rect 15476 -1964 15510 -1914
rect 15476 -2156 15510 -2140
rect 16058 -1913 16328 -1874
rect 16058 -1964 16092 -1913
rect 16058 -2156 16092 -2140
rect 16176 -1964 16210 -1948
rect 15122 -2233 15392 -2194
rect 16176 -2191 16210 -2140
rect 16294 -1964 16328 -1913
rect 16294 -2156 16328 -2140
rect 16412 -1964 16446 -1948
rect 16412 -2191 16446 -2140
rect 16499 -2156 16533 -2140
rect 16617 -1764 16651 -1748
rect 16176 -2230 16446 -2191
rect 16617 -2191 16651 -2140
rect 16735 -1764 16769 -1711
rect 16966 -1712 17236 -1673
rect 16735 -2156 16769 -2140
rect 16853 -1764 16887 -1748
rect 16853 -2191 16887 -2140
rect 16966 -1764 17000 -1712
rect 16966 -2156 17000 -2140
rect 17084 -1764 17118 -1748
rect 17084 -2191 17118 -2140
rect 17202 -1764 17236 -1712
rect 17438 -1712 17708 -1673
rect 17202 -2156 17236 -2140
rect 17320 -1764 17354 -1748
rect 17320 -2191 17354 -2140
rect 17438 -1764 17472 -1712
rect 17438 -2156 17472 -2140
rect 17556 -1764 17590 -1748
rect 17556 -2191 17590 -2140
rect 17674 -1764 17708 -1712
rect 17911 -1712 18181 -1673
rect 17674 -2156 17708 -2140
rect 17793 -1764 17827 -1748
rect 17793 -2191 17827 -2140
rect 17911 -1764 17945 -1712
rect 17911 -2156 17945 -2140
rect 18029 -1764 18063 -1748
rect 18029 -2191 18063 -2140
rect 18147 -1764 18181 -1712
rect 19631 -1707 19901 -1668
rect 19631 -1760 19665 -1707
rect 18384 -1914 18654 -1877
rect 18147 -2156 18181 -2140
rect 18266 -1964 18300 -1948
rect 16617 -2230 18063 -2191
rect 18266 -2194 18300 -2140
rect 18384 -1964 18418 -1914
rect 18384 -2156 18418 -2140
rect 18502 -1964 18536 -1948
rect 18502 -2194 18536 -2140
rect 18620 -1964 18654 -1914
rect 18620 -2156 18654 -2140
rect 19190 -1909 19460 -1870
rect 19190 -1960 19224 -1909
rect 19190 -2152 19224 -2136
rect 19308 -1960 19342 -1944
rect 18266 -2233 18536 -2194
rect 19308 -2187 19342 -2136
rect 19426 -1960 19460 -1909
rect 19426 -2152 19460 -2136
rect 19544 -1960 19578 -1944
rect 19544 -2187 19578 -2136
rect 19631 -2152 19665 -2136
rect 19749 -1760 19783 -1744
rect 19308 -2226 19578 -2187
rect 19749 -2187 19783 -2136
rect 19867 -1760 19901 -1707
rect 20098 -1708 20368 -1669
rect 19867 -2152 19901 -2136
rect 19985 -1760 20019 -1744
rect 19985 -2187 20019 -2136
rect 20098 -1760 20132 -1708
rect 20098 -2152 20132 -2136
rect 20216 -1760 20250 -1744
rect 20216 -2187 20250 -2136
rect 20334 -1760 20368 -1708
rect 20570 -1708 20840 -1669
rect 20334 -2152 20368 -2136
rect 20452 -1760 20486 -1744
rect 20452 -2187 20486 -2136
rect 20570 -1760 20604 -1708
rect 20570 -2152 20604 -2136
rect 20688 -1760 20722 -1744
rect 20688 -2187 20722 -2136
rect 20806 -1760 20840 -1708
rect 21043 -1708 21313 -1669
rect 20806 -2152 20840 -2136
rect 20925 -1760 20959 -1744
rect 20925 -2187 20959 -2136
rect 21043 -1760 21077 -1708
rect 21043 -2152 21077 -2136
rect 21161 -1760 21195 -1744
rect 21161 -2187 21195 -2136
rect 21279 -1760 21313 -1708
rect 22775 -1707 23045 -1668
rect 22775 -1760 22809 -1707
rect 21516 -1910 21786 -1873
rect 21279 -2152 21313 -2136
rect 21398 -1960 21432 -1944
rect 19749 -2226 21195 -2187
rect 21398 -2190 21432 -2136
rect 21516 -1960 21550 -1910
rect 21516 -2152 21550 -2136
rect 21634 -1960 21668 -1944
rect 21634 -2190 21668 -2136
rect 21752 -1960 21786 -1910
rect 21752 -2152 21786 -2136
rect 22334 -1909 22604 -1870
rect 22334 -1960 22368 -1909
rect 22334 -2152 22368 -2136
rect 22452 -1960 22486 -1944
rect 21398 -2229 21668 -2190
rect 22452 -2187 22486 -2136
rect 22570 -1960 22604 -1909
rect 22570 -2152 22604 -2136
rect 22688 -1960 22722 -1944
rect 22688 -2187 22722 -2136
rect 22775 -2152 22809 -2136
rect 22893 -1760 22927 -1744
rect 22452 -2226 22722 -2187
rect 22893 -2187 22927 -2136
rect 23011 -1760 23045 -1707
rect 23242 -1708 23512 -1669
rect 23011 -2152 23045 -2136
rect 23129 -1760 23163 -1744
rect 23129 -2187 23163 -2136
rect 23242 -1760 23276 -1708
rect 23242 -2152 23276 -2136
rect 23360 -1760 23394 -1744
rect 23360 -2187 23394 -2136
rect 23478 -1760 23512 -1708
rect 23714 -1708 23984 -1669
rect 23478 -2152 23512 -2136
rect 23596 -1760 23630 -1744
rect 23596 -2187 23630 -2136
rect 23714 -1760 23748 -1708
rect 23714 -2152 23748 -2136
rect 23832 -1760 23866 -1744
rect 23832 -2187 23866 -2136
rect 23950 -1760 23984 -1708
rect 24187 -1708 24457 -1669
rect 23950 -2152 23984 -2136
rect 24069 -1760 24103 -1744
rect 24069 -2187 24103 -2136
rect 24187 -1760 24221 -1708
rect 24187 -2152 24221 -2136
rect 24305 -1760 24339 -1744
rect 24305 -2187 24339 -2136
rect 24423 -1760 24457 -1708
rect 24660 -1910 24930 -1873
rect 24423 -2152 24457 -2136
rect 24542 -1960 24576 -1944
rect 22893 -2226 24339 -2187
rect 24542 -2190 24576 -2136
rect 24660 -1960 24694 -1910
rect 24660 -2152 24694 -2136
rect 24778 -1960 24812 -1944
rect 24778 -2190 24812 -2136
rect 24896 -1960 24930 -1910
rect 24896 -2152 24930 -2136
rect 24542 -2229 24812 -2190
rect 1378 -2355 1412 -2339
rect 2672 -2348 2688 -2314
rect 2722 -2348 2738 -2314
rect 1378 -2405 1412 -2389
rect 4522 -2355 4556 -2339
rect 5816 -2348 5832 -2314
rect 5866 -2348 5882 -2314
rect 4522 -2405 4556 -2389
rect 7654 -2351 7688 -2335
rect 8948 -2344 8964 -2310
rect 8998 -2344 9014 -2310
rect 7654 -2401 7688 -2385
rect 10798 -2351 10832 -2335
rect 12092 -2344 12108 -2310
rect 12142 -2344 12158 -2310
rect 10798 -2401 10832 -2385
rect 14000 -2355 14034 -2339
rect 15294 -2348 15310 -2314
rect 15344 -2348 15360 -2314
rect 14000 -2405 14034 -2389
rect 17144 -2355 17178 -2339
rect 18438 -2348 18454 -2314
rect 18488 -2348 18504 -2314
rect 17144 -2405 17178 -2389
rect 20276 -2351 20310 -2335
rect 21570 -2344 21586 -2310
rect 21620 -2344 21636 -2310
rect 20276 -2401 20310 -2385
rect 23420 -2351 23454 -2335
rect 24714 -2344 24730 -2310
rect 24764 -2344 24780 -2310
rect 23420 -2401 23454 -2385
rect 149 -2454 206 -2450
rect 149 -2514 153 -2454
rect 202 -2514 206 -2454
rect 149 -2518 206 -2514
rect 381 -2455 473 -2438
rect 381 -2510 397 -2455
rect 457 -2510 473 -2455
rect 381 -2523 473 -2510
rect 1466 -2454 1558 -2441
rect 1466 -2509 1482 -2454
rect 1542 -2509 1558 -2454
rect 1466 -2526 1558 -2509
rect 3293 -2454 3350 -2450
rect 3293 -2514 3297 -2454
rect 3346 -2514 3350 -2454
rect 3293 -2518 3350 -2514
rect 3525 -2455 3617 -2438
rect 3525 -2510 3541 -2455
rect 3601 -2510 3617 -2455
rect 3525 -2523 3617 -2510
rect 4610 -2454 4702 -2441
rect 4610 -2509 4626 -2454
rect 4686 -2509 4702 -2454
rect 4610 -2526 4702 -2509
rect 6425 -2450 6482 -2446
rect 6425 -2510 6429 -2450
rect 6478 -2510 6482 -2450
rect 6425 -2514 6482 -2510
rect 6657 -2451 6749 -2434
rect 6657 -2506 6673 -2451
rect 6733 -2506 6749 -2451
rect 6657 -2519 6749 -2506
rect 7742 -2450 7834 -2437
rect 7742 -2505 7758 -2450
rect 7818 -2505 7834 -2450
rect 7742 -2522 7834 -2505
rect 9569 -2450 9626 -2446
rect 9569 -2510 9573 -2450
rect 9622 -2510 9626 -2450
rect 9569 -2514 9626 -2510
rect 9801 -2451 9893 -2434
rect 9801 -2506 9817 -2451
rect 9877 -2506 9893 -2451
rect 9801 -2519 9893 -2506
rect 10886 -2450 10978 -2437
rect 10886 -2505 10902 -2450
rect 10962 -2505 10978 -2450
rect 10886 -2522 10978 -2505
rect 12771 -2454 12828 -2450
rect 12771 -2514 12775 -2454
rect 12824 -2514 12828 -2454
rect 12771 -2518 12828 -2514
rect 13003 -2455 13095 -2438
rect 13003 -2510 13019 -2455
rect 13079 -2510 13095 -2455
rect 13003 -2523 13095 -2510
rect 14088 -2454 14180 -2441
rect 14088 -2509 14104 -2454
rect 14164 -2509 14180 -2454
rect 14088 -2526 14180 -2509
rect 15915 -2454 15972 -2450
rect 15915 -2514 15919 -2454
rect 15968 -2514 15972 -2454
rect 15915 -2518 15972 -2514
rect 16147 -2455 16239 -2438
rect 16147 -2510 16163 -2455
rect 16223 -2510 16239 -2455
rect 16147 -2523 16239 -2510
rect 17232 -2454 17324 -2441
rect 17232 -2509 17248 -2454
rect 17308 -2509 17324 -2454
rect 17232 -2526 17324 -2509
rect 19047 -2450 19104 -2446
rect 19047 -2510 19051 -2450
rect 19100 -2510 19104 -2450
rect 19047 -2514 19104 -2510
rect 19279 -2451 19371 -2434
rect 19279 -2506 19295 -2451
rect 19355 -2506 19371 -2451
rect 19279 -2519 19371 -2506
rect 20364 -2450 20456 -2437
rect 20364 -2505 20380 -2450
rect 20440 -2505 20456 -2450
rect 20364 -2522 20456 -2505
rect 22191 -2450 22248 -2446
rect 22191 -2510 22195 -2450
rect 22244 -2510 22248 -2450
rect 22191 -2514 22248 -2510
rect 22423 -2451 22515 -2434
rect 22423 -2506 22439 -2451
rect 22499 -2506 22515 -2451
rect 22423 -2519 22515 -2506
rect 23508 -2450 23600 -2437
rect 23508 -2505 23524 -2450
rect 23584 -2505 23600 -2450
rect 23508 -2522 23600 -2505
rect 6425 -2566 6482 -2562
rect 149 -2570 206 -2566
rect 149 -2630 153 -2570
rect 202 -2630 206 -2570
rect 149 -2634 206 -2630
rect 1732 -2585 1766 -2569
rect 1732 -2635 1766 -2619
rect 3293 -2570 3350 -2566
rect 3293 -2630 3297 -2570
rect 3346 -2630 3350 -2570
rect 3293 -2634 3350 -2630
rect 4876 -2585 4910 -2569
rect 4876 -2635 4910 -2619
rect 6425 -2626 6429 -2566
rect 6478 -2626 6482 -2566
rect 6425 -2630 6482 -2626
rect 8008 -2581 8042 -2565
rect 8008 -2631 8042 -2615
rect 9569 -2566 9626 -2562
rect 9569 -2626 9573 -2566
rect 9622 -2626 9626 -2566
rect 9569 -2630 9626 -2626
rect 11152 -2581 11186 -2565
rect 19047 -2566 19104 -2562
rect 11152 -2631 11186 -2615
rect 12771 -2570 12828 -2566
rect 12771 -2630 12775 -2570
rect 12824 -2630 12828 -2570
rect 12771 -2634 12828 -2630
rect 14354 -2585 14388 -2569
rect 14354 -2635 14388 -2619
rect 15915 -2570 15972 -2566
rect 15915 -2630 15919 -2570
rect 15968 -2630 15972 -2570
rect 15915 -2634 15972 -2630
rect 17498 -2585 17532 -2569
rect 17498 -2635 17532 -2619
rect 19047 -2626 19051 -2566
rect 19100 -2626 19104 -2566
rect 19047 -2630 19104 -2626
rect 20630 -2581 20664 -2565
rect 20630 -2631 20664 -2615
rect 22191 -2566 22248 -2562
rect 22191 -2626 22195 -2566
rect 22244 -2626 22248 -2566
rect 22191 -2630 22248 -2626
rect 23774 -2581 23808 -2565
rect 23774 -2631 23808 -2615
rect 149 -2738 206 -2734
rect 149 -2798 153 -2738
rect 202 -2798 206 -2738
rect 149 -2802 206 -2798
rect 1348 -2739 1440 -2726
rect 1348 -2794 1364 -2739
rect 1424 -2794 1440 -2739
rect 1348 -2811 1440 -2794
rect 3293 -2738 3350 -2734
rect 3293 -2798 3297 -2738
rect 3346 -2798 3350 -2738
rect 3293 -2802 3350 -2798
rect 4492 -2739 4584 -2726
rect 4492 -2794 4508 -2739
rect 4568 -2794 4584 -2739
rect 4492 -2811 4584 -2794
rect 6425 -2734 6482 -2730
rect 6425 -2794 6429 -2734
rect 6478 -2794 6482 -2734
rect 6425 -2798 6482 -2794
rect 7624 -2735 7716 -2722
rect 7624 -2790 7640 -2735
rect 7700 -2790 7716 -2735
rect 7624 -2807 7716 -2790
rect 9569 -2734 9626 -2730
rect 9569 -2794 9573 -2734
rect 9622 -2794 9626 -2734
rect 9569 -2798 9626 -2794
rect 10768 -2735 10860 -2722
rect 10768 -2790 10784 -2735
rect 10844 -2790 10860 -2735
rect 10768 -2807 10860 -2790
rect 12771 -2738 12828 -2734
rect 12771 -2798 12775 -2738
rect 12824 -2798 12828 -2738
rect 12771 -2802 12828 -2798
rect 13970 -2739 14062 -2726
rect 13970 -2794 13986 -2739
rect 14046 -2794 14062 -2739
rect 13970 -2811 14062 -2794
rect 15915 -2738 15972 -2734
rect 15915 -2798 15919 -2738
rect 15968 -2798 15972 -2738
rect 15915 -2802 15972 -2798
rect 17114 -2739 17206 -2726
rect 17114 -2794 17130 -2739
rect 17190 -2794 17206 -2739
rect 17114 -2811 17206 -2794
rect 19047 -2734 19104 -2730
rect 19047 -2794 19051 -2734
rect 19100 -2794 19104 -2734
rect 19047 -2798 19104 -2794
rect 20246 -2735 20338 -2722
rect 20246 -2790 20262 -2735
rect 20322 -2790 20338 -2735
rect 20246 -2807 20338 -2790
rect 22191 -2734 22248 -2730
rect 22191 -2794 22195 -2734
rect 22244 -2794 22248 -2734
rect 22191 -2798 22248 -2794
rect 23390 -2735 23482 -2722
rect 23390 -2790 23406 -2735
rect 23466 -2790 23482 -2735
rect 23390 -2807 23482 -2790
rect 1613 -2975 1647 -2959
rect 1613 -3025 1647 -3009
rect 4757 -2975 4791 -2959
rect 4757 -3025 4791 -3009
rect 7889 -2971 7923 -2955
rect 7889 -3021 7923 -3005
rect 11033 -2971 11067 -2955
rect 11033 -3021 11067 -3005
rect 14235 -2975 14269 -2959
rect 14235 -3025 14269 -3009
rect 17379 -2975 17413 -2959
rect 17379 -3025 17413 -3009
rect 20511 -2971 20545 -2955
rect 20511 -3021 20545 -3005
rect 23655 -2971 23689 -2955
rect 23655 -3021 23689 -3005
rect 1126 -3097 1160 -3081
rect 1126 -3289 1160 -3273
rect 1244 -3085 1278 -3081
rect 1318 -3085 1352 -3081
rect 1244 -3097 1352 -3085
rect 1278 -3273 1318 -3097
rect 1244 -3285 1318 -3273
rect 1244 -3289 1278 -3285
rect 1318 -3489 1352 -3473
rect 1436 -3097 1470 -3081
rect 1436 -3489 1470 -3473
rect 1554 -3097 1588 -3081
rect 1554 -3489 1588 -3473
rect 1672 -3097 1706 -3081
rect 1672 -3489 1706 -3473
rect 1790 -3085 1824 -3081
rect 1868 -3085 1902 -3081
rect 1790 -3097 1902 -3085
rect 1824 -3273 1868 -3097
rect 1824 -3285 1902 -3273
rect 1868 -3289 1902 -3285
rect 1986 -3097 2020 -3081
rect 1986 -3289 2020 -3273
rect 4270 -3097 4304 -3081
rect 4270 -3289 4304 -3273
rect 4388 -3085 4422 -3081
rect 4462 -3085 4496 -3081
rect 4388 -3097 4496 -3085
rect 4422 -3273 4462 -3097
rect 4388 -3285 4462 -3273
rect 4388 -3289 4422 -3285
rect 1790 -3489 1824 -3473
rect 4462 -3489 4496 -3473
rect 4580 -3097 4614 -3081
rect 4580 -3489 4614 -3473
rect 4698 -3097 4732 -3081
rect 4698 -3489 4732 -3473
rect 4816 -3097 4850 -3081
rect 4816 -3489 4850 -3473
rect 4934 -3085 4968 -3081
rect 5012 -3085 5046 -3081
rect 4934 -3097 5046 -3085
rect 4968 -3273 5012 -3097
rect 4968 -3285 5046 -3273
rect 5012 -3289 5046 -3285
rect 5130 -3097 5164 -3081
rect 5130 -3289 5164 -3273
rect 7402 -3093 7436 -3077
rect 7402 -3285 7436 -3269
rect 7520 -3081 7554 -3077
rect 7594 -3081 7628 -3077
rect 7520 -3093 7628 -3081
rect 7554 -3269 7594 -3093
rect 7520 -3281 7594 -3269
rect 7520 -3285 7554 -3281
rect 4934 -3489 4968 -3473
rect 7594 -3485 7628 -3469
rect 7712 -3093 7746 -3077
rect 7712 -3485 7746 -3469
rect 7830 -3093 7864 -3077
rect 7830 -3485 7864 -3469
rect 7948 -3093 7982 -3077
rect 7948 -3485 7982 -3469
rect 8066 -3081 8100 -3077
rect 8144 -3081 8178 -3077
rect 8066 -3093 8178 -3081
rect 8100 -3269 8144 -3093
rect 8100 -3281 8178 -3269
rect 8144 -3285 8178 -3281
rect 8262 -3093 8296 -3077
rect 8262 -3285 8296 -3269
rect 10546 -3093 10580 -3077
rect 10546 -3285 10580 -3269
rect 10664 -3081 10698 -3077
rect 10738 -3081 10772 -3077
rect 10664 -3093 10772 -3081
rect 10698 -3269 10738 -3093
rect 10664 -3281 10738 -3269
rect 10664 -3285 10698 -3281
rect 8066 -3485 8100 -3469
rect 10738 -3485 10772 -3469
rect 10856 -3093 10890 -3077
rect 10856 -3485 10890 -3469
rect 10974 -3093 11008 -3077
rect 10974 -3485 11008 -3469
rect 11092 -3093 11126 -3077
rect 11092 -3485 11126 -3469
rect 11210 -3081 11244 -3077
rect 11288 -3081 11322 -3077
rect 11210 -3093 11322 -3081
rect 11244 -3269 11288 -3093
rect 11244 -3281 11322 -3269
rect 11288 -3285 11322 -3281
rect 11406 -3093 11440 -3077
rect 11406 -3285 11440 -3269
rect 13748 -3097 13782 -3081
rect 13748 -3289 13782 -3273
rect 13866 -3085 13900 -3081
rect 13940 -3085 13974 -3081
rect 13866 -3097 13974 -3085
rect 13900 -3273 13940 -3097
rect 13866 -3285 13940 -3273
rect 13866 -3289 13900 -3285
rect 11210 -3485 11244 -3469
rect 13940 -3489 13974 -3473
rect 14058 -3097 14092 -3081
rect 14058 -3489 14092 -3473
rect 14176 -3097 14210 -3081
rect 14176 -3489 14210 -3473
rect 14294 -3097 14328 -3081
rect 14294 -3489 14328 -3473
rect 14412 -3085 14446 -3081
rect 14490 -3085 14524 -3081
rect 14412 -3097 14524 -3085
rect 14446 -3273 14490 -3097
rect 14446 -3285 14524 -3273
rect 14490 -3289 14524 -3285
rect 14608 -3097 14642 -3081
rect 14608 -3289 14642 -3273
rect 16892 -3097 16926 -3081
rect 16892 -3289 16926 -3273
rect 17010 -3085 17044 -3081
rect 17084 -3085 17118 -3081
rect 17010 -3097 17118 -3085
rect 17044 -3273 17084 -3097
rect 17010 -3285 17084 -3273
rect 17010 -3289 17044 -3285
rect 14412 -3489 14446 -3473
rect 17084 -3489 17118 -3473
rect 17202 -3097 17236 -3081
rect 17202 -3489 17236 -3473
rect 17320 -3097 17354 -3081
rect 17320 -3489 17354 -3473
rect 17438 -3097 17472 -3081
rect 17438 -3489 17472 -3473
rect 17556 -3085 17590 -3081
rect 17634 -3085 17668 -3081
rect 17556 -3097 17668 -3085
rect 17590 -3273 17634 -3097
rect 17590 -3285 17668 -3273
rect 17634 -3289 17668 -3285
rect 17752 -3097 17786 -3081
rect 17752 -3289 17786 -3273
rect 20024 -3093 20058 -3077
rect 20024 -3285 20058 -3269
rect 20142 -3081 20176 -3077
rect 20216 -3081 20250 -3077
rect 20142 -3093 20250 -3081
rect 20176 -3269 20216 -3093
rect 20142 -3281 20216 -3269
rect 20142 -3285 20176 -3281
rect 17556 -3489 17590 -3473
rect 20216 -3485 20250 -3469
rect 20334 -3093 20368 -3077
rect 20334 -3485 20368 -3469
rect 20452 -3093 20486 -3077
rect 20452 -3485 20486 -3469
rect 20570 -3093 20604 -3077
rect 20570 -3485 20604 -3469
rect 20688 -3081 20722 -3077
rect 20766 -3081 20800 -3077
rect 20688 -3093 20800 -3081
rect 20722 -3269 20766 -3093
rect 20722 -3281 20800 -3269
rect 20766 -3285 20800 -3281
rect 20884 -3093 20918 -3077
rect 20884 -3285 20918 -3269
rect 23168 -3093 23202 -3077
rect 23168 -3285 23202 -3269
rect 23286 -3081 23320 -3077
rect 23360 -3081 23394 -3077
rect 23286 -3093 23394 -3081
rect 23320 -3269 23360 -3093
rect 23286 -3281 23360 -3269
rect 23286 -3285 23320 -3281
rect 20688 -3485 20722 -3469
rect 23360 -3485 23394 -3469
rect 23478 -3093 23512 -3077
rect 23478 -3485 23512 -3469
rect 23596 -3093 23630 -3077
rect 23596 -3485 23630 -3469
rect 23714 -3093 23748 -3077
rect 23714 -3485 23748 -3469
rect 23832 -3081 23866 -3077
rect 23910 -3081 23944 -3077
rect 23832 -3093 23944 -3081
rect 23866 -3269 23910 -3093
rect 23866 -3281 23944 -3269
rect 23910 -3285 23944 -3281
rect 24028 -3093 24062 -3077
rect 24028 -3285 24062 -3269
rect 23832 -3485 23866 -3469
rect 1539 -3608 1555 -3574
rect 1589 -3608 1605 -3574
rect 4683 -3608 4699 -3574
rect 4733 -3608 4749 -3574
rect 7815 -3604 7831 -3570
rect 7865 -3604 7881 -3570
rect 10959 -3604 10975 -3570
rect 11009 -3604 11025 -3570
rect 14161 -3608 14177 -3574
rect 14211 -3608 14227 -3574
rect 17305 -3608 17321 -3574
rect 17355 -3608 17371 -3574
rect 20437 -3604 20453 -3570
rect 20487 -3604 20503 -3570
rect 23581 -3604 23597 -3570
rect 23631 -3604 23647 -3570
rect 7796 -3722 7932 -3718
rect 1520 -3726 1656 -3722
rect 1520 -3740 1558 -3726
rect 1616 -3740 1656 -3726
rect 1520 -3786 1536 -3740
rect 1640 -3786 1656 -3740
rect 1520 -3808 1656 -3786
rect 4664 -3726 4800 -3722
rect 4664 -3740 4702 -3726
rect 4760 -3740 4800 -3726
rect 4664 -3786 4680 -3740
rect 4784 -3786 4800 -3740
rect 4664 -3808 4800 -3786
rect 7796 -3736 7834 -3722
rect 7892 -3736 7932 -3722
rect 7796 -3782 7812 -3736
rect 7916 -3782 7932 -3736
rect 7796 -3804 7932 -3782
rect 10940 -3722 11076 -3718
rect 20418 -3722 20554 -3718
rect 10940 -3736 10978 -3722
rect 11036 -3736 11076 -3722
rect 10940 -3782 10956 -3736
rect 11060 -3782 11076 -3736
rect 10940 -3804 11076 -3782
rect 14142 -3726 14278 -3722
rect 14142 -3740 14180 -3726
rect 14238 -3740 14278 -3726
rect 14142 -3786 14158 -3740
rect 14262 -3786 14278 -3740
rect 14142 -3808 14278 -3786
rect 17286 -3726 17422 -3722
rect 17286 -3740 17324 -3726
rect 17382 -3740 17422 -3726
rect 17286 -3786 17302 -3740
rect 17406 -3786 17422 -3740
rect 17286 -3808 17422 -3786
rect 20418 -3736 20456 -3722
rect 20514 -3736 20554 -3722
rect 20418 -3782 20434 -3736
rect 20538 -3782 20554 -3736
rect 20418 -3804 20554 -3782
rect 23562 -3722 23698 -3718
rect 23562 -3736 23600 -3722
rect 23658 -3736 23698 -3722
rect 23562 -3782 23578 -3736
rect 23682 -3782 23698 -3736
rect 23562 -3804 23698 -3782
<< viali >>
rect 1718 22176 1790 22230
rect 4862 22176 4934 22230
rect 7994 22180 8066 22234
rect 11138 22180 11210 22234
rect 14340 22176 14412 22230
rect 17484 22176 17556 22230
rect 20616 22180 20688 22234
rect 23760 22180 23832 22234
rect 466 21604 500 21780
rect 584 21604 618 21780
rect 702 21604 736 21780
rect 820 21604 854 21780
rect 907 21604 941 21980
rect 1025 21604 1059 21980
rect 1143 21604 1177 21980
rect 1261 21604 1295 21980
rect 1374 21604 1408 21980
rect 1492 21604 1526 21980
rect 1610 21604 1644 21980
rect 1728 21604 1762 21980
rect 1846 21604 1880 21980
rect 1964 21604 1998 21980
rect 2082 21604 2116 21980
rect 2201 21604 2235 21980
rect 2319 21604 2353 21980
rect 2437 21604 2471 21980
rect 2555 21604 2589 21980
rect 2674 21604 2708 21780
rect 2792 21604 2826 21780
rect 2910 21604 2944 21780
rect 3028 21604 3062 21780
rect 3610 21604 3644 21780
rect 3728 21604 3762 21780
rect 3846 21604 3880 21780
rect 3964 21604 3998 21780
rect 4051 21604 4085 21980
rect 4169 21604 4203 21980
rect 4287 21604 4321 21980
rect 4405 21604 4439 21980
rect 4518 21604 4552 21980
rect 4636 21604 4670 21980
rect 4754 21604 4788 21980
rect 4872 21604 4906 21980
rect 4990 21604 5024 21980
rect 5108 21604 5142 21980
rect 5226 21604 5260 21980
rect 5345 21604 5379 21980
rect 5463 21604 5497 21980
rect 5581 21604 5615 21980
rect 5699 21604 5733 21980
rect 5818 21604 5852 21780
rect 5936 21604 5970 21780
rect 6054 21604 6088 21780
rect 6172 21604 6206 21780
rect 6742 21608 6776 21784
rect 6860 21608 6894 21784
rect 6978 21608 7012 21784
rect 7096 21608 7130 21784
rect 7183 21608 7217 21984
rect 7301 21608 7335 21984
rect 7419 21608 7453 21984
rect 7537 21608 7571 21984
rect 7650 21608 7684 21984
rect 7768 21608 7802 21984
rect 7886 21608 7920 21984
rect 8004 21608 8038 21984
rect 8122 21608 8156 21984
rect 8240 21608 8274 21984
rect 8358 21608 8392 21984
rect 8477 21608 8511 21984
rect 8595 21608 8629 21984
rect 8713 21608 8747 21984
rect 8831 21608 8865 21984
rect 8950 21608 8984 21784
rect 9068 21608 9102 21784
rect 9186 21608 9220 21784
rect 9304 21608 9338 21784
rect 9886 21608 9920 21784
rect 10004 21608 10038 21784
rect 10122 21608 10156 21784
rect 10240 21608 10274 21784
rect 10327 21608 10361 21984
rect 10445 21608 10479 21984
rect 10563 21608 10597 21984
rect 10681 21608 10715 21984
rect 10794 21608 10828 21984
rect 10912 21608 10946 21984
rect 11030 21608 11064 21984
rect 11148 21608 11182 21984
rect 11266 21608 11300 21984
rect 11384 21608 11418 21984
rect 11502 21608 11536 21984
rect 11621 21608 11655 21984
rect 11739 21608 11773 21984
rect 11857 21608 11891 21984
rect 11975 21608 12009 21984
rect 12094 21608 12128 21784
rect 12212 21608 12246 21784
rect 12330 21608 12364 21784
rect 12448 21608 12482 21784
rect 13088 21604 13122 21780
rect 13206 21604 13240 21780
rect 13324 21604 13358 21780
rect 13442 21604 13476 21780
rect 13529 21604 13563 21980
rect 13647 21604 13681 21980
rect 13765 21604 13799 21980
rect 13883 21604 13917 21980
rect 13996 21604 14030 21980
rect 14114 21604 14148 21980
rect 14232 21604 14266 21980
rect 14350 21604 14384 21980
rect 14468 21604 14502 21980
rect 14586 21604 14620 21980
rect 14704 21604 14738 21980
rect 14823 21604 14857 21980
rect 14941 21604 14975 21980
rect 15059 21604 15093 21980
rect 15177 21604 15211 21980
rect 15296 21604 15330 21780
rect 15414 21604 15448 21780
rect 15532 21604 15566 21780
rect 15650 21604 15684 21780
rect 16232 21604 16266 21780
rect 16350 21604 16384 21780
rect 16468 21604 16502 21780
rect 16586 21604 16620 21780
rect 16673 21604 16707 21980
rect 16791 21604 16825 21980
rect 16909 21604 16943 21980
rect 17027 21604 17061 21980
rect 17140 21604 17174 21980
rect 17258 21604 17292 21980
rect 17376 21604 17410 21980
rect 17494 21604 17528 21980
rect 17612 21604 17646 21980
rect 17730 21604 17764 21980
rect 17848 21604 17882 21980
rect 17967 21604 18001 21980
rect 18085 21604 18119 21980
rect 18203 21604 18237 21980
rect 18321 21604 18355 21980
rect 18440 21604 18474 21780
rect 18558 21604 18592 21780
rect 18676 21604 18710 21780
rect 18794 21604 18828 21780
rect 19364 21608 19398 21784
rect 19482 21608 19516 21784
rect 19600 21608 19634 21784
rect 19718 21608 19752 21784
rect 19805 21608 19839 21984
rect 19923 21608 19957 21984
rect 20041 21608 20075 21984
rect 20159 21608 20193 21984
rect 20272 21608 20306 21984
rect 20390 21608 20424 21984
rect 20508 21608 20542 21984
rect 20626 21608 20660 21984
rect 20744 21608 20778 21984
rect 20862 21608 20896 21984
rect 20980 21608 21014 21984
rect 21099 21608 21133 21984
rect 21217 21608 21251 21984
rect 21335 21608 21369 21984
rect 21453 21608 21487 21984
rect 21572 21608 21606 21784
rect 21690 21608 21724 21784
rect 21808 21608 21842 21784
rect 21926 21608 21960 21784
rect 22508 21608 22542 21784
rect 22626 21608 22660 21784
rect 22744 21608 22778 21784
rect 22862 21608 22896 21784
rect 22949 21608 22983 21984
rect 23067 21608 23101 21984
rect 23185 21608 23219 21984
rect 23303 21608 23337 21984
rect 23416 21608 23450 21984
rect 23534 21608 23568 21984
rect 23652 21608 23686 21984
rect 23770 21608 23804 21984
rect 23888 21608 23922 21984
rect 24006 21608 24040 21984
rect 24124 21608 24158 21984
rect 24243 21608 24277 21984
rect 24361 21608 24395 21984
rect 24479 21608 24513 21984
rect 24597 21608 24631 21984
rect 24716 21608 24750 21784
rect 24834 21608 24868 21784
rect 24952 21608 24986 21784
rect 25070 21608 25104 21784
rect 2862 21396 2896 21430
rect 1552 21355 1586 21389
rect 6006 21396 6040 21430
rect 4696 21355 4730 21389
rect 9138 21400 9172 21434
rect 7828 21359 7862 21393
rect 12282 21400 12316 21434
rect 10972 21359 11006 21393
rect 15484 21396 15518 21430
rect 14174 21355 14208 21389
rect 18628 21396 18662 21430
rect 17318 21355 17352 21389
rect 21760 21400 21794 21434
rect 20450 21359 20484 21393
rect 24904 21400 24938 21434
rect 23594 21359 23628 21393
rect 327 21230 376 21290
rect 571 21234 629 21289
rect 629 21234 631 21289
rect 1656 21235 1658 21290
rect 1658 21235 1716 21290
rect 3715 21234 3773 21289
rect 3773 21234 3775 21289
rect 4800 21235 4802 21290
rect 4802 21235 4860 21290
rect 6847 21238 6905 21293
rect 6905 21238 6907 21293
rect 7932 21239 7934 21294
rect 7934 21239 7992 21294
rect 9991 21238 10049 21293
rect 10049 21238 10051 21293
rect 11076 21239 11078 21294
rect 11078 21239 11136 21294
rect 13193 21234 13251 21289
rect 13251 21234 13253 21289
rect 14278 21235 14280 21290
rect 14280 21235 14338 21290
rect 16337 21234 16395 21289
rect 16395 21234 16397 21289
rect 17422 21235 17424 21290
rect 17424 21235 17482 21290
rect 19469 21238 19527 21293
rect 19527 21238 19529 21293
rect 20554 21239 20556 21294
rect 20556 21239 20614 21294
rect 22613 21238 22671 21293
rect 22671 21238 22673 21293
rect 23698 21239 23700 21294
rect 23700 21239 23758 21294
rect 1906 21125 1940 21159
rect 3471 21114 3520 21174
rect 5050 21125 5084 21159
rect 8182 21129 8216 21163
rect 9747 21118 9796 21178
rect 11326 21129 11360 21163
rect 14528 21125 14562 21159
rect 16093 21114 16142 21174
rect 17672 21125 17706 21159
rect 327 20946 376 21006
rect 1538 20950 1540 21005
rect 1540 20950 1598 21005
rect 3471 20946 3520 21006
rect 4682 20950 4684 21005
rect 4684 20950 4742 21005
rect 6603 20950 6652 21010
rect 7814 20954 7816 21009
rect 7816 20954 7874 21009
rect 9747 20950 9796 21010
rect 10958 20954 10960 21009
rect 10960 20954 11018 21009
rect 12949 20946 12998 21006
rect 14160 20950 14162 21005
rect 14162 20950 14220 21005
rect 19225 21118 19274 21178
rect 20804 21129 20838 21163
rect 22369 21118 22418 21178
rect 23948 21129 23982 21163
rect 16093 20946 16142 21006
rect 17304 20950 17306 21005
rect 17306 20950 17364 21005
rect 19225 20950 19274 21010
rect 20436 20954 20438 21009
rect 20438 20954 20496 21009
rect 23580 20954 23582 21009
rect 23582 20954 23640 21009
rect 1787 20735 1821 20769
rect 4931 20735 4965 20769
rect 8063 20739 8097 20773
rect 11207 20739 11241 20773
rect 14409 20735 14443 20769
rect 17553 20735 17587 20769
rect 20685 20739 20719 20773
rect 23829 20739 23863 20773
rect 1300 20471 1334 20647
rect 1418 20471 1452 20647
rect 1492 20271 1526 20647
rect 1610 20271 1644 20647
rect 1728 20271 1762 20647
rect 1846 20271 1880 20647
rect 1964 20271 1998 20647
rect 2042 20471 2076 20647
rect 2160 20471 2194 20647
rect 4444 20471 4478 20647
rect 4562 20471 4596 20647
rect 4636 20271 4670 20647
rect 4754 20271 4788 20647
rect 4872 20271 4906 20647
rect 4990 20271 5024 20647
rect 5108 20271 5142 20647
rect 5186 20471 5220 20647
rect 5304 20471 5338 20647
rect 7576 20475 7610 20651
rect 7694 20475 7728 20651
rect 7768 20275 7802 20651
rect 7886 20275 7920 20651
rect 8004 20275 8038 20651
rect 8122 20275 8156 20651
rect 8240 20275 8274 20651
rect 8318 20475 8352 20651
rect 8436 20475 8470 20651
rect 10720 20475 10754 20651
rect 10838 20475 10872 20651
rect 10912 20275 10946 20651
rect 11030 20275 11064 20651
rect 11148 20275 11182 20651
rect 11266 20275 11300 20651
rect 11384 20275 11418 20651
rect 11462 20475 11496 20651
rect 11580 20475 11614 20651
rect 13922 20471 13956 20647
rect 14040 20471 14074 20647
rect 14114 20271 14148 20647
rect 14232 20271 14266 20647
rect 14350 20271 14384 20647
rect 14468 20271 14502 20647
rect 14586 20271 14620 20647
rect 14664 20471 14698 20647
rect 14782 20471 14816 20647
rect 17066 20471 17100 20647
rect 17184 20471 17218 20647
rect 17258 20271 17292 20647
rect 17376 20271 17410 20647
rect 17494 20271 17528 20647
rect 17612 20271 17646 20647
rect 17730 20271 17764 20647
rect 17808 20471 17842 20647
rect 17926 20471 17960 20647
rect 20198 20475 20232 20651
rect 20316 20475 20350 20651
rect 20390 20275 20424 20651
rect 20508 20275 20542 20651
rect 20626 20275 20660 20651
rect 20744 20275 20778 20651
rect 20862 20275 20896 20651
rect 20940 20475 20974 20651
rect 21058 20475 21092 20651
rect 23342 20475 23376 20651
rect 23460 20475 23494 20651
rect 23534 20275 23568 20651
rect 23652 20275 23686 20651
rect 23770 20275 23804 20651
rect 23888 20275 23922 20651
rect 24006 20275 24040 20651
rect 24084 20475 24118 20651
rect 24202 20475 24236 20651
rect 1729 20136 1763 20170
rect 4873 20136 4907 20170
rect 8005 20140 8039 20174
rect 11149 20140 11183 20174
rect 14351 20136 14385 20170
rect 17495 20136 17529 20170
rect 20627 20140 20661 20174
rect 23771 20140 23805 20174
rect 1732 20004 1790 20018
rect 1732 19972 1790 20004
rect 4876 20004 4934 20018
rect 4876 19972 4934 20004
rect 8008 20008 8066 20022
rect 8008 19976 8066 20008
rect 11152 20008 11210 20022
rect 11152 19976 11210 20008
rect 14354 20004 14412 20018
rect 14354 19972 14412 20004
rect 17498 20004 17556 20018
rect 17498 19972 17556 20004
rect 20630 20008 20688 20022
rect 20630 19976 20688 20008
rect 23774 20008 23832 20022
rect 23774 19976 23832 20008
rect 15230 16974 15310 17044
rect 15230 16972 15310 16974
rect 14582 16934 14616 16968
rect 16398 16974 16478 17044
rect 16398 16972 16478 16974
rect 15750 16934 15784 16968
rect 17566 16974 17646 17044
rect 17566 16972 17646 16974
rect 16918 16934 16952 16968
rect 18734 16974 18814 17044
rect 18734 16972 18814 16974
rect 18086 16934 18120 16968
rect 19908 16976 19988 17046
rect 19908 16974 19988 16976
rect 19260 16936 19294 16970
rect 21076 16976 21156 17046
rect 21076 16974 21156 16976
rect 20428 16936 20462 16970
rect 22244 16976 22324 17046
rect 22244 16974 22324 16976
rect 21596 16936 21630 16970
rect 23412 16976 23492 17046
rect 23412 16974 23492 16976
rect 22764 16936 22798 16970
rect 3250 16775 3310 16837
rect 4698 16775 4758 16837
rect 6196 16777 6256 16839
rect 7644 16777 7704 16839
rect 9164 16775 9224 16837
rect 10612 16775 10672 16837
rect 12110 16777 12170 16839
rect 13558 16777 13618 16839
rect 14582 16826 14616 16860
rect 15750 16826 15784 16860
rect 16918 16826 16952 16860
rect 18086 16826 18120 16860
rect 19260 16828 19294 16862
rect 20428 16828 20462 16862
rect 21596 16828 21630 16862
rect 22764 16828 22798 16862
rect 2909 16423 2943 16599
rect 3027 16423 3061 16599
rect 3145 16423 3179 16599
rect 3263 16423 3297 16599
rect 3381 16423 3415 16599
rect 3499 16423 3533 16599
rect 3617 16423 3651 16599
rect 3735 16423 3769 16599
rect 3853 16423 3887 16599
rect 3971 16423 4005 16599
rect 4357 16423 4391 16599
rect 4475 16423 4509 16599
rect 4593 16423 4627 16599
rect 4711 16423 4745 16599
rect 4829 16423 4863 16599
rect 4947 16423 4981 16599
rect 5065 16423 5099 16599
rect 5183 16423 5217 16599
rect 5301 16423 5335 16599
rect 5419 16423 5453 16599
rect 5855 16425 5889 16601
rect 5973 16425 6007 16601
rect 6091 16425 6125 16601
rect 6209 16425 6243 16601
rect 6327 16425 6361 16601
rect 6445 16425 6479 16601
rect 6563 16425 6597 16601
rect 6681 16425 6715 16601
rect 6799 16425 6833 16601
rect 6917 16425 6951 16601
rect 7303 16425 7337 16601
rect 7421 16425 7455 16601
rect 7539 16425 7573 16601
rect 7657 16425 7691 16601
rect 7775 16425 7809 16601
rect 7893 16425 7927 16601
rect 8011 16425 8045 16601
rect 8129 16425 8163 16601
rect 8247 16425 8281 16601
rect 8365 16425 8399 16601
rect 8823 16423 8857 16599
rect 8941 16423 8975 16599
rect 9059 16423 9093 16599
rect 9177 16423 9211 16599
rect 9295 16423 9329 16599
rect 9413 16423 9447 16599
rect 9531 16423 9565 16599
rect 9649 16423 9683 16599
rect 9767 16423 9801 16599
rect 9885 16423 9919 16599
rect 10271 16423 10305 16599
rect 10389 16423 10423 16599
rect 10507 16423 10541 16599
rect 10625 16423 10659 16599
rect 10743 16423 10777 16599
rect 10861 16423 10895 16599
rect 10979 16423 11013 16599
rect 11097 16423 11131 16599
rect 11215 16423 11249 16599
rect 11333 16423 11367 16599
rect 11769 16425 11803 16601
rect 11887 16425 11921 16601
rect 12005 16425 12039 16601
rect 12123 16425 12157 16601
rect 12241 16425 12275 16601
rect 12359 16425 12393 16601
rect 12477 16425 12511 16601
rect 12595 16425 12629 16601
rect 12713 16425 12747 16601
rect 12831 16425 12865 16601
rect 13217 16425 13251 16601
rect 13335 16425 13369 16601
rect 13453 16425 13487 16601
rect 13571 16425 13605 16601
rect 13689 16425 13723 16601
rect 13807 16425 13841 16601
rect 13925 16425 13959 16601
rect 14043 16425 14077 16601
rect 14161 16425 14195 16601
rect 14279 16425 14313 16601
rect 14672 16420 14706 16796
rect 14790 16420 14824 16796
rect 14908 16420 14942 16796
rect 15026 16420 15060 16796
rect 15144 16420 15178 16796
rect 15262 16420 15296 16796
rect 15380 16420 15414 16796
rect 15840 16420 15874 16796
rect 15958 16420 15992 16796
rect 16076 16420 16110 16796
rect 16194 16420 16228 16796
rect 16312 16420 16346 16796
rect 16430 16420 16464 16796
rect 16548 16420 16582 16796
rect 17008 16418 17042 16794
rect 17126 16418 17160 16794
rect 17244 16418 17278 16794
rect 17362 16418 17396 16794
rect 17480 16418 17514 16794
rect 17598 16418 17632 16794
rect 17716 16418 17750 16794
rect 18176 16420 18210 16796
rect 18294 16420 18328 16796
rect 18412 16420 18446 16796
rect 18530 16420 18564 16796
rect 18648 16420 18682 16796
rect 18766 16420 18800 16796
rect 18884 16420 18918 16796
rect 19350 16422 19384 16798
rect 19468 16422 19502 16798
rect 19586 16422 19620 16798
rect 19704 16422 19738 16798
rect 19822 16422 19856 16798
rect 19940 16422 19974 16798
rect 20058 16422 20092 16798
rect 20518 16420 20552 16796
rect 20636 16420 20670 16796
rect 20754 16420 20788 16796
rect 20872 16420 20906 16796
rect 20990 16420 21024 16796
rect 21108 16420 21142 16796
rect 21226 16420 21260 16796
rect 21686 16422 21720 16798
rect 21804 16422 21838 16798
rect 21922 16422 21956 16798
rect 22040 16422 22074 16798
rect 22158 16422 22192 16798
rect 22276 16422 22310 16798
rect 22394 16422 22428 16798
rect 22854 16420 22888 16796
rect 22972 16420 23006 16796
rect 23090 16420 23124 16796
rect 23208 16420 23242 16796
rect 23326 16420 23360 16796
rect 23444 16420 23478 16796
rect 23562 16420 23596 16796
rect 3676 16329 3710 16363
rect 5124 16329 5158 16363
rect 6622 16331 6656 16365
rect 8070 16331 8104 16365
rect 9590 16329 9624 16363
rect 11038 16329 11072 16363
rect 12536 16331 12570 16365
rect 13984 16331 14018 16365
rect 3558 16212 3592 16246
rect 5006 16212 5040 16246
rect 6504 16214 6538 16248
rect 7952 16214 7986 16248
rect 9472 16212 9506 16246
rect 10920 16212 10954 16246
rect 12418 16214 12452 16248
rect 13866 16214 13900 16248
rect 3146 15786 3180 16162
rect 3264 15786 3298 16162
rect 3382 15786 3416 16162
rect 3499 15986 3533 16162
rect 3617 15986 3651 16162
rect 4594 15786 4628 16162
rect 4712 15786 4746 16162
rect 4830 15786 4864 16162
rect 4947 15986 4981 16162
rect 5065 15986 5099 16162
rect 6092 15788 6126 16164
rect 6210 15788 6244 16164
rect 6328 15788 6362 16164
rect 6445 15988 6479 16164
rect 6563 15988 6597 16164
rect 7540 15788 7574 16164
rect 7658 15788 7692 16164
rect 7776 15788 7810 16164
rect 7893 15988 7927 16164
rect 8011 15988 8045 16164
rect 9060 15786 9094 16162
rect 9178 15786 9212 16162
rect 9296 15786 9330 16162
rect 9413 15986 9447 16162
rect 9531 15986 9565 16162
rect 10508 15786 10542 16162
rect 10626 15786 10660 16162
rect 10744 15786 10778 16162
rect 10861 15986 10895 16162
rect 10979 15986 11013 16162
rect 12006 15788 12040 16164
rect 12124 15788 12158 16164
rect 12242 15788 12276 16164
rect 12359 15988 12393 16164
rect 12477 15988 12511 16164
rect 13454 15788 13488 16164
rect 13572 15788 13606 16164
rect 13690 15788 13724 16164
rect 13807 15988 13841 16164
rect 13925 15988 13959 16164
rect 14877 16063 14911 16097
rect 16045 16063 16079 16097
rect 17213 16063 17247 16097
rect 14582 15834 14616 16010
rect 14700 15834 14734 16010
rect 14818 15834 14852 16010
rect 14936 15834 14970 16010
rect 15102 15830 15136 16006
rect 3205 15702 3239 15736
rect 3323 15702 3357 15736
rect 4653 15702 4687 15736
rect 4771 15702 4805 15736
rect 6151 15704 6185 15738
rect 6269 15704 6303 15738
rect 7599 15704 7633 15738
rect 7717 15704 7751 15738
rect 9119 15702 9153 15736
rect 9237 15702 9271 15736
rect 10567 15702 10601 15736
rect 10685 15702 10719 15736
rect 12065 15704 12099 15738
rect 12183 15704 12217 15738
rect 13513 15704 13547 15738
rect 13631 15704 13665 15738
rect 15220 15830 15254 16006
rect 15338 15830 15372 16006
rect 15456 15830 15490 16006
rect 15750 15836 15784 16012
rect 15868 15836 15902 16012
rect 15986 15836 16020 16012
rect 16104 15836 16138 16012
rect 16269 15836 16303 16012
rect 14766 15702 14832 15706
rect 3478 15579 3530 15625
rect 4926 15579 4978 15625
rect 6424 15581 6476 15627
rect 7872 15581 7924 15627
rect 9392 15579 9444 15625
rect 10840 15579 10892 15625
rect 12338 15581 12390 15627
rect 13786 15581 13838 15627
rect 14766 15636 14832 15702
rect 16387 15836 16421 16012
rect 16505 15836 16539 16012
rect 16623 15836 16657 16012
rect 16918 15836 16952 16012
rect 17036 15836 17070 16012
rect 17154 15836 17188 16012
rect 17272 15836 17306 16012
rect 17437 15836 17471 16012
rect 17555 15836 17589 16012
rect 17673 15836 17707 16012
rect 17791 15836 17825 16012
rect 15934 15702 16000 15706
rect 15934 15636 16000 15702
rect 17102 15702 17168 15706
rect 17102 15636 17168 15702
rect 4220 15038 4292 15092
rect 2968 14466 3002 14642
rect 3086 14466 3120 14642
rect 3204 14466 3238 14642
rect 3322 14466 3356 14642
rect 3409 14466 3443 14842
rect 3527 14466 3561 14842
rect 3645 14466 3679 14842
rect 3763 14466 3797 14842
rect 3876 14466 3910 14842
rect 3994 14466 4028 14842
rect 4112 14466 4146 14842
rect 4230 14466 4264 14842
rect 4348 14466 4382 14842
rect 4466 14466 4500 14842
rect 4584 14466 4618 14842
rect 4703 14466 4737 14842
rect 4821 14466 4855 14842
rect 4939 14466 4973 14842
rect 5057 14466 5091 14842
rect 5176 14466 5210 14642
rect 5294 14466 5328 14642
rect 5412 14466 5446 14642
rect 5530 14466 5564 14642
rect 5364 14258 5398 14292
rect 4054 14217 4088 14251
rect 3073 14096 3131 14151
rect 3131 14096 3133 14151
rect 4158 14097 4160 14152
rect 4160 14097 4218 14152
rect 2829 13976 2878 14036
rect 4408 13987 4442 14021
rect 2829 13808 2878 13868
rect 4040 13812 4042 13867
rect 4042 13812 4100 13867
rect 7364 15038 7436 15092
rect 6112 14466 6146 14642
rect 6230 14466 6264 14642
rect 6348 14466 6382 14642
rect 6466 14466 6500 14642
rect 6553 14466 6587 14842
rect 6671 14466 6705 14842
rect 6789 14466 6823 14842
rect 6907 14466 6941 14842
rect 7020 14466 7054 14842
rect 7138 14466 7172 14842
rect 7256 14466 7290 14842
rect 7374 14466 7408 14842
rect 7492 14466 7526 14842
rect 7610 14466 7644 14842
rect 7728 14466 7762 14842
rect 7847 14466 7881 14842
rect 7965 14466 7999 14842
rect 8083 14466 8117 14842
rect 8201 14466 8235 14842
rect 8320 14466 8354 14642
rect 8438 14466 8472 14642
rect 8556 14466 8590 14642
rect 8674 14466 8708 14642
rect 8508 14258 8542 14292
rect 7198 14217 7232 14251
rect 6217 14096 6275 14151
rect 6275 14096 6277 14151
rect 7302 14097 7304 14152
rect 7304 14097 7362 14152
rect 5973 13976 6022 14036
rect 7552 13987 7586 14021
rect 5973 13808 6022 13868
rect 7184 13812 7186 13867
rect 7186 13812 7244 13867
rect 18381 16063 18415 16097
rect 19555 16065 19589 16099
rect 20723 16065 20757 16099
rect 21891 16065 21925 16099
rect 23059 16065 23093 16099
rect 18086 15836 18120 16012
rect 18204 15836 18238 16012
rect 18322 15836 18356 16012
rect 18440 15836 18474 16012
rect 18606 15836 18640 16012
rect 18724 15836 18758 16012
rect 18842 15836 18876 16012
rect 18960 15836 18994 16012
rect 19260 15836 19294 16012
rect 19378 15836 19412 16012
rect 19496 15836 19530 16012
rect 19614 15836 19648 16012
rect 19778 15832 19812 16008
rect 19896 15832 19930 16008
rect 20014 15832 20048 16008
rect 20132 15832 20166 16008
rect 20428 15836 20462 16012
rect 20546 15836 20580 16012
rect 20664 15836 20698 16012
rect 20782 15836 20816 16012
rect 20947 15831 20981 16007
rect 18270 15702 18336 15706
rect 18270 15636 18336 15702
rect 19444 15704 19510 15708
rect 19444 15638 19510 15704
rect 21065 15831 21099 16007
rect 21183 15831 21217 16007
rect 21301 15831 21335 16007
rect 21596 15838 21630 16014
rect 21714 15838 21748 16014
rect 21832 15838 21866 16014
rect 21950 15838 21984 16014
rect 22115 15831 22149 16007
rect 22233 15831 22267 16007
rect 22351 15831 22385 16007
rect 22469 15831 22503 16007
rect 22764 15838 22798 16014
rect 22882 15838 22916 16014
rect 23000 15838 23034 16014
rect 23118 15838 23152 16014
rect 23283 15832 23317 16008
rect 20612 15704 20678 15708
rect 20612 15638 20678 15704
rect 10496 15042 10568 15096
rect 13640 15042 13712 15096
rect 9244 14470 9278 14646
rect 9362 14470 9396 14646
rect 9480 14470 9514 14646
rect 9598 14470 9632 14646
rect 9685 14470 9719 14846
rect 9803 14470 9837 14846
rect 9921 14470 9955 14846
rect 10039 14470 10073 14846
rect 10152 14470 10186 14846
rect 10270 14470 10304 14846
rect 10388 14470 10422 14846
rect 10506 14470 10540 14846
rect 10624 14470 10658 14846
rect 10742 14470 10776 14846
rect 10860 14470 10894 14846
rect 10979 14470 11013 14846
rect 11097 14470 11131 14846
rect 11215 14470 11249 14846
rect 11333 14470 11367 14846
rect 11452 14470 11486 14646
rect 11570 14470 11604 14646
rect 11688 14470 11722 14646
rect 11806 14470 11840 14646
rect 12388 14470 12422 14646
rect 12506 14470 12540 14646
rect 12624 14470 12658 14646
rect 12742 14470 12776 14646
rect 12829 14470 12863 14846
rect 12947 14470 12981 14846
rect 13065 14470 13099 14846
rect 13183 14470 13217 14846
rect 13296 14470 13330 14846
rect 13414 14470 13448 14846
rect 13532 14470 13566 14846
rect 13650 14470 13684 14846
rect 13768 14470 13802 14846
rect 13886 14470 13920 14846
rect 14004 14470 14038 14846
rect 14123 14470 14157 14846
rect 14241 14470 14275 14846
rect 14359 14470 14393 14846
rect 14477 14470 14511 14846
rect 14596 14470 14630 14646
rect 14714 14470 14748 14646
rect 14832 14470 14866 14646
rect 14950 14470 14984 14646
rect 11640 14262 11674 14296
rect 10330 14221 10364 14255
rect 14784 14262 14818 14296
rect 13474 14221 13508 14255
rect 9349 14100 9407 14155
rect 9407 14100 9409 14155
rect 10434 14101 10436 14156
rect 10436 14101 10494 14156
rect 12493 14100 12551 14155
rect 12551 14100 12553 14155
rect 13578 14101 13580 14156
rect 13580 14101 13638 14156
rect 9105 13980 9154 14040
rect 10684 13991 10718 14025
rect 12249 13980 12298 14040
rect 13828 13991 13862 14025
rect 9105 13812 9154 13872
rect 10316 13816 10318 13871
rect 10318 13816 10376 13871
rect 16842 15038 16914 15092
rect 15590 14466 15624 14642
rect 15708 14466 15742 14642
rect 15826 14466 15860 14642
rect 15944 14466 15978 14642
rect 16031 14466 16065 14842
rect 16149 14466 16183 14842
rect 16267 14466 16301 14842
rect 16385 14466 16419 14842
rect 16498 14466 16532 14842
rect 16616 14466 16650 14842
rect 16734 14466 16768 14842
rect 16852 14466 16886 14842
rect 16970 14466 17004 14842
rect 17088 14466 17122 14842
rect 17206 14466 17240 14842
rect 17325 14466 17359 14842
rect 17443 14466 17477 14842
rect 17561 14466 17595 14842
rect 17679 14466 17713 14842
rect 17798 14466 17832 14642
rect 17916 14466 17950 14642
rect 18034 14466 18068 14642
rect 18152 14466 18186 14642
rect 17986 14258 18020 14292
rect 16676 14217 16710 14251
rect 15695 14096 15753 14151
rect 15753 14096 15755 14151
rect 16780 14097 16782 14152
rect 16782 14097 16840 14152
rect 15451 13976 15500 14036
rect 17030 13987 17064 14021
rect 23401 15832 23435 16008
rect 23519 15832 23553 16008
rect 23637 15832 23671 16008
rect 21780 15704 21846 15708
rect 21780 15638 21846 15704
rect 22948 15704 23014 15708
rect 22948 15638 23014 15704
rect 19986 15038 20058 15092
rect 18734 14466 18768 14642
rect 18852 14466 18886 14642
rect 18970 14466 19004 14642
rect 19088 14466 19122 14642
rect 19175 14466 19209 14842
rect 19293 14466 19327 14842
rect 19411 14466 19445 14842
rect 19529 14466 19563 14842
rect 19642 14466 19676 14842
rect 19760 14466 19794 14842
rect 19878 14466 19912 14842
rect 19996 14466 20030 14842
rect 20114 14466 20148 14842
rect 20232 14466 20266 14842
rect 20350 14466 20384 14842
rect 20469 14466 20503 14842
rect 20587 14466 20621 14842
rect 20705 14466 20739 14842
rect 20823 14466 20857 14842
rect 20942 14466 20976 14642
rect 21060 14466 21094 14642
rect 21178 14466 21212 14642
rect 21296 14466 21330 14642
rect 21130 14258 21164 14292
rect 19820 14217 19854 14251
rect 23118 15042 23190 15096
rect 21866 14470 21900 14646
rect 21984 14470 22018 14646
rect 22102 14470 22136 14646
rect 22220 14470 22254 14646
rect 22307 14470 22341 14846
rect 22425 14470 22459 14846
rect 22543 14470 22577 14846
rect 22661 14470 22695 14846
rect 22774 14470 22808 14846
rect 22892 14470 22926 14846
rect 23010 14470 23044 14846
rect 23128 14470 23162 14846
rect 23246 14470 23280 14846
rect 23364 14470 23398 14846
rect 23482 14470 23516 14846
rect 23601 14470 23635 14846
rect 23719 14470 23753 14846
rect 23837 14470 23871 14846
rect 23955 14470 23989 14846
rect 24074 14470 24108 14646
rect 24192 14470 24226 14646
rect 24310 14470 24344 14646
rect 24428 14470 24462 14646
rect 24262 14262 24296 14296
rect 18839 14096 18897 14151
rect 18897 14096 18899 14151
rect 19924 14097 19926 14152
rect 19926 14097 19984 14152
rect 18595 13976 18644 14036
rect 20174 13987 20208 14021
rect 18595 13808 18644 13868
rect 19806 13812 19808 13867
rect 19808 13812 19866 13867
rect 22952 14221 22986 14255
rect 21971 14100 22029 14155
rect 22029 14100 22031 14155
rect 23056 14101 23058 14156
rect 23058 14101 23116 14156
rect 21727 13980 21776 14040
rect 23306 13991 23340 14025
rect 21727 13812 21776 13872
rect 22938 13816 22940 13871
rect 22940 13816 22998 13871
rect 26262 15042 26334 15096
rect 25010 14470 25044 14646
rect 25128 14470 25162 14646
rect 25246 14470 25280 14646
rect 25364 14470 25398 14646
rect 25451 14470 25485 14846
rect 25569 14470 25603 14846
rect 25687 14470 25721 14846
rect 25805 14470 25839 14846
rect 25918 14470 25952 14846
rect 26036 14470 26070 14846
rect 26154 14470 26188 14846
rect 26272 14470 26306 14846
rect 26390 14470 26424 14846
rect 26508 14470 26542 14846
rect 26626 14470 26660 14846
rect 26745 14470 26779 14846
rect 26863 14470 26897 14846
rect 26981 14470 27015 14846
rect 27099 14470 27133 14846
rect 27218 14470 27252 14646
rect 27336 14470 27370 14646
rect 27454 14470 27488 14646
rect 27572 14470 27606 14646
rect 27406 14262 27440 14296
rect 26096 14221 26130 14255
rect 25115 14100 25173 14155
rect 25173 14100 25175 14155
rect 26200 14101 26202 14156
rect 26202 14101 26260 14156
rect 24871 13980 24920 14040
rect 26450 13991 26484 14025
rect 24871 13812 24920 13872
rect 26082 13816 26084 13871
rect 26084 13816 26142 13871
rect 4289 13597 4323 13631
rect 7433 13597 7467 13631
rect 10565 13601 10599 13635
rect 13709 13601 13743 13635
rect 16911 13597 16945 13631
rect 20055 13597 20089 13631
rect 23187 13601 23221 13635
rect 26331 13601 26365 13635
rect 3802 13333 3836 13509
rect 3920 13333 3954 13509
rect 3994 13133 4028 13509
rect 4112 13133 4146 13509
rect 4230 13133 4264 13509
rect 4348 13133 4382 13509
rect 4466 13133 4500 13509
rect 4544 13333 4578 13509
rect 4662 13333 4696 13509
rect 6946 13333 6980 13509
rect 7064 13333 7098 13509
rect 7138 13133 7172 13509
rect 7256 13133 7290 13509
rect 7374 13133 7408 13509
rect 7492 13133 7526 13509
rect 7610 13133 7644 13509
rect 7688 13333 7722 13509
rect 7806 13333 7840 13509
rect 10078 13337 10112 13513
rect 10196 13337 10230 13513
rect 10270 13137 10304 13513
rect 10388 13137 10422 13513
rect 10506 13137 10540 13513
rect 10624 13137 10658 13513
rect 10742 13137 10776 13513
rect 10820 13337 10854 13513
rect 10938 13337 10972 13513
rect 13222 13337 13256 13513
rect 13340 13337 13374 13513
rect 13414 13137 13448 13513
rect 13532 13137 13566 13513
rect 13650 13137 13684 13513
rect 13768 13137 13802 13513
rect 13886 13137 13920 13513
rect 13964 13337 13998 13513
rect 14082 13337 14116 13513
rect 16424 13333 16458 13509
rect 16542 13333 16576 13509
rect 16616 13133 16650 13509
rect 16734 13133 16768 13509
rect 16852 13133 16886 13509
rect 16970 13133 17004 13509
rect 17088 13133 17122 13509
rect 17166 13333 17200 13509
rect 17284 13333 17318 13509
rect 19568 13333 19602 13509
rect 19686 13333 19720 13509
rect 19760 13133 19794 13509
rect 19878 13133 19912 13509
rect 19996 13133 20030 13509
rect 20114 13133 20148 13509
rect 20232 13133 20266 13509
rect 20310 13333 20344 13509
rect 20428 13333 20462 13509
rect 22700 13337 22734 13513
rect 22818 13337 22852 13513
rect 22892 13137 22926 13513
rect 23010 13137 23044 13513
rect 23128 13137 23162 13513
rect 23246 13137 23280 13513
rect 23364 13137 23398 13513
rect 23442 13337 23476 13513
rect 23560 13337 23594 13513
rect 25844 13337 25878 13513
rect 25962 13337 25996 13513
rect 26036 13137 26070 13513
rect 26154 13137 26188 13513
rect 26272 13137 26306 13513
rect 26390 13137 26424 13513
rect 26508 13137 26542 13513
rect 26586 13337 26620 13513
rect 26704 13337 26738 13513
rect 4231 12998 4265 13032
rect 7375 12998 7409 13032
rect 10507 13002 10541 13036
rect 13651 13002 13685 13036
rect 16853 12998 16887 13032
rect 19997 12998 20031 13032
rect 23129 13002 23163 13036
rect 26273 13002 26307 13036
rect 4234 12866 4292 12880
rect 4234 12834 4292 12866
rect 7378 12866 7436 12880
rect 7378 12834 7436 12866
rect 10510 12870 10568 12884
rect 10510 12838 10568 12870
rect 13654 12870 13712 12884
rect 13654 12838 13712 12870
rect 16856 12866 16914 12880
rect 16856 12834 16914 12866
rect 20000 12866 20058 12880
rect 20000 12834 20058 12866
rect 23132 12870 23190 12884
rect 23132 12838 23190 12870
rect 26276 12870 26334 12884
rect 26276 12838 26334 12870
rect 4220 12304 4292 12358
rect 7364 12304 7436 12358
rect 10496 12308 10568 12362
rect 13640 12308 13712 12362
rect 16842 12304 16914 12358
rect 19986 12304 20058 12358
rect 23118 12308 23190 12362
rect 26262 12308 26334 12362
rect 2968 11732 3002 11908
rect 3086 11732 3120 11908
rect 3204 11732 3238 11908
rect 3322 11732 3356 11908
rect 3409 11732 3443 12108
rect 3527 11732 3561 12108
rect 3645 11732 3679 12108
rect 3763 11732 3797 12108
rect 3876 11732 3910 12108
rect 3994 11732 4028 12108
rect 4112 11732 4146 12108
rect 4230 11732 4264 12108
rect 4348 11732 4382 12108
rect 4466 11732 4500 12108
rect 4584 11732 4618 12108
rect 4703 11732 4737 12108
rect 4821 11732 4855 12108
rect 4939 11732 4973 12108
rect 5057 11732 5091 12108
rect 5176 11732 5210 11908
rect 5294 11732 5328 11908
rect 5412 11732 5446 11908
rect 5530 11732 5564 11908
rect 6112 11732 6146 11908
rect 6230 11732 6264 11908
rect 6348 11732 6382 11908
rect 6466 11732 6500 11908
rect 6553 11732 6587 12108
rect 6671 11732 6705 12108
rect 6789 11732 6823 12108
rect 6907 11732 6941 12108
rect 7020 11732 7054 12108
rect 7138 11732 7172 12108
rect 7256 11732 7290 12108
rect 7374 11732 7408 12108
rect 7492 11732 7526 12108
rect 7610 11732 7644 12108
rect 7728 11732 7762 12108
rect 7847 11732 7881 12108
rect 7965 11732 7999 12108
rect 8083 11732 8117 12108
rect 8201 11732 8235 12108
rect 8320 11732 8354 11908
rect 8438 11732 8472 11908
rect 8556 11732 8590 11908
rect 8674 11732 8708 11908
rect 9244 11736 9278 11912
rect 9362 11736 9396 11912
rect 9480 11736 9514 11912
rect 9598 11736 9632 11912
rect 9685 11736 9719 12112
rect 9803 11736 9837 12112
rect 9921 11736 9955 12112
rect 10039 11736 10073 12112
rect 10152 11736 10186 12112
rect 10270 11736 10304 12112
rect 10388 11736 10422 12112
rect 10506 11736 10540 12112
rect 10624 11736 10658 12112
rect 10742 11736 10776 12112
rect 10860 11736 10894 12112
rect 10979 11736 11013 12112
rect 11097 11736 11131 12112
rect 11215 11736 11249 12112
rect 11333 11736 11367 12112
rect 11452 11736 11486 11912
rect 11570 11736 11604 11912
rect 11688 11736 11722 11912
rect 11806 11736 11840 11912
rect 12388 11736 12422 11912
rect 12506 11736 12540 11912
rect 12624 11736 12658 11912
rect 12742 11736 12776 11912
rect 12829 11736 12863 12112
rect 12947 11736 12981 12112
rect 13065 11736 13099 12112
rect 13183 11736 13217 12112
rect 13296 11736 13330 12112
rect 13414 11736 13448 12112
rect 13532 11736 13566 12112
rect 13650 11736 13684 12112
rect 13768 11736 13802 12112
rect 13886 11736 13920 12112
rect 14004 11736 14038 12112
rect 14123 11736 14157 12112
rect 14241 11736 14275 12112
rect 14359 11736 14393 12112
rect 14477 11736 14511 12112
rect 14596 11736 14630 11912
rect 14714 11736 14748 11912
rect 14832 11736 14866 11912
rect 14950 11736 14984 11912
rect 15590 11732 15624 11908
rect 15708 11732 15742 11908
rect 15826 11732 15860 11908
rect 15944 11732 15978 11908
rect 16031 11732 16065 12108
rect 16149 11732 16183 12108
rect 16267 11732 16301 12108
rect 16385 11732 16419 12108
rect 16498 11732 16532 12108
rect 16616 11732 16650 12108
rect 16734 11732 16768 12108
rect 16852 11732 16886 12108
rect 16970 11732 17004 12108
rect 17088 11732 17122 12108
rect 17206 11732 17240 12108
rect 17325 11732 17359 12108
rect 17443 11732 17477 12108
rect 17561 11732 17595 12108
rect 17679 11732 17713 12108
rect 17798 11732 17832 11908
rect 17916 11732 17950 11908
rect 18034 11732 18068 11908
rect 18152 11732 18186 11908
rect 18734 11732 18768 11908
rect 18852 11732 18886 11908
rect 18970 11732 19004 11908
rect 19088 11732 19122 11908
rect 19175 11732 19209 12108
rect 19293 11732 19327 12108
rect 19411 11732 19445 12108
rect 19529 11732 19563 12108
rect 19642 11732 19676 12108
rect 19760 11732 19794 12108
rect 19878 11732 19912 12108
rect 19996 11732 20030 12108
rect 20114 11732 20148 12108
rect 20232 11732 20266 12108
rect 20350 11732 20384 12108
rect 20469 11732 20503 12108
rect 20587 11732 20621 12108
rect 20705 11732 20739 12108
rect 20823 11732 20857 12108
rect 20942 11732 20976 11908
rect 21060 11732 21094 11908
rect 21178 11732 21212 11908
rect 21296 11732 21330 11908
rect 21866 11736 21900 11912
rect 21984 11736 22018 11912
rect 22102 11736 22136 11912
rect 22220 11736 22254 11912
rect 22307 11736 22341 12112
rect 22425 11736 22459 12112
rect 22543 11736 22577 12112
rect 22661 11736 22695 12112
rect 22774 11736 22808 12112
rect 22892 11736 22926 12112
rect 23010 11736 23044 12112
rect 23128 11736 23162 12112
rect 23246 11736 23280 12112
rect 23364 11736 23398 12112
rect 23482 11736 23516 12112
rect 23601 11736 23635 12112
rect 23719 11736 23753 12112
rect 23837 11736 23871 12112
rect 23955 11736 23989 12112
rect 24074 11736 24108 11912
rect 24192 11736 24226 11912
rect 24310 11736 24344 11912
rect 24428 11736 24462 11912
rect 25010 11736 25044 11912
rect 25128 11736 25162 11912
rect 25246 11736 25280 11912
rect 25364 11736 25398 11912
rect 25451 11736 25485 12112
rect 25569 11736 25603 12112
rect 25687 11736 25721 12112
rect 25805 11736 25839 12112
rect 25918 11736 25952 12112
rect 26036 11736 26070 12112
rect 26154 11736 26188 12112
rect 26272 11736 26306 12112
rect 26390 11736 26424 12112
rect 26508 11736 26542 12112
rect 26626 11736 26660 12112
rect 26745 11736 26779 12112
rect 26863 11736 26897 12112
rect 26981 11736 27015 12112
rect 27099 11736 27133 12112
rect 27218 11736 27252 11912
rect 27336 11736 27370 11912
rect 27454 11736 27488 11912
rect 27572 11736 27606 11912
rect 5364 11524 5398 11558
rect 4054 11483 4088 11517
rect 8508 11524 8542 11558
rect 7198 11483 7232 11517
rect 11640 11528 11674 11562
rect 10330 11487 10364 11521
rect 14784 11528 14818 11562
rect 13474 11487 13508 11521
rect 17986 11524 18020 11558
rect 16676 11483 16710 11517
rect 21130 11524 21164 11558
rect 19820 11483 19854 11517
rect 24262 11528 24296 11562
rect 22952 11487 22986 11521
rect 27406 11528 27440 11562
rect 26096 11487 26130 11521
rect 3073 11362 3131 11417
rect 3131 11362 3133 11417
rect 4158 11363 4160 11418
rect 4160 11363 4218 11418
rect 6217 11362 6275 11417
rect 6275 11362 6277 11417
rect 7302 11363 7304 11418
rect 7304 11363 7362 11418
rect 9349 11366 9407 11421
rect 9407 11366 9409 11421
rect 10434 11367 10436 11422
rect 10436 11367 10494 11422
rect 12493 11366 12551 11421
rect 12551 11366 12553 11421
rect 13578 11367 13580 11422
rect 13580 11367 13638 11422
rect 15695 11362 15753 11417
rect 15753 11362 15755 11417
rect 16780 11363 16782 11418
rect 16782 11363 16840 11418
rect 18595 11358 18644 11418
rect 18839 11362 18897 11417
rect 18897 11362 18899 11417
rect 19924 11363 19926 11418
rect 19926 11363 19984 11418
rect 21971 11366 22029 11421
rect 22029 11366 22031 11421
rect 23056 11367 23058 11422
rect 23058 11367 23116 11422
rect 25115 11366 25173 11421
rect 25173 11366 25175 11421
rect 26200 11367 26202 11422
rect 26202 11367 26260 11422
rect 2829 11242 2878 11302
rect 4408 11253 4442 11287
rect 5973 11242 6022 11302
rect 7552 11253 7586 11287
rect 9105 11246 9154 11306
rect 10684 11257 10718 11291
rect 12249 11246 12298 11306
rect 13828 11257 13862 11291
rect 15451 11242 15500 11302
rect 17030 11253 17064 11287
rect 18595 11242 18644 11302
rect 20174 11253 20208 11287
rect 21727 11246 21776 11306
rect 23306 11257 23340 11291
rect 24871 11246 24920 11306
rect 26450 11257 26484 11291
rect 2829 11074 2878 11134
rect 4040 11078 4042 11133
rect 4042 11078 4100 11133
rect 5973 11074 6022 11134
rect 7184 11078 7186 11133
rect 7186 11078 7244 11133
rect 9105 11078 9154 11138
rect 10316 11082 10318 11137
rect 10318 11082 10376 11137
rect 12249 11078 12298 11138
rect 13460 11082 13462 11137
rect 13462 11082 13520 11137
rect 15451 11074 15500 11134
rect 16662 11078 16664 11133
rect 16664 11078 16722 11133
rect 18595 11074 18644 11134
rect 19806 11078 19808 11133
rect 19808 11078 19866 11133
rect 21727 11078 21776 11138
rect 22938 11082 22940 11137
rect 22940 11082 22998 11137
rect 24871 11078 24920 11138
rect 26082 11082 26084 11137
rect 26084 11082 26142 11137
rect 4289 10863 4323 10897
rect 7433 10863 7467 10897
rect 10565 10867 10599 10901
rect 13709 10867 13743 10901
rect 16911 10863 16945 10897
rect 20055 10863 20089 10897
rect 23187 10867 23221 10901
rect 26331 10867 26365 10901
rect 3802 10599 3836 10775
rect 3920 10599 3954 10775
rect 3994 10399 4028 10775
rect 4112 10399 4146 10775
rect 4230 10399 4264 10775
rect 4348 10399 4382 10775
rect 4466 10399 4500 10775
rect 4544 10599 4578 10775
rect 4662 10599 4696 10775
rect 6946 10599 6980 10775
rect 7064 10599 7098 10775
rect 7138 10399 7172 10775
rect 7256 10399 7290 10775
rect 7374 10399 7408 10775
rect 7492 10399 7526 10775
rect 7610 10399 7644 10775
rect 7688 10599 7722 10775
rect 7806 10599 7840 10775
rect 10078 10603 10112 10779
rect 10196 10603 10230 10779
rect 10270 10403 10304 10779
rect 10388 10403 10422 10779
rect 10506 10403 10540 10779
rect 10624 10403 10658 10779
rect 10742 10403 10776 10779
rect 10820 10603 10854 10779
rect 10938 10603 10972 10779
rect 13222 10603 13256 10779
rect 13340 10603 13374 10779
rect 13414 10403 13448 10779
rect 13532 10403 13566 10779
rect 13650 10403 13684 10779
rect 13768 10403 13802 10779
rect 13886 10403 13920 10779
rect 13964 10603 13998 10779
rect 14082 10603 14116 10779
rect 16424 10599 16458 10775
rect 16542 10599 16576 10775
rect 16616 10399 16650 10775
rect 16734 10399 16768 10775
rect 16852 10399 16886 10775
rect 16970 10399 17004 10775
rect 17088 10399 17122 10775
rect 17166 10599 17200 10775
rect 17284 10599 17318 10775
rect 19568 10599 19602 10775
rect 19686 10599 19720 10775
rect 19760 10399 19794 10775
rect 19878 10399 19912 10775
rect 19996 10399 20030 10775
rect 20114 10399 20148 10775
rect 20232 10399 20266 10775
rect 20310 10599 20344 10775
rect 20428 10599 20462 10775
rect 22700 10603 22734 10779
rect 22818 10603 22852 10779
rect 22892 10403 22926 10779
rect 23010 10403 23044 10779
rect 23128 10403 23162 10779
rect 23246 10403 23280 10779
rect 23364 10403 23398 10779
rect 23442 10603 23476 10779
rect 23560 10603 23594 10779
rect 25844 10603 25878 10779
rect 25962 10603 25996 10779
rect 26036 10403 26070 10779
rect 26154 10403 26188 10779
rect 26272 10403 26306 10779
rect 26390 10403 26424 10779
rect 26508 10403 26542 10779
rect 26586 10603 26620 10779
rect 26704 10603 26738 10779
rect 4231 10264 4265 10298
rect 7375 10264 7409 10298
rect 10507 10268 10541 10302
rect 13651 10268 13685 10302
rect 16853 10264 16887 10298
rect 19997 10264 20031 10298
rect 23129 10268 23163 10302
rect 26273 10268 26307 10302
rect 4234 10132 4292 10146
rect 4234 10100 4292 10132
rect 7378 10132 7436 10146
rect 7378 10100 7436 10132
rect 10510 10136 10568 10150
rect 10510 10104 10568 10136
rect 13654 10136 13712 10150
rect 13654 10104 13712 10136
rect 16856 10132 16914 10146
rect 16856 10100 16914 10132
rect 20000 10132 20058 10146
rect 20000 10100 20058 10132
rect 23132 10136 23190 10150
rect 23132 10104 23190 10136
rect 26276 10136 26334 10150
rect 26276 10104 26334 10136
rect 4210 9572 4282 9626
rect 7354 9572 7426 9626
rect 10486 9576 10558 9630
rect 13630 9576 13702 9630
rect 16832 9572 16904 9626
rect 19976 9572 20048 9626
rect 23108 9576 23180 9630
rect 26252 9576 26324 9630
rect 2958 9000 2992 9176
rect 3076 9000 3110 9176
rect 3194 9000 3228 9176
rect 3312 9000 3346 9176
rect 3399 9000 3433 9376
rect 3517 9000 3551 9376
rect 3635 9000 3669 9376
rect 3753 9000 3787 9376
rect 3866 9000 3900 9376
rect 3984 9000 4018 9376
rect 4102 9000 4136 9376
rect 4220 9000 4254 9376
rect 4338 9000 4372 9376
rect 4456 9000 4490 9376
rect 4574 9000 4608 9376
rect 4693 9000 4727 9376
rect 4811 9000 4845 9376
rect 4929 9000 4963 9376
rect 5047 9000 5081 9376
rect 5166 9000 5200 9176
rect 5284 9000 5318 9176
rect 5402 9000 5436 9176
rect 5520 9000 5554 9176
rect 6102 9000 6136 9176
rect 6220 9000 6254 9176
rect 6338 9000 6372 9176
rect 6456 9000 6490 9176
rect 6543 9000 6577 9376
rect 6661 9000 6695 9376
rect 6779 9000 6813 9376
rect 6897 9000 6931 9376
rect 7010 9000 7044 9376
rect 7128 9000 7162 9376
rect 7246 9000 7280 9376
rect 7364 9000 7398 9376
rect 7482 9000 7516 9376
rect 7600 9000 7634 9376
rect 7718 9000 7752 9376
rect 7837 9000 7871 9376
rect 7955 9000 7989 9376
rect 8073 9000 8107 9376
rect 8191 9000 8225 9376
rect 8310 9000 8344 9176
rect 8428 9000 8462 9176
rect 8546 9000 8580 9176
rect 8664 9000 8698 9176
rect 9234 9004 9268 9180
rect 9352 9004 9386 9180
rect 9470 9004 9504 9180
rect 9588 9004 9622 9180
rect 9675 9004 9709 9380
rect 9793 9004 9827 9380
rect 9911 9004 9945 9380
rect 10029 9004 10063 9380
rect 10142 9004 10176 9380
rect 10260 9004 10294 9380
rect 10378 9004 10412 9380
rect 10496 9004 10530 9380
rect 10614 9004 10648 9380
rect 10732 9004 10766 9380
rect 10850 9004 10884 9380
rect 10969 9004 11003 9380
rect 11087 9004 11121 9380
rect 11205 9004 11239 9380
rect 11323 9004 11357 9380
rect 11442 9004 11476 9180
rect 11560 9004 11594 9180
rect 11678 9004 11712 9180
rect 11796 9004 11830 9180
rect 12378 9004 12412 9180
rect 12496 9004 12530 9180
rect 12614 9004 12648 9180
rect 12732 9004 12766 9180
rect 12819 9004 12853 9380
rect 12937 9004 12971 9380
rect 13055 9004 13089 9380
rect 13173 9004 13207 9380
rect 13286 9004 13320 9380
rect 13404 9004 13438 9380
rect 13522 9004 13556 9380
rect 13640 9004 13674 9380
rect 13758 9004 13792 9380
rect 13876 9004 13910 9380
rect 13994 9004 14028 9380
rect 14113 9004 14147 9380
rect 14231 9004 14265 9380
rect 14349 9004 14383 9380
rect 14467 9004 14501 9380
rect 14586 9004 14620 9180
rect 14704 9004 14738 9180
rect 14822 9004 14856 9180
rect 14940 9004 14974 9180
rect 15580 9000 15614 9176
rect 15698 9000 15732 9176
rect 15816 9000 15850 9176
rect 15934 9000 15968 9176
rect 16021 9000 16055 9376
rect 16139 9000 16173 9376
rect 16257 9000 16291 9376
rect 16375 9000 16409 9376
rect 16488 9000 16522 9376
rect 16606 9000 16640 9376
rect 16724 9000 16758 9376
rect 16842 9000 16876 9376
rect 16960 9000 16994 9376
rect 17078 9000 17112 9376
rect 17196 9000 17230 9376
rect 17315 9000 17349 9376
rect 17433 9000 17467 9376
rect 17551 9000 17585 9376
rect 17669 9000 17703 9376
rect 17788 9000 17822 9176
rect 17906 9000 17940 9176
rect 18024 9000 18058 9176
rect 18142 9000 18176 9176
rect 18724 9000 18758 9176
rect 18842 9000 18876 9176
rect 18960 9000 18994 9176
rect 19078 9000 19112 9176
rect 19165 9000 19199 9376
rect 19283 9000 19317 9376
rect 19401 9000 19435 9376
rect 19519 9000 19553 9376
rect 19632 9000 19666 9376
rect 19750 9000 19784 9376
rect 19868 9000 19902 9376
rect 19986 9000 20020 9376
rect 20104 9000 20138 9376
rect 20222 9000 20256 9376
rect 20340 9000 20374 9376
rect 20459 9000 20493 9376
rect 20577 9000 20611 9376
rect 20695 9000 20729 9376
rect 20813 9000 20847 9376
rect 20932 9000 20966 9176
rect 21050 9000 21084 9176
rect 21168 9000 21202 9176
rect 21286 9000 21320 9176
rect 21856 9004 21890 9180
rect 21974 9004 22008 9180
rect 22092 9004 22126 9180
rect 22210 9004 22244 9180
rect 22297 9004 22331 9380
rect 22415 9004 22449 9380
rect 22533 9004 22567 9380
rect 22651 9004 22685 9380
rect 22764 9004 22798 9380
rect 22882 9004 22916 9380
rect 23000 9004 23034 9380
rect 23118 9004 23152 9380
rect 23236 9004 23270 9380
rect 23354 9004 23388 9380
rect 23472 9004 23506 9380
rect 23591 9004 23625 9380
rect 23709 9004 23743 9380
rect 23827 9004 23861 9380
rect 23945 9004 23979 9380
rect 24064 9004 24098 9180
rect 24182 9004 24216 9180
rect 24300 9004 24334 9180
rect 24418 9004 24452 9180
rect 25000 9004 25034 9180
rect 25118 9004 25152 9180
rect 25236 9004 25270 9180
rect 25354 9004 25388 9180
rect 25441 9004 25475 9380
rect 25559 9004 25593 9380
rect 25677 9004 25711 9380
rect 25795 9004 25829 9380
rect 25908 9004 25942 9380
rect 26026 9004 26060 9380
rect 26144 9004 26178 9380
rect 26262 9004 26296 9380
rect 26380 9004 26414 9380
rect 26498 9004 26532 9380
rect 26616 9004 26650 9380
rect 26735 9004 26769 9380
rect 26853 9004 26887 9380
rect 26971 9004 27005 9380
rect 27089 9004 27123 9380
rect 27208 9004 27242 9180
rect 27326 9004 27360 9180
rect 27444 9004 27478 9180
rect 27562 9004 27596 9180
rect 5354 8792 5388 8826
rect 4044 8751 4078 8785
rect 8498 8792 8532 8826
rect 7188 8751 7222 8785
rect 11630 8796 11664 8830
rect 10320 8755 10354 8789
rect 14774 8796 14808 8830
rect 13464 8755 13498 8789
rect 17976 8792 18010 8826
rect 16666 8751 16700 8785
rect 21120 8792 21154 8826
rect 19810 8751 19844 8785
rect 24252 8796 24286 8830
rect 22942 8755 22976 8789
rect 27396 8796 27430 8830
rect 26086 8755 26120 8789
rect 2819 8626 2868 8686
rect 3063 8630 3121 8685
rect 3121 8630 3123 8685
rect 4148 8631 4150 8686
rect 4150 8631 4208 8686
rect 5963 8626 6012 8686
rect 6207 8630 6265 8685
rect 6265 8630 6267 8685
rect 7292 8631 7294 8686
rect 7294 8631 7352 8686
rect 9095 8630 9144 8690
rect 9339 8634 9397 8689
rect 9397 8634 9399 8689
rect 10424 8635 10426 8690
rect 10426 8635 10484 8690
rect 12239 8630 12288 8690
rect 12483 8634 12541 8689
rect 12541 8634 12543 8689
rect 13568 8635 13570 8690
rect 13570 8635 13628 8690
rect 15441 8626 15490 8686
rect 15685 8630 15743 8685
rect 15743 8630 15745 8685
rect 16770 8631 16772 8686
rect 16772 8631 16830 8686
rect 18585 8626 18634 8686
rect 18829 8630 18887 8685
rect 18887 8630 18889 8685
rect 19914 8631 19916 8686
rect 19916 8631 19974 8686
rect 21717 8630 21766 8690
rect 21961 8634 22019 8689
rect 22019 8634 22021 8689
rect 23046 8635 23048 8690
rect 23048 8635 23106 8690
rect 24861 8630 24910 8690
rect 25105 8634 25163 8689
rect 25163 8634 25165 8689
rect 26190 8635 26192 8690
rect 26192 8635 26250 8690
rect 2819 8510 2868 8570
rect 4398 8521 4432 8555
rect 5963 8510 6012 8570
rect 2819 8342 2868 8402
rect 4030 8346 4032 8401
rect 4032 8346 4090 8401
rect 4279 8131 4313 8165
rect 3792 7867 3826 8043
rect 3910 7867 3944 8043
rect 3984 7667 4018 8043
rect 4102 7667 4136 8043
rect 4220 7667 4254 8043
rect 4338 7667 4372 8043
rect 4456 7667 4490 8043
rect 4534 7867 4568 8043
rect 4652 7867 4686 8043
rect 4221 7532 4255 7566
rect 4224 7400 4282 7414
rect 4224 7368 4282 7400
rect 3532 6658 3570 6686
rect 3532 6648 3570 6658
rect 2695 6055 2729 6231
rect 2813 6055 2847 6231
rect 2931 6055 2965 6231
rect 3049 6055 3083 6231
rect 3179 6055 3213 6431
rect 3297 6055 3331 6431
rect 3415 6055 3449 6431
rect 3533 6055 3567 6431
rect 3651 6055 3685 6431
rect 3769 6055 3803 6431
rect 3887 6055 3921 6431
rect 4016 6055 4050 6231
rect 4134 6055 4168 6231
rect 4252 6055 4286 6231
rect 4370 6055 4404 6231
rect 4102 5876 4156 5886
rect 4102 5842 4112 5876
rect 4112 5842 4146 5876
rect 4146 5842 4156 5876
rect 4102 5832 4156 5842
rect 2702 5682 2768 5696
rect 2702 5648 2718 5682
rect 2718 5648 2752 5682
rect 2752 5648 2768 5682
rect 2702 5636 2768 5648
rect 3122 5362 3156 5738
rect 3240 5362 3274 5738
rect 3358 5362 3392 5738
rect 3476 5362 3510 5738
rect 3594 5362 3628 5738
rect 3712 5362 3746 5738
rect 3830 5362 3864 5738
rect 3152 5140 3186 5174
rect 2967 5073 3001 5107
rect 4334 5232 4436 5334
rect 7542 8521 7576 8555
rect 9095 8514 9144 8574
rect 5963 8342 6012 8402
rect 7174 8346 7176 8401
rect 7176 8346 7234 8401
rect 7423 8131 7457 8165
rect 10674 8525 10708 8559
rect 12239 8514 12288 8574
rect 9095 8346 9144 8406
rect 10306 8350 10308 8405
rect 10308 8350 10366 8405
rect 10555 8135 10589 8169
rect 6936 7867 6970 8043
rect 7054 7867 7088 8043
rect 7128 7667 7162 8043
rect 7246 7667 7280 8043
rect 7364 7667 7398 8043
rect 7482 7667 7516 8043
rect 7600 7667 7634 8043
rect 7678 7867 7712 8043
rect 7796 7867 7830 8043
rect 7365 7532 7399 7566
rect 7368 7400 7426 7414
rect 7368 7368 7426 7400
rect 5600 6660 5638 6688
rect 5600 6650 5638 6660
rect 4763 6057 4797 6233
rect 4881 6057 4915 6233
rect 4999 6057 5033 6233
rect 5117 6057 5151 6233
rect 5247 6057 5281 6433
rect 5365 6057 5399 6433
rect 5483 6057 5517 6433
rect 5601 6057 5635 6433
rect 5719 6057 5753 6433
rect 5837 6057 5871 6433
rect 5955 6057 5989 6433
rect 6084 6057 6118 6233
rect 6202 6057 6236 6233
rect 6320 6057 6354 6233
rect 6438 6057 6472 6233
rect 6170 5878 6224 5888
rect 6170 5844 6180 5878
rect 6180 5844 6214 5878
rect 6214 5844 6224 5878
rect 6170 5834 6224 5844
rect 4770 5684 4836 5698
rect 4770 5650 4786 5684
rect 4786 5650 4820 5684
rect 4820 5650 4836 5684
rect 4770 5638 4836 5650
rect 5190 5364 5224 5740
rect 5308 5364 5342 5740
rect 5426 5364 5460 5740
rect 5544 5364 5578 5740
rect 5662 5364 5696 5740
rect 5780 5364 5814 5740
rect 5898 5364 5932 5740
rect 3800 5140 3834 5174
rect 5220 5142 5254 5176
rect 3418 5056 3452 5090
rect 3536 5057 3570 5091
rect 4090 5072 4124 5106
rect 5035 5075 5069 5109
rect 6402 5234 6504 5336
rect 7669 6658 7707 6686
rect 7669 6648 7707 6658
rect 6832 6055 6866 6231
rect 6950 6055 6984 6231
rect 7068 6055 7102 6231
rect 7186 6055 7220 6231
rect 7316 6055 7350 6431
rect 7434 6055 7468 6431
rect 7552 6055 7586 6431
rect 7670 6055 7704 6431
rect 7788 6055 7822 6431
rect 7906 6055 7940 6431
rect 8024 6055 8058 6431
rect 8153 6055 8187 6231
rect 8271 6055 8305 6231
rect 8389 6055 8423 6231
rect 8507 6055 8541 6231
rect 8239 5876 8293 5886
rect 8239 5842 8249 5876
rect 8249 5842 8283 5876
rect 8283 5842 8293 5876
rect 8239 5832 8293 5842
rect 6839 5682 6905 5696
rect 6839 5648 6855 5682
rect 6855 5648 6889 5682
rect 6889 5648 6905 5682
rect 6839 5636 6905 5648
rect 7259 5362 7293 5738
rect 7377 5362 7411 5738
rect 7495 5362 7529 5738
rect 7613 5362 7647 5738
rect 7731 5362 7765 5738
rect 7849 5362 7883 5738
rect 7967 5362 8001 5738
rect 5868 5142 5902 5176
rect 7289 5140 7323 5174
rect 5486 5058 5520 5092
rect 5604 5059 5638 5093
rect 6158 5074 6192 5108
rect 7104 5073 7138 5107
rect 2820 4830 2854 5006
rect 2938 4830 2972 5006
rect 3240 4630 3274 5006
rect 3358 4630 3392 5006
rect 3476 4630 3510 5006
rect 3594 4630 3628 5006
rect 3712 4630 3746 5006
rect 4118 4830 4152 5006
rect 4236 4830 4270 5006
rect 4888 4832 4922 5008
rect 5006 4832 5040 5008
rect 5308 4632 5342 5008
rect 5426 4632 5460 5008
rect 5544 4632 5578 5008
rect 5662 4632 5696 5008
rect 5780 4632 5814 5008
rect 6186 4832 6220 5008
rect 8471 5232 8573 5334
rect 10068 7871 10102 8047
rect 10186 7871 10220 8047
rect 10260 7671 10294 8047
rect 10378 7671 10412 8047
rect 10496 7671 10530 8047
rect 10614 7671 10648 8047
rect 10732 7671 10766 8047
rect 10810 7871 10844 8047
rect 10928 7871 10962 8047
rect 10497 7536 10531 7570
rect 10500 7404 10558 7418
rect 10500 7372 10558 7404
rect 13818 8525 13852 8559
rect 15441 8510 15490 8570
rect 17020 8521 17054 8555
rect 12239 8346 12288 8406
rect 13450 8350 13452 8405
rect 13452 8350 13510 8405
rect 13699 8135 13733 8169
rect 13212 7871 13246 8047
rect 13330 7871 13364 8047
rect 13404 7671 13438 8047
rect 13522 7671 13556 8047
rect 13640 7671 13674 8047
rect 13758 7671 13792 8047
rect 13876 7671 13910 8047
rect 13954 7871 13988 8047
rect 14072 7871 14106 8047
rect 13641 7536 13675 7570
rect 13644 7404 13702 7418
rect 13644 7372 13702 7404
rect 18585 8510 18634 8570
rect 15441 8342 15490 8402
rect 16652 8346 16654 8401
rect 16654 8346 16712 8401
rect 16901 8131 16935 8165
rect 16414 7867 16448 8043
rect 16532 7867 16566 8043
rect 16606 7667 16640 8043
rect 16724 7667 16758 8043
rect 16842 7667 16876 8043
rect 16960 7667 16994 8043
rect 17078 7667 17112 8043
rect 17156 7867 17190 8043
rect 17274 7867 17308 8043
rect 16843 7532 16877 7566
rect 16846 7400 16904 7414
rect 16846 7368 16904 7400
rect 9737 6660 9775 6688
rect 9737 6650 9775 6660
rect 8900 6057 8934 6233
rect 9018 6057 9052 6233
rect 9136 6057 9170 6233
rect 9254 6057 9288 6233
rect 9384 6057 9418 6433
rect 9502 6057 9536 6433
rect 9620 6057 9654 6433
rect 9738 6057 9772 6433
rect 9856 6057 9890 6433
rect 9974 6057 10008 6433
rect 10092 6057 10126 6433
rect 10221 6057 10255 6233
rect 10339 6057 10373 6233
rect 10457 6057 10491 6233
rect 10575 6057 10609 6233
rect 10307 5878 10361 5888
rect 10307 5844 10317 5878
rect 10317 5844 10351 5878
rect 10351 5844 10361 5878
rect 10307 5834 10361 5844
rect 8907 5684 8973 5698
rect 8907 5650 8923 5684
rect 8923 5650 8957 5684
rect 8957 5650 8973 5684
rect 8907 5638 8973 5650
rect 9327 5364 9361 5740
rect 9445 5364 9479 5740
rect 9563 5364 9597 5740
rect 9681 5364 9715 5740
rect 9799 5364 9833 5740
rect 9917 5364 9951 5740
rect 10035 5364 10069 5740
rect 7937 5140 7971 5174
rect 9357 5142 9391 5176
rect 7555 5056 7589 5090
rect 7673 5057 7707 5091
rect 8227 5072 8261 5106
rect 9172 5075 9206 5109
rect 10539 5234 10641 5336
rect 11806 6660 11844 6688
rect 11806 6650 11844 6660
rect 10969 6057 11003 6233
rect 11087 6057 11121 6233
rect 11205 6057 11239 6233
rect 11323 6057 11357 6233
rect 11453 6057 11487 6433
rect 11571 6057 11605 6433
rect 11689 6057 11723 6433
rect 11807 6057 11841 6433
rect 11925 6057 11959 6433
rect 12043 6057 12077 6433
rect 12161 6057 12195 6433
rect 12290 6057 12324 6233
rect 12408 6057 12442 6233
rect 12526 6057 12560 6233
rect 12644 6057 12678 6233
rect 12376 5878 12430 5888
rect 12376 5844 12386 5878
rect 12386 5844 12420 5878
rect 12420 5844 12430 5878
rect 12376 5834 12430 5844
rect 10976 5684 11042 5698
rect 10976 5650 10992 5684
rect 10992 5650 11026 5684
rect 11026 5650 11042 5684
rect 10976 5638 11042 5650
rect 11396 5364 11430 5740
rect 11514 5364 11548 5740
rect 11632 5364 11666 5740
rect 11750 5364 11784 5740
rect 11868 5364 11902 5740
rect 11986 5364 12020 5740
rect 12104 5364 12138 5740
rect 10005 5142 10039 5176
rect 11426 5142 11460 5176
rect 9623 5058 9657 5092
rect 9741 5059 9775 5093
rect 10295 5074 10329 5108
rect 11241 5075 11275 5109
rect 12608 5234 12710 5336
rect 20164 8521 20198 8555
rect 21717 8514 21766 8574
rect 18585 8342 18634 8402
rect 19796 8346 19798 8401
rect 19798 8346 19856 8401
rect 20045 8131 20079 8165
rect 19558 7867 19592 8043
rect 19676 7867 19710 8043
rect 19750 7667 19784 8043
rect 19868 7667 19902 8043
rect 19986 7667 20020 8043
rect 20104 7667 20138 8043
rect 20222 7667 20256 8043
rect 20300 7867 20334 8043
rect 20418 7867 20452 8043
rect 19987 7532 20021 7566
rect 19990 7400 20048 7414
rect 19990 7368 20048 7400
rect 13874 6662 13912 6690
rect 13874 6652 13912 6662
rect 13037 6059 13071 6235
rect 13155 6059 13189 6235
rect 13273 6059 13307 6235
rect 13391 6059 13425 6235
rect 13521 6059 13555 6435
rect 13639 6059 13673 6435
rect 13757 6059 13791 6435
rect 13875 6059 13909 6435
rect 13993 6059 14027 6435
rect 14111 6059 14145 6435
rect 14229 6059 14263 6435
rect 14358 6059 14392 6235
rect 14476 6059 14510 6235
rect 14594 6059 14628 6235
rect 14712 6059 14746 6235
rect 14444 5880 14498 5890
rect 14444 5846 14454 5880
rect 14454 5846 14488 5880
rect 14488 5846 14498 5880
rect 14444 5836 14498 5846
rect 13044 5686 13110 5700
rect 13044 5652 13060 5686
rect 13060 5652 13094 5686
rect 13094 5652 13110 5686
rect 13044 5640 13110 5652
rect 13464 5366 13498 5742
rect 13582 5366 13616 5742
rect 13700 5366 13734 5742
rect 13818 5366 13852 5742
rect 13936 5366 13970 5742
rect 14054 5366 14088 5742
rect 14172 5366 14206 5742
rect 12074 5142 12108 5176
rect 13494 5144 13528 5178
rect 11692 5058 11726 5092
rect 11810 5059 11844 5093
rect 12364 5074 12398 5108
rect 13309 5077 13343 5111
rect 14676 5236 14778 5338
rect 23296 8525 23330 8559
rect 24861 8514 24910 8574
rect 26440 8525 26474 8559
rect 21717 8346 21766 8406
rect 22928 8350 22930 8405
rect 22930 8350 22988 8405
rect 23177 8135 23211 8169
rect 22690 7871 22724 8047
rect 22808 7871 22842 8047
rect 22882 7671 22916 8047
rect 23000 7671 23034 8047
rect 23118 7671 23152 8047
rect 23236 7671 23270 8047
rect 23354 7671 23388 8047
rect 23432 7871 23466 8047
rect 23550 7871 23584 8047
rect 23119 7536 23153 7570
rect 23122 7404 23180 7418
rect 23122 7372 23180 7404
rect 15943 6660 15981 6688
rect 15943 6650 15981 6660
rect 15106 6057 15140 6233
rect 15224 6057 15258 6233
rect 15342 6057 15376 6233
rect 15460 6057 15494 6233
rect 15590 6057 15624 6433
rect 15708 6057 15742 6433
rect 15826 6057 15860 6433
rect 15944 6057 15978 6433
rect 16062 6057 16096 6433
rect 16180 6057 16214 6433
rect 16298 6057 16332 6433
rect 16427 6057 16461 6233
rect 16545 6057 16579 6233
rect 16663 6057 16697 6233
rect 16781 6057 16815 6233
rect 16513 5878 16567 5888
rect 16513 5844 16523 5878
rect 16523 5844 16557 5878
rect 16557 5844 16567 5878
rect 16513 5834 16567 5844
rect 15113 5684 15179 5698
rect 15113 5650 15129 5684
rect 15129 5650 15163 5684
rect 15163 5650 15179 5684
rect 15113 5638 15179 5650
rect 15533 5364 15567 5740
rect 15651 5364 15685 5740
rect 15769 5364 15803 5740
rect 15887 5364 15921 5740
rect 16005 5364 16039 5740
rect 16123 5364 16157 5740
rect 16241 5364 16275 5740
rect 14142 5144 14176 5178
rect 15563 5142 15597 5176
rect 13760 5060 13794 5094
rect 13878 5061 13912 5095
rect 14432 5076 14466 5110
rect 15378 5075 15412 5109
rect 6304 4832 6338 5008
rect 6957 4830 6991 5006
rect 7075 4830 7109 5006
rect 7377 4630 7411 5006
rect 7495 4630 7529 5006
rect 7613 4630 7647 5006
rect 7731 4630 7765 5006
rect 7849 4630 7883 5006
rect 8255 4830 8289 5006
rect 8373 4830 8407 5006
rect 9025 4832 9059 5008
rect 9143 4832 9177 5008
rect 9445 4632 9479 5008
rect 9563 4632 9597 5008
rect 9681 4632 9715 5008
rect 9799 4632 9833 5008
rect 9917 4632 9951 5008
rect 10323 4832 10357 5008
rect 10441 4832 10475 5008
rect 11094 4832 11128 5008
rect 11212 4832 11246 5008
rect 11514 4632 11548 5008
rect 11632 4632 11666 5008
rect 11750 4632 11784 5008
rect 11868 4632 11902 5008
rect 11986 4632 12020 5008
rect 12392 4832 12426 5008
rect 12510 4832 12544 5008
rect 13162 4834 13196 5010
rect 13280 4834 13314 5010
rect 13582 4634 13616 5010
rect 13700 4634 13734 5010
rect 13818 4634 13852 5010
rect 13936 4634 13970 5010
rect 14054 4634 14088 5010
rect 14460 4834 14494 5010
rect 16745 5234 16847 5336
rect 24861 8346 24910 8406
rect 26072 8350 26074 8405
rect 26074 8350 26132 8405
rect 26321 8135 26355 8169
rect 25834 7871 25868 8047
rect 25952 7871 25986 8047
rect 26026 7671 26060 8047
rect 26144 7671 26178 8047
rect 26262 7671 26296 8047
rect 26380 7671 26414 8047
rect 26498 7671 26532 8047
rect 26576 7871 26610 8047
rect 26694 7871 26728 8047
rect 26263 7536 26297 7570
rect 26266 7404 26324 7418
rect 26266 7372 26324 7404
rect 18011 6662 18049 6690
rect 18011 6652 18049 6662
rect 17174 6059 17208 6235
rect 17292 6059 17326 6235
rect 17410 6059 17444 6235
rect 17528 6059 17562 6235
rect 17658 6059 17692 6435
rect 17776 6059 17810 6435
rect 17894 6059 17928 6435
rect 18012 6059 18046 6435
rect 18130 6059 18164 6435
rect 18248 6059 18282 6435
rect 18366 6059 18400 6435
rect 18495 6059 18529 6235
rect 18613 6059 18647 6235
rect 18731 6059 18765 6235
rect 18849 6059 18883 6235
rect 18581 5880 18635 5890
rect 18581 5846 18591 5880
rect 18591 5846 18625 5880
rect 18625 5846 18635 5880
rect 18581 5836 18635 5846
rect 17181 5686 17247 5700
rect 17181 5652 17197 5686
rect 17197 5652 17231 5686
rect 17231 5652 17247 5686
rect 17181 5640 17247 5652
rect 17601 5366 17635 5742
rect 17719 5366 17753 5742
rect 17837 5366 17871 5742
rect 17955 5366 17989 5742
rect 18073 5366 18107 5742
rect 18191 5366 18225 5742
rect 18309 5366 18343 5742
rect 16211 5142 16245 5176
rect 17631 5144 17665 5178
rect 15829 5058 15863 5092
rect 15947 5059 15981 5093
rect 16501 5074 16535 5108
rect 17446 5077 17480 5111
rect 18813 5236 18915 5338
rect 19571 6697 19667 6733
rect 20309 6695 20405 6731
rect 21047 6695 21143 6731
rect 21789 6695 21885 6731
rect 22529 6695 22625 6731
rect 23267 6695 23363 6731
rect 24005 6695 24101 6731
rect 24743 6695 24839 6731
rect 19427 6371 19461 6547
rect 19545 6371 19579 6547
rect 19663 6371 19697 6547
rect 19781 6371 19815 6547
rect 20165 6375 20199 6551
rect 20283 6375 20317 6551
rect 20401 6375 20435 6551
rect 20519 6375 20553 6551
rect 20903 6371 20937 6547
rect 21021 6371 21055 6547
rect 21139 6371 21173 6547
rect 21257 6371 21291 6547
rect 21645 6369 21679 6545
rect 21763 6369 21797 6545
rect 21881 6369 21915 6545
rect 21999 6369 22033 6545
rect 22385 6369 22419 6545
rect 22503 6369 22537 6545
rect 22621 6369 22655 6545
rect 22739 6369 22773 6545
rect 23123 6369 23157 6545
rect 23241 6369 23275 6545
rect 23359 6369 23393 6545
rect 23477 6369 23511 6545
rect 23861 6369 23895 6545
rect 23979 6369 24013 6545
rect 24097 6369 24131 6545
rect 24215 6369 24249 6545
rect 24599 6369 24633 6545
rect 24717 6369 24751 6545
rect 24835 6369 24869 6545
rect 24953 6369 24987 6545
rect 19603 6231 19637 6265
rect 18279 5144 18313 5178
rect 17897 5060 17931 5094
rect 18015 5061 18049 5095
rect 18569 5076 18603 5110
rect 14578 4834 14612 5010
rect 15231 4832 15265 5008
rect 15349 4832 15383 5008
rect 15651 4632 15685 5008
rect 15769 4632 15803 5008
rect 15887 4632 15921 5008
rect 16005 4632 16039 5008
rect 16123 4632 16157 5008
rect 16529 4832 16563 5008
rect 16647 4832 16681 5008
rect 17299 4834 17333 5010
rect 17417 4834 17451 5010
rect 17719 4634 17753 5010
rect 17837 4634 17871 5010
rect 17955 4634 17989 5010
rect 18073 4634 18107 5010
rect 18191 4634 18225 5010
rect 18597 4834 18631 5010
rect 18715 4834 18749 5010
rect 3470 4442 3520 4464
rect 3470 4422 3520 4442
rect 5538 4444 5588 4466
rect 5538 4424 5588 4444
rect 7607 4442 7657 4464
rect 7607 4422 7657 4442
rect 9675 4444 9725 4466
rect 9675 4424 9725 4444
rect 11744 4444 11794 4466
rect 11744 4424 11794 4444
rect 13812 4446 13862 4468
rect 13812 4426 13862 4446
rect 15881 4444 15931 4466
rect 15881 4424 15931 4444
rect 17949 4446 17999 4468
rect 17949 4426 17999 4446
rect 20341 6229 20375 6263
rect 21079 6229 21113 6263
rect 21821 6229 21855 6263
rect 22561 6229 22595 6263
rect 23299 6229 23333 6263
rect 19545 5985 19579 6161
rect 19663 5985 19697 6161
rect 19521 5811 19599 5865
rect 20283 5987 20317 6163
rect 20401 5987 20435 6163
rect 20259 5809 20337 5863
rect 4715 4004 4766 4055
rect 6750 3896 6797 3950
rect 21021 5983 21055 6159
rect 21139 5983 21173 6159
rect 20997 5809 21075 5863
rect 21763 5983 21797 6159
rect 21881 5983 21915 6159
rect 21739 5809 21817 5863
rect 8797 3793 8844 3847
rect 22503 5983 22537 6159
rect 22621 5983 22655 6159
rect 22479 5809 22557 5863
rect 10887 3686 10937 3737
rect 23854 6223 23890 6269
rect 24037 6229 24071 6263
rect 24591 6223 24629 6269
rect 24775 6229 24809 6263
rect 23241 5983 23275 6159
rect 23359 5983 23393 6159
rect 23217 5809 23295 5863
rect 12958 3589 13009 3642
rect 23979 5987 24013 6163
rect 24097 5987 24131 6163
rect 23955 5809 24033 5863
rect 24717 5987 24751 6163
rect 24835 5987 24869 6163
rect 24693 5809 24771 5863
rect 15061 3447 15105 3498
rect 17129 3349 17182 3403
rect 1512 2324 1584 2378
rect 4656 2324 4728 2378
rect 7788 2328 7860 2382
rect 10932 2328 11004 2382
rect 14134 2324 14206 2378
rect 17278 2324 17350 2378
rect 20410 2328 20482 2382
rect 23554 2328 23626 2382
rect 260 1752 294 1928
rect 378 1752 412 1928
rect 496 1752 530 1928
rect 614 1752 648 1928
rect 701 1752 735 2128
rect 819 1752 853 2128
rect 937 1752 971 2128
rect 1055 1752 1089 2128
rect 1168 1752 1202 2128
rect 1286 1752 1320 2128
rect 1404 1752 1438 2128
rect 1522 1752 1556 2128
rect 1640 1752 1674 2128
rect 1758 1752 1792 2128
rect 1876 1752 1910 2128
rect 1995 1752 2029 2128
rect 2113 1752 2147 2128
rect 2231 1752 2265 2128
rect 2349 1752 2383 2128
rect 2468 1752 2502 1928
rect 2586 1752 2620 1928
rect 2704 1752 2738 1928
rect 2822 1752 2856 1928
rect 3404 1752 3438 1928
rect 3522 1752 3556 1928
rect 3640 1752 3674 1928
rect 3758 1752 3792 1928
rect 3845 1752 3879 2128
rect 3963 1752 3997 2128
rect 4081 1752 4115 2128
rect 4199 1752 4233 2128
rect 4312 1752 4346 2128
rect 4430 1752 4464 2128
rect 4548 1752 4582 2128
rect 4666 1752 4700 2128
rect 4784 1752 4818 2128
rect 4902 1752 4936 2128
rect 5020 1752 5054 2128
rect 5139 1752 5173 2128
rect 5257 1752 5291 2128
rect 5375 1752 5409 2128
rect 5493 1752 5527 2128
rect 5612 1752 5646 1928
rect 5730 1752 5764 1928
rect 5848 1752 5882 1928
rect 5966 1752 6000 1928
rect 6536 1756 6570 1932
rect 6654 1756 6688 1932
rect 6772 1756 6806 1932
rect 6890 1756 6924 1932
rect 6977 1756 7011 2132
rect 7095 1756 7129 2132
rect 7213 1756 7247 2132
rect 7331 1756 7365 2132
rect 7444 1756 7478 2132
rect 7562 1756 7596 2132
rect 7680 1756 7714 2132
rect 7798 1756 7832 2132
rect 7916 1756 7950 2132
rect 8034 1756 8068 2132
rect 8152 1756 8186 2132
rect 8271 1756 8305 2132
rect 8389 1756 8423 2132
rect 8507 1756 8541 2132
rect 8625 1756 8659 2132
rect 8744 1756 8778 1932
rect 8862 1756 8896 1932
rect 8980 1756 9014 1932
rect 9098 1756 9132 1932
rect 9680 1756 9714 1932
rect 9798 1756 9832 1932
rect 9916 1756 9950 1932
rect 10034 1756 10068 1932
rect 10121 1756 10155 2132
rect 10239 1756 10273 2132
rect 10357 1756 10391 2132
rect 10475 1756 10509 2132
rect 10588 1756 10622 2132
rect 10706 1756 10740 2132
rect 10824 1756 10858 2132
rect 10942 1756 10976 2132
rect 11060 1756 11094 2132
rect 11178 1756 11212 2132
rect 11296 1756 11330 2132
rect 11415 1756 11449 2132
rect 11533 1756 11567 2132
rect 11651 1756 11685 2132
rect 11769 1756 11803 2132
rect 11888 1756 11922 1932
rect 12006 1756 12040 1932
rect 12124 1756 12158 1932
rect 12242 1756 12276 1932
rect 12882 1752 12916 1928
rect 13000 1752 13034 1928
rect 13118 1752 13152 1928
rect 13236 1752 13270 1928
rect 13323 1752 13357 2128
rect 13441 1752 13475 2128
rect 13559 1752 13593 2128
rect 13677 1752 13711 2128
rect 13790 1752 13824 2128
rect 13908 1752 13942 2128
rect 14026 1752 14060 2128
rect 14144 1752 14178 2128
rect 14262 1752 14296 2128
rect 14380 1752 14414 2128
rect 14498 1752 14532 2128
rect 14617 1752 14651 2128
rect 14735 1752 14769 2128
rect 14853 1752 14887 2128
rect 14971 1752 15005 2128
rect 15090 1752 15124 1928
rect 15208 1752 15242 1928
rect 15326 1752 15360 1928
rect 15444 1752 15478 1928
rect 16026 1752 16060 1928
rect 16144 1752 16178 1928
rect 16262 1752 16296 1928
rect 16380 1752 16414 1928
rect 16467 1752 16501 2128
rect 16585 1752 16619 2128
rect 16703 1752 16737 2128
rect 16821 1752 16855 2128
rect 16934 1752 16968 2128
rect 17052 1752 17086 2128
rect 17170 1752 17204 2128
rect 17288 1752 17322 2128
rect 17406 1752 17440 2128
rect 17524 1752 17558 2128
rect 17642 1752 17676 2128
rect 17761 1752 17795 2128
rect 17879 1752 17913 2128
rect 17997 1752 18031 2128
rect 18115 1752 18149 2128
rect 18234 1752 18268 1928
rect 18352 1752 18386 1928
rect 18470 1752 18504 1928
rect 18588 1752 18622 1928
rect 19158 1756 19192 1932
rect 19276 1756 19310 1932
rect 19394 1756 19428 1932
rect 19512 1756 19546 1932
rect 19599 1756 19633 2132
rect 19717 1756 19751 2132
rect 19835 1756 19869 2132
rect 19953 1756 19987 2132
rect 20066 1756 20100 2132
rect 20184 1756 20218 2132
rect 20302 1756 20336 2132
rect 20420 1756 20454 2132
rect 20538 1756 20572 2132
rect 20656 1756 20690 2132
rect 20774 1756 20808 2132
rect 20893 1756 20927 2132
rect 21011 1756 21045 2132
rect 21129 1756 21163 2132
rect 21247 1756 21281 2132
rect 21366 1756 21400 1932
rect 21484 1756 21518 1932
rect 21602 1756 21636 1932
rect 21720 1756 21754 1932
rect 22302 1756 22336 1932
rect 22420 1756 22454 1932
rect 22538 1756 22572 1932
rect 22656 1756 22690 1932
rect 22743 1756 22777 2132
rect 22861 1756 22895 2132
rect 22979 1756 23013 2132
rect 23097 1756 23131 2132
rect 23210 1756 23244 2132
rect 23328 1756 23362 2132
rect 23446 1756 23480 2132
rect 23564 1756 23598 2132
rect 23682 1756 23716 2132
rect 23800 1756 23834 2132
rect 23918 1756 23952 2132
rect 24037 1756 24071 2132
rect 24155 1756 24189 2132
rect 24273 1756 24307 2132
rect 24391 1756 24425 2132
rect 24510 1756 24544 1932
rect 24628 1756 24662 1932
rect 24746 1756 24780 1932
rect 24864 1756 24898 1932
rect 2656 1544 2690 1578
rect 1346 1503 1380 1537
rect 5800 1544 5834 1578
rect 4490 1503 4524 1537
rect 8932 1548 8966 1582
rect 7622 1507 7656 1541
rect 12076 1548 12110 1582
rect 10766 1507 10800 1541
rect 15278 1544 15312 1578
rect 13968 1503 14002 1537
rect 18422 1544 18456 1578
rect 17112 1503 17146 1537
rect 21554 1548 21588 1582
rect 20244 1507 20278 1541
rect 24698 1548 24732 1582
rect 23388 1507 23422 1541
rect 121 1378 170 1438
rect 365 1382 423 1437
rect 423 1382 425 1437
rect 1450 1383 1452 1438
rect 1452 1383 1510 1438
rect 3265 1378 3314 1438
rect 3509 1382 3567 1437
rect 3567 1382 3569 1437
rect 4594 1383 4596 1438
rect 4596 1383 4654 1438
rect 6397 1382 6446 1442
rect 6641 1386 6699 1441
rect 6699 1386 6701 1441
rect 7726 1387 7728 1442
rect 7728 1387 7786 1442
rect 9541 1382 9590 1442
rect 9785 1386 9843 1441
rect 9843 1386 9845 1441
rect 10870 1387 10872 1442
rect 10872 1387 10930 1442
rect 12743 1378 12792 1438
rect 12987 1382 13045 1437
rect 13045 1382 13047 1437
rect 14072 1383 14074 1438
rect 14074 1383 14132 1438
rect 15887 1378 15936 1438
rect 16131 1382 16189 1437
rect 16189 1382 16191 1437
rect 17216 1383 17218 1438
rect 17218 1383 17276 1438
rect 19019 1382 19068 1442
rect 19263 1386 19321 1441
rect 19321 1386 19323 1441
rect 20348 1387 20350 1442
rect 20350 1387 20408 1442
rect 22163 1382 22212 1442
rect 22407 1386 22465 1441
rect 22465 1386 22467 1441
rect 23492 1387 23494 1442
rect 23494 1387 23552 1442
rect 121 1262 170 1322
rect 1700 1273 1734 1307
rect 3265 1262 3314 1322
rect 4844 1273 4878 1307
rect 6397 1266 6446 1326
rect 7976 1277 8010 1311
rect 9541 1266 9590 1326
rect 11120 1277 11154 1311
rect 12743 1262 12792 1322
rect 14322 1273 14356 1307
rect 15887 1262 15936 1322
rect 17466 1273 17500 1307
rect 19019 1266 19068 1326
rect 20598 1277 20632 1311
rect 22163 1266 22212 1326
rect 23742 1277 23776 1311
rect 121 1094 170 1154
rect 1332 1098 1334 1153
rect 1334 1098 1392 1153
rect 3265 1094 3314 1154
rect 4476 1098 4478 1153
rect 4478 1098 4536 1153
rect 6397 1098 6446 1158
rect 7608 1102 7610 1157
rect 7610 1102 7668 1157
rect 9541 1098 9590 1158
rect 10752 1102 10754 1157
rect 10754 1102 10812 1157
rect 12743 1094 12792 1154
rect 13954 1098 13956 1153
rect 13956 1098 14014 1153
rect 15887 1094 15936 1154
rect 17098 1098 17100 1153
rect 17100 1098 17158 1153
rect 19019 1098 19068 1158
rect 20230 1102 20232 1157
rect 20232 1102 20290 1157
rect 22163 1098 22212 1158
rect 23374 1102 23376 1157
rect 23376 1102 23434 1157
rect 1581 883 1615 917
rect 4725 883 4759 917
rect 7857 887 7891 921
rect 11001 887 11035 921
rect 14203 883 14237 917
rect 17347 883 17381 917
rect 20479 887 20513 921
rect 23623 887 23657 921
rect 1094 619 1128 795
rect 1212 619 1246 795
rect 1286 419 1320 795
rect 1404 419 1438 795
rect 1522 419 1556 795
rect 1640 419 1674 795
rect 1758 419 1792 795
rect 1836 619 1870 795
rect 1954 619 1988 795
rect 4238 619 4272 795
rect 4356 619 4390 795
rect 4430 419 4464 795
rect 4548 419 4582 795
rect 4666 419 4700 795
rect 4784 419 4818 795
rect 4902 419 4936 795
rect 4980 619 5014 795
rect 5098 619 5132 795
rect 7370 623 7404 799
rect 7488 623 7522 799
rect 7562 423 7596 799
rect 7680 423 7714 799
rect 7798 423 7832 799
rect 7916 423 7950 799
rect 8034 423 8068 799
rect 8112 623 8146 799
rect 8230 623 8264 799
rect 10514 623 10548 799
rect 10632 623 10666 799
rect 10706 423 10740 799
rect 10824 423 10858 799
rect 10942 423 10976 799
rect 11060 423 11094 799
rect 11178 423 11212 799
rect 11256 623 11290 799
rect 11374 623 11408 799
rect 13716 619 13750 795
rect 13834 619 13868 795
rect 13908 419 13942 795
rect 14026 419 14060 795
rect 14144 419 14178 795
rect 14262 419 14296 795
rect 14380 419 14414 795
rect 14458 619 14492 795
rect 14576 619 14610 795
rect 16860 619 16894 795
rect 16978 619 17012 795
rect 17052 419 17086 795
rect 17170 419 17204 795
rect 17288 419 17322 795
rect 17406 419 17440 795
rect 17524 419 17558 795
rect 17602 619 17636 795
rect 17720 619 17754 795
rect 19992 623 20026 799
rect 20110 623 20144 799
rect 20184 423 20218 799
rect 20302 423 20336 799
rect 20420 423 20454 799
rect 20538 423 20572 799
rect 20656 423 20690 799
rect 20734 623 20768 799
rect 20852 623 20886 799
rect 23136 623 23170 799
rect 23254 623 23288 799
rect 23328 423 23362 799
rect 23446 423 23480 799
rect 23564 423 23598 799
rect 23682 423 23716 799
rect 23800 423 23834 799
rect 23878 623 23912 799
rect 23996 623 24030 799
rect 1523 284 1557 318
rect 4667 284 4701 318
rect 7799 288 7833 322
rect 10943 288 10977 322
rect 14145 284 14179 318
rect 17289 284 17323 318
rect 20421 288 20455 322
rect 23565 288 23599 322
rect 1526 152 1584 166
rect 1526 120 1584 152
rect 4670 152 4728 166
rect 4670 120 4728 152
rect 7802 156 7860 170
rect 7802 124 7860 156
rect 10946 156 11004 170
rect 10946 124 11004 156
rect 14148 152 14206 166
rect 14148 120 14206 152
rect 17292 152 17350 166
rect 17292 120 17350 152
rect 20424 156 20482 170
rect 20424 124 20482 156
rect 23568 156 23626 170
rect 23568 124 23626 156
rect 1544 -1568 1616 -1514
rect 4688 -1568 4760 -1514
rect 7820 -1564 7892 -1510
rect 10964 -1564 11036 -1510
rect 14166 -1568 14238 -1514
rect 17310 -1568 17382 -1514
rect 20442 -1564 20514 -1510
rect 23586 -1564 23658 -1510
rect 292 -2140 326 -1964
rect 410 -2140 444 -1964
rect 528 -2140 562 -1964
rect 646 -2140 680 -1964
rect 733 -2140 767 -1764
rect 851 -2140 885 -1764
rect 969 -2140 1003 -1764
rect 1087 -2140 1121 -1764
rect 1200 -2140 1234 -1764
rect 1318 -2140 1352 -1764
rect 1436 -2140 1470 -1764
rect 1554 -2140 1588 -1764
rect 1672 -2140 1706 -1764
rect 1790 -2140 1824 -1764
rect 1908 -2140 1942 -1764
rect 2027 -2140 2061 -1764
rect 2145 -2140 2179 -1764
rect 2263 -2140 2297 -1764
rect 2381 -2140 2415 -1764
rect 2500 -2140 2534 -1964
rect 2618 -2140 2652 -1964
rect 2736 -2140 2770 -1964
rect 2854 -2140 2888 -1964
rect 3436 -2140 3470 -1964
rect 3554 -2140 3588 -1964
rect 3672 -2140 3706 -1964
rect 3790 -2140 3824 -1964
rect 3877 -2140 3911 -1764
rect 3995 -2140 4029 -1764
rect 4113 -2140 4147 -1764
rect 4231 -2140 4265 -1764
rect 4344 -2140 4378 -1764
rect 4462 -2140 4496 -1764
rect 4580 -2140 4614 -1764
rect 4698 -2140 4732 -1764
rect 4816 -2140 4850 -1764
rect 4934 -2140 4968 -1764
rect 5052 -2140 5086 -1764
rect 5171 -2140 5205 -1764
rect 5289 -2140 5323 -1764
rect 5407 -2140 5441 -1764
rect 5525 -2140 5559 -1764
rect 5644 -2140 5678 -1964
rect 5762 -2140 5796 -1964
rect 5880 -2140 5914 -1964
rect 5998 -2140 6032 -1964
rect 6568 -2136 6602 -1960
rect 6686 -2136 6720 -1960
rect 6804 -2136 6838 -1960
rect 6922 -2136 6956 -1960
rect 7009 -2136 7043 -1760
rect 7127 -2136 7161 -1760
rect 7245 -2136 7279 -1760
rect 7363 -2136 7397 -1760
rect 7476 -2136 7510 -1760
rect 7594 -2136 7628 -1760
rect 7712 -2136 7746 -1760
rect 7830 -2136 7864 -1760
rect 7948 -2136 7982 -1760
rect 8066 -2136 8100 -1760
rect 8184 -2136 8218 -1760
rect 8303 -2136 8337 -1760
rect 8421 -2136 8455 -1760
rect 8539 -2136 8573 -1760
rect 8657 -2136 8691 -1760
rect 8776 -2136 8810 -1960
rect 8894 -2136 8928 -1960
rect 9012 -2136 9046 -1960
rect 9130 -2136 9164 -1960
rect 9712 -2136 9746 -1960
rect 9830 -2136 9864 -1960
rect 9948 -2136 9982 -1960
rect 10066 -2136 10100 -1960
rect 10153 -2136 10187 -1760
rect 10271 -2136 10305 -1760
rect 10389 -2136 10423 -1760
rect 10507 -2136 10541 -1760
rect 10620 -2136 10654 -1760
rect 10738 -2136 10772 -1760
rect 10856 -2136 10890 -1760
rect 10974 -2136 11008 -1760
rect 11092 -2136 11126 -1760
rect 11210 -2136 11244 -1760
rect 11328 -2136 11362 -1760
rect 11447 -2136 11481 -1760
rect 11565 -2136 11599 -1760
rect 11683 -2136 11717 -1760
rect 11801 -2136 11835 -1760
rect 11920 -2136 11954 -1960
rect 12038 -2136 12072 -1960
rect 12156 -2136 12190 -1960
rect 12274 -2136 12308 -1960
rect 12914 -2140 12948 -1964
rect 13032 -2140 13066 -1964
rect 13150 -2140 13184 -1964
rect 13268 -2140 13302 -1964
rect 13355 -2140 13389 -1764
rect 13473 -2140 13507 -1764
rect 13591 -2140 13625 -1764
rect 13709 -2140 13743 -1764
rect 13822 -2140 13856 -1764
rect 13940 -2140 13974 -1764
rect 14058 -2140 14092 -1764
rect 14176 -2140 14210 -1764
rect 14294 -2140 14328 -1764
rect 14412 -2140 14446 -1764
rect 14530 -2140 14564 -1764
rect 14649 -2140 14683 -1764
rect 14767 -2140 14801 -1764
rect 14885 -2140 14919 -1764
rect 15003 -2140 15037 -1764
rect 15122 -2140 15156 -1964
rect 15240 -2140 15274 -1964
rect 15358 -2140 15392 -1964
rect 15476 -2140 15510 -1964
rect 16058 -2140 16092 -1964
rect 16176 -2140 16210 -1964
rect 16294 -2140 16328 -1964
rect 16412 -2140 16446 -1964
rect 16499 -2140 16533 -1764
rect 16617 -2140 16651 -1764
rect 16735 -2140 16769 -1764
rect 16853 -2140 16887 -1764
rect 16966 -2140 17000 -1764
rect 17084 -2140 17118 -1764
rect 17202 -2140 17236 -1764
rect 17320 -2140 17354 -1764
rect 17438 -2140 17472 -1764
rect 17556 -2140 17590 -1764
rect 17674 -2140 17708 -1764
rect 17793 -2140 17827 -1764
rect 17911 -2140 17945 -1764
rect 18029 -2140 18063 -1764
rect 18147 -2140 18181 -1764
rect 18266 -2140 18300 -1964
rect 18384 -2140 18418 -1964
rect 18502 -2140 18536 -1964
rect 18620 -2140 18654 -1964
rect 19190 -2136 19224 -1960
rect 19308 -2136 19342 -1960
rect 19426 -2136 19460 -1960
rect 19544 -2136 19578 -1960
rect 19631 -2136 19665 -1760
rect 19749 -2136 19783 -1760
rect 19867 -2136 19901 -1760
rect 19985 -2136 20019 -1760
rect 20098 -2136 20132 -1760
rect 20216 -2136 20250 -1760
rect 20334 -2136 20368 -1760
rect 20452 -2136 20486 -1760
rect 20570 -2136 20604 -1760
rect 20688 -2136 20722 -1760
rect 20806 -2136 20840 -1760
rect 20925 -2136 20959 -1760
rect 21043 -2136 21077 -1760
rect 21161 -2136 21195 -1760
rect 21279 -2136 21313 -1760
rect 21398 -2136 21432 -1960
rect 21516 -2136 21550 -1960
rect 21634 -2136 21668 -1960
rect 21752 -2136 21786 -1960
rect 22334 -2136 22368 -1960
rect 22452 -2136 22486 -1960
rect 22570 -2136 22604 -1960
rect 22688 -2136 22722 -1960
rect 22775 -2136 22809 -1760
rect 22893 -2136 22927 -1760
rect 23011 -2136 23045 -1760
rect 23129 -2136 23163 -1760
rect 23242 -2136 23276 -1760
rect 23360 -2136 23394 -1760
rect 23478 -2136 23512 -1760
rect 23596 -2136 23630 -1760
rect 23714 -2136 23748 -1760
rect 23832 -2136 23866 -1760
rect 23950 -2136 23984 -1760
rect 24069 -2136 24103 -1760
rect 24187 -2136 24221 -1760
rect 24305 -2136 24339 -1760
rect 24423 -2136 24457 -1760
rect 24542 -2136 24576 -1960
rect 24660 -2136 24694 -1960
rect 24778 -2136 24812 -1960
rect 24896 -2136 24930 -1960
rect 2688 -2348 2722 -2314
rect 1378 -2389 1412 -2355
rect 5832 -2348 5866 -2314
rect 4522 -2389 4556 -2355
rect 8964 -2344 8998 -2310
rect 7654 -2385 7688 -2351
rect 12108 -2344 12142 -2310
rect 10798 -2385 10832 -2351
rect 15310 -2348 15344 -2314
rect 14000 -2389 14034 -2355
rect 18454 -2348 18488 -2314
rect 17144 -2389 17178 -2355
rect 21586 -2344 21620 -2310
rect 20276 -2385 20310 -2351
rect 24730 -2344 24764 -2310
rect 23420 -2385 23454 -2351
rect 153 -2514 202 -2454
rect 397 -2510 455 -2455
rect 455 -2510 457 -2455
rect 1482 -2509 1484 -2454
rect 1484 -2509 1542 -2454
rect 3297 -2514 3346 -2454
rect 3541 -2510 3599 -2455
rect 3599 -2510 3601 -2455
rect 4626 -2509 4628 -2454
rect 4628 -2509 4686 -2454
rect 6429 -2510 6478 -2450
rect 6673 -2506 6731 -2451
rect 6731 -2506 6733 -2451
rect 7758 -2505 7760 -2450
rect 7760 -2505 7818 -2450
rect 9573 -2510 9622 -2450
rect 9817 -2506 9875 -2451
rect 9875 -2506 9877 -2451
rect 10902 -2505 10904 -2450
rect 10904 -2505 10962 -2450
rect 12775 -2514 12824 -2454
rect 13019 -2510 13077 -2455
rect 13077 -2510 13079 -2455
rect 14104 -2509 14106 -2454
rect 14106 -2509 14164 -2454
rect 15919 -2514 15968 -2454
rect 16163 -2510 16221 -2455
rect 16221 -2510 16223 -2455
rect 17248 -2509 17250 -2454
rect 17250 -2509 17308 -2454
rect 19051 -2510 19100 -2450
rect 19295 -2506 19353 -2451
rect 19353 -2506 19355 -2451
rect 20380 -2505 20382 -2450
rect 20382 -2505 20440 -2450
rect 22195 -2510 22244 -2450
rect 22439 -2506 22497 -2451
rect 22497 -2506 22499 -2451
rect 23524 -2505 23526 -2450
rect 23526 -2505 23584 -2450
rect 153 -2630 202 -2570
rect 1732 -2619 1766 -2585
rect 3297 -2630 3346 -2570
rect 4876 -2619 4910 -2585
rect 6429 -2626 6478 -2566
rect 8008 -2615 8042 -2581
rect 9573 -2626 9622 -2566
rect 11152 -2615 11186 -2581
rect 12775 -2630 12824 -2570
rect 14354 -2619 14388 -2585
rect 15919 -2630 15968 -2570
rect 17498 -2619 17532 -2585
rect 19051 -2626 19100 -2566
rect 20630 -2615 20664 -2581
rect 22195 -2626 22244 -2566
rect 23774 -2615 23808 -2581
rect 153 -2798 202 -2738
rect 1364 -2794 1366 -2739
rect 1366 -2794 1424 -2739
rect 3297 -2798 3346 -2738
rect 4508 -2794 4510 -2739
rect 4510 -2794 4568 -2739
rect 6429 -2794 6478 -2734
rect 7640 -2790 7642 -2735
rect 7642 -2790 7700 -2735
rect 9573 -2794 9622 -2734
rect 10784 -2790 10786 -2735
rect 10786 -2790 10844 -2735
rect 12775 -2798 12824 -2738
rect 13986 -2794 13988 -2739
rect 13988 -2794 14046 -2739
rect 15919 -2798 15968 -2738
rect 17130 -2794 17132 -2739
rect 17132 -2794 17190 -2739
rect 19051 -2794 19100 -2734
rect 20262 -2790 20264 -2735
rect 20264 -2790 20322 -2735
rect 22195 -2794 22244 -2734
rect 23406 -2790 23408 -2735
rect 23408 -2790 23466 -2735
rect 1613 -3009 1647 -2975
rect 4757 -3009 4791 -2975
rect 7889 -3005 7923 -2971
rect 11033 -3005 11067 -2971
rect 14235 -3009 14269 -2975
rect 17379 -3009 17413 -2975
rect 20511 -3005 20545 -2971
rect 23655 -3005 23689 -2971
rect 1126 -3273 1160 -3097
rect 1244 -3273 1278 -3097
rect 1318 -3473 1352 -3097
rect 1436 -3473 1470 -3097
rect 1554 -3473 1588 -3097
rect 1672 -3473 1706 -3097
rect 1790 -3473 1824 -3097
rect 1868 -3273 1902 -3097
rect 1986 -3273 2020 -3097
rect 4270 -3273 4304 -3097
rect 4388 -3273 4422 -3097
rect 4462 -3473 4496 -3097
rect 4580 -3473 4614 -3097
rect 4698 -3473 4732 -3097
rect 4816 -3473 4850 -3097
rect 4934 -3473 4968 -3097
rect 5012 -3273 5046 -3097
rect 5130 -3273 5164 -3097
rect 7402 -3269 7436 -3093
rect 7520 -3269 7554 -3093
rect 7594 -3469 7628 -3093
rect 7712 -3469 7746 -3093
rect 7830 -3469 7864 -3093
rect 7948 -3469 7982 -3093
rect 8066 -3469 8100 -3093
rect 8144 -3269 8178 -3093
rect 8262 -3269 8296 -3093
rect 10546 -3269 10580 -3093
rect 10664 -3269 10698 -3093
rect 10738 -3469 10772 -3093
rect 10856 -3469 10890 -3093
rect 10974 -3469 11008 -3093
rect 11092 -3469 11126 -3093
rect 11210 -3469 11244 -3093
rect 11288 -3269 11322 -3093
rect 11406 -3269 11440 -3093
rect 13748 -3273 13782 -3097
rect 13866 -3273 13900 -3097
rect 13940 -3473 13974 -3097
rect 14058 -3473 14092 -3097
rect 14176 -3473 14210 -3097
rect 14294 -3473 14328 -3097
rect 14412 -3473 14446 -3097
rect 14490 -3273 14524 -3097
rect 14608 -3273 14642 -3097
rect 16892 -3273 16926 -3097
rect 17010 -3273 17044 -3097
rect 17084 -3473 17118 -3097
rect 17202 -3473 17236 -3097
rect 17320 -3473 17354 -3097
rect 17438 -3473 17472 -3097
rect 17556 -3473 17590 -3097
rect 17634 -3273 17668 -3097
rect 17752 -3273 17786 -3097
rect 20024 -3269 20058 -3093
rect 20142 -3269 20176 -3093
rect 20216 -3469 20250 -3093
rect 20334 -3469 20368 -3093
rect 20452 -3469 20486 -3093
rect 20570 -3469 20604 -3093
rect 20688 -3469 20722 -3093
rect 20766 -3269 20800 -3093
rect 20884 -3269 20918 -3093
rect 23168 -3269 23202 -3093
rect 23286 -3269 23320 -3093
rect 23360 -3469 23394 -3093
rect 23478 -3469 23512 -3093
rect 23596 -3469 23630 -3093
rect 23714 -3469 23748 -3093
rect 23832 -3469 23866 -3093
rect 23910 -3269 23944 -3093
rect 24028 -3269 24062 -3093
rect 1555 -3608 1589 -3574
rect 4699 -3608 4733 -3574
rect 7831 -3604 7865 -3570
rect 10975 -3604 11009 -3570
rect 14177 -3608 14211 -3574
rect 17321 -3608 17355 -3574
rect 20453 -3604 20487 -3570
rect 23597 -3604 23631 -3570
rect 1558 -3740 1616 -3726
rect 1558 -3772 1616 -3740
rect 4702 -3740 4760 -3726
rect 4702 -3772 4760 -3740
rect 7834 -3736 7892 -3722
rect 7834 -3768 7892 -3736
rect 10978 -3736 11036 -3722
rect 10978 -3768 11036 -3736
rect 14180 -3740 14238 -3726
rect 14180 -3772 14238 -3740
rect 17324 -3740 17382 -3726
rect 17324 -3772 17382 -3740
rect 20456 -3736 20514 -3722
rect 20456 -3768 20514 -3736
rect 23600 -3736 23658 -3722
rect 23600 -3768 23658 -3736
<< metal1 >>
rect 1704 22176 1714 22236
rect 1794 22176 1804 22236
rect 1704 22136 1804 22176
rect 4848 22176 4858 22236
rect 4938 22176 4948 22236
rect 4848 22136 4948 22176
rect 7980 22180 7990 22240
rect 8070 22180 8080 22240
rect 7980 22140 8080 22180
rect 11124 22180 11134 22240
rect 11214 22180 11224 22240
rect 11124 22140 11224 22180
rect 14326 22176 14336 22236
rect 14416 22176 14426 22236
rect 907 22079 2710 22136
rect 907 21992 941 22079
rect 2082 21992 2116 22079
rect 901 21980 947 21992
rect 901 21792 907 21980
rect 460 21780 506 21792
rect 460 21604 466 21780
rect 500 21604 506 21780
rect 460 21592 506 21604
rect 578 21780 624 21792
rect 578 21604 584 21780
rect 618 21604 624 21780
rect 578 21592 624 21604
rect 696 21780 742 21792
rect 696 21604 702 21780
rect 736 21604 742 21780
rect 696 21592 742 21604
rect 814 21780 907 21792
rect 814 21604 820 21780
rect 854 21604 907 21780
rect 941 21604 947 21980
rect 814 21592 947 21604
rect 1019 21980 1065 21992
rect 1019 21604 1025 21980
rect 1059 21604 1065 21980
rect 1019 21592 1065 21604
rect 1137 21980 1183 21992
rect 1137 21604 1143 21980
rect 1177 21604 1183 21980
rect 1137 21592 1183 21604
rect 1255 21980 1301 21992
rect 1255 21604 1261 21980
rect 1295 21604 1301 21980
rect 1255 21592 1301 21604
rect 1368 21980 1414 21992
rect 1368 21604 1374 21980
rect 1408 21604 1414 21980
rect 1368 21592 1414 21604
rect 1486 21980 1532 21992
rect 1486 21604 1492 21980
rect 1526 21604 1532 21980
rect 1486 21592 1532 21604
rect 1604 21980 1650 21992
rect 1604 21604 1610 21980
rect 1644 21604 1650 21980
rect 1604 21592 1650 21604
rect 1722 21980 1768 21992
rect 1722 21604 1728 21980
rect 1762 21604 1768 21980
rect 1722 21592 1768 21604
rect 1840 21980 1886 21992
rect 1840 21604 1846 21980
rect 1880 21604 1886 21980
rect 1840 21592 1886 21604
rect 1958 21980 2004 21992
rect 1958 21604 1964 21980
rect 1998 21604 2004 21980
rect 1958 21592 2004 21604
rect 2076 21980 2122 21992
rect 2076 21604 2082 21980
rect 2116 21604 2122 21980
rect 2076 21592 2122 21604
rect 2195 21980 2241 21992
rect 2195 21604 2201 21980
rect 2235 21604 2241 21980
rect 2195 21592 2241 21604
rect 2313 21980 2359 21992
rect 2313 21604 2319 21980
rect 2353 21604 2359 21980
rect 2313 21592 2359 21604
rect 2431 21980 2477 21992
rect 2431 21604 2437 21980
rect 2471 21604 2477 21980
rect 2431 21592 2477 21604
rect 2549 21980 2595 21992
rect 2549 21604 2555 21980
rect 2589 21604 2595 21980
rect 2673 21792 2710 22079
rect 4051 22079 5854 22136
rect 4051 21992 4085 22079
rect 5226 21992 5260 22079
rect 4045 21980 4091 21992
rect 4045 21792 4051 21980
rect 2549 21592 2595 21604
rect 2668 21780 2714 21792
rect 2668 21604 2674 21780
rect 2708 21604 2714 21780
rect 2668 21592 2714 21604
rect 2786 21780 2832 21792
rect 2786 21604 2792 21780
rect 2826 21604 2832 21780
rect 2786 21592 2832 21604
rect 2904 21780 2950 21792
rect 2904 21604 2910 21780
rect 2944 21604 2950 21780
rect 2904 21592 2950 21604
rect 3022 21780 3068 21792
rect 3022 21604 3028 21780
rect 3062 21604 3068 21780
rect 3022 21592 3068 21604
rect 3604 21780 3650 21792
rect 3604 21604 3610 21780
rect 3644 21604 3650 21780
rect 3604 21592 3650 21604
rect 3722 21780 3768 21792
rect 3722 21604 3728 21780
rect 3762 21604 3768 21780
rect 3722 21592 3768 21604
rect 3840 21780 3886 21792
rect 3840 21604 3846 21780
rect 3880 21604 3886 21780
rect 3840 21592 3886 21604
rect 3958 21780 4051 21792
rect 3958 21604 3964 21780
rect 3998 21604 4051 21780
rect 4085 21604 4091 21980
rect 3958 21592 4091 21604
rect 4163 21980 4209 21992
rect 4163 21604 4169 21980
rect 4203 21604 4209 21980
rect 4163 21592 4209 21604
rect 4281 21980 4327 21992
rect 4281 21604 4287 21980
rect 4321 21604 4327 21980
rect 4281 21592 4327 21604
rect 4399 21980 4445 21992
rect 4399 21604 4405 21980
rect 4439 21604 4445 21980
rect 4399 21592 4445 21604
rect 4512 21980 4558 21992
rect 4512 21604 4518 21980
rect 4552 21604 4558 21980
rect 4512 21592 4558 21604
rect 4630 21980 4676 21992
rect 4630 21604 4636 21980
rect 4670 21604 4676 21980
rect 4630 21592 4676 21604
rect 4748 21980 4794 21992
rect 4748 21604 4754 21980
rect 4788 21604 4794 21980
rect 4748 21592 4794 21604
rect 4866 21980 4912 21992
rect 4866 21604 4872 21980
rect 4906 21604 4912 21980
rect 4866 21592 4912 21604
rect 4984 21980 5030 21992
rect 4984 21604 4990 21980
rect 5024 21604 5030 21980
rect 4984 21592 5030 21604
rect 5102 21980 5148 21992
rect 5102 21604 5108 21980
rect 5142 21604 5148 21980
rect 5102 21592 5148 21604
rect 5220 21980 5266 21992
rect 5220 21604 5226 21980
rect 5260 21604 5266 21980
rect 5220 21592 5266 21604
rect 5339 21980 5385 21992
rect 5339 21604 5345 21980
rect 5379 21604 5385 21980
rect 5339 21592 5385 21604
rect 5457 21980 5503 21992
rect 5457 21604 5463 21980
rect 5497 21604 5503 21980
rect 5457 21592 5503 21604
rect 5575 21980 5621 21992
rect 5575 21604 5581 21980
rect 5615 21604 5621 21980
rect 5575 21592 5621 21604
rect 5693 21980 5739 21992
rect 5693 21604 5699 21980
rect 5733 21604 5739 21980
rect 5817 21792 5854 22079
rect 7183 22083 8986 22140
rect 7183 21996 7217 22083
rect 8358 21996 8392 22083
rect 7177 21984 7223 21996
rect 7177 21796 7183 21984
rect 5693 21592 5739 21604
rect 5812 21780 5858 21792
rect 5812 21604 5818 21780
rect 5852 21604 5858 21780
rect 5812 21592 5858 21604
rect 5930 21780 5976 21792
rect 5930 21604 5936 21780
rect 5970 21604 5976 21780
rect 5930 21592 5976 21604
rect 6048 21780 6094 21792
rect 6048 21604 6054 21780
rect 6088 21604 6094 21780
rect 6048 21592 6094 21604
rect 6166 21780 6212 21792
rect 6166 21604 6172 21780
rect 6206 21604 6212 21780
rect 6166 21592 6212 21604
rect 6736 21784 6782 21796
rect 6736 21608 6742 21784
rect 6776 21608 6782 21784
rect 6736 21596 6782 21608
rect 6854 21784 6900 21796
rect 6854 21608 6860 21784
rect 6894 21608 6900 21784
rect 6854 21596 6900 21608
rect 6972 21784 7018 21796
rect 6972 21608 6978 21784
rect 7012 21608 7018 21784
rect 6972 21596 7018 21608
rect 7090 21784 7183 21796
rect 7090 21608 7096 21784
rect 7130 21608 7183 21784
rect 7217 21608 7223 21984
rect 7090 21596 7223 21608
rect 7295 21984 7341 21996
rect 7295 21608 7301 21984
rect 7335 21608 7341 21984
rect 7295 21596 7341 21608
rect 7413 21984 7459 21996
rect 7413 21608 7419 21984
rect 7453 21608 7459 21984
rect 7413 21596 7459 21608
rect 7531 21984 7577 21996
rect 7531 21608 7537 21984
rect 7571 21608 7577 21984
rect 7531 21596 7577 21608
rect 7644 21984 7690 21996
rect 7644 21608 7650 21984
rect 7684 21608 7690 21984
rect 7644 21596 7690 21608
rect 7762 21984 7808 21996
rect 7762 21608 7768 21984
rect 7802 21608 7808 21984
rect 7762 21596 7808 21608
rect 7880 21984 7926 21996
rect 7880 21608 7886 21984
rect 7920 21608 7926 21984
rect 7880 21596 7926 21608
rect 7998 21984 8044 21996
rect 7998 21608 8004 21984
rect 8038 21608 8044 21984
rect 7998 21596 8044 21608
rect 8116 21984 8162 21996
rect 8116 21608 8122 21984
rect 8156 21608 8162 21984
rect 8116 21596 8162 21608
rect 8234 21984 8280 21996
rect 8234 21608 8240 21984
rect 8274 21608 8280 21984
rect 8234 21596 8280 21608
rect 8352 21984 8398 21996
rect 8352 21608 8358 21984
rect 8392 21608 8398 21984
rect 8352 21596 8398 21608
rect 8471 21984 8517 21996
rect 8471 21608 8477 21984
rect 8511 21608 8517 21984
rect 8471 21596 8517 21608
rect 8589 21984 8635 21996
rect 8589 21608 8595 21984
rect 8629 21608 8635 21984
rect 8589 21596 8635 21608
rect 8707 21984 8753 21996
rect 8707 21608 8713 21984
rect 8747 21608 8753 21984
rect 8707 21596 8753 21608
rect 8825 21984 8871 21996
rect 8825 21608 8831 21984
rect 8865 21608 8871 21984
rect 8949 21796 8986 22083
rect 10327 22083 12130 22140
rect 14326 22136 14426 22176
rect 17470 22176 17480 22236
rect 17560 22176 17570 22236
rect 17470 22136 17570 22176
rect 20602 22180 20612 22240
rect 20692 22180 20702 22240
rect 20602 22140 20702 22180
rect 23746 22180 23756 22240
rect 23836 22180 23846 22240
rect 23746 22140 23846 22180
rect 10327 21996 10361 22083
rect 11502 21996 11536 22083
rect 10321 21984 10367 21996
rect 10321 21796 10327 21984
rect 8825 21596 8871 21608
rect 8944 21784 8990 21796
rect 8944 21608 8950 21784
rect 8984 21608 8990 21784
rect 8944 21596 8990 21608
rect 9062 21784 9108 21796
rect 9062 21608 9068 21784
rect 9102 21608 9108 21784
rect 9062 21596 9108 21608
rect 9180 21784 9226 21796
rect 9180 21608 9186 21784
rect 9220 21608 9226 21784
rect 9180 21596 9226 21608
rect 9298 21784 9344 21796
rect 9298 21608 9304 21784
rect 9338 21608 9344 21784
rect 9298 21596 9344 21608
rect 9880 21784 9926 21796
rect 9880 21608 9886 21784
rect 9920 21608 9926 21784
rect 9880 21596 9926 21608
rect 9998 21784 10044 21796
rect 9998 21608 10004 21784
rect 10038 21608 10044 21784
rect 9998 21596 10044 21608
rect 10116 21784 10162 21796
rect 10116 21608 10122 21784
rect 10156 21608 10162 21784
rect 10116 21596 10162 21608
rect 10234 21784 10327 21796
rect 10234 21608 10240 21784
rect 10274 21608 10327 21784
rect 10361 21608 10367 21984
rect 10234 21596 10367 21608
rect 10439 21984 10485 21996
rect 10439 21608 10445 21984
rect 10479 21608 10485 21984
rect 10439 21596 10485 21608
rect 10557 21984 10603 21996
rect 10557 21608 10563 21984
rect 10597 21608 10603 21984
rect 10557 21596 10603 21608
rect 10675 21984 10721 21996
rect 10675 21608 10681 21984
rect 10715 21608 10721 21984
rect 10675 21596 10721 21608
rect 10788 21984 10834 21996
rect 10788 21608 10794 21984
rect 10828 21608 10834 21984
rect 10788 21596 10834 21608
rect 10906 21984 10952 21996
rect 10906 21608 10912 21984
rect 10946 21608 10952 21984
rect 10906 21596 10952 21608
rect 11024 21984 11070 21996
rect 11024 21608 11030 21984
rect 11064 21608 11070 21984
rect 11024 21596 11070 21608
rect 11142 21984 11188 21996
rect 11142 21608 11148 21984
rect 11182 21608 11188 21984
rect 11142 21596 11188 21608
rect 11260 21984 11306 21996
rect 11260 21608 11266 21984
rect 11300 21608 11306 21984
rect 11260 21596 11306 21608
rect 11378 21984 11424 21996
rect 11378 21608 11384 21984
rect 11418 21608 11424 21984
rect 11378 21596 11424 21608
rect 11496 21984 11542 21996
rect 11496 21608 11502 21984
rect 11536 21608 11542 21984
rect 11496 21596 11542 21608
rect 11615 21984 11661 21996
rect 11615 21608 11621 21984
rect 11655 21608 11661 21984
rect 11615 21596 11661 21608
rect 11733 21984 11779 21996
rect 11733 21608 11739 21984
rect 11773 21608 11779 21984
rect 11733 21596 11779 21608
rect 11851 21984 11897 21996
rect 11851 21608 11857 21984
rect 11891 21608 11897 21984
rect 11851 21596 11897 21608
rect 11969 21984 12015 21996
rect 11969 21608 11975 21984
rect 12009 21608 12015 21984
rect 12093 21796 12130 22083
rect 13529 22079 15332 22136
rect 13529 21992 13563 22079
rect 14704 21992 14738 22079
rect 13523 21980 13569 21992
rect 11969 21596 12015 21608
rect 12088 21784 12134 21796
rect 12088 21608 12094 21784
rect 12128 21608 12134 21784
rect 12088 21596 12134 21608
rect 12206 21784 12252 21796
rect 12206 21608 12212 21784
rect 12246 21608 12252 21784
rect 12206 21596 12252 21608
rect 12324 21784 12370 21796
rect 12324 21608 12330 21784
rect 12364 21608 12370 21784
rect 12324 21596 12370 21608
rect 12442 21784 12488 21796
rect 13523 21792 13529 21980
rect 12442 21608 12448 21784
rect 12482 21608 12488 21784
rect 12442 21596 12488 21608
rect 13082 21780 13128 21792
rect 13082 21604 13088 21780
rect 13122 21604 13128 21780
rect 61 21443 388 21444
rect 61 21381 324 21443
rect 378 21381 388 21443
rect 465 21406 500 21592
rect 1374 21508 1408 21592
rect 2555 21508 2589 21592
rect 1374 21466 2589 21508
rect 2555 21446 2589 21466
rect 2555 21430 2912 21446
rect 465 21389 1602 21406
rect 465 21355 1552 21389
rect 1586 21355 1602 21389
rect 2555 21396 2862 21430
rect 2896 21396 2912 21430
rect 2555 21380 2912 21396
rect 465 21339 1602 21355
rect 60 21294 382 21302
rect 60 21226 323 21294
rect 380 21226 390 21294
rect 60 21218 382 21226
rect 60 21018 225 21019
rect 60 21010 382 21018
rect 60 20942 323 21010
rect 380 20942 390 21010
rect 60 20934 382 20942
rect 60 20933 225 20934
rect 465 20829 500 21339
rect 555 21293 647 21306
rect 555 21230 567 21293
rect 638 21230 647 21293
rect 555 21221 647 21230
rect 1640 21293 1732 21303
rect 1640 21231 1652 21293
rect 1722 21231 1732 21293
rect 1640 21218 1732 21231
rect 3028 21238 3063 21592
rect 3609 21406 3644 21592
rect 4518 21508 4552 21592
rect 5699 21508 5733 21592
rect 4518 21466 5733 21508
rect 5699 21446 5733 21466
rect 5699 21430 6056 21446
rect 3342 21343 3352 21396
rect 3412 21343 3422 21396
rect 3609 21389 4746 21406
rect 3609 21355 4696 21389
rect 4730 21355 4746 21389
rect 5699 21396 6006 21430
rect 6040 21396 6056 21430
rect 5699 21380 6056 21396
rect 1887 21176 1952 21179
rect 1887 21173 1956 21176
rect 1887 21113 1893 21173
rect 1952 21113 1962 21173
rect 3028 21120 3209 21238
rect 3350 21186 3413 21343
rect 3609 21339 4746 21355
rect 3350 21178 3526 21186
rect 1887 21109 1956 21113
rect 1887 21107 1952 21109
rect 3028 21092 3210 21120
rect 3350 21110 3467 21178
rect 3524 21110 3534 21178
rect 3350 21102 3526 21110
rect 1522 21010 1614 21018
rect 1522 20945 1534 21010
rect 1602 20945 1614 21010
rect 1522 20933 1614 20945
rect 3028 20830 3063 21092
rect 465 20782 1837 20829
rect 2159 20783 3063 20830
rect 60 20768 387 20769
rect 60 20706 323 20768
rect 377 20706 387 20768
rect 1299 20659 1333 20782
rect 1771 20769 1837 20782
rect 1771 20735 1787 20769
rect 1821 20735 1837 20769
rect 1771 20719 1837 20735
rect 2160 20659 2194 20783
rect 1294 20647 1340 20659
rect 60 20633 387 20634
rect 60 20571 323 20633
rect 377 20571 387 20633
rect 62 20521 389 20522
rect 62 20459 325 20521
rect 379 20459 389 20521
rect 1294 20471 1300 20647
rect 1334 20471 1340 20647
rect 1294 20459 1340 20471
rect 1412 20647 1532 20659
rect 1412 20471 1418 20647
rect 1452 20471 1492 20647
rect 1412 20459 1492 20471
rect 62 20396 389 20397
rect 62 20334 325 20396
rect 379 20334 389 20396
rect 67 20155 394 20156
rect 67 20093 330 20155
rect 384 20093 394 20155
rect 1418 20092 1452 20459
rect 1486 20271 1492 20459
rect 1526 20271 1532 20647
rect 1486 20259 1532 20271
rect 1604 20647 1650 20659
rect 1604 20271 1610 20647
rect 1644 20271 1650 20647
rect 1604 20259 1650 20271
rect 1722 20647 1768 20659
rect 1722 20271 1728 20647
rect 1762 20271 1768 20647
rect 1722 20259 1768 20271
rect 1840 20647 1886 20659
rect 1840 20271 1846 20647
rect 1880 20271 1886 20647
rect 1840 20259 1886 20271
rect 1958 20647 2082 20659
rect 1958 20271 1964 20647
rect 1998 20471 2042 20647
rect 2076 20471 2082 20647
rect 1998 20459 2082 20471
rect 2154 20647 2200 20659
rect 2154 20471 2160 20647
rect 2194 20471 2200 20647
rect 2154 20459 2200 20471
rect 1998 20271 2004 20459
rect 1958 20259 2004 20271
rect 1728 20186 1762 20259
rect 1713 20170 1779 20186
rect 1713 20136 1729 20170
rect 1763 20136 1779 20170
rect 1713 20120 1779 20136
rect 2042 20092 2076 20459
rect 1418 20040 2076 20092
rect 1716 20018 1808 20040
rect 1716 19966 1728 20018
rect 1794 19966 1808 20018
rect 1716 19962 1808 19966
rect 64 19933 391 19934
rect 64 19871 327 19933
rect 381 19871 391 19933
rect 3149 19882 3210 21092
rect 3350 21010 3526 21018
rect 3350 20942 3467 21010
rect 3524 20942 3534 21010
rect 3350 20934 3526 20942
rect 3350 20772 3439 20934
rect 3609 20829 3644 21339
rect 3699 21293 3791 21306
rect 3699 21230 3711 21293
rect 3782 21230 3791 21293
rect 3699 21221 3791 21230
rect 4784 21293 4876 21303
rect 4784 21231 4796 21293
rect 4866 21231 4876 21293
rect 4784 21218 4876 21231
rect 6172 21238 6207 21592
rect 6741 21410 6776 21596
rect 7650 21512 7684 21596
rect 8831 21512 8865 21596
rect 7650 21470 8865 21512
rect 8831 21450 8865 21470
rect 8831 21434 9188 21450
rect 6741 21393 7878 21410
rect 6741 21359 7828 21393
rect 7862 21359 7878 21393
rect 8831 21400 9138 21434
rect 9172 21400 9188 21434
rect 8831 21384 9188 21400
rect 6741 21343 7878 21359
rect 5031 21176 5096 21179
rect 5031 21173 5100 21176
rect 5031 21113 5037 21173
rect 5096 21113 5106 21173
rect 5031 21109 5100 21113
rect 5031 21107 5096 21109
rect 6172 21092 6353 21238
rect 4666 21010 4758 21018
rect 4666 20945 4678 21010
rect 4746 20945 4758 21010
rect 4666 20933 4758 20945
rect 6172 20830 6207 21092
rect 3609 20782 4981 20829
rect 5303 20783 6207 20830
rect 3350 20712 3362 20772
rect 3432 20712 3442 20772
rect 3350 20705 3439 20712
rect 4443 20659 4477 20782
rect 4915 20769 4981 20782
rect 4915 20735 4931 20769
rect 4965 20735 4981 20769
rect 4915 20719 4981 20735
rect 5304 20659 5338 20783
rect 4438 20647 4484 20659
rect 4438 20471 4444 20647
rect 4478 20471 4484 20647
rect 4438 20459 4484 20471
rect 4556 20647 4676 20659
rect 4556 20471 4562 20647
rect 4596 20471 4636 20647
rect 4556 20459 4636 20471
rect 4562 20092 4596 20459
rect 4630 20271 4636 20459
rect 4670 20271 4676 20647
rect 4630 20259 4676 20271
rect 4748 20647 4794 20659
rect 4748 20271 4754 20647
rect 4788 20271 4794 20647
rect 4748 20259 4794 20271
rect 4866 20647 4912 20659
rect 4866 20271 4872 20647
rect 4906 20271 4912 20647
rect 4866 20259 4912 20271
rect 4984 20647 5030 20659
rect 4984 20271 4990 20647
rect 5024 20271 5030 20647
rect 4984 20259 5030 20271
rect 5102 20647 5226 20659
rect 5102 20271 5108 20647
rect 5142 20471 5186 20647
rect 5220 20471 5226 20647
rect 5142 20459 5226 20471
rect 5298 20647 5344 20659
rect 5298 20471 5304 20647
rect 5338 20471 5344 20647
rect 5298 20459 5344 20471
rect 5142 20271 5148 20459
rect 5102 20259 5148 20271
rect 4872 20186 4906 20259
rect 4857 20170 4923 20186
rect 4857 20136 4873 20170
rect 4907 20136 4923 20170
rect 4857 20120 4923 20136
rect 5186 20092 5220 20459
rect 6265 20162 6353 21092
rect 6482 21014 6658 21022
rect 6482 20946 6599 21014
rect 6656 20946 6666 21014
rect 6482 20938 6658 20946
rect 6502 20631 6579 20938
rect 6741 20833 6776 21343
rect 6831 21297 6923 21310
rect 6831 21234 6843 21297
rect 6914 21234 6923 21297
rect 6831 21225 6923 21234
rect 7916 21297 8008 21307
rect 7916 21235 7928 21297
rect 7998 21235 8008 21297
rect 7916 21222 8008 21235
rect 9304 21242 9339 21596
rect 9885 21410 9920 21596
rect 10794 21512 10828 21596
rect 11975 21512 12009 21596
rect 10794 21470 12009 21512
rect 11975 21450 12009 21470
rect 11975 21434 12332 21450
rect 9885 21393 11022 21410
rect 9885 21359 10972 21393
rect 11006 21359 11022 21393
rect 11975 21400 12282 21434
rect 12316 21400 12332 21434
rect 11975 21384 12332 21400
rect 9885 21343 11022 21359
rect 8163 21180 8228 21183
rect 8163 21177 8232 21180
rect 8163 21117 8169 21177
rect 8228 21117 8238 21177
rect 8163 21113 8232 21117
rect 8163 21111 8228 21113
rect 9304 21096 9485 21242
rect 9731 21182 9802 21190
rect 9731 21114 9743 21182
rect 9800 21114 9810 21182
rect 9731 21106 9802 21114
rect 7798 21014 7890 21022
rect 7798 20949 7810 21014
rect 7878 20949 7890 21014
rect 7798 20937 7890 20949
rect 9304 20834 9339 21096
rect 6741 20786 8113 20833
rect 8435 20787 9339 20834
rect 7575 20663 7609 20786
rect 8047 20773 8113 20786
rect 8047 20739 8063 20773
rect 8097 20739 8113 20773
rect 8047 20723 8113 20739
rect 8436 20663 8470 20787
rect 7570 20651 7616 20663
rect 6502 20574 6512 20631
rect 6576 20574 6586 20631
rect 6502 20570 6579 20574
rect 7570 20475 7576 20651
rect 7610 20475 7616 20651
rect 7570 20463 7616 20475
rect 7688 20651 7808 20663
rect 7688 20475 7694 20651
rect 7728 20475 7768 20651
rect 7688 20463 7768 20475
rect 6234 20096 6244 20162
rect 6303 20096 6353 20162
rect 7694 20096 7728 20463
rect 7762 20275 7768 20463
rect 7802 20275 7808 20651
rect 7762 20263 7808 20275
rect 7880 20651 7926 20663
rect 7880 20275 7886 20651
rect 7920 20275 7926 20651
rect 7880 20263 7926 20275
rect 7998 20651 8044 20663
rect 7998 20275 8004 20651
rect 8038 20275 8044 20651
rect 7998 20263 8044 20275
rect 8116 20651 8162 20663
rect 8116 20275 8122 20651
rect 8156 20275 8162 20651
rect 8116 20263 8162 20275
rect 8234 20651 8358 20663
rect 8234 20275 8240 20651
rect 8274 20475 8318 20651
rect 8352 20475 8358 20651
rect 8274 20463 8358 20475
rect 8430 20651 8476 20663
rect 8430 20475 8436 20651
rect 8470 20475 8476 20651
rect 8430 20463 8476 20475
rect 8274 20275 8280 20463
rect 8234 20263 8280 20275
rect 8004 20190 8038 20263
rect 7989 20174 8055 20190
rect 7989 20140 8005 20174
rect 8039 20140 8055 20174
rect 7989 20124 8055 20140
rect 8318 20096 8352 20463
rect 9388 20279 9485 21096
rect 9626 21014 9802 21022
rect 9626 20946 9743 21014
rect 9800 20946 9810 21014
rect 9626 20938 9802 20946
rect 9631 20526 9719 20938
rect 9885 20833 9920 21343
rect 9975 21297 10067 21310
rect 9975 21234 9987 21297
rect 10058 21234 10067 21297
rect 9975 21225 10067 21234
rect 11060 21297 11152 21307
rect 11060 21235 11072 21297
rect 11142 21235 11152 21297
rect 11060 21222 11152 21235
rect 12448 21242 12483 21596
rect 13082 21592 13128 21604
rect 13200 21780 13246 21792
rect 13200 21604 13206 21780
rect 13240 21604 13246 21780
rect 13200 21592 13246 21604
rect 13318 21780 13364 21792
rect 13318 21604 13324 21780
rect 13358 21604 13364 21780
rect 13318 21592 13364 21604
rect 13436 21780 13529 21792
rect 13436 21604 13442 21780
rect 13476 21604 13529 21780
rect 13563 21604 13569 21980
rect 13436 21592 13569 21604
rect 13641 21980 13687 21992
rect 13641 21604 13647 21980
rect 13681 21604 13687 21980
rect 13641 21592 13687 21604
rect 13759 21980 13805 21992
rect 13759 21604 13765 21980
rect 13799 21604 13805 21980
rect 13759 21592 13805 21604
rect 13877 21980 13923 21992
rect 13877 21604 13883 21980
rect 13917 21604 13923 21980
rect 13877 21592 13923 21604
rect 13990 21980 14036 21992
rect 13990 21604 13996 21980
rect 14030 21604 14036 21980
rect 13990 21592 14036 21604
rect 14108 21980 14154 21992
rect 14108 21604 14114 21980
rect 14148 21604 14154 21980
rect 14108 21592 14154 21604
rect 14226 21980 14272 21992
rect 14226 21604 14232 21980
rect 14266 21604 14272 21980
rect 14226 21592 14272 21604
rect 14344 21980 14390 21992
rect 14344 21604 14350 21980
rect 14384 21604 14390 21980
rect 14344 21592 14390 21604
rect 14462 21980 14508 21992
rect 14462 21604 14468 21980
rect 14502 21604 14508 21980
rect 14462 21592 14508 21604
rect 14580 21980 14626 21992
rect 14580 21604 14586 21980
rect 14620 21604 14626 21980
rect 14580 21592 14626 21604
rect 14698 21980 14744 21992
rect 14698 21604 14704 21980
rect 14738 21604 14744 21980
rect 14698 21592 14744 21604
rect 14817 21980 14863 21992
rect 14817 21604 14823 21980
rect 14857 21604 14863 21980
rect 14817 21592 14863 21604
rect 14935 21980 14981 21992
rect 14935 21604 14941 21980
rect 14975 21604 14981 21980
rect 14935 21592 14981 21604
rect 15053 21980 15099 21992
rect 15053 21604 15059 21980
rect 15093 21604 15099 21980
rect 15053 21592 15099 21604
rect 15171 21980 15217 21992
rect 15171 21604 15177 21980
rect 15211 21604 15217 21980
rect 15295 21792 15332 22079
rect 16673 22079 18476 22136
rect 16673 21992 16707 22079
rect 17848 21992 17882 22079
rect 16667 21980 16713 21992
rect 16667 21792 16673 21980
rect 15171 21592 15217 21604
rect 15290 21780 15336 21792
rect 15290 21604 15296 21780
rect 15330 21604 15336 21780
rect 15290 21592 15336 21604
rect 15408 21780 15454 21792
rect 15408 21604 15414 21780
rect 15448 21604 15454 21780
rect 15408 21592 15454 21604
rect 15526 21780 15572 21792
rect 15526 21604 15532 21780
rect 15566 21604 15572 21780
rect 15526 21592 15572 21604
rect 15644 21780 15690 21792
rect 15644 21604 15650 21780
rect 15684 21604 15690 21780
rect 15644 21592 15690 21604
rect 16226 21780 16272 21792
rect 16226 21604 16232 21780
rect 16266 21604 16272 21780
rect 16226 21592 16272 21604
rect 16344 21780 16390 21792
rect 16344 21604 16350 21780
rect 16384 21604 16390 21780
rect 16344 21592 16390 21604
rect 16462 21780 16508 21792
rect 16462 21604 16468 21780
rect 16502 21604 16508 21780
rect 16462 21592 16508 21604
rect 16580 21780 16673 21792
rect 16580 21604 16586 21780
rect 16620 21604 16673 21780
rect 16707 21604 16713 21980
rect 16580 21592 16713 21604
rect 16785 21980 16831 21992
rect 16785 21604 16791 21980
rect 16825 21604 16831 21980
rect 16785 21592 16831 21604
rect 16903 21980 16949 21992
rect 16903 21604 16909 21980
rect 16943 21604 16949 21980
rect 16903 21592 16949 21604
rect 17021 21980 17067 21992
rect 17021 21604 17027 21980
rect 17061 21604 17067 21980
rect 17021 21592 17067 21604
rect 17134 21980 17180 21992
rect 17134 21604 17140 21980
rect 17174 21604 17180 21980
rect 17134 21592 17180 21604
rect 17252 21980 17298 21992
rect 17252 21604 17258 21980
rect 17292 21604 17298 21980
rect 17252 21592 17298 21604
rect 17370 21980 17416 21992
rect 17370 21604 17376 21980
rect 17410 21604 17416 21980
rect 17370 21592 17416 21604
rect 17488 21980 17534 21992
rect 17488 21604 17494 21980
rect 17528 21604 17534 21980
rect 17488 21592 17534 21604
rect 17606 21980 17652 21992
rect 17606 21604 17612 21980
rect 17646 21604 17652 21980
rect 17606 21592 17652 21604
rect 17724 21980 17770 21992
rect 17724 21604 17730 21980
rect 17764 21604 17770 21980
rect 17724 21592 17770 21604
rect 17842 21980 17888 21992
rect 17842 21604 17848 21980
rect 17882 21604 17888 21980
rect 17842 21592 17888 21604
rect 17961 21980 18007 21992
rect 17961 21604 17967 21980
rect 18001 21604 18007 21980
rect 17961 21592 18007 21604
rect 18079 21980 18125 21992
rect 18079 21604 18085 21980
rect 18119 21604 18125 21980
rect 18079 21592 18125 21604
rect 18197 21980 18243 21992
rect 18197 21604 18203 21980
rect 18237 21604 18243 21980
rect 18197 21592 18243 21604
rect 18315 21980 18361 21992
rect 18315 21604 18321 21980
rect 18355 21604 18361 21980
rect 18439 21792 18476 22079
rect 19805 22083 21608 22140
rect 19805 21996 19839 22083
rect 20980 21996 21014 22083
rect 19799 21984 19845 21996
rect 19799 21796 19805 21984
rect 18315 21592 18361 21604
rect 18434 21780 18480 21792
rect 18434 21604 18440 21780
rect 18474 21604 18480 21780
rect 18434 21592 18480 21604
rect 18552 21780 18598 21792
rect 18552 21604 18558 21780
rect 18592 21604 18598 21780
rect 18552 21592 18598 21604
rect 18670 21780 18716 21792
rect 18670 21604 18676 21780
rect 18710 21604 18716 21780
rect 18670 21592 18716 21604
rect 18788 21780 18834 21792
rect 18788 21604 18794 21780
rect 18828 21604 18834 21780
rect 18788 21592 18834 21604
rect 19358 21784 19404 21796
rect 19358 21608 19364 21784
rect 19398 21608 19404 21784
rect 19358 21596 19404 21608
rect 19476 21784 19522 21796
rect 19476 21608 19482 21784
rect 19516 21608 19522 21784
rect 19476 21596 19522 21608
rect 19594 21784 19640 21796
rect 19594 21608 19600 21784
rect 19634 21608 19640 21784
rect 19594 21596 19640 21608
rect 19712 21784 19805 21796
rect 19712 21608 19718 21784
rect 19752 21608 19805 21784
rect 19839 21608 19845 21984
rect 19712 21596 19845 21608
rect 19917 21984 19963 21996
rect 19917 21608 19923 21984
rect 19957 21608 19963 21984
rect 19917 21596 19963 21608
rect 20035 21984 20081 21996
rect 20035 21608 20041 21984
rect 20075 21608 20081 21984
rect 20035 21596 20081 21608
rect 20153 21984 20199 21996
rect 20153 21608 20159 21984
rect 20193 21608 20199 21984
rect 20153 21596 20199 21608
rect 20266 21984 20312 21996
rect 20266 21608 20272 21984
rect 20306 21608 20312 21984
rect 20266 21596 20312 21608
rect 20384 21984 20430 21996
rect 20384 21608 20390 21984
rect 20424 21608 20430 21984
rect 20384 21596 20430 21608
rect 20502 21984 20548 21996
rect 20502 21608 20508 21984
rect 20542 21608 20548 21984
rect 20502 21596 20548 21608
rect 20620 21984 20666 21996
rect 20620 21608 20626 21984
rect 20660 21608 20666 21984
rect 20620 21596 20666 21608
rect 20738 21984 20784 21996
rect 20738 21608 20744 21984
rect 20778 21608 20784 21984
rect 20738 21596 20784 21608
rect 20856 21984 20902 21996
rect 20856 21608 20862 21984
rect 20896 21608 20902 21984
rect 20856 21596 20902 21608
rect 20974 21984 21020 21996
rect 20974 21608 20980 21984
rect 21014 21608 21020 21984
rect 20974 21596 21020 21608
rect 21093 21984 21139 21996
rect 21093 21608 21099 21984
rect 21133 21608 21139 21984
rect 21093 21596 21139 21608
rect 21211 21984 21257 21996
rect 21211 21608 21217 21984
rect 21251 21608 21257 21984
rect 21211 21596 21257 21608
rect 21329 21984 21375 21996
rect 21329 21608 21335 21984
rect 21369 21608 21375 21984
rect 21329 21596 21375 21608
rect 21447 21984 21493 21996
rect 21447 21608 21453 21984
rect 21487 21608 21493 21984
rect 21571 21796 21608 22083
rect 22949 22083 24752 22140
rect 22949 21996 22983 22083
rect 24124 21996 24158 22083
rect 22943 21984 22989 21996
rect 22943 21796 22949 21984
rect 21447 21596 21493 21608
rect 21566 21784 21612 21796
rect 21566 21608 21572 21784
rect 21606 21608 21612 21784
rect 21566 21596 21612 21608
rect 21684 21784 21730 21796
rect 21684 21608 21690 21784
rect 21724 21608 21730 21784
rect 21684 21596 21730 21608
rect 21802 21784 21848 21796
rect 21802 21608 21808 21784
rect 21842 21608 21848 21784
rect 21802 21596 21848 21608
rect 21920 21784 21966 21796
rect 21920 21608 21926 21784
rect 21960 21608 21966 21784
rect 21920 21596 21966 21608
rect 22502 21784 22548 21796
rect 22502 21608 22508 21784
rect 22542 21608 22548 21784
rect 22502 21596 22548 21608
rect 22620 21784 22666 21796
rect 22620 21608 22626 21784
rect 22660 21608 22666 21784
rect 22620 21596 22666 21608
rect 22738 21784 22784 21796
rect 22738 21608 22744 21784
rect 22778 21608 22784 21784
rect 22738 21596 22784 21608
rect 22856 21784 22949 21796
rect 22856 21608 22862 21784
rect 22896 21608 22949 21784
rect 22983 21608 22989 21984
rect 22856 21596 22989 21608
rect 23061 21984 23107 21996
rect 23061 21608 23067 21984
rect 23101 21608 23107 21984
rect 23061 21596 23107 21608
rect 23179 21984 23225 21996
rect 23179 21608 23185 21984
rect 23219 21608 23225 21984
rect 23179 21596 23225 21608
rect 23297 21984 23343 21996
rect 23297 21608 23303 21984
rect 23337 21608 23343 21984
rect 23297 21596 23343 21608
rect 23410 21984 23456 21996
rect 23410 21608 23416 21984
rect 23450 21608 23456 21984
rect 23410 21596 23456 21608
rect 23528 21984 23574 21996
rect 23528 21608 23534 21984
rect 23568 21608 23574 21984
rect 23528 21596 23574 21608
rect 23646 21984 23692 21996
rect 23646 21608 23652 21984
rect 23686 21608 23692 21984
rect 23646 21596 23692 21608
rect 23764 21984 23810 21996
rect 23764 21608 23770 21984
rect 23804 21608 23810 21984
rect 23764 21596 23810 21608
rect 23882 21984 23928 21996
rect 23882 21608 23888 21984
rect 23922 21608 23928 21984
rect 23882 21596 23928 21608
rect 24000 21984 24046 21996
rect 24000 21608 24006 21984
rect 24040 21608 24046 21984
rect 24000 21596 24046 21608
rect 24118 21984 24164 21996
rect 24118 21608 24124 21984
rect 24158 21608 24164 21984
rect 24118 21596 24164 21608
rect 24237 21984 24283 21996
rect 24237 21608 24243 21984
rect 24277 21608 24283 21984
rect 24237 21596 24283 21608
rect 24355 21984 24401 21996
rect 24355 21608 24361 21984
rect 24395 21608 24401 21984
rect 24355 21596 24401 21608
rect 24473 21984 24519 21996
rect 24473 21608 24479 21984
rect 24513 21608 24519 21984
rect 24473 21596 24519 21608
rect 24591 21984 24637 21996
rect 24591 21608 24597 21984
rect 24631 21608 24637 21984
rect 24715 21796 24752 22083
rect 24591 21596 24637 21608
rect 24710 21784 24756 21796
rect 24710 21608 24716 21784
rect 24750 21608 24756 21784
rect 24710 21596 24756 21608
rect 24828 21784 24874 21796
rect 24828 21608 24834 21784
rect 24868 21608 24874 21784
rect 24828 21596 24874 21608
rect 24946 21784 24992 21796
rect 24946 21608 24952 21784
rect 24986 21608 24992 21784
rect 24946 21596 24992 21608
rect 25064 21784 25110 21796
rect 25064 21608 25070 21784
rect 25104 21608 25110 21784
rect 25064 21596 25110 21608
rect 13087 21406 13122 21592
rect 13996 21508 14030 21592
rect 15177 21508 15211 21592
rect 13996 21466 15211 21508
rect 15177 21446 15211 21466
rect 15177 21430 15534 21446
rect 13087 21389 14224 21406
rect 13087 21355 14174 21389
rect 14208 21355 14224 21389
rect 15177 21396 15484 21430
rect 15518 21396 15534 21430
rect 15177 21380 15534 21396
rect 13087 21339 14224 21355
rect 11307 21180 11372 21183
rect 11307 21177 11376 21180
rect 11307 21117 11313 21177
rect 11372 21117 11382 21177
rect 11307 21113 11376 21117
rect 11307 21111 11372 21113
rect 12448 21096 12629 21242
rect 10942 21014 11034 21022
rect 10942 20949 10954 21014
rect 11022 20949 11034 21014
rect 10942 20937 11034 20949
rect 12448 20834 12483 21096
rect 9885 20786 11257 20833
rect 11579 20787 12483 20834
rect 10719 20663 10753 20786
rect 11191 20773 11257 20786
rect 11191 20739 11207 20773
rect 11241 20739 11257 20773
rect 11191 20723 11257 20739
rect 11580 20663 11614 20787
rect 9631 20468 9654 20526
rect 9708 20468 9719 20526
rect 9631 20458 9719 20468
rect 10714 20651 10760 20663
rect 10714 20475 10720 20651
rect 10754 20475 10760 20651
rect 10714 20463 10760 20475
rect 10832 20651 10952 20663
rect 10832 20475 10838 20651
rect 10872 20475 10912 20651
rect 10832 20463 10912 20475
rect 9360 20222 9370 20279
rect 9429 20222 9485 20279
rect 9360 20221 9485 20222
rect 4562 20040 5220 20092
rect 7694 20044 8352 20096
rect 10838 20096 10872 20463
rect 10906 20275 10912 20463
rect 10946 20275 10952 20651
rect 10906 20263 10952 20275
rect 11024 20651 11070 20663
rect 11024 20275 11030 20651
rect 11064 20275 11070 20651
rect 11024 20263 11070 20275
rect 11142 20651 11188 20663
rect 11142 20275 11148 20651
rect 11182 20275 11188 20651
rect 11142 20263 11188 20275
rect 11260 20651 11306 20663
rect 11260 20275 11266 20651
rect 11300 20275 11306 20651
rect 11260 20263 11306 20275
rect 11378 20651 11502 20663
rect 11378 20275 11384 20651
rect 11418 20475 11462 20651
rect 11496 20475 11502 20651
rect 11418 20463 11502 20475
rect 11574 20651 11620 20663
rect 11574 20475 11580 20651
rect 11614 20475 11620 20651
rect 11574 20463 11620 20475
rect 11418 20275 11424 20463
rect 11378 20263 11424 20275
rect 11148 20190 11182 20263
rect 11133 20174 11199 20190
rect 11133 20140 11149 20174
rect 11183 20140 11199 20174
rect 11133 20124 11199 20140
rect 11462 20096 11496 20463
rect 12535 20427 12628 21096
rect 12535 20359 12545 20427
rect 12607 20359 12628 20427
rect 12535 20354 12628 20359
rect 12828 21010 13004 21018
rect 12828 20942 12945 21010
rect 13002 20942 13012 21010
rect 12828 20934 13004 20942
rect 12828 20302 12894 20934
rect 13087 20829 13122 21339
rect 13177 21293 13269 21306
rect 13177 21230 13189 21293
rect 13260 21230 13269 21293
rect 13177 21221 13269 21230
rect 14262 21293 14354 21303
rect 14262 21231 14274 21293
rect 14344 21231 14354 21293
rect 14262 21218 14354 21231
rect 15650 21238 15685 21592
rect 16231 21406 16266 21592
rect 17140 21508 17174 21592
rect 18321 21508 18355 21592
rect 17140 21466 18355 21508
rect 18321 21446 18355 21466
rect 18321 21430 18678 21446
rect 16231 21389 17368 21406
rect 16231 21355 17318 21389
rect 17352 21355 17368 21389
rect 18321 21396 18628 21430
rect 18662 21396 18678 21430
rect 18321 21380 18678 21396
rect 16231 21339 17368 21355
rect 14509 21176 14574 21179
rect 14509 21173 14578 21176
rect 14509 21113 14515 21173
rect 14574 21113 14584 21173
rect 14509 21109 14578 21113
rect 14509 21107 14574 21109
rect 15650 21092 15831 21238
rect 16077 21178 16148 21183
rect 16077 21110 16089 21178
rect 16146 21110 16156 21178
rect 16077 21104 16148 21110
rect 14144 21010 14236 21018
rect 14144 20945 14156 21010
rect 14224 20945 14236 21010
rect 14144 20933 14236 20945
rect 15650 20830 15685 21092
rect 13087 20782 14459 20829
rect 14781 20783 15685 20830
rect 13921 20659 13955 20782
rect 14393 20769 14459 20782
rect 14393 20735 14409 20769
rect 14443 20735 14459 20769
rect 14393 20719 14459 20735
rect 14782 20659 14816 20783
rect 13916 20647 13962 20659
rect 13916 20471 13922 20647
rect 13956 20471 13962 20647
rect 13916 20459 13962 20471
rect 14034 20647 14154 20659
rect 14034 20471 14040 20647
rect 14074 20471 14114 20647
rect 14034 20459 14114 20471
rect 12814 20241 12824 20302
rect 12893 20241 12903 20302
rect 12814 20233 12903 20241
rect 10838 20044 11496 20096
rect 14040 20092 14074 20459
rect 14108 20271 14114 20459
rect 14148 20271 14154 20647
rect 14108 20259 14154 20271
rect 14226 20647 14272 20659
rect 14226 20271 14232 20647
rect 14266 20271 14272 20647
rect 14226 20259 14272 20271
rect 14344 20647 14390 20659
rect 14344 20271 14350 20647
rect 14384 20271 14390 20647
rect 14344 20259 14390 20271
rect 14462 20647 14508 20659
rect 14462 20271 14468 20647
rect 14502 20271 14508 20647
rect 14462 20259 14508 20271
rect 14580 20647 14704 20659
rect 14580 20271 14586 20647
rect 14620 20471 14664 20647
rect 14698 20471 14704 20647
rect 14620 20459 14704 20471
rect 14776 20647 14822 20659
rect 14776 20471 14782 20647
rect 14816 20471 14822 20647
rect 15761 20578 15831 21092
rect 15972 21010 16148 21018
rect 15972 20942 16089 21010
rect 16146 20942 16156 21010
rect 15972 20934 16148 20942
rect 15760 20509 15770 20578
rect 15826 20509 15836 20578
rect 15761 20503 15831 20509
rect 14776 20459 14822 20471
rect 14620 20271 14626 20459
rect 14580 20259 14626 20271
rect 14350 20186 14384 20259
rect 14335 20170 14401 20186
rect 14335 20136 14351 20170
rect 14385 20136 14401 20170
rect 14335 20120 14401 20136
rect 14664 20092 14698 20459
rect 15972 20167 16055 20934
rect 16231 20829 16266 21339
rect 16321 21293 16413 21306
rect 16321 21230 16333 21293
rect 16404 21230 16413 21293
rect 16321 21221 16413 21230
rect 17406 21293 17498 21303
rect 17406 21231 17418 21293
rect 17488 21231 17498 21293
rect 17406 21218 17498 21231
rect 18794 21238 18829 21592
rect 19363 21410 19398 21596
rect 20272 21512 20306 21596
rect 21453 21512 21487 21596
rect 20272 21470 21487 21512
rect 21453 21450 21487 21470
rect 21453 21434 21810 21450
rect 19363 21393 20500 21410
rect 19363 21359 20450 21393
rect 20484 21359 20500 21393
rect 21453 21400 21760 21434
rect 21794 21400 21810 21434
rect 21453 21384 21810 21400
rect 19363 21343 20500 21359
rect 17653 21176 17718 21179
rect 17653 21173 17722 21176
rect 17653 21113 17659 21173
rect 17718 21113 17728 21173
rect 17653 21109 17722 21113
rect 17653 21107 17718 21109
rect 18794 21092 18975 21238
rect 19210 21182 19280 21187
rect 19210 21114 19221 21182
rect 19278 21114 19288 21182
rect 19210 21108 19280 21114
rect 17288 21010 17380 21018
rect 17288 20945 17300 21010
rect 17368 20945 17380 21010
rect 17288 20933 17380 20945
rect 18794 20830 18829 21092
rect 16231 20782 17603 20829
rect 17925 20783 18829 20830
rect 17065 20659 17099 20782
rect 17537 20769 17603 20782
rect 17537 20735 17553 20769
rect 17587 20735 17603 20769
rect 17537 20719 17603 20735
rect 17926 20659 17960 20783
rect 18903 20731 18975 21092
rect 19104 21014 19280 21022
rect 19104 20946 19221 21014
rect 19278 20946 19288 21014
rect 19104 20938 19280 20946
rect 18896 20672 18906 20731
rect 18970 20672 18980 20731
rect 17060 20647 17106 20659
rect 17060 20471 17066 20647
rect 17100 20471 17106 20647
rect 17060 20459 17106 20471
rect 17178 20647 17298 20659
rect 17178 20471 17184 20647
rect 17218 20471 17258 20647
rect 17178 20459 17258 20471
rect 15965 20100 15975 20167
rect 16032 20103 16055 20167
rect 16032 20100 16042 20103
rect 4860 20018 4952 20040
rect 4860 19966 4872 20018
rect 4938 19966 4952 20018
rect 7992 20022 8084 20044
rect 7992 19970 8004 20022
rect 8070 19970 8084 20022
rect 7992 19966 8084 19970
rect 11136 20022 11228 20044
rect 14040 20040 14698 20092
rect 17184 20092 17218 20459
rect 17252 20271 17258 20459
rect 17292 20271 17298 20647
rect 17252 20259 17298 20271
rect 17370 20647 17416 20659
rect 17370 20271 17376 20647
rect 17410 20271 17416 20647
rect 17370 20259 17416 20271
rect 17488 20647 17534 20659
rect 17488 20271 17494 20647
rect 17528 20271 17534 20647
rect 17488 20259 17534 20271
rect 17606 20647 17652 20659
rect 17606 20271 17612 20647
rect 17646 20271 17652 20647
rect 17606 20259 17652 20271
rect 17724 20647 17848 20659
rect 17724 20271 17730 20647
rect 17764 20471 17808 20647
rect 17842 20471 17848 20647
rect 17764 20459 17848 20471
rect 17920 20647 17966 20659
rect 17920 20471 17926 20647
rect 17960 20471 17966 20647
rect 17920 20459 17966 20471
rect 17764 20271 17770 20459
rect 17724 20259 17770 20271
rect 17494 20186 17528 20259
rect 17479 20170 17545 20186
rect 17479 20136 17495 20170
rect 17529 20136 17545 20170
rect 17479 20120 17545 20136
rect 17808 20092 17842 20459
rect 17184 20040 17842 20092
rect 11136 19970 11148 20022
rect 11214 19970 11228 20022
rect 11136 19966 11228 19970
rect 14338 20018 14430 20040
rect 14338 19966 14350 20018
rect 14416 19966 14430 20018
rect 4860 19962 4952 19966
rect 14338 19962 14430 19966
rect 17482 20018 17574 20040
rect 17482 19966 17494 20018
rect 17560 19966 17574 20018
rect 17482 19962 17574 19966
rect 19104 19951 19177 20938
rect 19363 20833 19398 21343
rect 19453 21297 19545 21310
rect 19453 21234 19465 21297
rect 19536 21234 19545 21297
rect 19453 21225 19545 21234
rect 20538 21297 20630 21307
rect 20538 21235 20550 21297
rect 20620 21235 20630 21297
rect 20538 21222 20630 21235
rect 21926 21242 21961 21596
rect 22507 21410 22542 21596
rect 23416 21512 23450 21596
rect 24597 21512 24631 21596
rect 23416 21470 24631 21512
rect 24597 21450 24631 21470
rect 24597 21434 24954 21450
rect 22507 21393 23644 21410
rect 22507 21359 23594 21393
rect 23628 21359 23644 21393
rect 24597 21400 24904 21434
rect 24938 21400 24954 21434
rect 24597 21384 24954 21400
rect 22507 21343 23644 21359
rect 20785 21180 20850 21183
rect 20785 21177 20854 21180
rect 20785 21117 20791 21177
rect 20850 21117 20860 21177
rect 21926 21147 22107 21242
rect 22354 21182 22424 21187
rect 20785 21113 20854 21117
rect 20785 21111 20850 21113
rect 21926 21096 22108 21147
rect 22354 21114 22365 21182
rect 22422 21114 22432 21182
rect 22354 21108 22424 21114
rect 20420 21014 20512 21022
rect 20420 20949 20432 21014
rect 20500 20949 20512 21014
rect 20420 20937 20512 20949
rect 21926 20834 21961 21096
rect 19363 20786 20735 20833
rect 21057 20787 21961 20834
rect 22013 20858 22108 21096
rect 22013 20801 22051 20858
rect 22104 20801 22114 20858
rect 22507 20833 22542 21343
rect 22597 21297 22689 21310
rect 22597 21234 22609 21297
rect 22680 21234 22689 21297
rect 22597 21225 22689 21234
rect 23682 21297 23774 21307
rect 23682 21235 23694 21297
rect 23764 21235 23774 21297
rect 23682 21222 23774 21235
rect 25070 21242 25105 21596
rect 23929 21180 23994 21183
rect 23929 21177 23998 21180
rect 23929 21117 23935 21177
rect 23994 21117 24004 21177
rect 25070 21154 25684 21242
rect 23929 21113 23998 21117
rect 23929 21111 23994 21113
rect 23564 21014 23656 21022
rect 23564 20949 23576 21014
rect 23644 20949 23656 21014
rect 23564 20937 23656 20949
rect 25070 20834 25105 21154
rect 22013 20793 22108 20801
rect 20197 20663 20231 20786
rect 20669 20773 20735 20786
rect 20669 20739 20685 20773
rect 20719 20739 20735 20773
rect 20669 20723 20735 20739
rect 21058 20663 21092 20787
rect 22507 20786 23879 20833
rect 24201 20787 25105 20834
rect 25536 20866 25685 20878
rect 25536 20795 25549 20866
rect 25620 20795 25685 20866
rect 23341 20663 23375 20786
rect 23813 20773 23879 20786
rect 23813 20739 23829 20773
rect 23863 20739 23879 20773
rect 23813 20723 23879 20739
rect 24202 20663 24236 20787
rect 25536 20784 25685 20795
rect 25527 20730 25686 20741
rect 25527 20670 25537 20730
rect 25603 20670 25686 20730
rect 20192 20651 20238 20663
rect 20192 20475 20198 20651
rect 20232 20475 20238 20651
rect 20192 20463 20238 20475
rect 20310 20651 20430 20663
rect 20310 20475 20316 20651
rect 20350 20475 20390 20651
rect 20310 20463 20390 20475
rect 20316 20096 20350 20463
rect 20384 20275 20390 20463
rect 20424 20275 20430 20651
rect 20384 20263 20430 20275
rect 20502 20651 20548 20663
rect 20502 20275 20508 20651
rect 20542 20275 20548 20651
rect 20502 20263 20548 20275
rect 20620 20651 20666 20663
rect 20620 20275 20626 20651
rect 20660 20275 20666 20651
rect 20620 20263 20666 20275
rect 20738 20651 20784 20663
rect 20738 20275 20744 20651
rect 20778 20275 20784 20651
rect 20738 20263 20784 20275
rect 20856 20651 20980 20663
rect 20856 20275 20862 20651
rect 20896 20475 20940 20651
rect 20974 20475 20980 20651
rect 20896 20463 20980 20475
rect 21052 20651 21098 20663
rect 21052 20475 21058 20651
rect 21092 20475 21098 20651
rect 21052 20463 21098 20475
rect 23336 20651 23382 20663
rect 23336 20475 23342 20651
rect 23376 20475 23382 20651
rect 23336 20463 23382 20475
rect 23454 20651 23574 20663
rect 23454 20475 23460 20651
rect 23494 20475 23534 20651
rect 23454 20463 23534 20475
rect 20896 20275 20902 20463
rect 20856 20263 20902 20275
rect 20626 20190 20660 20263
rect 20611 20174 20677 20190
rect 20611 20140 20627 20174
rect 20661 20140 20677 20174
rect 20611 20124 20677 20140
rect 20940 20096 20974 20463
rect 20316 20044 20974 20096
rect 23460 20096 23494 20463
rect 23528 20275 23534 20463
rect 23568 20275 23574 20651
rect 23528 20263 23574 20275
rect 23646 20651 23692 20663
rect 23646 20275 23652 20651
rect 23686 20275 23692 20651
rect 23646 20263 23692 20275
rect 23764 20651 23810 20663
rect 23764 20275 23770 20651
rect 23804 20275 23810 20651
rect 23764 20263 23810 20275
rect 23882 20651 23928 20663
rect 23882 20275 23888 20651
rect 23922 20275 23928 20651
rect 23882 20263 23928 20275
rect 24000 20651 24124 20663
rect 24000 20275 24006 20651
rect 24040 20475 24084 20651
rect 24118 20475 24124 20651
rect 24040 20463 24124 20475
rect 24196 20651 24242 20663
rect 25527 20659 25686 20670
rect 24196 20475 24202 20651
rect 24236 20475 24242 20651
rect 25516 20572 25686 20583
rect 25516 20503 25527 20572
rect 25591 20503 25686 20572
rect 25516 20492 25686 20503
rect 24196 20463 24242 20475
rect 24040 20275 24046 20463
rect 24000 20263 24046 20275
rect 23770 20190 23804 20263
rect 23755 20174 23821 20190
rect 23755 20140 23771 20174
rect 23805 20140 23821 20174
rect 23755 20124 23821 20140
rect 24084 20096 24118 20463
rect 25516 20426 25686 20437
rect 25516 20357 25527 20426
rect 25591 20357 25686 20426
rect 25516 20346 25686 20357
rect 25516 20286 25686 20297
rect 25516 20217 25527 20286
rect 25591 20217 25686 20286
rect 25516 20206 25686 20217
rect 23460 20044 24118 20096
rect 25515 20147 25685 20158
rect 25515 20078 25526 20147
rect 25590 20078 25685 20147
rect 25515 20067 25685 20078
rect 20614 20022 20706 20044
rect 20614 19970 20626 20022
rect 20692 19970 20706 20022
rect 20614 19966 20706 19970
rect 23758 20022 23850 20044
rect 23758 19970 23770 20022
rect 23836 19970 23850 20022
rect 23758 19966 23850 19970
rect 3101 19801 3111 19882
rect 3184 19801 3210 19882
rect 19094 19875 19104 19951
rect 19174 19875 19184 19951
rect 25515 19879 25685 19890
rect 3149 19800 3210 19801
rect 25515 19810 25526 19879
rect 25590 19810 25685 19879
rect 25515 19799 25685 19810
rect 123 18577 230 18636
rect 290 18577 300 18636
rect 13002 18615 22814 18621
rect 13002 18561 13012 18615
rect 13066 18561 22814 18615
rect 13002 18557 22814 18561
rect 721 18527 13187 18528
rect 721 18522 22676 18527
rect 721 18468 13106 18522
rect 13160 18468 22676 18522
rect 721 18464 22676 18468
rect 123 18436 260 18439
rect 123 18374 227 18436
rect 287 18374 297 18436
rect 123 18246 250 18250
rect 123 18184 220 18246
rect 280 18184 290 18246
rect 123 17995 220 18064
rect 280 17995 290 18064
rect 123 17814 207 17877
rect 268 17814 278 17877
rect 123 17614 194 17686
rect 265 17614 275 17686
rect 123 15880 207 15881
rect 123 15825 211 15880
rect 265 15825 275 15880
rect 125 15451 182 15505
rect 238 15451 248 15505
rect 98 11425 203 11431
rect 98 11350 201 11425
rect 263 11350 273 11425
rect 99 11098 204 11104
rect 99 11023 202 11098
rect 264 11023 274 11098
rect 721 7157 800 18464
rect 13096 18463 22676 18464
rect 11467 18430 21646 18435
rect 11467 18376 11474 18430
rect 11528 18376 21646 18430
rect 11467 18371 21646 18376
rect 997 18342 1116 18343
rect 997 18341 2349 18342
rect 974 18335 21513 18341
rect 974 18281 11649 18335
rect 11703 18281 21513 18335
rect 974 18278 21513 18281
rect 405 7096 471 7157
rect 526 7096 536 7157
rect 717 7099 727 7157
rect 795 7099 805 7157
rect 405 6804 471 6865
rect 526 6804 536 6865
rect 405 6499 471 6560
rect 526 6499 536 6560
rect 405 6338 471 6399
rect 526 6338 536 6399
rect 405 6187 471 6248
rect 527 6187 537 6248
rect 405 6027 471 6088
rect 526 6027 536 6088
rect 405 5840 471 5901
rect 526 5840 536 5901
rect 405 5634 471 5695
rect 526 5634 536 5695
rect 721 3404 800 7099
rect 974 6863 1054 18278
rect 11339 18277 21513 18278
rect 10003 18245 20478 18249
rect 10003 18191 10013 18245
rect 10067 18191 20478 18245
rect 10003 18185 20478 18191
rect 974 6806 986 6863
rect 1042 6806 1054 6863
rect 974 3503 1054 6806
rect 1203 18155 10224 18157
rect 1203 18151 20350 18155
rect 1203 18097 10151 18151
rect 10205 18097 20350 18151
rect 1203 18093 20350 18097
rect 1203 6555 1267 18093
rect 10141 18091 20350 18093
rect 8501 18057 19310 18063
rect 8501 18003 8511 18057
rect 8565 18003 19310 18057
rect 8501 17999 19310 18003
rect 8677 17967 19160 17969
rect 1375 17963 19160 17967
rect 1375 17909 8690 17963
rect 8744 17909 19160 17963
rect 1194 6502 1204 6555
rect 1265 6502 1275 6555
rect 1203 3602 1267 6502
rect 1375 6398 1454 17909
rect 8677 17905 19160 17909
rect 7045 17873 18136 17877
rect 7045 17819 7055 17873
rect 7109 17819 18136 17873
rect 7045 17814 18136 17819
rect 13091 17813 18136 17814
rect 1578 17784 1652 17785
rect 1578 17783 12725 17784
rect 1578 17778 17962 17783
rect 1578 17724 7183 17778
rect 7237 17724 17962 17778
rect 1578 17720 17962 17724
rect 1369 6340 1379 6398
rect 1449 6340 1459 6398
rect 1375 3730 1454 6340
rect 1578 6248 1652 17720
rect 12998 17719 17962 17720
rect 5595 17691 12728 17692
rect 5595 17687 16968 17691
rect 5595 17633 5602 17687
rect 5656 17633 16968 17687
rect 5595 17628 16968 17633
rect 13174 17627 16968 17628
rect 1775 17597 12728 17598
rect 1775 17592 16791 17597
rect 1775 17543 5733 17592
rect 1571 6190 1581 6248
rect 1649 6190 1659 6248
rect 1578 3849 1652 6190
rect 1775 6085 1839 17543
rect 5724 17538 5733 17543
rect 5787 17538 16791 17592
rect 5724 17534 16791 17538
rect 13174 17533 16791 17534
rect 4157 17505 11596 17506
rect 4157 17501 15800 17505
rect 4147 17447 4157 17501
rect 4211 17447 15800 17501
rect 4157 17442 15800 17447
rect 13172 17441 15800 17442
rect 2014 17412 2540 17413
rect 2005 17411 11596 17412
rect 2005 17408 15644 17411
rect 2005 17354 4267 17408
rect 4321 17354 15644 17408
rect 2005 17348 15644 17354
rect 1767 6031 1777 6085
rect 1835 6031 1845 6085
rect 1775 3958 1839 6031
rect 2005 5901 2069 17348
rect 13172 17347 15644 17348
rect 2547 17255 14632 17319
rect 2547 16182 2610 17255
rect 2405 16181 2610 16182
rect 2405 16122 2415 16181
rect 2486 16122 2610 16181
rect 2547 15906 2610 16122
rect 2786 17161 14487 17225
rect 2786 16962 2849 17161
rect 2786 16107 2850 16962
rect 3214 16837 3350 16857
rect 3214 16775 3250 16837
rect 3310 16775 3350 16837
rect 3214 16747 3350 16775
rect 4662 16837 4798 16857
rect 4662 16775 4698 16837
rect 4758 16775 4798 16837
rect 4662 16747 4798 16775
rect 6160 16839 6296 16859
rect 6160 16777 6196 16839
rect 6256 16777 6296 16839
rect 6160 16749 6296 16777
rect 7608 16839 7744 16859
rect 7608 16777 7644 16839
rect 7704 16777 7744 16839
rect 7608 16749 7744 16777
rect 9128 16837 9264 16857
rect 9128 16775 9164 16837
rect 9224 16775 9264 16837
rect 2910 16717 3887 16747
rect 2910 16611 2942 16717
rect 3146 16611 3178 16717
rect 3382 16611 3414 16717
rect 3618 16611 3650 16717
rect 3853 16611 3887 16717
rect 4358 16717 5335 16747
rect 4358 16611 4390 16717
rect 4594 16611 4626 16717
rect 4830 16611 4862 16717
rect 5066 16611 5098 16717
rect 5301 16611 5335 16717
rect 5856 16719 6833 16749
rect 5856 16613 5888 16719
rect 6092 16613 6124 16719
rect 6328 16613 6360 16719
rect 6564 16613 6596 16719
rect 6799 16613 6833 16719
rect 7304 16719 8281 16749
rect 9128 16747 9264 16775
rect 10576 16837 10712 16857
rect 10576 16775 10612 16837
rect 10672 16775 10712 16837
rect 10576 16747 10712 16775
rect 12074 16839 12210 16859
rect 12074 16777 12110 16839
rect 12170 16777 12210 16839
rect 12074 16749 12210 16777
rect 13522 16839 13658 16859
rect 13522 16777 13558 16839
rect 13618 16777 13658 16839
rect 13522 16749 13658 16777
rect 14432 16797 14487 17161
rect 14568 17070 14632 17255
rect 14532 16968 14632 17070
rect 14532 16934 14582 16968
rect 14616 16934 14632 16968
rect 15218 17044 15322 17050
rect 15218 16972 15230 17044
rect 15310 16972 15322 17044
rect 15218 16966 15322 16972
rect 14532 16908 14632 16934
rect 15253 16910 15288 16966
rect 14532 16860 14632 16880
rect 14532 16826 14582 16860
rect 14616 16826 14632 16860
rect 14532 16797 14632 16826
rect 14790 16869 15060 16897
rect 14790 16808 14824 16869
rect 15026 16808 15060 16869
rect 15144 16869 15414 16910
rect 15144 16808 15178 16869
rect 15380 16808 15414 16869
rect 15580 16880 15644 17347
rect 15736 17070 15800 17441
rect 15700 16968 15800 17070
rect 15700 16934 15750 16968
rect 15784 16934 15800 16968
rect 16386 17044 16490 17050
rect 16386 16972 16398 17044
rect 16478 16972 16490 17044
rect 16386 16966 16490 16972
rect 15700 16908 15800 16934
rect 16421 16910 16456 16966
rect 15580 16860 15800 16880
rect 15580 16826 15750 16860
rect 15784 16826 15800 16860
rect 15580 16816 15800 16826
rect 7304 16613 7336 16719
rect 7540 16613 7572 16719
rect 7776 16613 7808 16719
rect 8012 16613 8044 16719
rect 8247 16613 8281 16719
rect 8824 16717 9801 16747
rect 2903 16599 2949 16611
rect 2903 16423 2909 16599
rect 2943 16423 2949 16599
rect 2903 16411 2949 16423
rect 3021 16599 3067 16611
rect 3021 16423 3027 16599
rect 3061 16423 3067 16599
rect 3021 16411 3067 16423
rect 3139 16599 3185 16611
rect 3139 16423 3145 16599
rect 3179 16423 3185 16599
rect 3139 16411 3185 16423
rect 3257 16599 3303 16611
rect 3257 16423 3263 16599
rect 3297 16423 3303 16599
rect 3257 16411 3303 16423
rect 3375 16599 3421 16611
rect 3375 16423 3381 16599
rect 3415 16423 3421 16599
rect 3375 16411 3421 16423
rect 3493 16599 3539 16611
rect 3493 16423 3499 16599
rect 3533 16423 3539 16599
rect 3493 16411 3539 16423
rect 3611 16599 3657 16611
rect 3611 16423 3617 16599
rect 3651 16423 3657 16599
rect 3611 16411 3657 16423
rect 3729 16599 3775 16611
rect 3729 16423 3735 16599
rect 3769 16423 3775 16599
rect 3729 16411 3775 16423
rect 3847 16599 3893 16611
rect 3847 16423 3853 16599
rect 3887 16423 3893 16599
rect 3847 16411 3893 16423
rect 3965 16599 4011 16611
rect 3965 16423 3971 16599
rect 4005 16423 4011 16599
rect 3965 16411 4011 16423
rect 4351 16599 4397 16611
rect 4351 16423 4357 16599
rect 4391 16423 4397 16599
rect 4351 16411 4397 16423
rect 4469 16599 4515 16611
rect 4469 16423 4475 16599
rect 4509 16423 4515 16599
rect 4469 16411 4515 16423
rect 4587 16599 4633 16611
rect 4587 16423 4593 16599
rect 4627 16423 4633 16599
rect 4587 16411 4633 16423
rect 4705 16599 4751 16611
rect 4705 16423 4711 16599
rect 4745 16423 4751 16599
rect 4705 16411 4751 16423
rect 4823 16599 4869 16611
rect 4823 16423 4829 16599
rect 4863 16423 4869 16599
rect 4823 16411 4869 16423
rect 4941 16599 4987 16611
rect 4941 16423 4947 16599
rect 4981 16423 4987 16599
rect 4941 16411 4987 16423
rect 5059 16599 5105 16611
rect 5059 16423 5065 16599
rect 5099 16423 5105 16599
rect 5059 16411 5105 16423
rect 5177 16599 5223 16611
rect 5177 16423 5183 16599
rect 5217 16423 5223 16599
rect 5177 16411 5223 16423
rect 5295 16599 5341 16611
rect 5295 16423 5301 16599
rect 5335 16423 5341 16599
rect 5295 16411 5341 16423
rect 5413 16599 5459 16611
rect 5413 16423 5419 16599
rect 5453 16423 5459 16599
rect 5413 16411 5459 16423
rect 5849 16601 5895 16613
rect 5849 16425 5855 16601
rect 5889 16425 5895 16601
rect 5849 16413 5895 16425
rect 5967 16601 6013 16613
rect 5967 16425 5973 16601
rect 6007 16425 6013 16601
rect 5967 16413 6013 16425
rect 6085 16601 6131 16613
rect 6085 16425 6091 16601
rect 6125 16425 6131 16601
rect 6085 16413 6131 16425
rect 6203 16601 6249 16613
rect 6203 16425 6209 16601
rect 6243 16425 6249 16601
rect 6203 16413 6249 16425
rect 6321 16601 6367 16613
rect 6321 16425 6327 16601
rect 6361 16425 6367 16601
rect 6321 16413 6367 16425
rect 6439 16601 6485 16613
rect 6439 16425 6445 16601
rect 6479 16425 6485 16601
rect 6439 16413 6485 16425
rect 6557 16601 6603 16613
rect 6557 16425 6563 16601
rect 6597 16425 6603 16601
rect 6557 16413 6603 16425
rect 6675 16601 6721 16613
rect 6675 16425 6681 16601
rect 6715 16425 6721 16601
rect 6675 16413 6721 16425
rect 6793 16601 6839 16613
rect 6793 16425 6799 16601
rect 6833 16425 6839 16601
rect 6793 16413 6839 16425
rect 6911 16601 6957 16613
rect 6911 16425 6917 16601
rect 6951 16425 6957 16601
rect 6911 16413 6957 16425
rect 7297 16601 7343 16613
rect 7297 16425 7303 16601
rect 7337 16425 7343 16601
rect 7297 16413 7343 16425
rect 7415 16601 7461 16613
rect 7415 16425 7421 16601
rect 7455 16425 7461 16601
rect 7415 16413 7461 16425
rect 7533 16601 7579 16613
rect 7533 16425 7539 16601
rect 7573 16425 7579 16601
rect 7533 16413 7579 16425
rect 7651 16601 7697 16613
rect 7651 16425 7657 16601
rect 7691 16425 7697 16601
rect 7651 16413 7697 16425
rect 7769 16601 7815 16613
rect 7769 16425 7775 16601
rect 7809 16425 7815 16601
rect 7769 16413 7815 16425
rect 7887 16601 7933 16613
rect 7887 16425 7893 16601
rect 7927 16425 7933 16601
rect 7887 16413 7933 16425
rect 8005 16601 8051 16613
rect 8005 16425 8011 16601
rect 8045 16425 8051 16601
rect 8005 16413 8051 16425
rect 8123 16601 8169 16613
rect 8123 16425 8129 16601
rect 8163 16425 8169 16601
rect 8123 16413 8169 16425
rect 8241 16601 8287 16613
rect 8241 16425 8247 16601
rect 8281 16425 8287 16601
rect 8241 16413 8287 16425
rect 8359 16601 8405 16613
rect 8824 16611 8856 16717
rect 9060 16611 9092 16717
rect 9296 16611 9328 16717
rect 9532 16611 9564 16717
rect 9767 16611 9801 16717
rect 10272 16717 11249 16747
rect 10272 16611 10304 16717
rect 10508 16611 10540 16717
rect 10744 16611 10776 16717
rect 10980 16611 11012 16717
rect 11215 16611 11249 16717
rect 11770 16719 12747 16749
rect 11770 16613 11802 16719
rect 12006 16613 12038 16719
rect 12242 16613 12274 16719
rect 12478 16613 12510 16719
rect 12713 16613 12747 16719
rect 13218 16719 14195 16749
rect 14432 16728 14632 16797
rect 14666 16796 14712 16808
rect 13218 16613 13250 16719
rect 13454 16613 13486 16719
rect 13690 16613 13722 16719
rect 13926 16613 13958 16719
rect 14161 16613 14195 16719
rect 8359 16425 8365 16601
rect 8399 16425 8405 16601
rect 8359 16413 8405 16425
rect 8817 16599 8863 16611
rect 8817 16423 8823 16599
rect 8857 16423 8863 16599
rect 3026 16317 3062 16411
rect 3262 16317 3298 16411
rect 3498 16318 3534 16411
rect 3660 16363 3726 16370
rect 3660 16329 3676 16363
rect 3710 16329 3726 16363
rect 3660 16318 3726 16329
rect 3498 16317 3726 16318
rect 3026 16288 3726 16317
rect 3026 16287 3608 16288
rect 3146 16174 3180 16287
rect 3542 16246 3608 16287
rect 3542 16212 3558 16246
rect 3592 16212 3608 16246
rect 3542 16205 3608 16212
rect 3970 16178 4005 16411
rect 4474 16317 4510 16411
rect 4710 16317 4746 16411
rect 4946 16318 4982 16411
rect 5108 16363 5174 16370
rect 5108 16329 5124 16363
rect 5158 16329 5174 16363
rect 5108 16318 5174 16329
rect 4946 16317 5174 16318
rect 4474 16288 5174 16317
rect 4474 16287 5056 16288
rect 3616 16174 4005 16178
rect 4594 16174 4628 16287
rect 4990 16246 5056 16287
rect 4990 16212 5006 16246
rect 5040 16212 5056 16246
rect 4990 16205 5056 16212
rect 5418 16178 5453 16411
rect 5972 16319 6008 16413
rect 6208 16319 6244 16413
rect 6444 16320 6480 16413
rect 6606 16365 6672 16372
rect 6606 16331 6622 16365
rect 6656 16331 6672 16365
rect 6606 16320 6672 16331
rect 6444 16319 6672 16320
rect 5972 16290 6672 16319
rect 5972 16289 6554 16290
rect 5064 16174 5453 16178
rect 6092 16176 6126 16289
rect 6488 16248 6554 16289
rect 6488 16214 6504 16248
rect 6538 16214 6554 16248
rect 6488 16207 6554 16214
rect 6916 16180 6951 16413
rect 7420 16319 7456 16413
rect 7656 16319 7692 16413
rect 7892 16320 7928 16413
rect 8054 16365 8120 16372
rect 8054 16331 8070 16365
rect 8104 16331 8120 16365
rect 8054 16320 8120 16331
rect 7892 16319 8120 16320
rect 7420 16290 8120 16319
rect 7420 16289 8002 16290
rect 6562 16176 6951 16180
rect 7540 16176 7574 16289
rect 7936 16248 8002 16289
rect 7936 16214 7952 16248
rect 7986 16214 8002 16248
rect 7936 16207 8002 16214
rect 8364 16180 8399 16413
rect 8817 16411 8863 16423
rect 8935 16599 8981 16611
rect 8935 16423 8941 16599
rect 8975 16423 8981 16599
rect 8935 16411 8981 16423
rect 9053 16599 9099 16611
rect 9053 16423 9059 16599
rect 9093 16423 9099 16599
rect 9053 16411 9099 16423
rect 9171 16599 9217 16611
rect 9171 16423 9177 16599
rect 9211 16423 9217 16599
rect 9171 16411 9217 16423
rect 9289 16599 9335 16611
rect 9289 16423 9295 16599
rect 9329 16423 9335 16599
rect 9289 16411 9335 16423
rect 9407 16599 9453 16611
rect 9407 16423 9413 16599
rect 9447 16423 9453 16599
rect 9407 16411 9453 16423
rect 9525 16599 9571 16611
rect 9525 16423 9531 16599
rect 9565 16423 9571 16599
rect 9525 16411 9571 16423
rect 9643 16599 9689 16611
rect 9643 16423 9649 16599
rect 9683 16423 9689 16599
rect 9643 16411 9689 16423
rect 9761 16599 9807 16611
rect 9761 16423 9767 16599
rect 9801 16423 9807 16599
rect 9761 16411 9807 16423
rect 9879 16599 9925 16611
rect 9879 16423 9885 16599
rect 9919 16423 9925 16599
rect 9879 16411 9925 16423
rect 10265 16599 10311 16611
rect 10265 16423 10271 16599
rect 10305 16423 10311 16599
rect 10265 16411 10311 16423
rect 10383 16599 10429 16611
rect 10383 16423 10389 16599
rect 10423 16423 10429 16599
rect 10383 16411 10429 16423
rect 10501 16599 10547 16611
rect 10501 16423 10507 16599
rect 10541 16423 10547 16599
rect 10501 16411 10547 16423
rect 10619 16599 10665 16611
rect 10619 16423 10625 16599
rect 10659 16423 10665 16599
rect 10619 16411 10665 16423
rect 10737 16599 10783 16611
rect 10737 16423 10743 16599
rect 10777 16423 10783 16599
rect 10737 16411 10783 16423
rect 10855 16599 10901 16611
rect 10855 16423 10861 16599
rect 10895 16423 10901 16599
rect 10855 16411 10901 16423
rect 10973 16599 11019 16611
rect 10973 16423 10979 16599
rect 11013 16423 11019 16599
rect 10973 16411 11019 16423
rect 11091 16599 11137 16611
rect 11091 16423 11097 16599
rect 11131 16423 11137 16599
rect 11091 16411 11137 16423
rect 11209 16599 11255 16611
rect 11209 16423 11215 16599
rect 11249 16423 11255 16599
rect 11209 16411 11255 16423
rect 11327 16599 11373 16611
rect 11327 16423 11333 16599
rect 11367 16423 11373 16599
rect 11327 16411 11373 16423
rect 11763 16601 11809 16613
rect 11763 16425 11769 16601
rect 11803 16425 11809 16601
rect 11763 16413 11809 16425
rect 11881 16601 11927 16613
rect 11881 16425 11887 16601
rect 11921 16425 11927 16601
rect 11881 16413 11927 16425
rect 11999 16601 12045 16613
rect 11999 16425 12005 16601
rect 12039 16425 12045 16601
rect 11999 16413 12045 16425
rect 12117 16601 12163 16613
rect 12117 16425 12123 16601
rect 12157 16425 12163 16601
rect 12117 16413 12163 16425
rect 12235 16601 12281 16613
rect 12235 16425 12241 16601
rect 12275 16425 12281 16601
rect 12235 16413 12281 16425
rect 12353 16601 12399 16613
rect 12353 16425 12359 16601
rect 12393 16425 12399 16601
rect 12353 16413 12399 16425
rect 12471 16601 12517 16613
rect 12471 16425 12477 16601
rect 12511 16425 12517 16601
rect 12471 16413 12517 16425
rect 12589 16601 12635 16613
rect 12589 16425 12595 16601
rect 12629 16425 12635 16601
rect 12589 16413 12635 16425
rect 12707 16601 12753 16613
rect 12707 16425 12713 16601
rect 12747 16425 12753 16601
rect 12707 16413 12753 16425
rect 12825 16601 12871 16613
rect 12825 16425 12831 16601
rect 12865 16425 12871 16601
rect 12825 16413 12871 16425
rect 13211 16601 13257 16613
rect 13211 16425 13217 16601
rect 13251 16425 13257 16601
rect 13211 16413 13257 16425
rect 13329 16601 13375 16613
rect 13329 16425 13335 16601
rect 13369 16425 13375 16601
rect 13329 16413 13375 16425
rect 13447 16601 13493 16613
rect 13447 16425 13453 16601
rect 13487 16425 13493 16601
rect 13447 16413 13493 16425
rect 13565 16601 13611 16613
rect 13565 16425 13571 16601
rect 13605 16425 13611 16601
rect 13565 16413 13611 16425
rect 13683 16601 13729 16613
rect 13683 16425 13689 16601
rect 13723 16425 13729 16601
rect 13683 16413 13729 16425
rect 13801 16601 13847 16613
rect 13801 16425 13807 16601
rect 13841 16425 13847 16601
rect 13801 16413 13847 16425
rect 13919 16601 13965 16613
rect 13919 16425 13925 16601
rect 13959 16425 13965 16601
rect 13919 16413 13965 16425
rect 14037 16601 14083 16613
rect 14037 16425 14043 16601
rect 14077 16425 14083 16601
rect 14037 16413 14083 16425
rect 14155 16601 14201 16613
rect 14155 16425 14161 16601
rect 14195 16425 14201 16601
rect 14155 16413 14201 16425
rect 14273 16601 14319 16613
rect 14273 16425 14279 16601
rect 14313 16425 14319 16601
rect 14273 16413 14319 16425
rect 14666 16420 14672 16796
rect 14706 16420 14712 16796
rect 8940 16317 8976 16411
rect 9176 16317 9212 16411
rect 9412 16318 9448 16411
rect 9574 16363 9640 16370
rect 9574 16329 9590 16363
rect 9624 16329 9640 16363
rect 9574 16318 9640 16329
rect 9412 16317 9640 16318
rect 8940 16288 9640 16317
rect 8940 16287 9522 16288
rect 8010 16176 8399 16180
rect 2691 16085 2850 16107
rect 2691 16021 2701 16085
rect 2770 16034 2850 16085
rect 3140 16162 3186 16174
rect 2770 16021 3100 16034
rect 2691 16010 3100 16021
rect 2786 15934 3100 16010
rect 2547 15806 2988 15906
rect 2910 15657 2964 15806
rect 3024 15742 3078 15934
rect 3140 15786 3146 16162
rect 3180 15786 3186 16162
rect 3140 15774 3186 15786
rect 3258 16162 3304 16174
rect 3258 15786 3264 16162
rect 3298 15786 3304 16162
rect 3258 15774 3304 15786
rect 3376 16162 3422 16174
rect 3376 15786 3382 16162
rect 3416 15813 3422 16162
rect 3493 16162 3539 16174
rect 3493 15986 3499 16162
rect 3533 15986 3539 16162
rect 3493 15979 3539 15986
rect 3611 16162 4005 16174
rect 3611 15986 3617 16162
rect 3651 16156 4005 16162
rect 4588 16162 4634 16174
rect 3651 16149 4006 16156
rect 3651 15986 3657 16149
rect 3898 16016 4006 16149
rect 3898 15994 4007 16016
rect 3493 15974 3542 15979
rect 3611 15974 3657 15986
rect 3499 15813 3542 15974
rect 3416 15786 3542 15813
rect 3376 15774 3542 15786
rect 3382 15770 3542 15774
rect 3024 15736 3255 15742
rect 3024 15702 3205 15736
rect 3239 15702 3255 15736
rect 3024 15686 3255 15702
rect 3307 15736 3373 15742
rect 3307 15702 3323 15736
rect 3357 15702 3373 15736
rect 3307 15657 3373 15702
rect 2910 15649 3373 15657
rect 2910 15617 3374 15649
rect 3466 15633 3542 15770
rect 3462 15573 3472 15633
rect 3534 15573 3544 15633
rect 3899 15467 4007 15994
rect 4448 16012 4548 16034
rect 4448 15958 4474 16012
rect 4528 15958 4548 16012
rect 4448 15934 4548 15958
rect 4336 15881 4436 15906
rect 4336 15826 4359 15881
rect 4413 15826 4436 15881
rect 4336 15806 4436 15826
rect 4358 15657 4412 15806
rect 4472 15742 4526 15934
rect 4588 15786 4594 16162
rect 4628 15786 4634 16162
rect 4588 15774 4634 15786
rect 4706 16162 4752 16174
rect 4706 15786 4712 16162
rect 4746 15786 4752 16162
rect 4706 15774 4752 15786
rect 4824 16162 4870 16174
rect 4824 15786 4830 16162
rect 4864 15813 4870 16162
rect 4941 16162 4987 16174
rect 4941 15986 4947 16162
rect 4981 15986 4987 16162
rect 4941 15979 4987 15986
rect 5059 16162 5453 16174
rect 5059 15986 5065 16162
rect 5099 16149 5453 16162
rect 5099 15986 5105 16149
rect 4941 15974 4990 15979
rect 5059 15974 5105 15986
rect 4947 15813 4990 15974
rect 4864 15786 4990 15813
rect 4824 15774 4990 15786
rect 4830 15770 4990 15774
rect 4472 15736 4703 15742
rect 4472 15702 4653 15736
rect 4687 15702 4703 15736
rect 4472 15686 4703 15702
rect 4755 15736 4821 15742
rect 4755 15702 4771 15736
rect 4805 15702 4821 15736
rect 4755 15657 4821 15702
rect 4358 15649 4821 15657
rect 4358 15617 4822 15649
rect 4914 15633 4990 15770
rect 4910 15573 4920 15633
rect 4982 15573 4992 15633
rect 3899 15338 4005 15467
rect 2707 15292 4005 15338
rect 5349 15338 5453 16149
rect 6086 16164 6132 16176
rect 5946 16011 6046 16036
rect 5946 15957 5968 16011
rect 6022 15957 6046 16011
rect 5946 15936 6046 15957
rect 5834 15879 5934 15908
rect 5834 15825 5857 15879
rect 5911 15825 5934 15879
rect 5834 15808 5934 15825
rect 5856 15659 5910 15808
rect 5970 15744 6024 15936
rect 6086 15788 6092 16164
rect 6126 15788 6132 16164
rect 6086 15776 6132 15788
rect 6204 16164 6250 16176
rect 6204 15788 6210 16164
rect 6244 15788 6250 16164
rect 6204 15776 6250 15788
rect 6322 16164 6368 16176
rect 6322 15788 6328 16164
rect 6362 15815 6368 16164
rect 6439 16164 6485 16176
rect 6439 15988 6445 16164
rect 6479 15988 6485 16164
rect 6439 15981 6485 15988
rect 6557 16164 6951 16176
rect 6557 15988 6563 16164
rect 6597 16151 6951 16164
rect 6597 15988 6603 16151
rect 6439 15976 6488 15981
rect 6557 15976 6603 15988
rect 6445 15815 6488 15976
rect 6362 15788 6488 15815
rect 6322 15776 6488 15788
rect 6328 15772 6488 15776
rect 5970 15738 6201 15744
rect 5970 15704 6151 15738
rect 6185 15704 6201 15738
rect 5970 15688 6201 15704
rect 6253 15738 6319 15744
rect 6253 15704 6269 15738
rect 6303 15704 6319 15738
rect 6253 15659 6319 15704
rect 5856 15651 6319 15659
rect 5856 15619 6320 15651
rect 6412 15635 6488 15772
rect 6408 15575 6418 15635
rect 6480 15575 6490 15635
rect 2707 15245 4004 15292
rect 5349 15245 5939 15338
rect 2189 14158 2299 14165
rect 2189 14070 2205 14158
rect 2288 14080 2299 14158
rect 2288 14070 2298 14080
rect 2189 11247 2298 14070
rect 2707 14048 2794 15245
rect 3868 15244 4004 15245
rect 4206 15038 4216 15098
rect 4296 15038 4306 15098
rect 4206 14998 4306 15038
rect 3409 14941 5212 14998
rect 3409 14854 3443 14941
rect 4584 14854 4618 14941
rect 3403 14842 3449 14854
rect 3403 14654 3409 14842
rect 2962 14642 3008 14654
rect 2962 14466 2968 14642
rect 3002 14466 3008 14642
rect 2962 14454 3008 14466
rect 3080 14642 3126 14654
rect 3080 14466 3086 14642
rect 3120 14466 3126 14642
rect 3080 14454 3126 14466
rect 3198 14642 3244 14654
rect 3198 14466 3204 14642
rect 3238 14466 3244 14642
rect 3198 14454 3244 14466
rect 3316 14642 3409 14654
rect 3316 14466 3322 14642
rect 3356 14466 3409 14642
rect 3443 14466 3449 14842
rect 3316 14454 3449 14466
rect 3521 14842 3567 14854
rect 3521 14466 3527 14842
rect 3561 14466 3567 14842
rect 3521 14454 3567 14466
rect 3639 14842 3685 14854
rect 3639 14466 3645 14842
rect 3679 14466 3685 14842
rect 3639 14454 3685 14466
rect 3757 14842 3803 14854
rect 3757 14466 3763 14842
rect 3797 14466 3803 14842
rect 3757 14454 3803 14466
rect 3870 14842 3916 14854
rect 3870 14466 3876 14842
rect 3910 14466 3916 14842
rect 3870 14454 3916 14466
rect 3988 14842 4034 14854
rect 3988 14466 3994 14842
rect 4028 14466 4034 14842
rect 3988 14454 4034 14466
rect 4106 14842 4152 14854
rect 4106 14466 4112 14842
rect 4146 14466 4152 14842
rect 4106 14454 4152 14466
rect 4224 14842 4270 14854
rect 4224 14466 4230 14842
rect 4264 14466 4270 14842
rect 4224 14454 4270 14466
rect 4342 14842 4388 14854
rect 4342 14466 4348 14842
rect 4382 14466 4388 14842
rect 4342 14454 4388 14466
rect 4460 14842 4506 14854
rect 4460 14466 4466 14842
rect 4500 14466 4506 14842
rect 4460 14454 4506 14466
rect 4578 14842 4624 14854
rect 4578 14466 4584 14842
rect 4618 14466 4624 14842
rect 4578 14454 4624 14466
rect 4697 14842 4743 14854
rect 4697 14466 4703 14842
rect 4737 14466 4743 14842
rect 4697 14454 4743 14466
rect 4815 14842 4861 14854
rect 4815 14466 4821 14842
rect 4855 14466 4861 14842
rect 4815 14454 4861 14466
rect 4933 14842 4979 14854
rect 4933 14466 4939 14842
rect 4973 14466 4979 14842
rect 4933 14454 4979 14466
rect 5051 14842 5097 14854
rect 5051 14466 5057 14842
rect 5091 14466 5097 14842
rect 5175 14654 5212 14941
rect 5051 14454 5097 14466
rect 5170 14642 5216 14654
rect 5170 14466 5176 14642
rect 5210 14466 5216 14642
rect 5170 14454 5216 14466
rect 5288 14642 5334 14654
rect 5288 14466 5294 14642
rect 5328 14466 5334 14642
rect 5288 14454 5334 14466
rect 5406 14642 5452 14654
rect 5406 14466 5412 14642
rect 5446 14466 5452 14642
rect 5406 14454 5452 14466
rect 5524 14642 5570 14654
rect 5524 14466 5530 14642
rect 5564 14466 5570 14642
rect 5524 14454 5570 14466
rect 2967 14268 3002 14454
rect 3876 14370 3910 14454
rect 5057 14370 5091 14454
rect 3876 14328 5091 14370
rect 5057 14308 5091 14328
rect 5057 14292 5414 14308
rect 2967 14251 4104 14268
rect 2967 14217 4054 14251
rect 4088 14217 4104 14251
rect 5057 14258 5364 14292
rect 5398 14258 5414 14292
rect 5057 14242 5414 14258
rect 2967 14201 4104 14217
rect 2707 14040 2884 14048
rect 2707 13972 2825 14040
rect 2882 13972 2892 14040
rect 2707 13964 2884 13972
rect 2811 13872 2884 13880
rect 2811 13804 2825 13872
rect 2882 13804 2892 13872
rect 2811 13796 2884 13804
rect 2967 13691 3002 14201
rect 3057 14155 3149 14168
rect 3057 14092 3069 14155
rect 3140 14092 3149 14155
rect 3057 14083 3149 14092
rect 4142 14155 4234 14165
rect 4142 14093 4154 14155
rect 4224 14093 4234 14155
rect 4142 14080 4234 14093
rect 5530 14100 5565 14454
rect 4389 14038 4454 14041
rect 4389 14035 4458 14038
rect 4389 13975 4395 14035
rect 4454 13975 4464 14035
rect 4389 13971 4458 13975
rect 4389 13969 4454 13971
rect 5530 13954 5711 14100
rect 5852 14048 5939 15245
rect 6847 15302 6951 16151
rect 7534 16164 7580 16176
rect 7394 16014 7494 16036
rect 7394 15960 7418 16014
rect 7472 15960 7494 16014
rect 7394 15936 7494 15960
rect 7282 15884 7382 15908
rect 7282 15830 7305 15884
rect 7359 15830 7382 15884
rect 7282 15808 7382 15830
rect 7304 15659 7358 15808
rect 7418 15744 7472 15936
rect 7534 15788 7540 16164
rect 7574 15788 7580 16164
rect 7534 15776 7580 15788
rect 7652 16164 7698 16176
rect 7652 15788 7658 16164
rect 7692 15788 7698 16164
rect 7652 15776 7698 15788
rect 7770 16164 7816 16176
rect 7770 15788 7776 16164
rect 7810 15815 7816 16164
rect 7887 16164 7933 16176
rect 7887 15988 7893 16164
rect 7927 15988 7933 16164
rect 7887 15981 7933 15988
rect 8005 16164 8399 16176
rect 9060 16174 9094 16287
rect 9456 16246 9522 16287
rect 9456 16212 9472 16246
rect 9506 16212 9522 16246
rect 9456 16205 9522 16212
rect 9884 16178 9919 16411
rect 10388 16317 10424 16411
rect 10624 16317 10660 16411
rect 10860 16318 10896 16411
rect 11022 16363 11088 16370
rect 11022 16329 11038 16363
rect 11072 16329 11088 16363
rect 11022 16318 11088 16329
rect 10860 16317 11088 16318
rect 10388 16288 11088 16317
rect 10388 16287 10970 16288
rect 9530 16174 9919 16178
rect 10508 16174 10542 16287
rect 10904 16246 10970 16287
rect 10904 16212 10920 16246
rect 10954 16212 10970 16246
rect 10904 16205 10970 16212
rect 11332 16178 11367 16411
rect 11886 16319 11922 16413
rect 12122 16319 12158 16413
rect 12358 16320 12394 16413
rect 12520 16365 12586 16372
rect 12520 16331 12536 16365
rect 12570 16331 12586 16365
rect 12520 16320 12586 16331
rect 12358 16319 12586 16320
rect 11886 16290 12586 16319
rect 11886 16289 12468 16290
rect 10978 16174 11367 16178
rect 12006 16176 12040 16289
rect 12402 16248 12468 16289
rect 12402 16214 12418 16248
rect 12452 16214 12468 16248
rect 12402 16207 12468 16214
rect 12830 16180 12865 16413
rect 13334 16319 13370 16413
rect 13570 16319 13606 16413
rect 13806 16320 13842 16413
rect 13968 16365 14034 16372
rect 13968 16331 13984 16365
rect 14018 16331 14034 16365
rect 13968 16320 14034 16331
rect 13806 16319 14034 16320
rect 13334 16290 14034 16319
rect 13334 16289 13916 16290
rect 12476 16176 12865 16180
rect 13454 16176 13488 16289
rect 13850 16248 13916 16289
rect 13850 16214 13866 16248
rect 13900 16214 13916 16248
rect 13850 16207 13916 16214
rect 14278 16180 14313 16413
rect 14666 16408 14712 16420
rect 14784 16796 14830 16808
rect 14784 16420 14790 16796
rect 14824 16420 14830 16796
rect 14784 16408 14830 16420
rect 14902 16796 14948 16808
rect 14902 16420 14908 16796
rect 14942 16420 14948 16796
rect 14902 16408 14948 16420
rect 15020 16796 15066 16808
rect 15020 16420 15026 16796
rect 15060 16420 15066 16796
rect 15020 16408 15066 16420
rect 15138 16796 15184 16808
rect 15138 16420 15144 16796
rect 15178 16420 15184 16796
rect 15138 16408 15184 16420
rect 15256 16796 15302 16808
rect 15256 16420 15262 16796
rect 15296 16420 15302 16796
rect 15256 16408 15302 16420
rect 15374 16796 15420 16808
rect 15374 16420 15380 16796
rect 15414 16420 15420 16796
rect 15700 16728 15800 16816
rect 15958 16869 16228 16897
rect 15958 16808 15992 16869
rect 16194 16808 16228 16869
rect 16312 16869 16582 16910
rect 16312 16808 16346 16869
rect 16548 16808 16582 16869
rect 16727 16880 16791 17533
rect 16904 17070 16968 17627
rect 16868 16968 16968 17070
rect 16868 16934 16918 16968
rect 16952 16934 16968 16968
rect 17554 17044 17658 17050
rect 17554 16972 17566 17044
rect 17646 16972 17658 17044
rect 17554 16966 17658 16972
rect 16868 16908 16968 16934
rect 17589 16910 17624 16966
rect 16727 16860 16968 16880
rect 16727 16826 16918 16860
rect 16952 16826 16968 16860
rect 16727 16816 16968 16826
rect 15834 16796 15880 16808
rect 15374 16408 15420 16420
rect 15834 16420 15840 16796
rect 15874 16420 15880 16796
rect 15834 16408 15880 16420
rect 15952 16796 15998 16808
rect 15952 16420 15958 16796
rect 15992 16420 15998 16796
rect 15952 16408 15998 16420
rect 16070 16796 16116 16808
rect 16070 16420 16076 16796
rect 16110 16420 16116 16796
rect 16070 16408 16116 16420
rect 16188 16796 16234 16808
rect 16188 16420 16194 16796
rect 16228 16420 16234 16796
rect 16188 16408 16234 16420
rect 16306 16796 16352 16808
rect 16306 16420 16312 16796
rect 16346 16420 16352 16796
rect 16306 16408 16352 16420
rect 16424 16796 16470 16808
rect 16424 16420 16430 16796
rect 16464 16420 16470 16796
rect 16424 16408 16470 16420
rect 16542 16796 16588 16808
rect 16542 16420 16548 16796
rect 16582 16420 16588 16796
rect 16868 16728 16968 16816
rect 17126 16869 17396 16897
rect 17126 16806 17160 16869
rect 17362 16806 17396 16869
rect 17480 16869 17750 16910
rect 17480 16806 17514 16869
rect 17716 16806 17750 16869
rect 17898 16880 17962 17719
rect 18072 17070 18136 17813
rect 18036 16968 18136 17070
rect 18036 16934 18086 16968
rect 18120 16934 18136 16968
rect 18722 17044 18826 17050
rect 18722 16972 18734 17044
rect 18814 16972 18826 17044
rect 18722 16966 18826 16972
rect 18036 16908 18136 16934
rect 18757 16910 18792 16966
rect 17898 16860 18136 16880
rect 17898 16826 18086 16860
rect 18120 16826 18136 16860
rect 17898 16816 18136 16826
rect 17002 16794 17048 16806
rect 16542 16408 16588 16420
rect 17002 16418 17008 16794
rect 17042 16418 17048 16794
rect 14672 16365 14706 16408
rect 14908 16365 14942 16408
rect 14672 16337 14942 16365
rect 15026 16366 15060 16408
rect 15262 16366 15296 16408
rect 15026 16337 15296 16366
rect 14672 16289 14706 16337
rect 14672 16259 14735 16289
rect 13924 16176 14313 16180
rect 8005 15988 8011 16164
rect 8045 16151 8399 16164
rect 8045 15988 8051 16151
rect 7887 15976 7936 15981
rect 8005 15976 8051 15988
rect 7893 15815 7936 15976
rect 7810 15788 7936 15815
rect 7770 15776 7936 15788
rect 7776 15772 7936 15776
rect 7418 15738 7649 15744
rect 7418 15704 7599 15738
rect 7633 15704 7649 15738
rect 7418 15688 7649 15704
rect 7701 15738 7767 15744
rect 7701 15704 7717 15738
rect 7751 15704 7767 15738
rect 7701 15659 7767 15704
rect 7304 15651 7767 15659
rect 7304 15619 7768 15651
rect 7860 15635 7936 15772
rect 7856 15575 7866 15635
rect 7928 15575 7938 15635
rect 8295 15402 8399 16151
rect 9054 16162 9100 16174
rect 8914 16009 9014 16034
rect 8914 15955 8937 16009
rect 8991 15955 9014 16009
rect 8914 15934 9014 15955
rect 8802 15884 8902 15906
rect 8802 15830 8821 15884
rect 8875 15830 8902 15884
rect 8802 15806 8902 15830
rect 8824 15657 8878 15806
rect 8938 15742 8992 15934
rect 9054 15786 9060 16162
rect 9094 15786 9100 16162
rect 9054 15774 9100 15786
rect 9172 16162 9218 16174
rect 9172 15786 9178 16162
rect 9212 15786 9218 16162
rect 9172 15774 9218 15786
rect 9290 16162 9336 16174
rect 9290 15786 9296 16162
rect 9330 15813 9336 16162
rect 9407 16162 9453 16174
rect 9407 15986 9413 16162
rect 9447 15986 9453 16162
rect 9407 15979 9453 15986
rect 9525 16162 9919 16174
rect 9525 15986 9531 16162
rect 9565 16149 9919 16162
rect 9565 15986 9571 16149
rect 9407 15974 9456 15979
rect 9525 15974 9571 15986
rect 9413 15813 9456 15974
rect 9330 15786 9456 15813
rect 9290 15774 9456 15786
rect 9296 15770 9456 15774
rect 8938 15736 9169 15742
rect 8938 15702 9119 15736
rect 9153 15702 9169 15736
rect 8938 15686 9169 15702
rect 9221 15736 9287 15742
rect 9221 15702 9237 15736
rect 9271 15702 9287 15736
rect 9221 15657 9287 15702
rect 8824 15649 9287 15657
rect 8824 15617 9288 15649
rect 9380 15633 9456 15770
rect 9376 15573 9386 15633
rect 9448 15573 9458 15633
rect 9815 15407 9919 16149
rect 10502 16162 10548 16174
rect 10362 16016 10462 16034
rect 10362 15962 10385 16016
rect 10439 15962 10462 16016
rect 10362 15934 10462 15962
rect 10250 15878 10350 15906
rect 10250 15824 10273 15878
rect 10327 15824 10350 15878
rect 10250 15806 10350 15824
rect 10272 15657 10326 15806
rect 10386 15742 10440 15934
rect 10502 15786 10508 16162
rect 10542 15786 10548 16162
rect 10502 15774 10548 15786
rect 10620 16162 10666 16174
rect 10620 15786 10626 16162
rect 10660 15786 10666 16162
rect 10620 15774 10666 15786
rect 10738 16162 10784 16174
rect 10738 15786 10744 16162
rect 10778 15813 10784 16162
rect 10855 16162 10901 16174
rect 10855 15986 10861 16162
rect 10895 15986 10901 16162
rect 10855 15979 10901 15986
rect 10973 16162 11367 16174
rect 10973 15986 10979 16162
rect 11013 16149 11367 16162
rect 11013 15986 11019 16149
rect 10855 15974 10904 15979
rect 10973 15974 11019 15986
rect 10861 15813 10904 15974
rect 10778 15786 10904 15813
rect 10738 15774 10904 15786
rect 10744 15770 10904 15774
rect 10386 15736 10617 15742
rect 10386 15702 10567 15736
rect 10601 15702 10617 15736
rect 10386 15686 10617 15702
rect 10669 15736 10735 15742
rect 10669 15702 10685 15736
rect 10719 15702 10735 15736
rect 10669 15657 10735 15702
rect 10272 15649 10735 15657
rect 10272 15617 10736 15649
rect 10828 15633 10904 15770
rect 10824 15573 10834 15633
rect 10896 15573 10906 15633
rect 11263 15496 11367 16149
rect 12000 16164 12046 16176
rect 11860 16014 11960 16036
rect 11860 15960 11882 16014
rect 11936 15960 11960 16014
rect 11860 15936 11960 15960
rect 11748 15884 11848 15908
rect 11748 15830 11770 15884
rect 11824 15830 11848 15884
rect 11748 15808 11848 15830
rect 11770 15659 11824 15808
rect 11884 15744 11938 15936
rect 12000 15788 12006 16164
rect 12040 15788 12046 16164
rect 12000 15776 12046 15788
rect 12118 16164 12164 16176
rect 12118 15788 12124 16164
rect 12158 15788 12164 16164
rect 12118 15776 12164 15788
rect 12236 16164 12282 16176
rect 12236 15788 12242 16164
rect 12276 15815 12282 16164
rect 12353 16164 12399 16176
rect 12353 15988 12359 16164
rect 12393 15988 12399 16164
rect 12353 15981 12399 15988
rect 12471 16164 12865 16176
rect 12471 15988 12477 16164
rect 12511 16151 12865 16164
rect 12511 15988 12517 16151
rect 12353 15976 12402 15981
rect 12471 15976 12517 15988
rect 12359 15815 12402 15976
rect 12276 15788 12402 15815
rect 12236 15776 12402 15788
rect 12242 15772 12402 15776
rect 11884 15738 12115 15744
rect 11884 15704 12065 15738
rect 12099 15704 12115 15738
rect 11884 15688 12115 15704
rect 12167 15738 12233 15744
rect 12167 15704 12183 15738
rect 12217 15704 12233 15738
rect 12167 15659 12233 15704
rect 11770 15651 12233 15659
rect 11770 15619 12234 15651
rect 12326 15635 12402 15772
rect 12322 15575 12332 15635
rect 12394 15575 12404 15635
rect 11263 15436 12430 15496
rect 12761 15486 12865 16151
rect 13448 16164 13494 16176
rect 13308 16030 13408 16036
rect 13304 15942 13314 16030
rect 13400 15942 13410 16030
rect 13308 15936 13408 15942
rect 13196 15901 13296 15908
rect 13190 15813 13200 15901
rect 13286 15813 13296 15901
rect 13196 15808 13296 15813
rect 13218 15659 13272 15808
rect 13332 15744 13386 15936
rect 13448 15788 13454 16164
rect 13488 15788 13494 16164
rect 13448 15776 13494 15788
rect 13566 16164 13612 16176
rect 13566 15788 13572 16164
rect 13606 15788 13612 16164
rect 13566 15776 13612 15788
rect 13684 16164 13730 16176
rect 13684 15788 13690 16164
rect 13724 15815 13730 16164
rect 13801 16164 13847 16176
rect 13801 15988 13807 16164
rect 13841 15988 13847 16164
rect 13801 15981 13847 15988
rect 13919 16164 14313 16176
rect 13919 15988 13925 16164
rect 13959 16151 14313 16164
rect 13959 15988 13965 16151
rect 13801 15976 13850 15981
rect 13919 15976 13965 15988
rect 13807 15815 13850 15976
rect 13724 15788 13850 15815
rect 13684 15776 13850 15788
rect 13690 15772 13850 15776
rect 13332 15738 13563 15744
rect 13332 15704 13513 15738
rect 13547 15704 13563 15738
rect 13332 15688 13563 15704
rect 13615 15738 13681 15744
rect 13615 15704 13631 15738
rect 13665 15704 13681 15738
rect 13615 15659 13681 15704
rect 13218 15651 13681 15659
rect 13218 15619 13682 15651
rect 13774 15635 13850 15772
rect 13770 15575 13780 15635
rect 13842 15575 13852 15635
rect 14209 15562 14313 16151
rect 14700 16167 14735 16259
rect 15380 16224 15414 16408
rect 15840 16365 15874 16408
rect 16076 16365 16110 16408
rect 15840 16337 16110 16365
rect 16194 16366 16228 16408
rect 16430 16366 16464 16408
rect 16194 16337 16464 16366
rect 15840 16289 15874 16337
rect 15840 16259 15903 16289
rect 15380 16170 15489 16224
rect 14700 16131 14927 16167
rect 14700 16022 14735 16131
rect 14861 16097 14927 16131
rect 14861 16063 14877 16097
rect 14911 16063 14927 16097
rect 14861 16057 14927 16063
rect 14576 16010 14622 16022
rect 14576 15834 14582 16010
rect 14616 15834 14622 16010
rect 14576 15822 14622 15834
rect 14694 16010 14740 16022
rect 14694 15834 14700 16010
rect 14734 15834 14740 16010
rect 14694 15822 14740 15834
rect 14812 16010 14858 16022
rect 14812 15834 14818 16010
rect 14852 15834 14858 16010
rect 14812 15822 14858 15834
rect 14930 16010 14976 16022
rect 15338 16018 15371 16049
rect 15455 16018 15489 16170
rect 15868 16167 15903 16259
rect 16548 16224 16582 16408
rect 17002 16406 17048 16418
rect 17120 16794 17166 16806
rect 17120 16418 17126 16794
rect 17160 16418 17166 16794
rect 17120 16406 17166 16418
rect 17238 16794 17284 16806
rect 17238 16418 17244 16794
rect 17278 16418 17284 16794
rect 17238 16406 17284 16418
rect 17356 16794 17402 16806
rect 17356 16418 17362 16794
rect 17396 16418 17402 16794
rect 17356 16406 17402 16418
rect 17474 16794 17520 16806
rect 17474 16418 17480 16794
rect 17514 16418 17520 16794
rect 17474 16406 17520 16418
rect 17592 16794 17638 16806
rect 17592 16418 17598 16794
rect 17632 16418 17638 16794
rect 17592 16406 17638 16418
rect 17710 16794 17756 16806
rect 17710 16418 17716 16794
rect 17750 16418 17756 16794
rect 18036 16728 18136 16816
rect 18294 16869 18564 16897
rect 18294 16808 18328 16869
rect 18530 16808 18564 16869
rect 18648 16869 18918 16910
rect 18648 16808 18682 16869
rect 18884 16808 18918 16869
rect 19096 16882 19160 17905
rect 19246 17072 19310 17999
rect 19210 16970 19310 17072
rect 19210 16936 19260 16970
rect 19294 16936 19310 16970
rect 19896 17046 20000 17052
rect 19896 16974 19908 17046
rect 19988 16974 20000 17046
rect 19896 16968 20000 16974
rect 19210 16910 19310 16936
rect 19931 16912 19966 16968
rect 19096 16862 19310 16882
rect 19096 16828 19260 16862
rect 19294 16828 19310 16862
rect 19096 16818 19310 16828
rect 18170 16796 18216 16808
rect 17710 16406 17756 16418
rect 18170 16420 18176 16796
rect 18210 16420 18216 16796
rect 18170 16408 18216 16420
rect 18288 16796 18334 16808
rect 18288 16420 18294 16796
rect 18328 16420 18334 16796
rect 18288 16408 18334 16420
rect 18406 16796 18452 16808
rect 18406 16420 18412 16796
rect 18446 16420 18452 16796
rect 18406 16408 18452 16420
rect 18524 16796 18570 16808
rect 18524 16420 18530 16796
rect 18564 16420 18570 16796
rect 18524 16408 18570 16420
rect 18642 16796 18688 16808
rect 18642 16420 18648 16796
rect 18682 16420 18688 16796
rect 18642 16408 18688 16420
rect 18760 16796 18806 16808
rect 18760 16420 18766 16796
rect 18800 16420 18806 16796
rect 18760 16408 18806 16420
rect 18878 16796 18924 16808
rect 18878 16420 18884 16796
rect 18918 16420 18924 16796
rect 19210 16730 19310 16818
rect 19468 16871 19738 16899
rect 19468 16810 19502 16871
rect 19704 16810 19738 16871
rect 19822 16871 20092 16912
rect 19822 16810 19856 16871
rect 20058 16810 20092 16871
rect 20286 16882 20350 18091
rect 20378 16970 20478 18185
rect 20378 16936 20428 16970
rect 20462 16936 20478 16970
rect 21064 17046 21168 17052
rect 21064 16974 21076 17046
rect 21156 16974 21168 17046
rect 21064 16968 21168 16974
rect 20378 16910 20478 16936
rect 21099 16912 21134 16968
rect 20286 16862 20478 16882
rect 20286 16828 20428 16862
rect 20462 16828 20478 16862
rect 20286 16818 20478 16828
rect 19344 16798 19390 16810
rect 18878 16408 18924 16420
rect 19344 16422 19350 16798
rect 19384 16422 19390 16798
rect 19344 16410 19390 16422
rect 19462 16798 19508 16810
rect 19462 16422 19468 16798
rect 19502 16422 19508 16798
rect 19462 16410 19508 16422
rect 19580 16798 19626 16810
rect 19580 16422 19586 16798
rect 19620 16422 19626 16798
rect 19580 16410 19626 16422
rect 19698 16798 19744 16810
rect 19698 16422 19704 16798
rect 19738 16422 19744 16798
rect 19698 16410 19744 16422
rect 19816 16798 19862 16810
rect 19816 16422 19822 16798
rect 19856 16422 19862 16798
rect 19816 16410 19862 16422
rect 19934 16798 19980 16810
rect 19934 16422 19940 16798
rect 19974 16422 19980 16798
rect 19934 16410 19980 16422
rect 20052 16798 20098 16810
rect 20052 16422 20058 16798
rect 20092 16422 20098 16798
rect 20378 16730 20478 16818
rect 20636 16871 20906 16899
rect 20636 16808 20670 16871
rect 20872 16808 20906 16871
rect 20990 16871 21260 16912
rect 20990 16808 21024 16871
rect 21226 16808 21260 16871
rect 21449 16882 21513 18277
rect 21546 16970 21646 18371
rect 21546 16936 21596 16970
rect 21630 16936 21646 16970
rect 22232 17046 22336 17052
rect 22232 16974 22244 17046
rect 22324 16974 22336 17046
rect 22232 16968 22336 16974
rect 21546 16910 21646 16936
rect 22267 16912 22302 16968
rect 21449 16862 21646 16882
rect 21449 16828 21596 16862
rect 21630 16828 21646 16862
rect 21449 16818 21646 16828
rect 20512 16796 20558 16808
rect 20052 16410 20098 16422
rect 20512 16420 20518 16796
rect 20552 16420 20558 16796
rect 17008 16365 17042 16406
rect 17244 16365 17278 16406
rect 17008 16337 17278 16365
rect 17362 16366 17396 16406
rect 17598 16366 17632 16406
rect 17362 16337 17632 16366
rect 17008 16289 17042 16337
rect 17008 16259 17071 16289
rect 16548 16170 16657 16224
rect 15868 16131 16095 16167
rect 15868 16024 15903 16131
rect 16029 16097 16095 16131
rect 16029 16063 16045 16097
rect 16079 16063 16095 16097
rect 16029 16057 16095 16063
rect 16270 16024 16303 16028
rect 16506 16024 16539 16028
rect 16623 16024 16657 16170
rect 17036 16167 17071 16259
rect 17716 16224 17750 16406
rect 18176 16365 18210 16408
rect 18412 16365 18446 16408
rect 18176 16337 18446 16365
rect 18530 16366 18564 16408
rect 18766 16366 18800 16408
rect 18530 16337 18800 16366
rect 18176 16289 18210 16337
rect 18176 16259 18239 16289
rect 17716 16170 17825 16224
rect 17036 16131 17263 16167
rect 17036 16024 17071 16131
rect 17197 16097 17263 16131
rect 17197 16063 17213 16097
rect 17247 16063 17263 16097
rect 17197 16057 17263 16063
rect 17438 16024 17471 16028
rect 17674 16024 17707 16028
rect 17791 16024 17825 16170
rect 18204 16167 18239 16259
rect 18884 16224 18918 16408
rect 19350 16367 19384 16410
rect 19586 16367 19620 16410
rect 19350 16339 19620 16367
rect 19704 16368 19738 16410
rect 19940 16368 19974 16410
rect 19704 16339 19974 16368
rect 19350 16291 19384 16339
rect 19350 16261 19413 16291
rect 18884 16170 18993 16224
rect 18204 16131 18431 16167
rect 18204 16024 18239 16131
rect 18365 16097 18431 16131
rect 18365 16063 18381 16097
rect 18415 16063 18431 16097
rect 18365 16057 18431 16063
rect 18606 16024 18639 16028
rect 18842 16024 18875 16028
rect 18959 16024 18993 16170
rect 19378 16169 19413 16261
rect 20058 16226 20092 16410
rect 20512 16408 20558 16420
rect 20630 16796 20676 16808
rect 20630 16420 20636 16796
rect 20670 16420 20676 16796
rect 20630 16408 20676 16420
rect 20748 16796 20794 16808
rect 20748 16420 20754 16796
rect 20788 16420 20794 16796
rect 20748 16408 20794 16420
rect 20866 16796 20912 16808
rect 20866 16420 20872 16796
rect 20906 16420 20912 16796
rect 20866 16408 20912 16420
rect 20984 16796 21030 16808
rect 20984 16420 20990 16796
rect 21024 16420 21030 16796
rect 20984 16408 21030 16420
rect 21102 16796 21148 16808
rect 21102 16420 21108 16796
rect 21142 16420 21148 16796
rect 21102 16408 21148 16420
rect 21220 16796 21266 16808
rect 21220 16420 21226 16796
rect 21260 16420 21266 16796
rect 21546 16730 21646 16818
rect 21804 16871 22074 16899
rect 21804 16810 21838 16871
rect 22040 16810 22074 16871
rect 22158 16871 22428 16912
rect 22158 16810 22192 16871
rect 22394 16810 22428 16871
rect 22612 16883 22676 18463
rect 22714 16970 22814 18557
rect 22714 16936 22764 16970
rect 22798 16936 22814 16970
rect 23400 17046 23504 17052
rect 23400 16974 23412 17046
rect 23492 16974 23504 17046
rect 23400 16968 23504 16974
rect 22714 16911 22814 16936
rect 23435 16912 23470 16968
rect 22612 16862 22814 16883
rect 22612 16828 22764 16862
rect 22798 16828 22814 16862
rect 22612 16811 22814 16828
rect 22972 16871 23242 16899
rect 21680 16798 21726 16810
rect 21220 16408 21266 16420
rect 21680 16422 21686 16798
rect 21720 16422 21726 16798
rect 21680 16410 21726 16422
rect 21798 16798 21844 16810
rect 21798 16422 21804 16798
rect 21838 16422 21844 16798
rect 21798 16410 21844 16422
rect 21916 16798 21962 16810
rect 21916 16422 21922 16798
rect 21956 16422 21962 16798
rect 21916 16410 21962 16422
rect 22034 16798 22080 16810
rect 22034 16422 22040 16798
rect 22074 16422 22080 16798
rect 22034 16410 22080 16422
rect 22152 16798 22198 16810
rect 22152 16422 22158 16798
rect 22192 16422 22198 16798
rect 22152 16410 22198 16422
rect 22270 16798 22316 16810
rect 22270 16422 22276 16798
rect 22310 16422 22316 16798
rect 22270 16410 22316 16422
rect 22388 16798 22434 16810
rect 22972 16808 23006 16871
rect 23208 16808 23242 16871
rect 23326 16871 23596 16912
rect 23326 16808 23360 16871
rect 23562 16808 23596 16871
rect 22388 16422 22394 16798
rect 22428 16422 22434 16798
rect 22388 16410 22434 16422
rect 22848 16796 22894 16808
rect 22848 16420 22854 16796
rect 22888 16420 22894 16796
rect 20518 16367 20552 16408
rect 20754 16367 20788 16408
rect 20518 16339 20788 16367
rect 20872 16368 20906 16408
rect 21108 16368 21142 16408
rect 20872 16339 21142 16368
rect 20518 16291 20552 16339
rect 20518 16261 20581 16291
rect 20058 16172 20167 16226
rect 19378 16133 19605 16169
rect 19378 16024 19413 16133
rect 19539 16099 19605 16133
rect 19539 16065 19555 16099
rect 19589 16065 19605 16099
rect 19539 16059 19605 16065
rect 14930 15834 14936 16010
rect 14970 15957 14976 16010
rect 15096 16006 15142 16018
rect 15096 15957 15102 16006
rect 14970 15869 15102 15957
rect 14970 15834 14976 15869
rect 14930 15822 14976 15834
rect 15096 15830 15102 15869
rect 15136 15830 15142 16006
rect 14582 15785 14616 15822
rect 14818 15785 14852 15822
rect 15096 15818 15142 15830
rect 15214 16006 15260 16018
rect 15214 15830 15220 16006
rect 15254 15830 15260 16006
rect 15214 15818 15260 15830
rect 15332 16006 15378 16018
rect 15332 15830 15338 16006
rect 15372 15830 15378 16006
rect 15332 15818 15378 15830
rect 15450 16006 15496 16018
rect 15450 15830 15456 16006
rect 15490 15830 15496 16006
rect 15450 15818 15496 15830
rect 15744 16012 15790 16024
rect 15744 15836 15750 16012
rect 15784 15836 15790 16012
rect 15744 15824 15790 15836
rect 15862 16012 15908 16024
rect 15862 15836 15868 16012
rect 15902 15836 15908 16012
rect 15862 15824 15908 15836
rect 15980 16012 16026 16024
rect 15980 15836 15986 16012
rect 16020 15836 16026 16012
rect 15980 15824 16026 15836
rect 16098 16012 16144 16024
rect 16098 15836 16104 16012
rect 16138 15957 16144 16012
rect 16263 16012 16309 16024
rect 16263 15957 16269 16012
rect 16138 15869 16269 15957
rect 16138 15836 16144 15869
rect 16098 15824 16144 15836
rect 16263 15836 16269 15869
rect 16303 15836 16309 16012
rect 16263 15824 16309 15836
rect 16381 16012 16427 16024
rect 16381 15836 16387 16012
rect 16421 15836 16427 16012
rect 16381 15824 16427 15836
rect 16499 16012 16545 16024
rect 16499 15836 16505 16012
rect 16539 15836 16545 16012
rect 16499 15824 16545 15836
rect 16617 16012 16663 16024
rect 16617 15836 16623 16012
rect 16657 15836 16663 16012
rect 16617 15824 16663 15836
rect 16912 16012 16958 16024
rect 16912 15836 16918 16012
rect 16952 15836 16958 16012
rect 16912 15824 16958 15836
rect 17030 16012 17076 16024
rect 17030 15836 17036 16012
rect 17070 15836 17076 16012
rect 17030 15824 17076 15836
rect 17148 16012 17194 16024
rect 17148 15836 17154 16012
rect 17188 15836 17194 16012
rect 17148 15824 17194 15836
rect 17266 16012 17312 16024
rect 17266 15836 17272 16012
rect 17306 15957 17312 16012
rect 17431 16012 17477 16024
rect 17431 15957 17437 16012
rect 17306 15869 17437 15957
rect 17306 15836 17312 15869
rect 17266 15824 17312 15836
rect 17431 15836 17437 15869
rect 17471 15836 17477 16012
rect 17431 15824 17477 15836
rect 17549 16012 17595 16024
rect 17549 15836 17555 16012
rect 17589 15836 17595 16012
rect 17549 15824 17595 15836
rect 17667 16012 17713 16024
rect 17667 15836 17673 16012
rect 17707 15836 17713 16012
rect 17667 15824 17713 15836
rect 17785 16012 17831 16024
rect 17785 15836 17791 16012
rect 17825 15836 17831 16012
rect 17785 15824 17831 15836
rect 18080 16012 18126 16024
rect 18080 15836 18086 16012
rect 18120 15836 18126 16012
rect 18080 15824 18126 15836
rect 18198 16012 18244 16024
rect 18198 15836 18204 16012
rect 18238 15836 18244 16012
rect 18198 15824 18244 15836
rect 18316 16012 18362 16024
rect 18316 15836 18322 16012
rect 18356 15836 18362 16012
rect 18316 15824 18362 15836
rect 18434 16012 18480 16024
rect 18434 15836 18440 16012
rect 18474 15957 18480 16012
rect 18600 16012 18646 16024
rect 18600 15957 18606 16012
rect 18474 15869 18606 15957
rect 18474 15836 18480 15869
rect 18434 15824 18480 15836
rect 18600 15836 18606 15869
rect 18640 15836 18646 16012
rect 18600 15824 18646 15836
rect 18718 16012 18764 16024
rect 18718 15836 18724 16012
rect 18758 15836 18764 16012
rect 18718 15824 18764 15836
rect 18836 16012 18882 16024
rect 18836 15836 18842 16012
rect 18876 15836 18882 16012
rect 18836 15824 18882 15836
rect 18954 16012 19000 16024
rect 18954 15836 18960 16012
rect 18994 15836 19000 16012
rect 18954 15824 19000 15836
rect 19254 16012 19300 16024
rect 19254 15836 19260 16012
rect 19294 15836 19300 16012
rect 19254 15824 19300 15836
rect 19372 16012 19418 16024
rect 19372 15836 19378 16012
rect 19412 15836 19418 16012
rect 19372 15824 19418 15836
rect 19490 16012 19536 16024
rect 19490 15836 19496 16012
rect 19530 15836 19536 16012
rect 19490 15824 19536 15836
rect 19608 16012 19654 16024
rect 19780 16020 19813 16024
rect 20016 16020 20049 16024
rect 20133 16020 20167 16172
rect 20546 16169 20581 16261
rect 21226 16226 21260 16408
rect 21686 16367 21720 16410
rect 21922 16367 21956 16410
rect 21686 16339 21956 16367
rect 22040 16368 22074 16410
rect 22276 16368 22310 16410
rect 22040 16339 22310 16368
rect 21686 16291 21720 16339
rect 21686 16261 21749 16291
rect 21226 16172 21335 16226
rect 20546 16133 20773 16169
rect 20546 16024 20581 16133
rect 20707 16099 20773 16133
rect 20707 16065 20723 16099
rect 20757 16065 20773 16099
rect 20707 16059 20773 16065
rect 19608 15836 19614 16012
rect 19648 15959 19654 16012
rect 19772 16008 19818 16020
rect 19772 15959 19778 16008
rect 19648 15871 19778 15959
rect 19648 15836 19654 15871
rect 19608 15824 19654 15836
rect 19772 15832 19778 15871
rect 19812 15832 19818 16008
rect 14582 15746 14852 15785
rect 15219 15786 15252 15818
rect 15455 15786 15488 15818
rect 15219 15750 15488 15786
rect 15750 15785 15784 15824
rect 15986 15785 16020 15824
rect 15750 15746 16020 15785
rect 16387 15786 16420 15824
rect 16623 15786 16656 15824
rect 16387 15750 16656 15786
rect 16918 15785 16952 15824
rect 17154 15785 17188 15824
rect 16918 15746 17188 15785
rect 17555 15786 17588 15824
rect 17791 15786 17824 15824
rect 17555 15750 17824 15786
rect 18086 15785 18120 15824
rect 18322 15785 18356 15824
rect 18086 15746 18356 15785
rect 18723 15786 18756 15824
rect 18959 15786 18992 15824
rect 18723 15750 18992 15786
rect 19260 15787 19294 15824
rect 19496 15787 19530 15824
rect 19772 15820 19818 15832
rect 19890 16008 19936 16020
rect 19890 15832 19896 16008
rect 19930 15832 19936 16008
rect 19890 15820 19936 15832
rect 20008 16008 20054 16020
rect 20008 15832 20014 16008
rect 20048 15832 20054 16008
rect 20008 15820 20054 15832
rect 20126 16008 20172 16020
rect 20126 15832 20132 16008
rect 20166 15832 20172 16008
rect 20126 15820 20172 15832
rect 20422 16012 20468 16024
rect 20422 15836 20428 16012
rect 20462 15836 20468 16012
rect 20422 15824 20468 15836
rect 20540 16012 20586 16024
rect 20540 15836 20546 16012
rect 20580 15836 20586 16012
rect 20540 15824 20586 15836
rect 20658 16012 20704 16024
rect 20658 15836 20664 16012
rect 20698 15836 20704 16012
rect 20658 15824 20704 15836
rect 20776 16012 20822 16024
rect 20948 16019 20981 16023
rect 21184 16019 21217 16024
rect 21301 16019 21335 16172
rect 21714 16169 21749 16261
rect 22394 16226 22428 16410
rect 22848 16408 22894 16420
rect 22966 16796 23012 16808
rect 22966 16420 22972 16796
rect 23006 16420 23012 16796
rect 22966 16408 23012 16420
rect 23084 16796 23130 16808
rect 23084 16420 23090 16796
rect 23124 16420 23130 16796
rect 23084 16408 23130 16420
rect 23202 16796 23248 16808
rect 23202 16420 23208 16796
rect 23242 16420 23248 16796
rect 23202 16408 23248 16420
rect 23320 16796 23366 16808
rect 23320 16420 23326 16796
rect 23360 16420 23366 16796
rect 23320 16408 23366 16420
rect 23438 16796 23484 16808
rect 23438 16420 23444 16796
rect 23478 16420 23484 16796
rect 23438 16408 23484 16420
rect 23556 16796 23602 16808
rect 23556 16420 23562 16796
rect 23596 16420 23602 16796
rect 23556 16408 23602 16420
rect 22854 16367 22888 16408
rect 23090 16367 23124 16408
rect 22854 16339 23124 16367
rect 23208 16368 23242 16408
rect 23444 16368 23478 16408
rect 23208 16339 23478 16368
rect 22854 16291 22888 16339
rect 22854 16261 22917 16291
rect 22394 16172 22503 16226
rect 21714 16133 21941 16169
rect 21714 16026 21749 16133
rect 21875 16099 21941 16133
rect 21875 16065 21891 16099
rect 21925 16065 21941 16099
rect 21875 16059 21941 16065
rect 20776 15836 20782 16012
rect 20816 15959 20822 16012
rect 20941 16007 20987 16019
rect 20941 15959 20947 16007
rect 20816 15871 20947 15959
rect 20816 15836 20822 15871
rect 20776 15824 20822 15836
rect 20941 15831 20947 15871
rect 20981 15831 20987 16007
rect 19260 15748 19530 15787
rect 19897 15788 19930 15820
rect 20133 15788 20166 15820
rect 19897 15752 20166 15788
rect 20428 15787 20462 15824
rect 20664 15787 20698 15824
rect 20941 15819 20987 15831
rect 21059 16007 21105 16019
rect 21059 15831 21065 16007
rect 21099 15831 21105 16007
rect 21059 15819 21105 15831
rect 21177 16007 21223 16019
rect 21177 15831 21183 16007
rect 21217 15831 21223 16007
rect 21177 15819 21223 15831
rect 21295 16007 21341 16019
rect 21295 15831 21301 16007
rect 21335 15831 21341 16007
rect 21295 15819 21341 15831
rect 21590 16014 21636 16026
rect 21590 15838 21596 16014
rect 21630 15838 21636 16014
rect 21590 15826 21636 15838
rect 21708 16014 21754 16026
rect 21708 15838 21714 16014
rect 21748 15838 21754 16014
rect 21708 15826 21754 15838
rect 21826 16014 21872 16026
rect 21826 15838 21832 16014
rect 21866 15838 21872 16014
rect 21826 15826 21872 15838
rect 21944 16014 21990 16026
rect 22116 16019 22149 16023
rect 22352 16019 22385 16023
rect 22469 16019 22503 16172
rect 22882 16169 22917 16261
rect 23562 16226 23596 16408
rect 23562 16215 23671 16226
rect 23563 16172 23671 16215
rect 22882 16133 23109 16169
rect 22882 16026 22917 16133
rect 23043 16099 23109 16133
rect 23043 16065 23059 16099
rect 23093 16065 23109 16099
rect 23043 16059 23109 16065
rect 21944 15838 21950 16014
rect 21984 15959 21990 16014
rect 22109 16007 22155 16019
rect 22109 15959 22115 16007
rect 21984 15871 22115 15959
rect 21984 15838 21990 15871
rect 21944 15826 21990 15838
rect 22109 15831 22115 15871
rect 22149 15831 22155 16007
rect 20428 15748 20698 15787
rect 21065 15788 21098 15819
rect 21301 15788 21334 15819
rect 21065 15752 21334 15788
rect 21596 15787 21630 15826
rect 21832 15787 21866 15826
rect 22109 15819 22155 15831
rect 22227 16007 22273 16019
rect 22227 15831 22233 16007
rect 22267 15831 22273 16007
rect 22227 15819 22273 15831
rect 22345 16007 22391 16019
rect 22345 15831 22351 16007
rect 22385 15831 22391 16007
rect 22345 15819 22391 15831
rect 22463 16007 22509 16019
rect 22463 15831 22469 16007
rect 22503 15831 22509 16007
rect 22463 15819 22509 15831
rect 22758 16014 22804 16026
rect 22758 15838 22764 16014
rect 22798 15838 22804 16014
rect 22758 15826 22804 15838
rect 22876 16014 22922 16026
rect 22876 15838 22882 16014
rect 22916 15838 22922 16014
rect 22876 15826 22922 15838
rect 22994 16014 23040 16026
rect 22994 15838 23000 16014
rect 23034 15838 23040 16014
rect 22994 15826 23040 15838
rect 23112 16014 23158 16026
rect 23284 16020 23317 16024
rect 23520 16020 23553 16025
rect 23637 16020 23671 16172
rect 23112 15838 23118 16014
rect 23152 15959 23158 16014
rect 23277 16008 23323 16020
rect 23277 15959 23283 16008
rect 23152 15871 23283 15959
rect 23152 15838 23158 15871
rect 23112 15826 23158 15838
rect 23277 15832 23283 15871
rect 23317 15832 23323 16008
rect 21596 15748 21866 15787
rect 22233 15788 22266 15819
rect 22469 15788 22502 15819
rect 22233 15752 22502 15788
rect 22764 15787 22798 15826
rect 23000 15787 23034 15826
rect 23277 15820 23323 15832
rect 23395 16008 23441 16020
rect 23395 15832 23401 16008
rect 23435 15832 23441 16008
rect 23395 15820 23441 15832
rect 23513 16008 23559 16020
rect 23513 15832 23519 16008
rect 23553 15832 23559 16008
rect 23513 15820 23559 15832
rect 23631 16008 23677 16020
rect 23631 15832 23637 16008
rect 23671 15832 23677 16008
rect 23631 15820 23677 15832
rect 22764 15748 23034 15787
rect 23401 15788 23434 15820
rect 23637 15788 23670 15820
rect 23401 15752 23670 15788
rect 14782 15718 14816 15746
rect 15950 15718 15984 15746
rect 17118 15718 17152 15746
rect 18286 15718 18320 15746
rect 19460 15720 19494 15748
rect 20628 15720 20662 15748
rect 21796 15720 21830 15748
rect 22964 15720 22998 15748
rect 14760 15706 14838 15718
rect 14760 15636 14766 15706
rect 14832 15636 14838 15706
rect 14760 15624 14838 15636
rect 15928 15706 16006 15718
rect 15928 15636 15934 15706
rect 16000 15636 16006 15706
rect 15928 15624 16006 15636
rect 17096 15706 17174 15718
rect 17096 15636 17102 15706
rect 17168 15636 17174 15706
rect 17096 15624 17174 15636
rect 18264 15706 18342 15718
rect 18264 15636 18270 15706
rect 18336 15636 18342 15706
rect 18264 15624 18342 15636
rect 19438 15708 19516 15720
rect 19438 15638 19444 15708
rect 19510 15638 19516 15708
rect 19438 15626 19516 15638
rect 20606 15708 20684 15720
rect 20606 15638 20612 15708
rect 20678 15638 20684 15708
rect 20606 15626 20684 15638
rect 21774 15708 21852 15720
rect 21774 15638 21780 15708
rect 21846 15638 21852 15708
rect 21774 15626 21852 15638
rect 22942 15708 23020 15720
rect 22942 15638 22948 15708
rect 23014 15638 23020 15708
rect 22942 15626 23020 15638
rect 14209 15514 15709 15562
rect 15671 15509 15709 15514
rect 12761 15438 15639 15486
rect 12371 15409 12430 15436
rect 15592 15409 15639 15438
rect 15671 15437 18829 15509
rect 8295 15330 9240 15402
rect 9815 15334 12339 15407
rect 12371 15336 15564 15409
rect 15592 15336 18719 15409
rect 9161 15306 9240 15330
rect 12265 15307 12339 15334
rect 15478 15307 15564 15336
rect 18640 15307 18719 15336
rect 18757 15407 18829 15437
rect 18757 15335 21810 15407
rect 21738 15307 21810 15335
rect 6847 15234 9088 15302
rect 9161 15234 12232 15306
rect 12265 15234 15432 15307
rect 15478 15234 18578 15307
rect 18640 15235 21709 15307
rect 21738 15235 24853 15307
rect 7350 15038 7360 15098
rect 7440 15038 7450 15098
rect 7350 14998 7450 15038
rect 6553 14941 8356 14998
rect 6553 14854 6587 14941
rect 7728 14854 7762 14941
rect 6547 14842 6593 14854
rect 6547 14654 6553 14842
rect 6106 14642 6152 14654
rect 6106 14466 6112 14642
rect 6146 14466 6152 14642
rect 6106 14454 6152 14466
rect 6224 14642 6270 14654
rect 6224 14466 6230 14642
rect 6264 14466 6270 14642
rect 6224 14454 6270 14466
rect 6342 14642 6388 14654
rect 6342 14466 6348 14642
rect 6382 14466 6388 14642
rect 6342 14454 6388 14466
rect 6460 14642 6553 14654
rect 6460 14466 6466 14642
rect 6500 14466 6553 14642
rect 6587 14466 6593 14842
rect 6460 14454 6593 14466
rect 6665 14842 6711 14854
rect 6665 14466 6671 14842
rect 6705 14466 6711 14842
rect 6665 14454 6711 14466
rect 6783 14842 6829 14854
rect 6783 14466 6789 14842
rect 6823 14466 6829 14842
rect 6783 14454 6829 14466
rect 6901 14842 6947 14854
rect 6901 14466 6907 14842
rect 6941 14466 6947 14842
rect 6901 14454 6947 14466
rect 7014 14842 7060 14854
rect 7014 14466 7020 14842
rect 7054 14466 7060 14842
rect 7014 14454 7060 14466
rect 7132 14842 7178 14854
rect 7132 14466 7138 14842
rect 7172 14466 7178 14842
rect 7132 14454 7178 14466
rect 7250 14842 7296 14854
rect 7250 14466 7256 14842
rect 7290 14466 7296 14842
rect 7250 14454 7296 14466
rect 7368 14842 7414 14854
rect 7368 14466 7374 14842
rect 7408 14466 7414 14842
rect 7368 14454 7414 14466
rect 7486 14842 7532 14854
rect 7486 14466 7492 14842
rect 7526 14466 7532 14842
rect 7486 14454 7532 14466
rect 7604 14842 7650 14854
rect 7604 14466 7610 14842
rect 7644 14466 7650 14842
rect 7604 14454 7650 14466
rect 7722 14842 7768 14854
rect 7722 14466 7728 14842
rect 7762 14466 7768 14842
rect 7722 14454 7768 14466
rect 7841 14842 7887 14854
rect 7841 14466 7847 14842
rect 7881 14466 7887 14842
rect 7841 14454 7887 14466
rect 7959 14842 8005 14854
rect 7959 14466 7965 14842
rect 7999 14466 8005 14842
rect 7959 14454 8005 14466
rect 8077 14842 8123 14854
rect 8077 14466 8083 14842
rect 8117 14466 8123 14842
rect 8077 14454 8123 14466
rect 8195 14842 8241 14854
rect 8195 14466 8201 14842
rect 8235 14466 8241 14842
rect 8319 14654 8356 14941
rect 8195 14454 8241 14466
rect 8314 14642 8360 14654
rect 8314 14466 8320 14642
rect 8354 14466 8360 14642
rect 8314 14454 8360 14466
rect 8432 14642 8478 14654
rect 8432 14466 8438 14642
rect 8472 14466 8478 14642
rect 8432 14454 8478 14466
rect 8550 14642 8596 14654
rect 8550 14466 8556 14642
rect 8590 14466 8596 14642
rect 8550 14454 8596 14466
rect 8668 14642 8714 14654
rect 8668 14466 8674 14642
rect 8708 14466 8714 14642
rect 8668 14454 8714 14466
rect 6111 14268 6146 14454
rect 7020 14370 7054 14454
rect 8201 14370 8235 14454
rect 7020 14328 8235 14370
rect 8201 14308 8235 14328
rect 8201 14292 8558 14308
rect 6111 14251 7248 14268
rect 6111 14217 7198 14251
rect 7232 14217 7248 14251
rect 8201 14258 8508 14292
rect 8542 14258 8558 14292
rect 8201 14242 8558 14258
rect 6111 14201 7248 14217
rect 5852 14040 6028 14048
rect 5852 13972 5969 14040
rect 6026 13972 6036 14040
rect 5852 13964 6028 13972
rect 4024 13872 4116 13880
rect 4024 13807 4036 13872
rect 4104 13807 4116 13872
rect 4024 13795 4116 13807
rect 5530 13692 5565 13954
rect 2967 13644 4339 13691
rect 4661 13645 5565 13692
rect 3801 13521 3835 13644
rect 4273 13631 4339 13644
rect 4273 13597 4289 13631
rect 4323 13597 4339 13631
rect 4273 13581 4339 13597
rect 4662 13521 4696 13645
rect 3796 13509 3842 13521
rect 3796 13333 3802 13509
rect 3836 13333 3842 13509
rect 3796 13321 3842 13333
rect 3914 13509 4034 13521
rect 3914 13333 3920 13509
rect 3954 13333 3994 13509
rect 3914 13321 3994 13333
rect 3920 12954 3954 13321
rect 3988 13133 3994 13321
rect 4028 13133 4034 13509
rect 3988 13121 4034 13133
rect 4106 13509 4152 13521
rect 4106 13133 4112 13509
rect 4146 13133 4152 13509
rect 4106 13121 4152 13133
rect 4224 13509 4270 13521
rect 4224 13133 4230 13509
rect 4264 13133 4270 13509
rect 4224 13121 4270 13133
rect 4342 13509 4388 13521
rect 4342 13133 4348 13509
rect 4382 13133 4388 13509
rect 4342 13121 4388 13133
rect 4460 13509 4584 13521
rect 4460 13133 4466 13509
rect 4500 13333 4544 13509
rect 4578 13333 4584 13509
rect 4500 13321 4584 13333
rect 4656 13509 4702 13521
rect 4656 13333 4662 13509
rect 4696 13333 4702 13509
rect 4656 13321 4702 13333
rect 4500 13133 4506 13321
rect 4460 13121 4506 13133
rect 4230 13048 4264 13121
rect 4215 13032 4281 13048
rect 4215 12998 4231 13032
rect 4265 12998 4281 13032
rect 4215 12982 4281 12998
rect 4544 12954 4578 13321
rect 3920 12902 4578 12954
rect 4218 12880 4310 12902
rect 4218 12828 4230 12880
rect 4296 12828 4310 12880
rect 4218 12824 4310 12828
rect 5638 12700 5710 13954
rect 5958 13872 6028 13880
rect 5958 13804 5969 13872
rect 6026 13804 6036 13872
rect 5958 13796 6028 13804
rect 6111 13691 6146 14201
rect 6201 14155 6293 14168
rect 6201 14092 6213 14155
rect 6284 14092 6293 14155
rect 6201 14083 6293 14092
rect 7286 14155 7378 14165
rect 7286 14093 7298 14155
rect 7368 14093 7378 14155
rect 7286 14080 7378 14093
rect 8674 14100 8709 14454
rect 7533 14038 7598 14041
rect 7533 14035 7602 14038
rect 7533 13975 7539 14035
rect 7598 13975 7608 14035
rect 7533 13971 7602 13975
rect 7533 13969 7598 13971
rect 8674 13954 8855 14100
rect 9001 14052 9088 15234
rect 10482 15042 10492 15102
rect 10572 15042 10582 15102
rect 10482 15002 10582 15042
rect 9685 14945 11488 15002
rect 9685 14858 9719 14945
rect 10860 14858 10894 14945
rect 9679 14846 9725 14858
rect 9679 14658 9685 14846
rect 9238 14646 9284 14658
rect 9238 14470 9244 14646
rect 9278 14470 9284 14646
rect 9238 14458 9284 14470
rect 9356 14646 9402 14658
rect 9356 14470 9362 14646
rect 9396 14470 9402 14646
rect 9356 14458 9402 14470
rect 9474 14646 9520 14658
rect 9474 14470 9480 14646
rect 9514 14470 9520 14646
rect 9474 14458 9520 14470
rect 9592 14646 9685 14658
rect 9592 14470 9598 14646
rect 9632 14470 9685 14646
rect 9719 14470 9725 14846
rect 9592 14458 9725 14470
rect 9797 14846 9843 14858
rect 9797 14470 9803 14846
rect 9837 14470 9843 14846
rect 9797 14458 9843 14470
rect 9915 14846 9961 14858
rect 9915 14470 9921 14846
rect 9955 14470 9961 14846
rect 9915 14458 9961 14470
rect 10033 14846 10079 14858
rect 10033 14470 10039 14846
rect 10073 14470 10079 14846
rect 10033 14458 10079 14470
rect 10146 14846 10192 14858
rect 10146 14470 10152 14846
rect 10186 14470 10192 14846
rect 10146 14458 10192 14470
rect 10264 14846 10310 14858
rect 10264 14470 10270 14846
rect 10304 14470 10310 14846
rect 10264 14458 10310 14470
rect 10382 14846 10428 14858
rect 10382 14470 10388 14846
rect 10422 14470 10428 14846
rect 10382 14458 10428 14470
rect 10500 14846 10546 14858
rect 10500 14470 10506 14846
rect 10540 14470 10546 14846
rect 10500 14458 10546 14470
rect 10618 14846 10664 14858
rect 10618 14470 10624 14846
rect 10658 14470 10664 14846
rect 10618 14458 10664 14470
rect 10736 14846 10782 14858
rect 10736 14470 10742 14846
rect 10776 14470 10782 14846
rect 10736 14458 10782 14470
rect 10854 14846 10900 14858
rect 10854 14470 10860 14846
rect 10894 14470 10900 14846
rect 10854 14458 10900 14470
rect 10973 14846 11019 14858
rect 10973 14470 10979 14846
rect 11013 14470 11019 14846
rect 10973 14458 11019 14470
rect 11091 14846 11137 14858
rect 11091 14470 11097 14846
rect 11131 14470 11137 14846
rect 11091 14458 11137 14470
rect 11209 14846 11255 14858
rect 11209 14470 11215 14846
rect 11249 14470 11255 14846
rect 11209 14458 11255 14470
rect 11327 14846 11373 14858
rect 11327 14470 11333 14846
rect 11367 14470 11373 14846
rect 11451 14658 11488 14945
rect 11327 14458 11373 14470
rect 11446 14646 11492 14658
rect 11446 14470 11452 14646
rect 11486 14470 11492 14646
rect 11446 14458 11492 14470
rect 11564 14646 11610 14658
rect 11564 14470 11570 14646
rect 11604 14470 11610 14646
rect 11564 14458 11610 14470
rect 11682 14646 11728 14658
rect 11682 14470 11688 14646
rect 11722 14470 11728 14646
rect 11682 14458 11728 14470
rect 11800 14646 11846 14658
rect 11800 14470 11806 14646
rect 11840 14470 11846 14646
rect 11800 14458 11846 14470
rect 9243 14272 9278 14458
rect 10152 14374 10186 14458
rect 11333 14374 11367 14458
rect 10152 14332 11367 14374
rect 11333 14312 11367 14332
rect 11333 14296 11690 14312
rect 9243 14255 10380 14272
rect 9243 14221 10330 14255
rect 10364 14221 10380 14255
rect 11333 14262 11640 14296
rect 11674 14262 11690 14296
rect 11333 14246 11690 14262
rect 9243 14205 10380 14221
rect 9001 14044 9160 14052
rect 9001 13976 9101 14044
rect 9158 13976 9168 14044
rect 9001 13968 9160 13976
rect 7168 13872 7260 13880
rect 7168 13807 7180 13872
rect 7248 13807 7260 13872
rect 7168 13795 7260 13807
rect 8674 13692 8709 13954
rect 6111 13644 7483 13691
rect 7805 13645 8709 13692
rect 6945 13521 6979 13644
rect 7417 13631 7483 13644
rect 7417 13597 7433 13631
rect 7467 13597 7483 13631
rect 7417 13581 7483 13597
rect 7806 13521 7840 13645
rect 6940 13509 6986 13521
rect 6940 13333 6946 13509
rect 6980 13333 6986 13509
rect 6940 13321 6986 13333
rect 7058 13509 7178 13521
rect 7058 13333 7064 13509
rect 7098 13333 7138 13509
rect 7058 13321 7138 13333
rect 7064 12954 7098 13321
rect 7132 13133 7138 13321
rect 7172 13133 7178 13509
rect 7132 13121 7178 13133
rect 7250 13509 7296 13521
rect 7250 13133 7256 13509
rect 7290 13133 7296 13509
rect 7250 13121 7296 13133
rect 7368 13509 7414 13521
rect 7368 13133 7374 13509
rect 7408 13133 7414 13509
rect 7368 13121 7414 13133
rect 7486 13509 7532 13521
rect 7486 13133 7492 13509
rect 7526 13133 7532 13509
rect 7486 13121 7532 13133
rect 7604 13509 7728 13521
rect 7604 13133 7610 13509
rect 7644 13333 7688 13509
rect 7722 13333 7728 13509
rect 7644 13321 7728 13333
rect 7800 13509 7846 13521
rect 7800 13333 7806 13509
rect 7840 13333 7846 13509
rect 7800 13321 7846 13333
rect 7644 13133 7650 13321
rect 7604 13121 7650 13133
rect 7374 13048 7408 13121
rect 7359 13032 7425 13048
rect 7359 12998 7375 13032
rect 7409 12998 7425 13032
rect 7359 12982 7425 12998
rect 7688 12954 7722 13321
rect 7064 12902 7722 12954
rect 7362 12880 7454 12902
rect 7362 12828 7374 12880
rect 7440 12828 7454 12880
rect 7362 12824 7454 12828
rect 8781 12701 8853 13954
rect 9088 13876 9160 13884
rect 9088 13808 9101 13876
rect 9158 13808 9168 13876
rect 9088 13800 9160 13808
rect 9243 13695 9278 14205
rect 9333 14159 9425 14172
rect 9333 14096 9345 14159
rect 9416 14096 9425 14159
rect 9333 14087 9425 14096
rect 10418 14159 10510 14169
rect 10418 14097 10430 14159
rect 10500 14097 10510 14159
rect 10418 14084 10510 14097
rect 11806 14104 11841 14458
rect 10665 14042 10730 14045
rect 10665 14039 10734 14042
rect 10665 13979 10671 14039
rect 10730 13979 10740 14039
rect 10665 13975 10734 13979
rect 10665 13973 10730 13975
rect 11806 13958 11986 14104
rect 12145 14052 12232 15234
rect 13626 15042 13636 15102
rect 13716 15042 13726 15102
rect 13626 15002 13726 15042
rect 12829 14945 14632 15002
rect 12829 14858 12863 14945
rect 14004 14858 14038 14945
rect 12823 14846 12869 14858
rect 12823 14658 12829 14846
rect 12382 14646 12428 14658
rect 12382 14470 12388 14646
rect 12422 14470 12428 14646
rect 12382 14458 12428 14470
rect 12500 14646 12546 14658
rect 12500 14470 12506 14646
rect 12540 14470 12546 14646
rect 12500 14458 12546 14470
rect 12618 14646 12664 14658
rect 12618 14470 12624 14646
rect 12658 14470 12664 14646
rect 12618 14458 12664 14470
rect 12736 14646 12829 14658
rect 12736 14470 12742 14646
rect 12776 14470 12829 14646
rect 12863 14470 12869 14846
rect 12736 14458 12869 14470
rect 12941 14846 12987 14858
rect 12941 14470 12947 14846
rect 12981 14470 12987 14846
rect 12941 14458 12987 14470
rect 13059 14846 13105 14858
rect 13059 14470 13065 14846
rect 13099 14470 13105 14846
rect 13059 14458 13105 14470
rect 13177 14846 13223 14858
rect 13177 14470 13183 14846
rect 13217 14470 13223 14846
rect 13177 14458 13223 14470
rect 13290 14846 13336 14858
rect 13290 14470 13296 14846
rect 13330 14470 13336 14846
rect 13290 14458 13336 14470
rect 13408 14846 13454 14858
rect 13408 14470 13414 14846
rect 13448 14470 13454 14846
rect 13408 14458 13454 14470
rect 13526 14846 13572 14858
rect 13526 14470 13532 14846
rect 13566 14470 13572 14846
rect 13526 14458 13572 14470
rect 13644 14846 13690 14858
rect 13644 14470 13650 14846
rect 13684 14470 13690 14846
rect 13644 14458 13690 14470
rect 13762 14846 13808 14858
rect 13762 14470 13768 14846
rect 13802 14470 13808 14846
rect 13762 14458 13808 14470
rect 13880 14846 13926 14858
rect 13880 14470 13886 14846
rect 13920 14470 13926 14846
rect 13880 14458 13926 14470
rect 13998 14846 14044 14858
rect 13998 14470 14004 14846
rect 14038 14470 14044 14846
rect 13998 14458 14044 14470
rect 14117 14846 14163 14858
rect 14117 14470 14123 14846
rect 14157 14470 14163 14846
rect 14117 14458 14163 14470
rect 14235 14846 14281 14858
rect 14235 14470 14241 14846
rect 14275 14470 14281 14846
rect 14235 14458 14281 14470
rect 14353 14846 14399 14858
rect 14353 14470 14359 14846
rect 14393 14470 14399 14846
rect 14353 14458 14399 14470
rect 14471 14846 14517 14858
rect 14471 14470 14477 14846
rect 14511 14470 14517 14846
rect 14595 14658 14632 14945
rect 14471 14458 14517 14470
rect 14590 14646 14636 14658
rect 14590 14470 14596 14646
rect 14630 14470 14636 14646
rect 14590 14458 14636 14470
rect 14708 14646 14754 14658
rect 14708 14470 14714 14646
rect 14748 14470 14754 14646
rect 14708 14458 14754 14470
rect 14826 14646 14872 14658
rect 14826 14470 14832 14646
rect 14866 14470 14872 14646
rect 14826 14458 14872 14470
rect 14944 14646 14990 14658
rect 14944 14470 14950 14646
rect 14984 14470 14990 14646
rect 14944 14458 14990 14470
rect 12387 14272 12422 14458
rect 13296 14374 13330 14458
rect 14477 14374 14511 14458
rect 13296 14332 14511 14374
rect 14477 14312 14511 14332
rect 14477 14296 14834 14312
rect 12387 14255 13524 14272
rect 12387 14221 13474 14255
rect 13508 14221 13524 14255
rect 14477 14262 14784 14296
rect 14818 14262 14834 14296
rect 14477 14246 14834 14262
rect 12387 14205 13524 14221
rect 12145 14044 12304 14052
rect 12145 13976 12245 14044
rect 12302 13976 12312 14044
rect 12145 13968 12304 13976
rect 10300 13876 10392 13884
rect 10300 13811 10312 13876
rect 10380 13811 10392 13876
rect 10300 13799 10392 13811
rect 11806 13696 11841 13958
rect 9243 13648 10615 13695
rect 10937 13649 11841 13696
rect 10077 13525 10111 13648
rect 10549 13635 10615 13648
rect 10549 13601 10565 13635
rect 10599 13601 10615 13635
rect 10549 13585 10615 13601
rect 10938 13525 10972 13649
rect 10072 13513 10118 13525
rect 10072 13337 10078 13513
rect 10112 13337 10118 13513
rect 10072 13325 10118 13337
rect 10190 13513 10310 13525
rect 10190 13337 10196 13513
rect 10230 13337 10270 13513
rect 10190 13325 10270 13337
rect 10196 12958 10230 13325
rect 10264 13137 10270 13325
rect 10304 13137 10310 13513
rect 10264 13125 10310 13137
rect 10382 13513 10428 13525
rect 10382 13137 10388 13513
rect 10422 13137 10428 13513
rect 10382 13125 10428 13137
rect 10500 13513 10546 13525
rect 10500 13137 10506 13513
rect 10540 13137 10546 13513
rect 10500 13125 10546 13137
rect 10618 13513 10664 13525
rect 10618 13137 10624 13513
rect 10658 13137 10664 13513
rect 10618 13125 10664 13137
rect 10736 13513 10860 13525
rect 10736 13137 10742 13513
rect 10776 13337 10820 13513
rect 10854 13337 10860 13513
rect 10776 13325 10860 13337
rect 10932 13513 10978 13525
rect 10932 13337 10938 13513
rect 10972 13337 10978 13513
rect 10932 13325 10978 13337
rect 10776 13137 10782 13325
rect 10736 13125 10782 13137
rect 10506 13052 10540 13125
rect 10491 13036 10557 13052
rect 10491 13002 10507 13036
rect 10541 13002 10557 13036
rect 10491 12986 10557 13002
rect 10820 12958 10854 13325
rect 10196 12906 10854 12958
rect 10494 12884 10586 12906
rect 10494 12832 10506 12884
rect 10572 12832 10586 12884
rect 10494 12828 10586 12832
rect 11914 12701 11986 13958
rect 12387 13695 12422 14205
rect 12477 14159 12569 14172
rect 12477 14096 12489 14159
rect 12560 14096 12569 14159
rect 12477 14087 12569 14096
rect 13562 14159 13654 14169
rect 13562 14097 13574 14159
rect 13644 14097 13654 14159
rect 13562 14084 13654 14097
rect 14950 14104 14985 14458
rect 13809 14042 13874 14045
rect 13809 14039 13878 14042
rect 13809 13979 13815 14039
rect 13874 13979 13884 14039
rect 13809 13975 13878 13979
rect 13809 13973 13874 13975
rect 14950 13958 15126 14104
rect 15345 14048 15432 15234
rect 16828 15038 16838 15098
rect 16918 15038 16928 15098
rect 16828 14998 16928 15038
rect 16031 14941 17834 14998
rect 16031 14854 16065 14941
rect 17206 14854 17240 14941
rect 16025 14842 16071 14854
rect 16025 14654 16031 14842
rect 15584 14642 15630 14654
rect 15584 14466 15590 14642
rect 15624 14466 15630 14642
rect 15584 14454 15630 14466
rect 15702 14642 15748 14654
rect 15702 14466 15708 14642
rect 15742 14466 15748 14642
rect 15702 14454 15748 14466
rect 15820 14642 15866 14654
rect 15820 14466 15826 14642
rect 15860 14466 15866 14642
rect 15820 14454 15866 14466
rect 15938 14642 16031 14654
rect 15938 14466 15944 14642
rect 15978 14466 16031 14642
rect 16065 14466 16071 14842
rect 15938 14454 16071 14466
rect 16143 14842 16189 14854
rect 16143 14466 16149 14842
rect 16183 14466 16189 14842
rect 16143 14454 16189 14466
rect 16261 14842 16307 14854
rect 16261 14466 16267 14842
rect 16301 14466 16307 14842
rect 16261 14454 16307 14466
rect 16379 14842 16425 14854
rect 16379 14466 16385 14842
rect 16419 14466 16425 14842
rect 16379 14454 16425 14466
rect 16492 14842 16538 14854
rect 16492 14466 16498 14842
rect 16532 14466 16538 14842
rect 16492 14454 16538 14466
rect 16610 14842 16656 14854
rect 16610 14466 16616 14842
rect 16650 14466 16656 14842
rect 16610 14454 16656 14466
rect 16728 14842 16774 14854
rect 16728 14466 16734 14842
rect 16768 14466 16774 14842
rect 16728 14454 16774 14466
rect 16846 14842 16892 14854
rect 16846 14466 16852 14842
rect 16886 14466 16892 14842
rect 16846 14454 16892 14466
rect 16964 14842 17010 14854
rect 16964 14466 16970 14842
rect 17004 14466 17010 14842
rect 16964 14454 17010 14466
rect 17082 14842 17128 14854
rect 17082 14466 17088 14842
rect 17122 14466 17128 14842
rect 17082 14454 17128 14466
rect 17200 14842 17246 14854
rect 17200 14466 17206 14842
rect 17240 14466 17246 14842
rect 17200 14454 17246 14466
rect 17319 14842 17365 14854
rect 17319 14466 17325 14842
rect 17359 14466 17365 14842
rect 17319 14454 17365 14466
rect 17437 14842 17483 14854
rect 17437 14466 17443 14842
rect 17477 14466 17483 14842
rect 17437 14454 17483 14466
rect 17555 14842 17601 14854
rect 17555 14466 17561 14842
rect 17595 14466 17601 14842
rect 17555 14454 17601 14466
rect 17673 14842 17719 14854
rect 17673 14466 17679 14842
rect 17713 14466 17719 14842
rect 17797 14654 17834 14941
rect 17673 14454 17719 14466
rect 17792 14642 17838 14654
rect 17792 14466 17798 14642
rect 17832 14466 17838 14642
rect 17792 14454 17838 14466
rect 17910 14642 17956 14654
rect 17910 14466 17916 14642
rect 17950 14466 17956 14642
rect 17910 14454 17956 14466
rect 18028 14642 18074 14654
rect 18028 14466 18034 14642
rect 18068 14466 18074 14642
rect 18028 14454 18074 14466
rect 18146 14642 18192 14654
rect 18146 14466 18152 14642
rect 18186 14466 18192 14642
rect 18146 14454 18192 14466
rect 15589 14268 15624 14454
rect 16498 14370 16532 14454
rect 17679 14370 17713 14454
rect 16498 14328 17713 14370
rect 17679 14308 17713 14328
rect 17679 14292 18036 14308
rect 15589 14251 16726 14268
rect 15589 14217 16676 14251
rect 16710 14217 16726 14251
rect 17679 14258 17986 14292
rect 18020 14258 18036 14292
rect 17679 14242 18036 14258
rect 15589 14201 16726 14217
rect 15345 14040 15506 14048
rect 15345 13972 15447 14040
rect 15504 13972 15514 14040
rect 15345 13964 15506 13972
rect 14950 13696 14985 13958
rect 12387 13648 13759 13695
rect 14081 13649 14985 13696
rect 13221 13525 13255 13648
rect 13693 13635 13759 13648
rect 13693 13601 13709 13635
rect 13743 13601 13759 13635
rect 13693 13585 13759 13601
rect 14082 13525 14116 13649
rect 13216 13513 13262 13525
rect 13216 13337 13222 13513
rect 13256 13337 13262 13513
rect 13216 13325 13262 13337
rect 13334 13513 13454 13525
rect 13334 13337 13340 13513
rect 13374 13337 13414 13513
rect 13334 13325 13414 13337
rect 13340 12958 13374 13325
rect 13408 13137 13414 13325
rect 13448 13137 13454 13513
rect 13408 13125 13454 13137
rect 13526 13513 13572 13525
rect 13526 13137 13532 13513
rect 13566 13137 13572 13513
rect 13526 13125 13572 13137
rect 13644 13513 13690 13525
rect 13644 13137 13650 13513
rect 13684 13137 13690 13513
rect 13644 13125 13690 13137
rect 13762 13513 13808 13525
rect 13762 13137 13768 13513
rect 13802 13137 13808 13513
rect 13762 13125 13808 13137
rect 13880 13513 14004 13525
rect 13880 13137 13886 13513
rect 13920 13337 13964 13513
rect 13998 13337 14004 13513
rect 13920 13325 14004 13337
rect 14076 13513 14122 13525
rect 14076 13337 14082 13513
rect 14116 13337 14122 13513
rect 14076 13325 14122 13337
rect 13920 13137 13926 13325
rect 13880 13125 13926 13137
rect 13650 13052 13684 13125
rect 13635 13036 13701 13052
rect 13635 13002 13651 13036
rect 13685 13002 13701 13036
rect 13635 12986 13701 13002
rect 13964 12958 13998 13325
rect 13340 12906 13998 12958
rect 13638 12884 13730 12906
rect 13638 12832 13650 12884
rect 13716 12832 13730 12884
rect 13638 12828 13730 12832
rect 15054 12704 15126 13958
rect 15589 13691 15624 14201
rect 15679 14155 15771 14168
rect 15679 14092 15691 14155
rect 15762 14092 15771 14155
rect 15679 14083 15771 14092
rect 16764 14155 16856 14165
rect 16764 14093 16776 14155
rect 16846 14093 16856 14155
rect 16764 14080 16856 14093
rect 18152 14100 18187 14454
rect 17011 14038 17076 14041
rect 17011 14035 17080 14038
rect 17011 13975 17017 14035
rect 17076 13975 17086 14035
rect 17011 13971 17080 13975
rect 17011 13969 17076 13971
rect 18152 13954 18333 14100
rect 18491 14048 18578 15234
rect 19972 15038 19982 15098
rect 20062 15038 20072 15098
rect 19972 14998 20072 15038
rect 19175 14941 20978 14998
rect 19175 14854 19209 14941
rect 20350 14854 20384 14941
rect 19169 14842 19215 14854
rect 19169 14654 19175 14842
rect 18728 14642 18774 14654
rect 18728 14466 18734 14642
rect 18768 14466 18774 14642
rect 18728 14454 18774 14466
rect 18846 14642 18892 14654
rect 18846 14466 18852 14642
rect 18886 14466 18892 14642
rect 18846 14454 18892 14466
rect 18964 14642 19010 14654
rect 18964 14466 18970 14642
rect 19004 14466 19010 14642
rect 18964 14454 19010 14466
rect 19082 14642 19175 14654
rect 19082 14466 19088 14642
rect 19122 14466 19175 14642
rect 19209 14466 19215 14842
rect 19082 14454 19215 14466
rect 19287 14842 19333 14854
rect 19287 14466 19293 14842
rect 19327 14466 19333 14842
rect 19287 14454 19333 14466
rect 19405 14842 19451 14854
rect 19405 14466 19411 14842
rect 19445 14466 19451 14842
rect 19405 14454 19451 14466
rect 19523 14842 19569 14854
rect 19523 14466 19529 14842
rect 19563 14466 19569 14842
rect 19523 14454 19569 14466
rect 19636 14842 19682 14854
rect 19636 14466 19642 14842
rect 19676 14466 19682 14842
rect 19636 14454 19682 14466
rect 19754 14842 19800 14854
rect 19754 14466 19760 14842
rect 19794 14466 19800 14842
rect 19754 14454 19800 14466
rect 19872 14842 19918 14854
rect 19872 14466 19878 14842
rect 19912 14466 19918 14842
rect 19872 14454 19918 14466
rect 19990 14842 20036 14854
rect 19990 14466 19996 14842
rect 20030 14466 20036 14842
rect 19990 14454 20036 14466
rect 20108 14842 20154 14854
rect 20108 14466 20114 14842
rect 20148 14466 20154 14842
rect 20108 14454 20154 14466
rect 20226 14842 20272 14854
rect 20226 14466 20232 14842
rect 20266 14466 20272 14842
rect 20226 14454 20272 14466
rect 20344 14842 20390 14854
rect 20344 14466 20350 14842
rect 20384 14466 20390 14842
rect 20344 14454 20390 14466
rect 20463 14842 20509 14854
rect 20463 14466 20469 14842
rect 20503 14466 20509 14842
rect 20463 14454 20509 14466
rect 20581 14842 20627 14854
rect 20581 14466 20587 14842
rect 20621 14466 20627 14842
rect 20581 14454 20627 14466
rect 20699 14842 20745 14854
rect 20699 14466 20705 14842
rect 20739 14466 20745 14842
rect 20699 14454 20745 14466
rect 20817 14842 20863 14854
rect 20817 14466 20823 14842
rect 20857 14466 20863 14842
rect 20941 14654 20978 14941
rect 20817 14454 20863 14466
rect 20936 14642 20982 14654
rect 20936 14466 20942 14642
rect 20976 14466 20982 14642
rect 20936 14454 20982 14466
rect 21054 14642 21100 14654
rect 21054 14466 21060 14642
rect 21094 14466 21100 14642
rect 21054 14454 21100 14466
rect 21172 14642 21218 14654
rect 21172 14466 21178 14642
rect 21212 14466 21218 14642
rect 21172 14454 21218 14466
rect 21290 14642 21336 14654
rect 21290 14466 21296 14642
rect 21330 14466 21336 14642
rect 21290 14454 21336 14466
rect 18733 14268 18768 14454
rect 19642 14370 19676 14454
rect 20823 14370 20857 14454
rect 19642 14328 20857 14370
rect 20823 14308 20857 14328
rect 20823 14292 21180 14308
rect 18733 14251 19870 14268
rect 18733 14217 19820 14251
rect 19854 14217 19870 14251
rect 20823 14258 21130 14292
rect 21164 14258 21180 14292
rect 20823 14242 21180 14258
rect 18733 14201 19870 14217
rect 18491 14040 18650 14048
rect 18491 13972 18591 14040
rect 18648 13972 18658 14040
rect 18491 13964 18650 13972
rect 18152 13692 18187 13954
rect 15589 13644 16961 13691
rect 17283 13645 18187 13692
rect 16423 13521 16457 13644
rect 16895 13631 16961 13644
rect 16895 13597 16911 13631
rect 16945 13597 16961 13631
rect 16895 13581 16961 13597
rect 17284 13521 17318 13645
rect 16418 13509 16464 13521
rect 16418 13333 16424 13509
rect 16458 13333 16464 13509
rect 16418 13321 16464 13333
rect 16536 13509 16656 13521
rect 16536 13333 16542 13509
rect 16576 13333 16616 13509
rect 16536 13321 16616 13333
rect 16542 12954 16576 13321
rect 16610 13133 16616 13321
rect 16650 13133 16656 13509
rect 16610 13121 16656 13133
rect 16728 13509 16774 13521
rect 16728 13133 16734 13509
rect 16768 13133 16774 13509
rect 16728 13121 16774 13133
rect 16846 13509 16892 13521
rect 16846 13133 16852 13509
rect 16886 13133 16892 13509
rect 16846 13121 16892 13133
rect 16964 13509 17010 13521
rect 16964 13133 16970 13509
rect 17004 13133 17010 13509
rect 16964 13121 17010 13133
rect 17082 13509 17206 13521
rect 17082 13133 17088 13509
rect 17122 13333 17166 13509
rect 17200 13333 17206 13509
rect 17122 13321 17206 13333
rect 17278 13509 17324 13521
rect 17278 13333 17284 13509
rect 17318 13333 17324 13509
rect 17278 13321 17324 13333
rect 17122 13133 17128 13321
rect 17082 13121 17128 13133
rect 16852 13048 16886 13121
rect 16837 13032 16903 13048
rect 16837 12998 16853 13032
rect 16887 12998 16903 13032
rect 16837 12982 16903 12998
rect 17166 12954 17200 13321
rect 16542 12902 17200 12954
rect 16840 12880 16932 12902
rect 16840 12828 16852 12880
rect 16918 12828 16932 12880
rect 16840 12824 16932 12828
rect 18246 12704 18333 13954
rect 18580 13872 18650 13880
rect 18580 13804 18591 13872
rect 18648 13804 18658 13872
rect 18580 13796 18650 13804
rect 18733 13691 18768 14201
rect 18823 14155 18915 14168
rect 18823 14092 18835 14155
rect 18906 14092 18915 14155
rect 18823 14083 18915 14092
rect 19908 14155 20000 14165
rect 19908 14093 19920 14155
rect 19990 14093 20000 14155
rect 19908 14080 20000 14093
rect 21296 14100 21331 14454
rect 20155 14038 20220 14041
rect 20155 14035 20224 14038
rect 20155 13975 20161 14035
rect 20220 13975 20230 14035
rect 20155 13971 20224 13975
rect 20155 13969 20220 13971
rect 21296 13967 21477 14100
rect 21622 14052 21709 15235
rect 23104 15042 23114 15102
rect 23194 15042 23204 15102
rect 23104 15002 23204 15042
rect 22307 14945 24110 15002
rect 22307 14858 22341 14945
rect 23482 14858 23516 14945
rect 22301 14846 22347 14858
rect 22301 14658 22307 14846
rect 21860 14646 21906 14658
rect 21860 14470 21866 14646
rect 21900 14470 21906 14646
rect 21860 14458 21906 14470
rect 21978 14646 22024 14658
rect 21978 14470 21984 14646
rect 22018 14470 22024 14646
rect 21978 14458 22024 14470
rect 22096 14646 22142 14658
rect 22096 14470 22102 14646
rect 22136 14470 22142 14646
rect 22096 14458 22142 14470
rect 22214 14646 22307 14658
rect 22214 14470 22220 14646
rect 22254 14470 22307 14646
rect 22341 14470 22347 14846
rect 22214 14458 22347 14470
rect 22419 14846 22465 14858
rect 22419 14470 22425 14846
rect 22459 14470 22465 14846
rect 22419 14458 22465 14470
rect 22537 14846 22583 14858
rect 22537 14470 22543 14846
rect 22577 14470 22583 14846
rect 22537 14458 22583 14470
rect 22655 14846 22701 14858
rect 22655 14470 22661 14846
rect 22695 14470 22701 14846
rect 22655 14458 22701 14470
rect 22768 14846 22814 14858
rect 22768 14470 22774 14846
rect 22808 14470 22814 14846
rect 22768 14458 22814 14470
rect 22886 14846 22932 14858
rect 22886 14470 22892 14846
rect 22926 14470 22932 14846
rect 22886 14458 22932 14470
rect 23004 14846 23050 14858
rect 23004 14470 23010 14846
rect 23044 14470 23050 14846
rect 23004 14458 23050 14470
rect 23122 14846 23168 14858
rect 23122 14470 23128 14846
rect 23162 14470 23168 14846
rect 23122 14458 23168 14470
rect 23240 14846 23286 14858
rect 23240 14470 23246 14846
rect 23280 14470 23286 14846
rect 23240 14458 23286 14470
rect 23358 14846 23404 14858
rect 23358 14470 23364 14846
rect 23398 14470 23404 14846
rect 23358 14458 23404 14470
rect 23476 14846 23522 14858
rect 23476 14470 23482 14846
rect 23516 14470 23522 14846
rect 23476 14458 23522 14470
rect 23595 14846 23641 14858
rect 23595 14470 23601 14846
rect 23635 14470 23641 14846
rect 23595 14458 23641 14470
rect 23713 14846 23759 14858
rect 23713 14470 23719 14846
rect 23753 14470 23759 14846
rect 23713 14458 23759 14470
rect 23831 14846 23877 14858
rect 23831 14470 23837 14846
rect 23871 14470 23877 14846
rect 23831 14458 23877 14470
rect 23949 14846 23995 14858
rect 23949 14470 23955 14846
rect 23989 14470 23995 14846
rect 24073 14658 24110 14945
rect 23949 14458 23995 14470
rect 24068 14646 24114 14658
rect 24068 14470 24074 14646
rect 24108 14470 24114 14646
rect 24068 14458 24114 14470
rect 24186 14646 24232 14658
rect 24186 14470 24192 14646
rect 24226 14470 24232 14646
rect 24186 14458 24232 14470
rect 24304 14646 24350 14658
rect 24304 14470 24310 14646
rect 24344 14470 24350 14646
rect 24304 14458 24350 14470
rect 24422 14646 24468 14658
rect 24422 14470 24428 14646
rect 24462 14470 24468 14646
rect 24422 14458 24468 14470
rect 21865 14272 21900 14458
rect 22774 14374 22808 14458
rect 23955 14374 23989 14458
rect 22774 14332 23989 14374
rect 23955 14312 23989 14332
rect 23955 14296 24312 14312
rect 21865 14255 23002 14272
rect 21865 14221 22952 14255
rect 22986 14221 23002 14255
rect 23955 14262 24262 14296
rect 24296 14262 24312 14296
rect 23955 14246 24312 14262
rect 21865 14205 23002 14221
rect 21622 14044 21782 14052
rect 21622 13976 21723 14044
rect 21780 13976 21790 14044
rect 21622 13968 21782 13976
rect 21296 13954 21478 13967
rect 19790 13872 19882 13880
rect 19790 13807 19802 13872
rect 19870 13807 19882 13872
rect 19790 13795 19882 13807
rect 21296 13692 21331 13954
rect 18733 13644 20105 13691
rect 20427 13645 21331 13692
rect 19567 13521 19601 13644
rect 20039 13631 20105 13644
rect 20039 13597 20055 13631
rect 20089 13597 20105 13631
rect 20039 13581 20105 13597
rect 20428 13521 20462 13645
rect 19562 13509 19608 13521
rect 19562 13333 19568 13509
rect 19602 13333 19608 13509
rect 19562 13321 19608 13333
rect 19680 13509 19800 13521
rect 19680 13333 19686 13509
rect 19720 13333 19760 13509
rect 19680 13321 19760 13333
rect 19686 12954 19720 13321
rect 19754 13133 19760 13321
rect 19794 13133 19800 13509
rect 19754 13121 19800 13133
rect 19872 13509 19918 13521
rect 19872 13133 19878 13509
rect 19912 13133 19918 13509
rect 19872 13121 19918 13133
rect 19990 13509 20036 13521
rect 19990 13133 19996 13509
rect 20030 13133 20036 13509
rect 19990 13121 20036 13133
rect 20108 13509 20154 13521
rect 20108 13133 20114 13509
rect 20148 13133 20154 13509
rect 20108 13121 20154 13133
rect 20226 13509 20350 13521
rect 20226 13133 20232 13509
rect 20266 13333 20310 13509
rect 20344 13333 20350 13509
rect 20266 13321 20350 13333
rect 20422 13509 20468 13521
rect 20422 13333 20428 13509
rect 20462 13333 20468 13509
rect 20422 13321 20468 13333
rect 20266 13133 20272 13321
rect 20226 13121 20272 13133
rect 19996 13048 20030 13121
rect 19981 13032 20047 13048
rect 19981 12998 19997 13032
rect 20031 12998 20047 13032
rect 19981 12982 20047 12998
rect 20310 12954 20344 13321
rect 19686 12902 20344 12954
rect 19984 12880 20076 12902
rect 19984 12828 19996 12880
rect 20062 12828 20076 12880
rect 19984 12824 20076 12828
rect 21375 12704 21478 13954
rect 21711 13876 21782 13884
rect 21711 13808 21723 13876
rect 21780 13808 21790 13876
rect 21711 13800 21782 13808
rect 21865 13695 21900 14205
rect 21955 14159 22047 14172
rect 21955 14096 21967 14159
rect 22038 14096 22047 14159
rect 21955 14087 22047 14096
rect 23040 14159 23132 14169
rect 23040 14097 23052 14159
rect 23122 14097 23132 14159
rect 23040 14084 23132 14097
rect 24428 14104 24463 14458
rect 23287 14042 23352 14045
rect 23287 14039 23356 14042
rect 23287 13979 23293 14039
rect 23352 13979 23362 14039
rect 23287 13975 23356 13979
rect 23287 13973 23352 13975
rect 24428 13958 24607 14104
rect 24766 14052 24853 15235
rect 26248 15042 26258 15102
rect 26338 15042 26348 15102
rect 26248 15002 26348 15042
rect 25451 14945 27254 15002
rect 25451 14858 25485 14945
rect 26626 14858 26660 14945
rect 25445 14846 25491 14858
rect 25445 14658 25451 14846
rect 25004 14646 25050 14658
rect 25004 14470 25010 14646
rect 25044 14470 25050 14646
rect 25004 14458 25050 14470
rect 25122 14646 25168 14658
rect 25122 14470 25128 14646
rect 25162 14470 25168 14646
rect 25122 14458 25168 14470
rect 25240 14646 25286 14658
rect 25240 14470 25246 14646
rect 25280 14470 25286 14646
rect 25240 14458 25286 14470
rect 25358 14646 25451 14658
rect 25358 14470 25364 14646
rect 25398 14470 25451 14646
rect 25485 14470 25491 14846
rect 25358 14458 25491 14470
rect 25563 14846 25609 14858
rect 25563 14470 25569 14846
rect 25603 14470 25609 14846
rect 25563 14458 25609 14470
rect 25681 14846 25727 14858
rect 25681 14470 25687 14846
rect 25721 14470 25727 14846
rect 25681 14458 25727 14470
rect 25799 14846 25845 14858
rect 25799 14470 25805 14846
rect 25839 14470 25845 14846
rect 25799 14458 25845 14470
rect 25912 14846 25958 14858
rect 25912 14470 25918 14846
rect 25952 14470 25958 14846
rect 25912 14458 25958 14470
rect 26030 14846 26076 14858
rect 26030 14470 26036 14846
rect 26070 14470 26076 14846
rect 26030 14458 26076 14470
rect 26148 14846 26194 14858
rect 26148 14470 26154 14846
rect 26188 14470 26194 14846
rect 26148 14458 26194 14470
rect 26266 14846 26312 14858
rect 26266 14470 26272 14846
rect 26306 14470 26312 14846
rect 26266 14458 26312 14470
rect 26384 14846 26430 14858
rect 26384 14470 26390 14846
rect 26424 14470 26430 14846
rect 26384 14458 26430 14470
rect 26502 14846 26548 14858
rect 26502 14470 26508 14846
rect 26542 14470 26548 14846
rect 26502 14458 26548 14470
rect 26620 14846 26666 14858
rect 26620 14470 26626 14846
rect 26660 14470 26666 14846
rect 26620 14458 26666 14470
rect 26739 14846 26785 14858
rect 26739 14470 26745 14846
rect 26779 14470 26785 14846
rect 26739 14458 26785 14470
rect 26857 14846 26903 14858
rect 26857 14470 26863 14846
rect 26897 14470 26903 14846
rect 26857 14458 26903 14470
rect 26975 14846 27021 14858
rect 26975 14470 26981 14846
rect 27015 14470 27021 14846
rect 26975 14458 27021 14470
rect 27093 14846 27139 14858
rect 27093 14470 27099 14846
rect 27133 14470 27139 14846
rect 27217 14658 27254 14945
rect 27093 14458 27139 14470
rect 27212 14646 27258 14658
rect 27212 14470 27218 14646
rect 27252 14470 27258 14646
rect 27212 14458 27258 14470
rect 27330 14646 27376 14658
rect 27330 14470 27336 14646
rect 27370 14470 27376 14646
rect 27330 14458 27376 14470
rect 27448 14646 27494 14658
rect 27448 14470 27454 14646
rect 27488 14470 27494 14646
rect 27448 14458 27494 14470
rect 27566 14646 27612 14658
rect 27566 14470 27572 14646
rect 27606 14470 27612 14646
rect 27566 14458 27612 14470
rect 25009 14272 25044 14458
rect 25918 14374 25952 14458
rect 27099 14374 27133 14458
rect 25918 14332 27133 14374
rect 27099 14312 27133 14332
rect 27099 14296 27456 14312
rect 25009 14255 26146 14272
rect 25009 14221 26096 14255
rect 26130 14221 26146 14255
rect 27099 14262 27406 14296
rect 27440 14262 27456 14296
rect 27099 14246 27456 14262
rect 25009 14205 26146 14221
rect 24766 14044 24926 14052
rect 24766 13976 24867 14044
rect 24924 13976 24934 14044
rect 24766 13968 24926 13976
rect 22922 13876 23014 13884
rect 22922 13811 22934 13876
rect 23002 13811 23014 13876
rect 22922 13799 23014 13811
rect 24428 13696 24463 13958
rect 21865 13648 23237 13695
rect 23559 13649 24463 13696
rect 22699 13525 22733 13648
rect 23171 13635 23237 13648
rect 23171 13601 23187 13635
rect 23221 13601 23237 13635
rect 23171 13585 23237 13601
rect 23560 13525 23594 13649
rect 22694 13513 22740 13525
rect 22694 13337 22700 13513
rect 22734 13337 22740 13513
rect 22694 13325 22740 13337
rect 22812 13513 22932 13525
rect 22812 13337 22818 13513
rect 22852 13337 22892 13513
rect 22812 13325 22892 13337
rect 22818 12958 22852 13325
rect 22886 13137 22892 13325
rect 22926 13137 22932 13513
rect 22886 13125 22932 13137
rect 23004 13513 23050 13525
rect 23004 13137 23010 13513
rect 23044 13137 23050 13513
rect 23004 13125 23050 13137
rect 23122 13513 23168 13525
rect 23122 13137 23128 13513
rect 23162 13137 23168 13513
rect 23122 13125 23168 13137
rect 23240 13513 23286 13525
rect 23240 13137 23246 13513
rect 23280 13137 23286 13513
rect 23240 13125 23286 13137
rect 23358 13513 23482 13525
rect 23358 13137 23364 13513
rect 23398 13337 23442 13513
rect 23476 13337 23482 13513
rect 23398 13325 23482 13337
rect 23554 13513 23600 13525
rect 23554 13337 23560 13513
rect 23594 13337 23600 13513
rect 23554 13325 23600 13337
rect 23398 13137 23404 13325
rect 23358 13125 23404 13137
rect 23128 13052 23162 13125
rect 23113 13036 23179 13052
rect 23113 13002 23129 13036
rect 23163 13002 23179 13036
rect 23113 12986 23179 13002
rect 23442 12958 23476 13325
rect 22818 12906 23476 12958
rect 23116 12884 23208 12906
rect 23116 12832 23128 12884
rect 23194 12832 23208 12884
rect 23116 12828 23208 12832
rect 24516 12704 24607 13958
rect 24856 13876 24926 13884
rect 24856 13808 24867 13876
rect 24924 13808 24934 13876
rect 24856 13800 24926 13808
rect 25009 13695 25044 14205
rect 25099 14159 25191 14172
rect 25099 14096 25111 14159
rect 25182 14096 25191 14159
rect 25099 14087 25191 14096
rect 26184 14159 26276 14169
rect 26184 14097 26196 14159
rect 26266 14097 26276 14159
rect 26184 14084 26276 14097
rect 27572 14104 27607 14458
rect 26431 14042 26496 14045
rect 26431 14039 26500 14042
rect 26431 13979 26437 14039
rect 26496 13979 26506 14039
rect 26431 13975 26500 13979
rect 26431 13973 26496 13975
rect 27572 13958 27753 14104
rect 26066 13876 26158 13884
rect 26066 13811 26078 13876
rect 26146 13811 26158 13876
rect 26066 13799 26158 13811
rect 27572 13696 27607 13958
rect 25009 13648 26381 13695
rect 26703 13649 27607 13696
rect 25843 13525 25877 13648
rect 26315 13635 26381 13648
rect 26315 13601 26331 13635
rect 26365 13601 26381 13635
rect 26315 13585 26381 13601
rect 26704 13525 26738 13649
rect 25838 13513 25884 13525
rect 25838 13337 25844 13513
rect 25878 13337 25884 13513
rect 25838 13325 25884 13337
rect 25956 13513 26076 13525
rect 25956 13337 25962 13513
rect 25996 13337 26036 13513
rect 25956 13325 26036 13337
rect 25962 12958 25996 13325
rect 26030 13137 26036 13325
rect 26070 13137 26076 13513
rect 26030 13125 26076 13137
rect 26148 13513 26194 13525
rect 26148 13137 26154 13513
rect 26188 13137 26194 13513
rect 26148 13125 26194 13137
rect 26266 13513 26312 13525
rect 26266 13137 26272 13513
rect 26306 13137 26312 13513
rect 26266 13125 26312 13137
rect 26384 13513 26430 13525
rect 26384 13137 26390 13513
rect 26424 13137 26430 13513
rect 26384 13125 26430 13137
rect 26502 13513 26626 13525
rect 26502 13137 26508 13513
rect 26542 13337 26586 13513
rect 26620 13337 26626 13513
rect 26542 13325 26626 13337
rect 26698 13513 26744 13525
rect 26698 13337 26704 13513
rect 26738 13337 26744 13513
rect 26698 13325 26744 13337
rect 26542 13137 26548 13325
rect 26502 13125 26548 13137
rect 26272 13052 26306 13125
rect 26257 13036 26323 13052
rect 26257 13002 26273 13036
rect 26307 13002 26323 13036
rect 26257 12986 26323 13002
rect 26586 12958 26620 13325
rect 25962 12906 26620 12958
rect 26260 12884 26352 12906
rect 26260 12832 26272 12884
rect 26338 12832 26352 12884
rect 26260 12828 26352 12832
rect 27673 12705 27753 13958
rect 2708 12636 5710 12700
rect 5852 12636 8853 12701
rect 8984 12636 11986 12701
rect 12128 12636 15126 12704
rect 15330 12636 18333 12704
rect 18474 12636 21478 12704
rect 21606 12636 24607 12704
rect 24750 12637 27753 12705
rect 2708 11314 2780 12636
rect 4206 12304 4216 12364
rect 4296 12304 4306 12364
rect 4206 12264 4306 12304
rect 3409 12207 5212 12264
rect 3409 12120 3443 12207
rect 4584 12120 4618 12207
rect 3403 12108 3449 12120
rect 3403 11920 3409 12108
rect 2962 11908 3008 11920
rect 2962 11732 2968 11908
rect 3002 11732 3008 11908
rect 2962 11720 3008 11732
rect 3080 11908 3126 11920
rect 3080 11732 3086 11908
rect 3120 11732 3126 11908
rect 3080 11720 3126 11732
rect 3198 11908 3244 11920
rect 3198 11732 3204 11908
rect 3238 11732 3244 11908
rect 3198 11720 3244 11732
rect 3316 11908 3409 11920
rect 3316 11732 3322 11908
rect 3356 11732 3409 11908
rect 3443 11732 3449 12108
rect 3316 11720 3449 11732
rect 3521 12108 3567 12120
rect 3521 11732 3527 12108
rect 3561 11732 3567 12108
rect 3521 11720 3567 11732
rect 3639 12108 3685 12120
rect 3639 11732 3645 12108
rect 3679 11732 3685 12108
rect 3639 11720 3685 11732
rect 3757 12108 3803 12120
rect 3757 11732 3763 12108
rect 3797 11732 3803 12108
rect 3757 11720 3803 11732
rect 3870 12108 3916 12120
rect 3870 11732 3876 12108
rect 3910 11732 3916 12108
rect 3870 11720 3916 11732
rect 3988 12108 4034 12120
rect 3988 11732 3994 12108
rect 4028 11732 4034 12108
rect 3988 11720 4034 11732
rect 4106 12108 4152 12120
rect 4106 11732 4112 12108
rect 4146 11732 4152 12108
rect 4106 11720 4152 11732
rect 4224 12108 4270 12120
rect 4224 11732 4230 12108
rect 4264 11732 4270 12108
rect 4224 11720 4270 11732
rect 4342 12108 4388 12120
rect 4342 11732 4348 12108
rect 4382 11732 4388 12108
rect 4342 11720 4388 11732
rect 4460 12108 4506 12120
rect 4460 11732 4466 12108
rect 4500 11732 4506 12108
rect 4460 11720 4506 11732
rect 4578 12108 4624 12120
rect 4578 11732 4584 12108
rect 4618 11732 4624 12108
rect 4578 11720 4624 11732
rect 4697 12108 4743 12120
rect 4697 11732 4703 12108
rect 4737 11732 4743 12108
rect 4697 11720 4743 11732
rect 4815 12108 4861 12120
rect 4815 11732 4821 12108
rect 4855 11732 4861 12108
rect 4815 11720 4861 11732
rect 4933 12108 4979 12120
rect 4933 11732 4939 12108
rect 4973 11732 4979 12108
rect 4933 11720 4979 11732
rect 5051 12108 5097 12120
rect 5051 11732 5057 12108
rect 5091 11732 5097 12108
rect 5175 11920 5212 12207
rect 5051 11720 5097 11732
rect 5170 11908 5216 11920
rect 5170 11732 5176 11908
rect 5210 11732 5216 11908
rect 5170 11720 5216 11732
rect 5288 11908 5334 11920
rect 5288 11732 5294 11908
rect 5328 11732 5334 11908
rect 5288 11720 5334 11732
rect 5406 11908 5452 11920
rect 5406 11732 5412 11908
rect 5446 11732 5452 11908
rect 5406 11720 5452 11732
rect 5524 11908 5570 11920
rect 5524 11732 5530 11908
rect 5564 11732 5570 11908
rect 5524 11720 5570 11732
rect 2967 11534 3002 11720
rect 3876 11636 3910 11720
rect 5057 11636 5091 11720
rect 3876 11594 5091 11636
rect 5057 11574 5091 11594
rect 5057 11558 5414 11574
rect 2967 11517 4104 11534
rect 2967 11483 4054 11517
rect 4088 11483 4104 11517
rect 5057 11524 5364 11558
rect 5398 11524 5414 11558
rect 5057 11508 5414 11524
rect 2967 11467 4104 11483
rect 2708 11306 2884 11314
rect 2189 11099 2299 11247
rect 2708 11238 2825 11306
rect 2882 11238 2892 11306
rect 2708 11230 2884 11238
rect 2189 11029 2212 11099
rect 2279 11029 2299 11099
rect 2189 8698 2299 11029
rect 2708 11138 2884 11146
rect 2708 11070 2825 11138
rect 2882 11070 2892 11138
rect 2708 11062 2884 11070
rect 2708 9874 2792 11062
rect 2967 10957 3002 11467
rect 3057 11421 3149 11434
rect 3057 11358 3069 11421
rect 3140 11358 3149 11421
rect 3057 11349 3149 11358
rect 4142 11421 4234 11431
rect 4142 11359 4154 11421
rect 4224 11359 4234 11421
rect 4142 11346 4234 11359
rect 5530 11366 5565 11720
rect 4389 11304 4454 11307
rect 4389 11301 4458 11304
rect 4389 11241 4395 11301
rect 4454 11241 4464 11301
rect 4389 11237 4458 11241
rect 4389 11235 4454 11237
rect 5530 11220 5711 11366
rect 5852 11314 5923 12636
rect 7350 12304 7360 12364
rect 7440 12304 7450 12364
rect 7350 12264 7450 12304
rect 6553 12207 8356 12264
rect 6553 12120 6587 12207
rect 7728 12120 7762 12207
rect 6547 12108 6593 12120
rect 6547 11920 6553 12108
rect 6106 11908 6152 11920
rect 6106 11732 6112 11908
rect 6146 11732 6152 11908
rect 6106 11720 6152 11732
rect 6224 11908 6270 11920
rect 6224 11732 6230 11908
rect 6264 11732 6270 11908
rect 6224 11720 6270 11732
rect 6342 11908 6388 11920
rect 6342 11732 6348 11908
rect 6382 11732 6388 11908
rect 6342 11720 6388 11732
rect 6460 11908 6553 11920
rect 6460 11732 6466 11908
rect 6500 11732 6553 11908
rect 6587 11732 6593 12108
rect 6460 11720 6593 11732
rect 6665 12108 6711 12120
rect 6665 11732 6671 12108
rect 6705 11732 6711 12108
rect 6665 11720 6711 11732
rect 6783 12108 6829 12120
rect 6783 11732 6789 12108
rect 6823 11732 6829 12108
rect 6783 11720 6829 11732
rect 6901 12108 6947 12120
rect 6901 11732 6907 12108
rect 6941 11732 6947 12108
rect 6901 11720 6947 11732
rect 7014 12108 7060 12120
rect 7014 11732 7020 12108
rect 7054 11732 7060 12108
rect 7014 11720 7060 11732
rect 7132 12108 7178 12120
rect 7132 11732 7138 12108
rect 7172 11732 7178 12108
rect 7132 11720 7178 11732
rect 7250 12108 7296 12120
rect 7250 11732 7256 12108
rect 7290 11732 7296 12108
rect 7250 11720 7296 11732
rect 7368 12108 7414 12120
rect 7368 11732 7374 12108
rect 7408 11732 7414 12108
rect 7368 11720 7414 11732
rect 7486 12108 7532 12120
rect 7486 11732 7492 12108
rect 7526 11732 7532 12108
rect 7486 11720 7532 11732
rect 7604 12108 7650 12120
rect 7604 11732 7610 12108
rect 7644 11732 7650 12108
rect 7604 11720 7650 11732
rect 7722 12108 7768 12120
rect 7722 11732 7728 12108
rect 7762 11732 7768 12108
rect 7722 11720 7768 11732
rect 7841 12108 7887 12120
rect 7841 11732 7847 12108
rect 7881 11732 7887 12108
rect 7841 11720 7887 11732
rect 7959 12108 8005 12120
rect 7959 11732 7965 12108
rect 7999 11732 8005 12108
rect 7959 11720 8005 11732
rect 8077 12108 8123 12120
rect 8077 11732 8083 12108
rect 8117 11732 8123 12108
rect 8077 11720 8123 11732
rect 8195 12108 8241 12120
rect 8195 11732 8201 12108
rect 8235 11732 8241 12108
rect 8319 11920 8356 12207
rect 8195 11720 8241 11732
rect 8314 11908 8360 11920
rect 8314 11732 8320 11908
rect 8354 11732 8360 11908
rect 8314 11720 8360 11732
rect 8432 11908 8478 11920
rect 8432 11732 8438 11908
rect 8472 11732 8478 11908
rect 8432 11720 8478 11732
rect 8550 11908 8596 11920
rect 8550 11732 8556 11908
rect 8590 11732 8596 11908
rect 8550 11720 8596 11732
rect 8668 11908 8714 11920
rect 8668 11732 8674 11908
rect 8708 11732 8714 11908
rect 8668 11720 8714 11732
rect 6111 11534 6146 11720
rect 7020 11636 7054 11720
rect 8201 11636 8235 11720
rect 7020 11594 8235 11636
rect 8201 11574 8235 11594
rect 8201 11558 8558 11574
rect 6111 11517 7248 11534
rect 6111 11483 7198 11517
rect 7232 11483 7248 11517
rect 8201 11524 8508 11558
rect 8542 11524 8558 11558
rect 8201 11508 8558 11524
rect 6111 11467 7248 11483
rect 5852 11306 6028 11314
rect 5852 11238 5969 11306
rect 6026 11238 6036 11306
rect 5852 11230 6028 11238
rect 4024 11138 4116 11146
rect 4024 11073 4036 11138
rect 4104 11073 4116 11138
rect 4024 11061 4116 11073
rect 5530 10958 5565 11220
rect 2967 10910 4339 10957
rect 4661 10911 5565 10958
rect 3801 10787 3835 10910
rect 4273 10897 4339 10910
rect 4273 10863 4289 10897
rect 4323 10863 4339 10897
rect 4273 10847 4339 10863
rect 4662 10787 4696 10911
rect 3796 10775 3842 10787
rect 3796 10599 3802 10775
rect 3836 10599 3842 10775
rect 3796 10587 3842 10599
rect 3914 10775 4034 10787
rect 3914 10599 3920 10775
rect 3954 10599 3994 10775
rect 3914 10587 3994 10599
rect 3920 10220 3954 10587
rect 3988 10399 3994 10587
rect 4028 10399 4034 10775
rect 3988 10387 4034 10399
rect 4106 10775 4152 10787
rect 4106 10399 4112 10775
rect 4146 10399 4152 10775
rect 4106 10387 4152 10399
rect 4224 10775 4270 10787
rect 4224 10399 4230 10775
rect 4264 10399 4270 10775
rect 4224 10387 4270 10399
rect 4342 10775 4388 10787
rect 4342 10399 4348 10775
rect 4382 10399 4388 10775
rect 4342 10387 4388 10399
rect 4460 10775 4584 10787
rect 4460 10399 4466 10775
rect 4500 10599 4544 10775
rect 4578 10599 4584 10775
rect 4500 10587 4584 10599
rect 4656 10775 4702 10787
rect 4656 10599 4662 10775
rect 4696 10599 4702 10775
rect 4656 10587 4702 10599
rect 4500 10399 4506 10587
rect 4460 10387 4506 10399
rect 4230 10314 4264 10387
rect 4215 10298 4281 10314
rect 4215 10264 4231 10298
rect 4265 10264 4281 10298
rect 4215 10248 4281 10264
rect 4544 10220 4578 10587
rect 3920 10168 4578 10220
rect 5638 10177 5711 11220
rect 5852 11138 6028 11146
rect 5852 11070 5969 11138
rect 6026 11070 6036 11138
rect 5852 11065 6028 11070
rect 5851 11062 6028 11065
rect 4218 10146 4310 10168
rect 4218 10094 4230 10146
rect 4296 10094 4310 10146
rect 5634 10100 5644 10177
rect 5708 10100 5718 10177
rect 5638 10099 5711 10100
rect 4218 10090 4310 10094
rect 5851 9875 5926 11062
rect 6111 10957 6146 11467
rect 6201 11421 6293 11434
rect 6201 11358 6213 11421
rect 6284 11358 6293 11421
rect 6201 11349 6293 11358
rect 7286 11421 7378 11431
rect 7286 11359 7298 11421
rect 7368 11359 7378 11421
rect 7286 11346 7378 11359
rect 8674 11366 8709 11720
rect 7533 11304 7598 11307
rect 7533 11301 7602 11304
rect 7533 11241 7539 11301
rect 7598 11241 7608 11301
rect 7533 11237 7602 11241
rect 8674 11238 8855 11366
rect 8984 11318 9055 12636
rect 10482 12308 10492 12368
rect 10572 12308 10582 12368
rect 10482 12268 10582 12308
rect 9685 12211 11488 12268
rect 9685 12124 9719 12211
rect 10860 12124 10894 12211
rect 9679 12112 9725 12124
rect 9679 11924 9685 12112
rect 9238 11912 9284 11924
rect 9238 11736 9244 11912
rect 9278 11736 9284 11912
rect 9238 11724 9284 11736
rect 9356 11912 9402 11924
rect 9356 11736 9362 11912
rect 9396 11736 9402 11912
rect 9356 11724 9402 11736
rect 9474 11912 9520 11924
rect 9474 11736 9480 11912
rect 9514 11736 9520 11912
rect 9474 11724 9520 11736
rect 9592 11912 9685 11924
rect 9592 11736 9598 11912
rect 9632 11736 9685 11912
rect 9719 11736 9725 12112
rect 9592 11724 9725 11736
rect 9797 12112 9843 12124
rect 9797 11736 9803 12112
rect 9837 11736 9843 12112
rect 9797 11724 9843 11736
rect 9915 12112 9961 12124
rect 9915 11736 9921 12112
rect 9955 11736 9961 12112
rect 9915 11724 9961 11736
rect 10033 12112 10079 12124
rect 10033 11736 10039 12112
rect 10073 11736 10079 12112
rect 10033 11724 10079 11736
rect 10146 12112 10192 12124
rect 10146 11736 10152 12112
rect 10186 11736 10192 12112
rect 10146 11724 10192 11736
rect 10264 12112 10310 12124
rect 10264 11736 10270 12112
rect 10304 11736 10310 12112
rect 10264 11724 10310 11736
rect 10382 12112 10428 12124
rect 10382 11736 10388 12112
rect 10422 11736 10428 12112
rect 10382 11724 10428 11736
rect 10500 12112 10546 12124
rect 10500 11736 10506 12112
rect 10540 11736 10546 12112
rect 10500 11724 10546 11736
rect 10618 12112 10664 12124
rect 10618 11736 10624 12112
rect 10658 11736 10664 12112
rect 10618 11724 10664 11736
rect 10736 12112 10782 12124
rect 10736 11736 10742 12112
rect 10776 11736 10782 12112
rect 10736 11724 10782 11736
rect 10854 12112 10900 12124
rect 10854 11736 10860 12112
rect 10894 11736 10900 12112
rect 10854 11724 10900 11736
rect 10973 12112 11019 12124
rect 10973 11736 10979 12112
rect 11013 11736 11019 12112
rect 10973 11724 11019 11736
rect 11091 12112 11137 12124
rect 11091 11736 11097 12112
rect 11131 11736 11137 12112
rect 11091 11724 11137 11736
rect 11209 12112 11255 12124
rect 11209 11736 11215 12112
rect 11249 11736 11255 12112
rect 11209 11724 11255 11736
rect 11327 12112 11373 12124
rect 11327 11736 11333 12112
rect 11367 11736 11373 12112
rect 11451 11924 11488 12211
rect 11327 11724 11373 11736
rect 11446 11912 11492 11924
rect 11446 11736 11452 11912
rect 11486 11736 11492 11912
rect 11446 11724 11492 11736
rect 11564 11912 11610 11924
rect 11564 11736 11570 11912
rect 11604 11736 11610 11912
rect 11564 11724 11610 11736
rect 11682 11912 11728 11924
rect 11682 11736 11688 11912
rect 11722 11736 11728 11912
rect 11682 11724 11728 11736
rect 11800 11912 11846 11924
rect 11800 11736 11806 11912
rect 11840 11736 11846 11912
rect 11800 11724 11846 11736
rect 9243 11538 9278 11724
rect 10152 11640 10186 11724
rect 11333 11640 11367 11724
rect 10152 11598 11367 11640
rect 11333 11578 11367 11598
rect 11333 11562 11690 11578
rect 9243 11521 10380 11538
rect 9243 11487 10330 11521
rect 10364 11487 10380 11521
rect 11333 11528 11640 11562
rect 11674 11528 11690 11562
rect 11333 11512 11690 11528
rect 9243 11471 10380 11487
rect 8984 11310 9160 11318
rect 8984 11242 9101 11310
rect 9158 11242 9168 11310
rect 7533 11235 7598 11237
rect 8674 11220 8856 11238
rect 8984 11234 9160 11242
rect 7168 11138 7260 11146
rect 7168 11073 7180 11138
rect 7248 11073 7260 11138
rect 7168 11061 7260 11073
rect 8674 10958 8709 11220
rect 6111 10910 7483 10957
rect 7805 10911 8709 10958
rect 6945 10787 6979 10910
rect 7417 10897 7483 10910
rect 7417 10863 7433 10897
rect 7467 10863 7483 10897
rect 7417 10847 7483 10863
rect 7806 10787 7840 10911
rect 6940 10775 6986 10787
rect 6940 10599 6946 10775
rect 6980 10599 6986 10775
rect 6940 10587 6986 10599
rect 7058 10775 7178 10787
rect 7058 10599 7064 10775
rect 7098 10599 7138 10775
rect 7058 10587 7138 10599
rect 7064 10220 7098 10587
rect 7132 10399 7138 10587
rect 7172 10399 7178 10775
rect 7132 10387 7178 10399
rect 7250 10775 7296 10787
rect 7250 10399 7256 10775
rect 7290 10399 7296 10775
rect 7250 10387 7296 10399
rect 7368 10775 7414 10787
rect 7368 10399 7374 10775
rect 7408 10399 7414 10775
rect 7368 10387 7414 10399
rect 7486 10775 7532 10787
rect 7486 10399 7492 10775
rect 7526 10399 7532 10775
rect 7486 10387 7532 10399
rect 7604 10775 7728 10787
rect 7604 10399 7610 10775
rect 7644 10599 7688 10775
rect 7722 10599 7728 10775
rect 7644 10587 7728 10599
rect 7800 10775 7846 10787
rect 7800 10599 7806 10775
rect 7840 10599 7846 10775
rect 7800 10587 7846 10599
rect 7644 10399 7650 10587
rect 7604 10387 7650 10399
rect 7374 10314 7408 10387
rect 7359 10298 7425 10314
rect 7359 10264 7375 10298
rect 7409 10264 7425 10298
rect 7359 10248 7425 10264
rect 7688 10220 7722 10587
rect 7064 10168 7722 10220
rect 7362 10146 7454 10168
rect 7362 10094 7374 10146
rect 7440 10094 7454 10146
rect 8758 10118 8856 11220
rect 7362 10090 7454 10094
rect 8744 10046 8754 10118
rect 8822 10068 8856 10118
rect 9001 11142 9160 11150
rect 9001 11074 9101 11142
rect 9158 11074 9168 11142
rect 9001 11066 9160 11074
rect 8822 10046 8832 10068
rect 9001 9875 9050 11066
rect 9243 10961 9278 11471
rect 9333 11425 9425 11438
rect 9333 11362 9345 11425
rect 9416 11362 9425 11425
rect 9333 11353 9425 11362
rect 10418 11425 10510 11435
rect 10418 11363 10430 11425
rect 10500 11363 10510 11425
rect 10418 11350 10510 11363
rect 11806 11370 11841 11724
rect 10665 11308 10730 11311
rect 10665 11305 10734 11308
rect 10665 11245 10671 11305
rect 10730 11245 10740 11305
rect 10665 11241 10734 11245
rect 10665 11239 10730 11241
rect 11806 11224 11987 11370
rect 12128 11318 12199 12636
rect 13626 12308 13636 12368
rect 13716 12308 13726 12368
rect 13626 12268 13726 12308
rect 12829 12211 14632 12268
rect 12829 12124 12863 12211
rect 14004 12124 14038 12211
rect 12823 12112 12869 12124
rect 12823 11924 12829 12112
rect 12382 11912 12428 11924
rect 12382 11736 12388 11912
rect 12422 11736 12428 11912
rect 12382 11724 12428 11736
rect 12500 11912 12546 11924
rect 12500 11736 12506 11912
rect 12540 11736 12546 11912
rect 12500 11724 12546 11736
rect 12618 11912 12664 11924
rect 12618 11736 12624 11912
rect 12658 11736 12664 11912
rect 12618 11724 12664 11736
rect 12736 11912 12829 11924
rect 12736 11736 12742 11912
rect 12776 11736 12829 11912
rect 12863 11736 12869 12112
rect 12736 11724 12869 11736
rect 12941 12112 12987 12124
rect 12941 11736 12947 12112
rect 12981 11736 12987 12112
rect 12941 11724 12987 11736
rect 13059 12112 13105 12124
rect 13059 11736 13065 12112
rect 13099 11736 13105 12112
rect 13059 11724 13105 11736
rect 13177 12112 13223 12124
rect 13177 11736 13183 12112
rect 13217 11736 13223 12112
rect 13177 11724 13223 11736
rect 13290 12112 13336 12124
rect 13290 11736 13296 12112
rect 13330 11736 13336 12112
rect 13290 11724 13336 11736
rect 13408 12112 13454 12124
rect 13408 11736 13414 12112
rect 13448 11736 13454 12112
rect 13408 11724 13454 11736
rect 13526 12112 13572 12124
rect 13526 11736 13532 12112
rect 13566 11736 13572 12112
rect 13526 11724 13572 11736
rect 13644 12112 13690 12124
rect 13644 11736 13650 12112
rect 13684 11736 13690 12112
rect 13644 11724 13690 11736
rect 13762 12112 13808 12124
rect 13762 11736 13768 12112
rect 13802 11736 13808 12112
rect 13762 11724 13808 11736
rect 13880 12112 13926 12124
rect 13880 11736 13886 12112
rect 13920 11736 13926 12112
rect 13880 11724 13926 11736
rect 13998 12112 14044 12124
rect 13998 11736 14004 12112
rect 14038 11736 14044 12112
rect 13998 11724 14044 11736
rect 14117 12112 14163 12124
rect 14117 11736 14123 12112
rect 14157 11736 14163 12112
rect 14117 11724 14163 11736
rect 14235 12112 14281 12124
rect 14235 11736 14241 12112
rect 14275 11736 14281 12112
rect 14235 11724 14281 11736
rect 14353 12112 14399 12124
rect 14353 11736 14359 12112
rect 14393 11736 14399 12112
rect 14353 11724 14399 11736
rect 14471 12112 14517 12124
rect 14471 11736 14477 12112
rect 14511 11736 14517 12112
rect 14595 11924 14632 12211
rect 14471 11724 14517 11736
rect 14590 11912 14636 11924
rect 14590 11736 14596 11912
rect 14630 11736 14636 11912
rect 14590 11724 14636 11736
rect 14708 11912 14754 11924
rect 14708 11736 14714 11912
rect 14748 11736 14754 11912
rect 14708 11724 14754 11736
rect 14826 11912 14872 11924
rect 14826 11736 14832 11912
rect 14866 11736 14872 11912
rect 14826 11724 14872 11736
rect 14944 11912 14990 11924
rect 14944 11736 14950 11912
rect 14984 11736 14990 11912
rect 14944 11724 14990 11736
rect 12387 11538 12422 11724
rect 13296 11640 13330 11724
rect 14477 11640 14511 11724
rect 13296 11598 14511 11640
rect 14477 11578 14511 11598
rect 14477 11562 14834 11578
rect 12387 11521 13524 11538
rect 12387 11487 13474 11521
rect 13508 11487 13524 11521
rect 14477 11528 14784 11562
rect 14818 11528 14834 11562
rect 14477 11512 14834 11528
rect 12387 11471 13524 11487
rect 12128 11310 12304 11318
rect 12128 11242 12245 11310
rect 12302 11242 12312 11310
rect 12128 11234 12304 11242
rect 10300 11142 10392 11150
rect 10300 11077 10312 11142
rect 10380 11077 10392 11142
rect 10300 11065 10392 11077
rect 11806 10962 11841 11224
rect 9243 10914 10615 10961
rect 10937 10915 11841 10962
rect 10077 10791 10111 10914
rect 10549 10901 10615 10914
rect 10549 10867 10565 10901
rect 10599 10867 10615 10901
rect 10549 10851 10615 10867
rect 10938 10791 10972 10915
rect 10072 10779 10118 10791
rect 10072 10603 10078 10779
rect 10112 10603 10118 10779
rect 10072 10591 10118 10603
rect 10190 10779 10310 10791
rect 10190 10603 10196 10779
rect 10230 10603 10270 10779
rect 10190 10591 10270 10603
rect 10196 10224 10230 10591
rect 10264 10403 10270 10591
rect 10304 10403 10310 10779
rect 10264 10391 10310 10403
rect 10382 10779 10428 10791
rect 10382 10403 10388 10779
rect 10422 10403 10428 10779
rect 10382 10391 10428 10403
rect 10500 10779 10546 10791
rect 10500 10403 10506 10779
rect 10540 10403 10546 10779
rect 10500 10391 10546 10403
rect 10618 10779 10664 10791
rect 10618 10403 10624 10779
rect 10658 10403 10664 10779
rect 10618 10391 10664 10403
rect 10736 10779 10860 10791
rect 10736 10403 10742 10779
rect 10776 10603 10820 10779
rect 10854 10603 10860 10779
rect 10776 10591 10860 10603
rect 10932 10779 10978 10791
rect 10932 10603 10938 10779
rect 10972 10603 10978 10779
rect 10932 10591 10978 10603
rect 10776 10403 10782 10591
rect 10736 10391 10782 10403
rect 10506 10318 10540 10391
rect 10491 10302 10557 10318
rect 10491 10268 10507 10302
rect 10541 10268 10557 10302
rect 10491 10252 10557 10268
rect 10820 10224 10854 10591
rect 10196 10172 10854 10224
rect 10494 10150 10586 10172
rect 10494 10098 10506 10150
rect 10572 10098 10586 10150
rect 10494 10094 10586 10098
rect 11896 9992 11987 11224
rect 11880 9924 11890 9992
rect 11957 9926 11987 9992
rect 12152 11142 12304 11150
rect 12152 11074 12245 11142
rect 12302 11074 12312 11142
rect 12152 11066 12304 11074
rect 11957 9924 11967 9926
rect 12152 9875 12213 11066
rect 12387 10961 12422 11471
rect 12477 11425 12569 11438
rect 12477 11362 12489 11425
rect 12560 11362 12569 11425
rect 12477 11353 12569 11362
rect 13562 11425 13654 11435
rect 13562 11363 13574 11425
rect 13644 11363 13654 11425
rect 13562 11350 13654 11363
rect 14950 11370 14985 11724
rect 13809 11308 13874 11311
rect 13809 11305 13878 11308
rect 13809 11245 13815 11305
rect 13874 11245 13884 11305
rect 13809 11241 13878 11245
rect 13809 11239 13874 11241
rect 14950 11224 15131 11370
rect 15330 11314 15401 12636
rect 16828 12304 16838 12364
rect 16918 12304 16928 12364
rect 16828 12264 16928 12304
rect 16031 12207 17834 12264
rect 16031 12120 16065 12207
rect 17206 12120 17240 12207
rect 16025 12108 16071 12120
rect 16025 11920 16031 12108
rect 15584 11908 15630 11920
rect 15584 11732 15590 11908
rect 15624 11732 15630 11908
rect 15584 11720 15630 11732
rect 15702 11908 15748 11920
rect 15702 11732 15708 11908
rect 15742 11732 15748 11908
rect 15702 11720 15748 11732
rect 15820 11908 15866 11920
rect 15820 11732 15826 11908
rect 15860 11732 15866 11908
rect 15820 11720 15866 11732
rect 15938 11908 16031 11920
rect 15938 11732 15944 11908
rect 15978 11732 16031 11908
rect 16065 11732 16071 12108
rect 15938 11720 16071 11732
rect 16143 12108 16189 12120
rect 16143 11732 16149 12108
rect 16183 11732 16189 12108
rect 16143 11720 16189 11732
rect 16261 12108 16307 12120
rect 16261 11732 16267 12108
rect 16301 11732 16307 12108
rect 16261 11720 16307 11732
rect 16379 12108 16425 12120
rect 16379 11732 16385 12108
rect 16419 11732 16425 12108
rect 16379 11720 16425 11732
rect 16492 12108 16538 12120
rect 16492 11732 16498 12108
rect 16532 11732 16538 12108
rect 16492 11720 16538 11732
rect 16610 12108 16656 12120
rect 16610 11732 16616 12108
rect 16650 11732 16656 12108
rect 16610 11720 16656 11732
rect 16728 12108 16774 12120
rect 16728 11732 16734 12108
rect 16768 11732 16774 12108
rect 16728 11720 16774 11732
rect 16846 12108 16892 12120
rect 16846 11732 16852 12108
rect 16886 11732 16892 12108
rect 16846 11720 16892 11732
rect 16964 12108 17010 12120
rect 16964 11732 16970 12108
rect 17004 11732 17010 12108
rect 16964 11720 17010 11732
rect 17082 12108 17128 12120
rect 17082 11732 17088 12108
rect 17122 11732 17128 12108
rect 17082 11720 17128 11732
rect 17200 12108 17246 12120
rect 17200 11732 17206 12108
rect 17240 11732 17246 12108
rect 17200 11720 17246 11732
rect 17319 12108 17365 12120
rect 17319 11732 17325 12108
rect 17359 11732 17365 12108
rect 17319 11720 17365 11732
rect 17437 12108 17483 12120
rect 17437 11732 17443 12108
rect 17477 11732 17483 12108
rect 17437 11720 17483 11732
rect 17555 12108 17601 12120
rect 17555 11732 17561 12108
rect 17595 11732 17601 12108
rect 17555 11720 17601 11732
rect 17673 12108 17719 12120
rect 17673 11732 17679 12108
rect 17713 11732 17719 12108
rect 17797 11920 17834 12207
rect 17673 11720 17719 11732
rect 17792 11908 17838 11920
rect 17792 11732 17798 11908
rect 17832 11732 17838 11908
rect 17792 11720 17838 11732
rect 17910 11908 17956 11920
rect 17910 11732 17916 11908
rect 17950 11732 17956 11908
rect 17910 11720 17956 11732
rect 18028 11908 18074 11920
rect 18028 11732 18034 11908
rect 18068 11732 18074 11908
rect 18028 11720 18074 11732
rect 18146 11908 18192 11920
rect 18146 11732 18152 11908
rect 18186 11732 18192 11908
rect 18146 11720 18192 11732
rect 15589 11534 15624 11720
rect 16498 11636 16532 11720
rect 17679 11636 17713 11720
rect 16498 11594 17713 11636
rect 17679 11574 17713 11594
rect 17679 11558 18036 11574
rect 15589 11517 16726 11534
rect 15589 11483 16676 11517
rect 16710 11483 16726 11517
rect 17679 11524 17986 11558
rect 18020 11524 18036 11558
rect 17679 11508 18036 11524
rect 15589 11467 16726 11483
rect 15330 11306 15506 11314
rect 15330 11238 15447 11306
rect 15504 11238 15514 11306
rect 15330 11230 15506 11238
rect 13444 11142 13536 11150
rect 13444 11077 13456 11142
rect 13524 11077 13536 11142
rect 13444 11065 13536 11077
rect 14950 10962 14985 11224
rect 12387 10914 13759 10961
rect 14081 10915 14985 10962
rect 13221 10791 13255 10914
rect 13693 10901 13759 10914
rect 13693 10867 13709 10901
rect 13743 10867 13759 10901
rect 13693 10851 13759 10867
rect 14082 10791 14116 10915
rect 13216 10779 13262 10791
rect 13216 10603 13222 10779
rect 13256 10603 13262 10779
rect 13216 10591 13262 10603
rect 13334 10779 13454 10791
rect 13334 10603 13340 10779
rect 13374 10603 13414 10779
rect 13334 10591 13414 10603
rect 13340 10224 13374 10591
rect 13408 10403 13414 10591
rect 13448 10403 13454 10779
rect 13408 10391 13454 10403
rect 13526 10779 13572 10791
rect 13526 10403 13532 10779
rect 13566 10403 13572 10779
rect 13526 10391 13572 10403
rect 13644 10779 13690 10791
rect 13644 10403 13650 10779
rect 13684 10403 13690 10779
rect 13644 10391 13690 10403
rect 13762 10779 13808 10791
rect 13762 10403 13768 10779
rect 13802 10403 13808 10779
rect 13762 10391 13808 10403
rect 13880 10779 14004 10791
rect 13880 10403 13886 10779
rect 13920 10603 13964 10779
rect 13998 10603 14004 10779
rect 13920 10591 14004 10603
rect 14076 10779 14122 10791
rect 14076 10603 14082 10779
rect 14116 10603 14122 10779
rect 14076 10591 14122 10603
rect 13920 10403 13926 10591
rect 13880 10391 13926 10403
rect 13650 10318 13684 10391
rect 13635 10302 13701 10318
rect 13635 10268 13651 10302
rect 13685 10268 13701 10302
rect 13635 10252 13701 10268
rect 13964 10224 13998 10591
rect 15037 10336 15130 11224
rect 15027 10267 15037 10336
rect 15115 10267 15130 10336
rect 15330 11138 15506 11146
rect 15330 11070 15447 11138
rect 15504 11070 15514 11138
rect 15330 11062 15506 11070
rect 13340 10172 13998 10224
rect 13638 10150 13730 10172
rect 13638 10098 13650 10150
rect 13716 10098 13730 10150
rect 13638 10094 13730 10098
rect 15330 9876 15406 11062
rect 15589 10957 15624 11467
rect 15679 11421 15771 11434
rect 15679 11358 15691 11421
rect 15762 11358 15771 11421
rect 15679 11349 15771 11358
rect 16764 11421 16856 11431
rect 16764 11359 16776 11421
rect 16846 11359 16856 11421
rect 16764 11346 16856 11359
rect 18152 11366 18187 11720
rect 17011 11304 17076 11307
rect 17011 11301 17080 11304
rect 17011 11241 17017 11301
rect 17076 11241 17086 11301
rect 18152 11269 18333 11366
rect 18474 11314 18545 12636
rect 19972 12304 19982 12364
rect 20062 12304 20072 12364
rect 19972 12264 20072 12304
rect 19175 12207 20978 12264
rect 19175 12120 19209 12207
rect 20350 12120 20384 12207
rect 19169 12108 19215 12120
rect 19169 11920 19175 12108
rect 18728 11908 18774 11920
rect 18728 11732 18734 11908
rect 18768 11732 18774 11908
rect 18728 11720 18774 11732
rect 18846 11908 18892 11920
rect 18846 11732 18852 11908
rect 18886 11732 18892 11908
rect 18846 11720 18892 11732
rect 18964 11908 19010 11920
rect 18964 11732 18970 11908
rect 19004 11732 19010 11908
rect 18964 11720 19010 11732
rect 19082 11908 19175 11920
rect 19082 11732 19088 11908
rect 19122 11732 19175 11908
rect 19209 11732 19215 12108
rect 19082 11720 19215 11732
rect 19287 12108 19333 12120
rect 19287 11732 19293 12108
rect 19327 11732 19333 12108
rect 19287 11720 19333 11732
rect 19405 12108 19451 12120
rect 19405 11732 19411 12108
rect 19445 11732 19451 12108
rect 19405 11720 19451 11732
rect 19523 12108 19569 12120
rect 19523 11732 19529 12108
rect 19563 11732 19569 12108
rect 19523 11720 19569 11732
rect 19636 12108 19682 12120
rect 19636 11732 19642 12108
rect 19676 11732 19682 12108
rect 19636 11720 19682 11732
rect 19754 12108 19800 12120
rect 19754 11732 19760 12108
rect 19794 11732 19800 12108
rect 19754 11720 19800 11732
rect 19872 12108 19918 12120
rect 19872 11732 19878 12108
rect 19912 11732 19918 12108
rect 19872 11720 19918 11732
rect 19990 12108 20036 12120
rect 19990 11732 19996 12108
rect 20030 11732 20036 12108
rect 19990 11720 20036 11732
rect 20108 12108 20154 12120
rect 20108 11732 20114 12108
rect 20148 11732 20154 12108
rect 20108 11720 20154 11732
rect 20226 12108 20272 12120
rect 20226 11732 20232 12108
rect 20266 11732 20272 12108
rect 20226 11720 20272 11732
rect 20344 12108 20390 12120
rect 20344 11732 20350 12108
rect 20384 11732 20390 12108
rect 20344 11720 20390 11732
rect 20463 12108 20509 12120
rect 20463 11732 20469 12108
rect 20503 11732 20509 12108
rect 20463 11720 20509 11732
rect 20581 12108 20627 12120
rect 20581 11732 20587 12108
rect 20621 11732 20627 12108
rect 20581 11720 20627 11732
rect 20699 12108 20745 12120
rect 20699 11732 20705 12108
rect 20739 11732 20745 12108
rect 20699 11720 20745 11732
rect 20817 12108 20863 12120
rect 20817 11732 20823 12108
rect 20857 11732 20863 12108
rect 20941 11920 20978 12207
rect 20817 11720 20863 11732
rect 20936 11908 20982 11920
rect 20936 11732 20942 11908
rect 20976 11732 20982 11908
rect 20936 11720 20982 11732
rect 21054 11908 21100 11920
rect 21054 11732 21060 11908
rect 21094 11732 21100 11908
rect 21054 11720 21100 11732
rect 21172 11908 21218 11920
rect 21172 11732 21178 11908
rect 21212 11732 21218 11908
rect 21172 11720 21218 11732
rect 21290 11908 21336 11920
rect 21290 11732 21296 11908
rect 21330 11732 21336 11908
rect 21290 11720 21336 11732
rect 18733 11534 18768 11720
rect 19642 11636 19676 11720
rect 20823 11636 20857 11720
rect 19642 11594 20857 11636
rect 20823 11574 20857 11594
rect 20823 11558 21180 11574
rect 18733 11517 19870 11534
rect 18733 11483 19820 11517
rect 19854 11483 19870 11517
rect 20823 11524 21130 11558
rect 21164 11524 21180 11558
rect 20823 11508 21180 11524
rect 18733 11467 19870 11483
rect 18584 11422 18650 11430
rect 18584 11354 18591 11422
rect 18648 11354 18658 11422
rect 18584 11346 18650 11354
rect 18474 11306 18650 11314
rect 17011 11237 17080 11241
rect 17011 11235 17076 11237
rect 18152 11220 18335 11269
rect 18474 11238 18591 11306
rect 18648 11238 18658 11306
rect 18474 11230 18650 11238
rect 16646 11138 16738 11146
rect 16646 11073 16658 11138
rect 16726 11073 16738 11138
rect 16646 11061 16738 11073
rect 18152 10958 18187 11220
rect 15589 10910 16961 10957
rect 17283 10911 18187 10958
rect 16423 10787 16457 10910
rect 16895 10897 16961 10910
rect 16895 10863 16911 10897
rect 16945 10863 16961 10897
rect 16895 10847 16961 10863
rect 17284 10787 17318 10911
rect 16418 10775 16464 10787
rect 16418 10599 16424 10775
rect 16458 10599 16464 10775
rect 16418 10587 16464 10599
rect 16536 10775 16656 10787
rect 16536 10599 16542 10775
rect 16576 10599 16616 10775
rect 16536 10587 16616 10599
rect 16542 10220 16576 10587
rect 16610 10399 16616 10587
rect 16650 10399 16656 10775
rect 16610 10387 16656 10399
rect 16728 10775 16774 10787
rect 16728 10399 16734 10775
rect 16768 10399 16774 10775
rect 16728 10387 16774 10399
rect 16846 10775 16892 10787
rect 16846 10399 16852 10775
rect 16886 10399 16892 10775
rect 16846 10387 16892 10399
rect 16964 10775 17010 10787
rect 16964 10399 16970 10775
rect 17004 10399 17010 10775
rect 16964 10387 17010 10399
rect 17082 10775 17206 10787
rect 17082 10399 17088 10775
rect 17122 10599 17166 10775
rect 17200 10599 17206 10775
rect 17122 10587 17206 10599
rect 17278 10775 17324 10787
rect 17278 10599 17284 10775
rect 17318 10599 17324 10775
rect 17278 10587 17324 10599
rect 17122 10399 17128 10587
rect 17082 10387 17128 10399
rect 16852 10314 16886 10387
rect 16837 10298 16903 10314
rect 16837 10264 16853 10298
rect 16887 10264 16903 10298
rect 16837 10248 16903 10264
rect 17166 10220 17200 10587
rect 18237 10540 18335 11220
rect 18498 11138 18650 11146
rect 18498 11070 18591 11138
rect 18648 11070 18658 11138
rect 18498 11062 18650 11070
rect 18227 10445 18237 10540
rect 18333 10445 18343 10540
rect 16542 10168 17200 10220
rect 16840 10146 16932 10168
rect 16840 10094 16852 10146
rect 16918 10094 16932 10146
rect 16840 10090 16932 10094
rect 18498 9876 18555 11062
rect 18733 10957 18768 11467
rect 18823 11421 18915 11434
rect 18823 11358 18835 11421
rect 18906 11358 18915 11421
rect 18823 11349 18915 11358
rect 19908 11421 20000 11431
rect 19908 11359 19920 11421
rect 19990 11359 20000 11421
rect 19908 11346 20000 11359
rect 21296 11366 21331 11720
rect 20155 11304 20220 11307
rect 20155 11301 20224 11304
rect 20155 11241 20161 11301
rect 20220 11241 20230 11301
rect 20155 11237 20224 11241
rect 20155 11235 20220 11237
rect 21296 11220 21477 11366
rect 21606 11318 21677 12636
rect 23104 12308 23114 12368
rect 23194 12308 23204 12368
rect 23104 12268 23204 12308
rect 22307 12211 24110 12268
rect 22307 12124 22341 12211
rect 23482 12124 23516 12211
rect 22301 12112 22347 12124
rect 22301 11924 22307 12112
rect 21860 11912 21906 11924
rect 21860 11736 21866 11912
rect 21900 11736 21906 11912
rect 21860 11724 21906 11736
rect 21978 11912 22024 11924
rect 21978 11736 21984 11912
rect 22018 11736 22024 11912
rect 21978 11724 22024 11736
rect 22096 11912 22142 11924
rect 22096 11736 22102 11912
rect 22136 11736 22142 11912
rect 22096 11724 22142 11736
rect 22214 11912 22307 11924
rect 22214 11736 22220 11912
rect 22254 11736 22307 11912
rect 22341 11736 22347 12112
rect 22214 11724 22347 11736
rect 22419 12112 22465 12124
rect 22419 11736 22425 12112
rect 22459 11736 22465 12112
rect 22419 11724 22465 11736
rect 22537 12112 22583 12124
rect 22537 11736 22543 12112
rect 22577 11736 22583 12112
rect 22537 11724 22583 11736
rect 22655 12112 22701 12124
rect 22655 11736 22661 12112
rect 22695 11736 22701 12112
rect 22655 11724 22701 11736
rect 22768 12112 22814 12124
rect 22768 11736 22774 12112
rect 22808 11736 22814 12112
rect 22768 11724 22814 11736
rect 22886 12112 22932 12124
rect 22886 11736 22892 12112
rect 22926 11736 22932 12112
rect 22886 11724 22932 11736
rect 23004 12112 23050 12124
rect 23004 11736 23010 12112
rect 23044 11736 23050 12112
rect 23004 11724 23050 11736
rect 23122 12112 23168 12124
rect 23122 11736 23128 12112
rect 23162 11736 23168 12112
rect 23122 11724 23168 11736
rect 23240 12112 23286 12124
rect 23240 11736 23246 12112
rect 23280 11736 23286 12112
rect 23240 11724 23286 11736
rect 23358 12112 23404 12124
rect 23358 11736 23364 12112
rect 23398 11736 23404 12112
rect 23358 11724 23404 11736
rect 23476 12112 23522 12124
rect 23476 11736 23482 12112
rect 23516 11736 23522 12112
rect 23476 11724 23522 11736
rect 23595 12112 23641 12124
rect 23595 11736 23601 12112
rect 23635 11736 23641 12112
rect 23595 11724 23641 11736
rect 23713 12112 23759 12124
rect 23713 11736 23719 12112
rect 23753 11736 23759 12112
rect 23713 11724 23759 11736
rect 23831 12112 23877 12124
rect 23831 11736 23837 12112
rect 23871 11736 23877 12112
rect 23831 11724 23877 11736
rect 23949 12112 23995 12124
rect 23949 11736 23955 12112
rect 23989 11736 23995 12112
rect 24073 11924 24110 12211
rect 23949 11724 23995 11736
rect 24068 11912 24114 11924
rect 24068 11736 24074 11912
rect 24108 11736 24114 11912
rect 24068 11724 24114 11736
rect 24186 11912 24232 11924
rect 24186 11736 24192 11912
rect 24226 11736 24232 11912
rect 24186 11724 24232 11736
rect 24304 11912 24350 11924
rect 24304 11736 24310 11912
rect 24344 11736 24350 11912
rect 24304 11724 24350 11736
rect 24422 11912 24468 11924
rect 24422 11736 24428 11912
rect 24462 11736 24468 11912
rect 24422 11724 24468 11736
rect 21865 11538 21900 11724
rect 22774 11640 22808 11724
rect 23955 11640 23989 11724
rect 22774 11598 23989 11640
rect 23955 11578 23989 11598
rect 23955 11562 24312 11578
rect 21865 11521 23002 11538
rect 21865 11487 22952 11521
rect 22986 11487 23002 11521
rect 23955 11528 24262 11562
rect 24296 11528 24312 11562
rect 23955 11512 24312 11528
rect 21865 11471 23002 11487
rect 21606 11310 21782 11318
rect 21606 11242 21723 11310
rect 21780 11242 21790 11310
rect 21606 11234 21782 11242
rect 19790 11138 19882 11146
rect 19790 11073 19802 11138
rect 19870 11073 19882 11138
rect 19790 11061 19882 11073
rect 21296 10958 21331 11220
rect 18733 10910 20105 10957
rect 20427 10911 21331 10958
rect 19567 10787 19601 10910
rect 20039 10897 20105 10910
rect 20039 10863 20055 10897
rect 20089 10863 20105 10897
rect 20039 10847 20105 10863
rect 20428 10787 20462 10911
rect 19562 10775 19608 10787
rect 19562 10599 19568 10775
rect 19602 10599 19608 10775
rect 19562 10587 19608 10599
rect 19680 10775 19800 10787
rect 19680 10599 19686 10775
rect 19720 10599 19760 10775
rect 19680 10587 19760 10599
rect 19686 10220 19720 10587
rect 19754 10399 19760 10587
rect 19794 10399 19800 10775
rect 19754 10387 19800 10399
rect 19872 10775 19918 10787
rect 19872 10399 19878 10775
rect 19912 10399 19918 10775
rect 19872 10387 19918 10399
rect 19990 10775 20036 10787
rect 19990 10399 19996 10775
rect 20030 10399 20036 10775
rect 19990 10387 20036 10399
rect 20108 10775 20154 10787
rect 20108 10399 20114 10775
rect 20148 10399 20154 10775
rect 20108 10387 20154 10399
rect 20226 10775 20350 10787
rect 20226 10399 20232 10775
rect 20266 10599 20310 10775
rect 20344 10599 20350 10775
rect 20266 10587 20350 10599
rect 20422 10775 20468 10787
rect 20422 10599 20428 10775
rect 20462 10599 20468 10775
rect 21387 10771 21477 11220
rect 21386 10678 21396 10771
rect 21466 10678 21477 10771
rect 21387 10670 21477 10678
rect 21614 11142 21782 11150
rect 21614 11074 21723 11142
rect 21780 11074 21790 11142
rect 21614 11066 21782 11074
rect 20422 10587 20468 10599
rect 20266 10399 20272 10587
rect 20226 10387 20272 10399
rect 19996 10314 20030 10387
rect 19981 10298 20047 10314
rect 19981 10264 19997 10298
rect 20031 10264 20047 10298
rect 19981 10248 20047 10264
rect 20310 10220 20344 10587
rect 19686 10168 20344 10220
rect 19984 10146 20076 10168
rect 19984 10094 19996 10146
rect 20062 10094 20076 10146
rect 19984 10090 20076 10094
rect 2708 9814 5702 9874
rect 5851 9814 8845 9875
rect 4196 9572 4206 9632
rect 4286 9572 4296 9632
rect 4196 9532 4296 9572
rect 3399 9475 5202 9532
rect 3399 9388 3433 9475
rect 4574 9388 4608 9475
rect 3393 9376 3439 9388
rect 3393 9188 3399 9376
rect 2952 9176 2998 9188
rect 2952 9000 2958 9176
rect 2992 9000 2998 9176
rect 2952 8988 2998 9000
rect 3070 9176 3116 9188
rect 3070 9000 3076 9176
rect 3110 9000 3116 9176
rect 3070 8988 3116 9000
rect 3188 9176 3234 9188
rect 3188 9000 3194 9176
rect 3228 9000 3234 9176
rect 3188 8988 3234 9000
rect 3306 9176 3399 9188
rect 3306 9000 3312 9176
rect 3346 9000 3399 9176
rect 3433 9000 3439 9376
rect 3306 8988 3439 9000
rect 3511 9376 3557 9388
rect 3511 9000 3517 9376
rect 3551 9000 3557 9376
rect 3511 8988 3557 9000
rect 3629 9376 3675 9388
rect 3629 9000 3635 9376
rect 3669 9000 3675 9376
rect 3629 8988 3675 9000
rect 3747 9376 3793 9388
rect 3747 9000 3753 9376
rect 3787 9000 3793 9376
rect 3747 8988 3793 9000
rect 3860 9376 3906 9388
rect 3860 9000 3866 9376
rect 3900 9000 3906 9376
rect 3860 8988 3906 9000
rect 3978 9376 4024 9388
rect 3978 9000 3984 9376
rect 4018 9000 4024 9376
rect 3978 8988 4024 9000
rect 4096 9376 4142 9388
rect 4096 9000 4102 9376
rect 4136 9000 4142 9376
rect 4096 8988 4142 9000
rect 4214 9376 4260 9388
rect 4214 9000 4220 9376
rect 4254 9000 4260 9376
rect 4214 8988 4260 9000
rect 4332 9376 4378 9388
rect 4332 9000 4338 9376
rect 4372 9000 4378 9376
rect 4332 8988 4378 9000
rect 4450 9376 4496 9388
rect 4450 9000 4456 9376
rect 4490 9000 4496 9376
rect 4450 8988 4496 9000
rect 4568 9376 4614 9388
rect 4568 9000 4574 9376
rect 4608 9000 4614 9376
rect 4568 8988 4614 9000
rect 4687 9376 4733 9388
rect 4687 9000 4693 9376
rect 4727 9000 4733 9376
rect 4687 8988 4733 9000
rect 4805 9376 4851 9388
rect 4805 9000 4811 9376
rect 4845 9000 4851 9376
rect 4805 8988 4851 9000
rect 4923 9376 4969 9388
rect 4923 9000 4929 9376
rect 4963 9000 4969 9376
rect 4923 8988 4969 9000
rect 5041 9376 5087 9388
rect 5041 9000 5047 9376
rect 5081 9000 5087 9376
rect 5165 9188 5202 9475
rect 5041 8988 5087 9000
rect 5160 9176 5206 9188
rect 5160 9000 5166 9176
rect 5200 9000 5206 9176
rect 5160 8988 5206 9000
rect 5278 9176 5324 9188
rect 5278 9000 5284 9176
rect 5318 9000 5324 9176
rect 5278 8988 5324 9000
rect 5396 9176 5442 9188
rect 5396 9000 5402 9176
rect 5436 9000 5442 9176
rect 5396 8988 5442 9000
rect 5514 9176 5560 9188
rect 5514 9000 5520 9176
rect 5554 9000 5560 9176
rect 5514 8988 5560 9000
rect 2957 8802 2992 8988
rect 3866 8904 3900 8988
rect 5047 8904 5081 8988
rect 3866 8862 5081 8904
rect 5047 8842 5081 8862
rect 5047 8826 5404 8842
rect 2957 8785 4094 8802
rect 2957 8751 4044 8785
rect 4078 8751 4094 8785
rect 5047 8792 5354 8826
rect 5388 8792 5404 8826
rect 5047 8776 5404 8792
rect 2957 8735 4094 8751
rect 2189 8690 2874 8698
rect 2189 8622 2815 8690
rect 2872 8622 2882 8690
rect 2189 8614 2874 8622
rect 2799 8574 2874 8582
rect 2799 8506 2815 8574
rect 2872 8506 2882 8574
rect 2799 8498 2874 8506
rect 2740 8406 2874 8414
rect 2740 8338 2815 8406
rect 2872 8338 2882 8406
rect 2740 8330 2874 8338
rect 2740 6899 2804 8330
rect 2957 8225 2992 8735
rect 3047 8689 3139 8702
rect 3047 8626 3059 8689
rect 3130 8626 3139 8689
rect 3047 8617 3139 8626
rect 4132 8689 4224 8699
rect 4132 8627 4144 8689
rect 4214 8627 4224 8689
rect 4132 8614 4224 8627
rect 5520 8634 5555 8988
rect 5630 8634 5702 9814
rect 7340 9572 7350 9632
rect 7430 9572 7440 9632
rect 7340 9532 7440 9572
rect 6543 9475 8346 9532
rect 6543 9388 6577 9475
rect 7718 9388 7752 9475
rect 6537 9376 6583 9388
rect 6537 9188 6543 9376
rect 6096 9176 6142 9188
rect 6096 9000 6102 9176
rect 6136 9000 6142 9176
rect 6096 8988 6142 9000
rect 6214 9176 6260 9188
rect 6214 9000 6220 9176
rect 6254 9000 6260 9176
rect 6214 8988 6260 9000
rect 6332 9176 6378 9188
rect 6332 9000 6338 9176
rect 6372 9000 6378 9176
rect 6332 8988 6378 9000
rect 6450 9176 6543 9188
rect 6450 9000 6456 9176
rect 6490 9000 6543 9176
rect 6577 9000 6583 9376
rect 6450 8988 6583 9000
rect 6655 9376 6701 9388
rect 6655 9000 6661 9376
rect 6695 9000 6701 9376
rect 6655 8988 6701 9000
rect 6773 9376 6819 9388
rect 6773 9000 6779 9376
rect 6813 9000 6819 9376
rect 6773 8988 6819 9000
rect 6891 9376 6937 9388
rect 6891 9000 6897 9376
rect 6931 9000 6937 9376
rect 6891 8988 6937 9000
rect 7004 9376 7050 9388
rect 7004 9000 7010 9376
rect 7044 9000 7050 9376
rect 7004 8988 7050 9000
rect 7122 9376 7168 9388
rect 7122 9000 7128 9376
rect 7162 9000 7168 9376
rect 7122 8988 7168 9000
rect 7240 9376 7286 9388
rect 7240 9000 7246 9376
rect 7280 9000 7286 9376
rect 7240 8988 7286 9000
rect 7358 9376 7404 9388
rect 7358 9000 7364 9376
rect 7398 9000 7404 9376
rect 7358 8988 7404 9000
rect 7476 9376 7522 9388
rect 7476 9000 7482 9376
rect 7516 9000 7522 9376
rect 7476 8988 7522 9000
rect 7594 9376 7640 9388
rect 7594 9000 7600 9376
rect 7634 9000 7640 9376
rect 7594 8988 7640 9000
rect 7712 9376 7758 9388
rect 7712 9000 7718 9376
rect 7752 9000 7758 9376
rect 7712 8988 7758 9000
rect 7831 9376 7877 9388
rect 7831 9000 7837 9376
rect 7871 9000 7877 9376
rect 7831 8988 7877 9000
rect 7949 9376 7995 9388
rect 7949 9000 7955 9376
rect 7989 9000 7995 9376
rect 7949 8988 7995 9000
rect 8067 9376 8113 9388
rect 8067 9000 8073 9376
rect 8107 9000 8113 9376
rect 8067 8988 8113 9000
rect 8185 9376 8231 9388
rect 8185 9000 8191 9376
rect 8225 9000 8231 9376
rect 8309 9188 8346 9475
rect 8185 8988 8231 9000
rect 8304 9176 8350 9188
rect 8304 9000 8310 9176
rect 8344 9000 8350 9176
rect 8304 8988 8350 9000
rect 8422 9176 8468 9188
rect 8422 9000 8428 9176
rect 8462 9000 8468 9176
rect 8422 8988 8468 9000
rect 8540 9176 8586 9188
rect 8540 9000 8546 9176
rect 8580 9000 8586 9176
rect 8540 8988 8586 9000
rect 8658 9176 8704 9188
rect 8658 9000 8664 9176
rect 8698 9000 8704 9176
rect 8658 8988 8704 9000
rect 6101 8802 6136 8988
rect 7010 8904 7044 8988
rect 8191 8904 8225 8988
rect 7010 8862 8225 8904
rect 8191 8842 8225 8862
rect 8191 8826 8548 8842
rect 6101 8785 7238 8802
rect 6101 8751 7188 8785
rect 7222 8751 7238 8785
rect 8191 8792 8498 8826
rect 8532 8792 8548 8826
rect 8191 8776 8548 8792
rect 6101 8735 7238 8751
rect 5520 8626 5702 8634
rect 5842 8690 6018 8698
rect 4379 8572 4444 8575
rect 4379 8569 4448 8572
rect 4379 8509 4385 8569
rect 4444 8509 4454 8569
rect 4379 8505 4448 8509
rect 4379 8503 4444 8505
rect 5520 8488 5701 8626
rect 5842 8622 5959 8690
rect 6016 8622 6026 8690
rect 5842 8614 6018 8622
rect 5947 8574 6018 8582
rect 5947 8506 5959 8574
rect 6016 8506 6026 8574
rect 5947 8498 6018 8506
rect 4014 8406 4106 8414
rect 4014 8341 4026 8406
rect 4094 8341 4106 8406
rect 4014 8329 4106 8341
rect 5520 8226 5555 8488
rect 2957 8178 4329 8225
rect 4651 8179 5555 8226
rect 5884 8406 6018 8414
rect 5884 8338 5959 8406
rect 6016 8338 6026 8406
rect 5884 8330 6018 8338
rect 3791 8055 3825 8178
rect 4263 8165 4329 8178
rect 4263 8131 4279 8165
rect 4313 8131 4329 8165
rect 4263 8115 4329 8131
rect 4652 8055 4686 8179
rect 3786 8043 3832 8055
rect 3786 7867 3792 8043
rect 3826 7867 3832 8043
rect 3786 7855 3832 7867
rect 3904 8043 4024 8055
rect 3904 7867 3910 8043
rect 3944 7867 3984 8043
rect 3904 7855 3984 7867
rect 3910 7488 3944 7855
rect 3978 7667 3984 7855
rect 4018 7667 4024 8043
rect 3978 7655 4024 7667
rect 4096 8043 4142 8055
rect 4096 7667 4102 8043
rect 4136 7667 4142 8043
rect 4096 7655 4142 7667
rect 4214 8043 4260 8055
rect 4214 7667 4220 8043
rect 4254 7667 4260 8043
rect 4214 7655 4260 7667
rect 4332 8043 4378 8055
rect 4332 7667 4338 8043
rect 4372 7667 4378 8043
rect 4332 7655 4378 7667
rect 4450 8043 4574 8055
rect 4450 7667 4456 8043
rect 4490 7867 4534 8043
rect 4568 7867 4574 8043
rect 4490 7855 4574 7867
rect 4646 8043 4692 8055
rect 4646 7867 4652 8043
rect 4686 7867 4692 8043
rect 4646 7855 4692 7867
rect 4490 7667 4496 7855
rect 4450 7655 4496 7667
rect 4220 7582 4254 7655
rect 4205 7566 4271 7582
rect 4205 7532 4221 7566
rect 4255 7532 4271 7566
rect 4205 7516 4271 7532
rect 4534 7488 4568 7855
rect 3910 7436 4568 7488
rect 4208 7414 4300 7436
rect 4208 7362 4220 7414
rect 4286 7362 4300 7414
rect 4208 7358 4300 7362
rect 5884 7008 5948 8330
rect 6101 8225 6136 8735
rect 6191 8689 6283 8702
rect 6191 8626 6203 8689
rect 6274 8626 6283 8689
rect 6191 8617 6283 8626
rect 7276 8689 7368 8699
rect 7276 8627 7288 8689
rect 7358 8627 7368 8689
rect 7276 8614 7368 8627
rect 8664 8634 8699 8988
rect 8774 8634 8845 9814
rect 9001 9814 11977 9875
rect 12152 9814 15122 9875
rect 15330 9815 18182 9876
rect 18498 9815 21467 9876
rect 9001 9812 9050 9814
rect 10472 9576 10482 9636
rect 10562 9576 10572 9636
rect 10472 9536 10572 9576
rect 9675 9479 11478 9536
rect 9675 9392 9709 9479
rect 10850 9392 10884 9479
rect 9669 9380 9715 9392
rect 9669 9192 9675 9380
rect 9228 9180 9274 9192
rect 9228 9004 9234 9180
rect 9268 9004 9274 9180
rect 9228 8992 9274 9004
rect 9346 9180 9392 9192
rect 9346 9004 9352 9180
rect 9386 9004 9392 9180
rect 9346 8992 9392 9004
rect 9464 9180 9510 9192
rect 9464 9004 9470 9180
rect 9504 9004 9510 9180
rect 9464 8992 9510 9004
rect 9582 9180 9675 9192
rect 9582 9004 9588 9180
rect 9622 9004 9675 9180
rect 9709 9004 9715 9380
rect 9582 8992 9715 9004
rect 9787 9380 9833 9392
rect 9787 9004 9793 9380
rect 9827 9004 9833 9380
rect 9787 8992 9833 9004
rect 9905 9380 9951 9392
rect 9905 9004 9911 9380
rect 9945 9004 9951 9380
rect 9905 8992 9951 9004
rect 10023 9380 10069 9392
rect 10023 9004 10029 9380
rect 10063 9004 10069 9380
rect 10023 8992 10069 9004
rect 10136 9380 10182 9392
rect 10136 9004 10142 9380
rect 10176 9004 10182 9380
rect 10136 8992 10182 9004
rect 10254 9380 10300 9392
rect 10254 9004 10260 9380
rect 10294 9004 10300 9380
rect 10254 8992 10300 9004
rect 10372 9380 10418 9392
rect 10372 9004 10378 9380
rect 10412 9004 10418 9380
rect 10372 8992 10418 9004
rect 10490 9380 10536 9392
rect 10490 9004 10496 9380
rect 10530 9004 10536 9380
rect 10490 8992 10536 9004
rect 10608 9380 10654 9392
rect 10608 9004 10614 9380
rect 10648 9004 10654 9380
rect 10608 8992 10654 9004
rect 10726 9380 10772 9392
rect 10726 9004 10732 9380
rect 10766 9004 10772 9380
rect 10726 8992 10772 9004
rect 10844 9380 10890 9392
rect 10844 9004 10850 9380
rect 10884 9004 10890 9380
rect 10844 8992 10890 9004
rect 10963 9380 11009 9392
rect 10963 9004 10969 9380
rect 11003 9004 11009 9380
rect 10963 8992 11009 9004
rect 11081 9380 11127 9392
rect 11081 9004 11087 9380
rect 11121 9004 11127 9380
rect 11081 8992 11127 9004
rect 11199 9380 11245 9392
rect 11199 9004 11205 9380
rect 11239 9004 11245 9380
rect 11199 8992 11245 9004
rect 11317 9380 11363 9392
rect 11317 9004 11323 9380
rect 11357 9004 11363 9380
rect 11441 9192 11478 9479
rect 11317 8992 11363 9004
rect 11436 9180 11482 9192
rect 11436 9004 11442 9180
rect 11476 9004 11482 9180
rect 11436 8992 11482 9004
rect 11554 9180 11600 9192
rect 11554 9004 11560 9180
rect 11594 9004 11600 9180
rect 11554 8992 11600 9004
rect 11672 9180 11718 9192
rect 11672 9004 11678 9180
rect 11712 9004 11718 9180
rect 11672 8992 11718 9004
rect 11790 9180 11836 9192
rect 11790 9004 11796 9180
rect 11830 9004 11836 9180
rect 11790 8992 11836 9004
rect 9233 8806 9268 8992
rect 10142 8908 10176 8992
rect 11323 8908 11357 8992
rect 10142 8866 11357 8908
rect 11323 8846 11357 8866
rect 11323 8830 11680 8846
rect 9233 8789 10370 8806
rect 9233 8755 10320 8789
rect 10354 8755 10370 8789
rect 11323 8796 11630 8830
rect 11664 8796 11680 8830
rect 11323 8780 11680 8796
rect 9233 8739 10370 8755
rect 7523 8572 7588 8575
rect 7523 8569 7592 8572
rect 7523 8509 7529 8569
rect 7588 8509 7598 8569
rect 7523 8505 7592 8509
rect 7523 8503 7588 8505
rect 8664 8488 8845 8634
rect 8974 8694 9150 8702
rect 8974 8626 9091 8694
rect 9148 8626 9158 8694
rect 8974 8618 9150 8626
rect 9079 8578 9150 8586
rect 9079 8510 9091 8578
rect 9148 8510 9158 8578
rect 9079 8502 9150 8510
rect 7158 8406 7250 8414
rect 7158 8341 7170 8406
rect 7238 8341 7250 8406
rect 7158 8329 7250 8341
rect 8664 8226 8699 8488
rect 8974 8410 9150 8418
rect 8974 8342 9091 8410
rect 9148 8342 9158 8410
rect 8974 8334 9150 8342
rect 6101 8178 7473 8225
rect 7795 8179 8699 8226
rect 6935 8055 6969 8178
rect 7407 8165 7473 8178
rect 7407 8131 7423 8165
rect 7457 8131 7473 8165
rect 7407 8115 7473 8131
rect 7796 8055 7830 8179
rect 6930 8043 6976 8055
rect 6930 7867 6936 8043
rect 6970 7867 6976 8043
rect 6930 7855 6976 7867
rect 7048 8043 7168 8055
rect 7048 7867 7054 8043
rect 7088 7867 7128 8043
rect 7048 7855 7128 7867
rect 7054 7488 7088 7855
rect 7122 7667 7128 7855
rect 7162 7667 7168 8043
rect 7122 7655 7168 7667
rect 7240 8043 7286 8055
rect 7240 7667 7246 8043
rect 7280 7667 7286 8043
rect 7240 7655 7286 7667
rect 7358 8043 7404 8055
rect 7358 7667 7364 8043
rect 7398 7667 7404 8043
rect 7358 7655 7404 7667
rect 7476 8043 7522 8055
rect 7476 7667 7482 8043
rect 7516 7667 7522 8043
rect 7476 7655 7522 7667
rect 7594 8043 7718 8055
rect 7594 7667 7600 8043
rect 7634 7867 7678 8043
rect 7712 7867 7718 8043
rect 7634 7855 7718 7867
rect 7790 8043 7836 8055
rect 7790 7867 7796 8043
rect 7830 7867 7836 8043
rect 7790 7855 7836 7867
rect 7634 7667 7640 7855
rect 7594 7655 7640 7667
rect 7364 7582 7398 7655
rect 7349 7566 7415 7582
rect 7349 7532 7365 7566
rect 7399 7532 7415 7566
rect 7349 7516 7415 7532
rect 7678 7488 7712 7855
rect 7054 7436 7712 7488
rect 7352 7414 7444 7436
rect 7352 7362 7364 7414
rect 7430 7362 7444 7414
rect 7352 7358 7444 7362
rect 9016 7244 9079 8334
rect 9233 8229 9268 8739
rect 9323 8693 9415 8706
rect 9323 8630 9335 8693
rect 9406 8630 9415 8693
rect 9323 8621 9415 8630
rect 10408 8693 10500 8703
rect 10408 8631 10420 8693
rect 10490 8631 10500 8693
rect 10408 8618 10500 8631
rect 11796 8638 11831 8992
rect 11906 8638 11977 9814
rect 13616 9576 13626 9636
rect 13706 9576 13716 9636
rect 13616 9536 13716 9576
rect 12819 9479 14622 9536
rect 12819 9392 12853 9479
rect 13994 9392 14028 9479
rect 12813 9380 12859 9392
rect 12813 9192 12819 9380
rect 12372 9180 12418 9192
rect 12372 9004 12378 9180
rect 12412 9004 12418 9180
rect 12372 8992 12418 9004
rect 12490 9180 12536 9192
rect 12490 9004 12496 9180
rect 12530 9004 12536 9180
rect 12490 8992 12536 9004
rect 12608 9180 12654 9192
rect 12608 9004 12614 9180
rect 12648 9004 12654 9180
rect 12608 8992 12654 9004
rect 12726 9180 12819 9192
rect 12726 9004 12732 9180
rect 12766 9004 12819 9180
rect 12853 9004 12859 9380
rect 12726 8992 12859 9004
rect 12931 9380 12977 9392
rect 12931 9004 12937 9380
rect 12971 9004 12977 9380
rect 12931 8992 12977 9004
rect 13049 9380 13095 9392
rect 13049 9004 13055 9380
rect 13089 9004 13095 9380
rect 13049 8992 13095 9004
rect 13167 9380 13213 9392
rect 13167 9004 13173 9380
rect 13207 9004 13213 9380
rect 13167 8992 13213 9004
rect 13280 9380 13326 9392
rect 13280 9004 13286 9380
rect 13320 9004 13326 9380
rect 13280 8992 13326 9004
rect 13398 9380 13444 9392
rect 13398 9004 13404 9380
rect 13438 9004 13444 9380
rect 13398 8992 13444 9004
rect 13516 9380 13562 9392
rect 13516 9004 13522 9380
rect 13556 9004 13562 9380
rect 13516 8992 13562 9004
rect 13634 9380 13680 9392
rect 13634 9004 13640 9380
rect 13674 9004 13680 9380
rect 13634 8992 13680 9004
rect 13752 9380 13798 9392
rect 13752 9004 13758 9380
rect 13792 9004 13798 9380
rect 13752 8992 13798 9004
rect 13870 9380 13916 9392
rect 13870 9004 13876 9380
rect 13910 9004 13916 9380
rect 13870 8992 13916 9004
rect 13988 9380 14034 9392
rect 13988 9004 13994 9380
rect 14028 9004 14034 9380
rect 13988 8992 14034 9004
rect 14107 9380 14153 9392
rect 14107 9004 14113 9380
rect 14147 9004 14153 9380
rect 14107 8992 14153 9004
rect 14225 9380 14271 9392
rect 14225 9004 14231 9380
rect 14265 9004 14271 9380
rect 14225 8992 14271 9004
rect 14343 9380 14389 9392
rect 14343 9004 14349 9380
rect 14383 9004 14389 9380
rect 14343 8992 14389 9004
rect 14461 9380 14507 9392
rect 14461 9004 14467 9380
rect 14501 9004 14507 9380
rect 14585 9192 14622 9479
rect 14461 8992 14507 9004
rect 14580 9180 14626 9192
rect 14580 9004 14586 9180
rect 14620 9004 14626 9180
rect 14580 8992 14626 9004
rect 14698 9180 14744 9192
rect 14698 9004 14704 9180
rect 14738 9004 14744 9180
rect 14698 8992 14744 9004
rect 14816 9180 14862 9192
rect 14816 9004 14822 9180
rect 14856 9004 14862 9180
rect 14816 8992 14862 9004
rect 14934 9180 14980 9192
rect 14934 9004 14940 9180
rect 14974 9004 14980 9180
rect 14934 8992 14980 9004
rect 12377 8806 12412 8992
rect 13286 8908 13320 8992
rect 14467 8908 14501 8992
rect 13286 8866 14501 8908
rect 14467 8846 14501 8866
rect 14467 8830 14824 8846
rect 12377 8789 13514 8806
rect 12377 8755 13464 8789
rect 13498 8755 13514 8789
rect 14467 8796 14774 8830
rect 14808 8796 14824 8830
rect 14467 8780 14824 8796
rect 12377 8739 13514 8755
rect 10655 8576 10720 8579
rect 10655 8573 10724 8576
rect 10655 8513 10661 8573
rect 10720 8513 10730 8573
rect 10655 8509 10724 8513
rect 10655 8507 10720 8509
rect 11796 8500 11977 8638
rect 12118 8694 12294 8702
rect 12118 8626 12235 8694
rect 12292 8626 12302 8694
rect 12118 8618 12294 8626
rect 12224 8578 12294 8586
rect 12224 8510 12235 8578
rect 12292 8510 12302 8578
rect 12224 8502 12294 8510
rect 10290 8410 10382 8418
rect 10290 8345 10302 8410
rect 10370 8345 10382 8410
rect 10290 8333 10382 8345
rect 11796 8230 11831 8500
rect 9233 8182 10605 8229
rect 10927 8183 11831 8230
rect 12176 8410 12294 8418
rect 12176 8342 12235 8410
rect 12292 8342 12302 8410
rect 12176 8334 12294 8342
rect 10067 8059 10101 8182
rect 10539 8169 10605 8182
rect 10539 8135 10555 8169
rect 10589 8135 10605 8169
rect 10539 8119 10605 8135
rect 10928 8059 10962 8183
rect 10062 8047 10108 8059
rect 10062 7871 10068 8047
rect 10102 7871 10108 8047
rect 10062 7859 10108 7871
rect 10180 8047 10300 8059
rect 10180 7871 10186 8047
rect 10220 7871 10260 8047
rect 10180 7859 10260 7871
rect 10186 7492 10220 7859
rect 10254 7671 10260 7859
rect 10294 7671 10300 8047
rect 10254 7659 10300 7671
rect 10372 8047 10418 8059
rect 10372 7671 10378 8047
rect 10412 7671 10418 8047
rect 10372 7659 10418 7671
rect 10490 8047 10536 8059
rect 10490 7671 10496 8047
rect 10530 7671 10536 8047
rect 10490 7659 10536 7671
rect 10608 8047 10654 8059
rect 10608 7671 10614 8047
rect 10648 7671 10654 8047
rect 10608 7659 10654 7671
rect 10726 8047 10850 8059
rect 10726 7671 10732 8047
rect 10766 7871 10810 8047
rect 10844 7871 10850 8047
rect 10766 7859 10850 7871
rect 10922 8047 10968 8059
rect 10922 7871 10928 8047
rect 10962 7871 10968 8047
rect 10922 7859 10968 7871
rect 10766 7671 10772 7859
rect 10726 7659 10772 7671
rect 10496 7586 10530 7659
rect 10481 7570 10547 7586
rect 10481 7536 10497 7570
rect 10531 7536 10547 7570
rect 10481 7520 10547 7536
rect 10810 7492 10844 7859
rect 10186 7440 10844 7492
rect 10484 7418 10576 7440
rect 10484 7366 10496 7418
rect 10562 7366 10576 7418
rect 10484 7362 10576 7366
rect 12176 7320 12224 8334
rect 12377 8229 12412 8739
rect 12467 8693 12559 8706
rect 12467 8630 12479 8693
rect 12550 8630 12559 8693
rect 12467 8621 12559 8630
rect 13552 8693 13644 8703
rect 13552 8631 13564 8693
rect 13634 8631 13644 8693
rect 13552 8618 13644 8631
rect 14940 8638 14975 8992
rect 15051 8638 15122 9814
rect 16818 9572 16828 9632
rect 16908 9572 16918 9632
rect 16818 9532 16918 9572
rect 16021 9475 17824 9532
rect 16021 9388 16055 9475
rect 17196 9388 17230 9475
rect 16015 9376 16061 9388
rect 16015 9188 16021 9376
rect 15574 9176 15620 9188
rect 15574 9000 15580 9176
rect 15614 9000 15620 9176
rect 15574 8988 15620 9000
rect 15692 9176 15738 9188
rect 15692 9000 15698 9176
rect 15732 9000 15738 9176
rect 15692 8988 15738 9000
rect 15810 9176 15856 9188
rect 15810 9000 15816 9176
rect 15850 9000 15856 9176
rect 15810 8988 15856 9000
rect 15928 9176 16021 9188
rect 15928 9000 15934 9176
rect 15968 9000 16021 9176
rect 16055 9000 16061 9376
rect 15928 8988 16061 9000
rect 16133 9376 16179 9388
rect 16133 9000 16139 9376
rect 16173 9000 16179 9376
rect 16133 8988 16179 9000
rect 16251 9376 16297 9388
rect 16251 9000 16257 9376
rect 16291 9000 16297 9376
rect 16251 8988 16297 9000
rect 16369 9376 16415 9388
rect 16369 9000 16375 9376
rect 16409 9000 16415 9376
rect 16369 8988 16415 9000
rect 16482 9376 16528 9388
rect 16482 9000 16488 9376
rect 16522 9000 16528 9376
rect 16482 8988 16528 9000
rect 16600 9376 16646 9388
rect 16600 9000 16606 9376
rect 16640 9000 16646 9376
rect 16600 8988 16646 9000
rect 16718 9376 16764 9388
rect 16718 9000 16724 9376
rect 16758 9000 16764 9376
rect 16718 8988 16764 9000
rect 16836 9376 16882 9388
rect 16836 9000 16842 9376
rect 16876 9000 16882 9376
rect 16836 8988 16882 9000
rect 16954 9376 17000 9388
rect 16954 9000 16960 9376
rect 16994 9000 17000 9376
rect 16954 8988 17000 9000
rect 17072 9376 17118 9388
rect 17072 9000 17078 9376
rect 17112 9000 17118 9376
rect 17072 8988 17118 9000
rect 17190 9376 17236 9388
rect 17190 9000 17196 9376
rect 17230 9000 17236 9376
rect 17190 8988 17236 9000
rect 17309 9376 17355 9388
rect 17309 9000 17315 9376
rect 17349 9000 17355 9376
rect 17309 8988 17355 9000
rect 17427 9376 17473 9388
rect 17427 9000 17433 9376
rect 17467 9000 17473 9376
rect 17427 8988 17473 9000
rect 17545 9376 17591 9388
rect 17545 9000 17551 9376
rect 17585 9000 17591 9376
rect 17545 8988 17591 9000
rect 17663 9376 17709 9388
rect 17663 9000 17669 9376
rect 17703 9000 17709 9376
rect 17787 9188 17824 9475
rect 17663 8988 17709 9000
rect 17782 9176 17828 9188
rect 17782 9000 17788 9176
rect 17822 9000 17828 9176
rect 17782 8988 17828 9000
rect 17900 9176 17946 9188
rect 17900 9000 17906 9176
rect 17940 9000 17946 9176
rect 17900 8988 17946 9000
rect 18018 9176 18064 9188
rect 18018 9000 18024 9176
rect 18058 9000 18064 9176
rect 18018 8988 18064 9000
rect 18136 9176 18182 9815
rect 19962 9572 19972 9632
rect 20052 9572 20062 9632
rect 19962 9532 20062 9572
rect 19165 9475 20968 9532
rect 19165 9388 19199 9475
rect 20340 9388 20374 9475
rect 19159 9376 19205 9388
rect 19159 9188 19165 9376
rect 18136 9000 18142 9176
rect 18176 9000 18182 9176
rect 18136 8988 18182 9000
rect 18718 9176 18764 9188
rect 18718 9000 18724 9176
rect 18758 9000 18764 9176
rect 18718 8988 18764 9000
rect 18836 9176 18882 9188
rect 18836 9000 18842 9176
rect 18876 9000 18882 9176
rect 18836 8988 18882 9000
rect 18954 9176 19000 9188
rect 18954 9000 18960 9176
rect 18994 9000 19000 9176
rect 18954 8988 19000 9000
rect 19072 9176 19165 9188
rect 19072 9000 19078 9176
rect 19112 9000 19165 9176
rect 19199 9000 19205 9376
rect 19072 8988 19205 9000
rect 19277 9376 19323 9388
rect 19277 9000 19283 9376
rect 19317 9000 19323 9376
rect 19277 8988 19323 9000
rect 19395 9376 19441 9388
rect 19395 9000 19401 9376
rect 19435 9000 19441 9376
rect 19395 8988 19441 9000
rect 19513 9376 19559 9388
rect 19513 9000 19519 9376
rect 19553 9000 19559 9376
rect 19513 8988 19559 9000
rect 19626 9376 19672 9388
rect 19626 9000 19632 9376
rect 19666 9000 19672 9376
rect 19626 8988 19672 9000
rect 19744 9376 19790 9388
rect 19744 9000 19750 9376
rect 19784 9000 19790 9376
rect 19744 8988 19790 9000
rect 19862 9376 19908 9388
rect 19862 9000 19868 9376
rect 19902 9000 19908 9376
rect 19862 8988 19908 9000
rect 19980 9376 20026 9388
rect 19980 9000 19986 9376
rect 20020 9000 20026 9376
rect 19980 8988 20026 9000
rect 20098 9376 20144 9388
rect 20098 9000 20104 9376
rect 20138 9000 20144 9376
rect 20098 8988 20144 9000
rect 20216 9376 20262 9388
rect 20216 9000 20222 9376
rect 20256 9000 20262 9376
rect 20216 8988 20262 9000
rect 20334 9376 20380 9388
rect 20334 9000 20340 9376
rect 20374 9000 20380 9376
rect 20334 8988 20380 9000
rect 20453 9376 20499 9388
rect 20453 9000 20459 9376
rect 20493 9000 20499 9376
rect 20453 8988 20499 9000
rect 20571 9376 20617 9388
rect 20571 9000 20577 9376
rect 20611 9000 20617 9376
rect 20571 8988 20617 9000
rect 20689 9376 20735 9388
rect 20689 9000 20695 9376
rect 20729 9000 20735 9376
rect 20689 8988 20735 9000
rect 20807 9376 20853 9388
rect 20807 9000 20813 9376
rect 20847 9000 20853 9376
rect 20931 9188 20968 9475
rect 20807 8988 20853 9000
rect 20926 9176 20972 9188
rect 20926 9000 20932 9176
rect 20966 9000 20972 9176
rect 20926 8988 20972 9000
rect 21044 9176 21090 9188
rect 21044 9000 21050 9176
rect 21084 9000 21090 9176
rect 21044 8988 21090 9000
rect 21162 9176 21208 9188
rect 21162 9000 21168 9176
rect 21202 9000 21208 9176
rect 21162 8988 21208 9000
rect 21280 9176 21326 9188
rect 21280 9000 21286 9176
rect 21320 9000 21326 9176
rect 21280 8988 21326 9000
rect 15579 8802 15614 8988
rect 16488 8904 16522 8988
rect 17669 8904 17703 8988
rect 16488 8862 17703 8904
rect 17669 8842 17703 8862
rect 17669 8826 18026 8842
rect 15579 8785 16716 8802
rect 15579 8751 16666 8785
rect 16700 8751 16716 8785
rect 17669 8792 17976 8826
rect 18010 8792 18026 8826
rect 17669 8776 18026 8792
rect 15579 8735 16716 8751
rect 15320 8690 15496 8698
rect 13799 8576 13864 8579
rect 13799 8573 13868 8576
rect 13799 8513 13805 8573
rect 13864 8513 13874 8573
rect 13799 8509 13868 8513
rect 13799 8507 13864 8509
rect 14940 8492 15121 8638
rect 15320 8622 15437 8690
rect 15494 8622 15504 8690
rect 15320 8614 15496 8622
rect 15426 8574 15496 8582
rect 15426 8506 15437 8574
rect 15494 8506 15504 8574
rect 15426 8498 15496 8506
rect 13434 8410 13526 8418
rect 13434 8345 13446 8410
rect 13514 8345 13526 8410
rect 13434 8333 13526 8345
rect 14940 8230 14975 8492
rect 12377 8182 13749 8229
rect 14071 8183 14975 8230
rect 15380 8406 15496 8414
rect 15380 8338 15437 8406
rect 15494 8338 15504 8406
rect 15380 8330 15496 8338
rect 13211 8059 13245 8182
rect 13683 8169 13749 8182
rect 13683 8135 13699 8169
rect 13733 8135 13749 8169
rect 13683 8119 13749 8135
rect 14072 8059 14106 8183
rect 13206 8047 13252 8059
rect 13206 7871 13212 8047
rect 13246 7871 13252 8047
rect 13206 7859 13252 7871
rect 13324 8047 13444 8059
rect 13324 7871 13330 8047
rect 13364 7871 13404 8047
rect 13324 7859 13404 7871
rect 13330 7492 13364 7859
rect 13398 7671 13404 7859
rect 13438 7671 13444 8047
rect 13398 7659 13444 7671
rect 13516 8047 13562 8059
rect 13516 7671 13522 8047
rect 13556 7671 13562 8047
rect 13516 7659 13562 7671
rect 13634 8047 13680 8059
rect 13634 7671 13640 8047
rect 13674 7671 13680 8047
rect 13634 7659 13680 7671
rect 13752 8047 13798 8059
rect 13752 7671 13758 8047
rect 13792 7671 13798 8047
rect 13752 7659 13798 7671
rect 13870 8047 13994 8059
rect 13870 7671 13876 8047
rect 13910 7871 13954 8047
rect 13988 7871 13994 8047
rect 13910 7859 13994 7871
rect 14066 8047 14112 8059
rect 14066 7871 14072 8047
rect 14106 7871 14112 8047
rect 14066 7859 14112 7871
rect 13910 7671 13916 7859
rect 13870 7659 13916 7671
rect 13640 7586 13674 7659
rect 13625 7570 13691 7586
rect 13625 7536 13641 7570
rect 13675 7536 13691 7570
rect 13625 7520 13691 7536
rect 13954 7492 13988 7859
rect 13330 7440 13988 7492
rect 13628 7418 13720 7440
rect 13628 7366 13640 7418
rect 13706 7366 13720 7418
rect 13628 7362 13720 7366
rect 15380 7323 15428 8330
rect 15579 8225 15614 8735
rect 15669 8689 15761 8702
rect 15669 8626 15681 8689
rect 15752 8626 15761 8689
rect 15669 8617 15761 8626
rect 16754 8689 16846 8699
rect 16754 8627 16766 8689
rect 16836 8627 16846 8689
rect 16754 8614 16846 8627
rect 17001 8572 17066 8575
rect 17001 8569 17070 8572
rect 17001 8509 17007 8569
rect 17066 8509 17076 8569
rect 17001 8505 17070 8509
rect 17001 8503 17066 8505
rect 16636 8406 16728 8414
rect 16636 8341 16648 8406
rect 16716 8341 16728 8406
rect 16636 8329 16728 8341
rect 18142 8226 18177 8988
rect 18723 8802 18758 8988
rect 19632 8904 19666 8988
rect 20813 8904 20847 8988
rect 19632 8862 20847 8904
rect 20813 8842 20847 8862
rect 20813 8826 21170 8842
rect 18723 8785 19860 8802
rect 18723 8751 19810 8785
rect 19844 8751 19860 8785
rect 20813 8792 21120 8826
rect 21154 8792 21170 8826
rect 20813 8776 21170 8792
rect 18723 8735 19860 8751
rect 18464 8690 18640 8698
rect 18464 8622 18581 8690
rect 18638 8622 18648 8690
rect 18464 8614 18640 8622
rect 18569 8574 18640 8582
rect 18569 8506 18581 8574
rect 18638 8506 18648 8574
rect 18569 8498 18640 8506
rect 18522 8414 18570 8415
rect 18521 8406 18640 8414
rect 18521 8338 18581 8406
rect 18638 8338 18648 8406
rect 18521 8330 18640 8338
rect 15579 8178 16951 8225
rect 17273 8179 18177 8226
rect 16413 8055 16447 8178
rect 16885 8165 16951 8178
rect 16885 8131 16901 8165
rect 16935 8131 16951 8165
rect 16885 8115 16951 8131
rect 17274 8055 17308 8179
rect 16408 8043 16454 8055
rect 16408 7867 16414 8043
rect 16448 7867 16454 8043
rect 16408 7855 16454 7867
rect 16526 8043 16646 8055
rect 16526 7867 16532 8043
rect 16566 7867 16606 8043
rect 16526 7855 16606 7867
rect 16532 7488 16566 7855
rect 16600 7667 16606 7855
rect 16640 7667 16646 8043
rect 16600 7655 16646 7667
rect 16718 8043 16764 8055
rect 16718 7667 16724 8043
rect 16758 7667 16764 8043
rect 16718 7655 16764 7667
rect 16836 8043 16882 8055
rect 16836 7667 16842 8043
rect 16876 7667 16882 8043
rect 16836 7655 16882 7667
rect 16954 8043 17000 8055
rect 16954 7667 16960 8043
rect 16994 7667 17000 8043
rect 16954 7655 17000 7667
rect 17072 8043 17196 8055
rect 17072 7667 17078 8043
rect 17112 7867 17156 8043
rect 17190 7867 17196 8043
rect 17112 7855 17196 7867
rect 17268 8043 17314 8055
rect 17268 7867 17274 8043
rect 17308 7867 17314 8043
rect 17268 7855 17314 7867
rect 17112 7667 17118 7855
rect 17072 7655 17118 7667
rect 16842 7582 16876 7655
rect 16827 7566 16893 7582
rect 16827 7532 16843 7566
rect 16877 7532 16893 7566
rect 16827 7516 16893 7532
rect 17156 7488 17190 7855
rect 16532 7436 17190 7488
rect 16830 7414 16922 7436
rect 16830 7362 16842 7414
rect 16908 7362 16922 7414
rect 16830 7358 16922 7362
rect 18522 7323 18570 8330
rect 18723 8225 18758 8735
rect 18813 8689 18905 8702
rect 18813 8626 18825 8689
rect 18896 8626 18905 8689
rect 18813 8617 18905 8626
rect 19898 8689 19990 8699
rect 19898 8627 19910 8689
rect 19980 8627 19990 8689
rect 19898 8614 19990 8627
rect 21286 8634 21321 8988
rect 21396 8634 21467 9815
rect 21614 9875 21694 11066
rect 21865 10961 21900 11471
rect 21955 11425 22047 11438
rect 21955 11362 21967 11425
rect 22038 11362 22047 11425
rect 21955 11353 22047 11362
rect 23040 11425 23132 11435
rect 23040 11363 23052 11425
rect 23122 11363 23132 11425
rect 23040 11350 23132 11363
rect 24428 11370 24463 11724
rect 23287 11308 23352 11311
rect 23287 11305 23356 11308
rect 23287 11245 23293 11305
rect 23352 11245 23362 11305
rect 23287 11241 23356 11245
rect 23287 11239 23352 11241
rect 24428 11224 24609 11370
rect 24750 11318 24821 12637
rect 26248 12308 26258 12368
rect 26338 12308 26348 12368
rect 26248 12268 26348 12308
rect 25451 12211 27254 12268
rect 25451 12124 25485 12211
rect 26626 12124 26660 12211
rect 25445 12112 25491 12124
rect 25445 11924 25451 12112
rect 25004 11912 25050 11924
rect 25004 11736 25010 11912
rect 25044 11736 25050 11912
rect 25004 11724 25050 11736
rect 25122 11912 25168 11924
rect 25122 11736 25128 11912
rect 25162 11736 25168 11912
rect 25122 11724 25168 11736
rect 25240 11912 25286 11924
rect 25240 11736 25246 11912
rect 25280 11736 25286 11912
rect 25240 11724 25286 11736
rect 25358 11912 25451 11924
rect 25358 11736 25364 11912
rect 25398 11736 25451 11912
rect 25485 11736 25491 12112
rect 25358 11724 25491 11736
rect 25563 12112 25609 12124
rect 25563 11736 25569 12112
rect 25603 11736 25609 12112
rect 25563 11724 25609 11736
rect 25681 12112 25727 12124
rect 25681 11736 25687 12112
rect 25721 11736 25727 12112
rect 25681 11724 25727 11736
rect 25799 12112 25845 12124
rect 25799 11736 25805 12112
rect 25839 11736 25845 12112
rect 25799 11724 25845 11736
rect 25912 12112 25958 12124
rect 25912 11736 25918 12112
rect 25952 11736 25958 12112
rect 25912 11724 25958 11736
rect 26030 12112 26076 12124
rect 26030 11736 26036 12112
rect 26070 11736 26076 12112
rect 26030 11724 26076 11736
rect 26148 12112 26194 12124
rect 26148 11736 26154 12112
rect 26188 11736 26194 12112
rect 26148 11724 26194 11736
rect 26266 12112 26312 12124
rect 26266 11736 26272 12112
rect 26306 11736 26312 12112
rect 26266 11724 26312 11736
rect 26384 12112 26430 12124
rect 26384 11736 26390 12112
rect 26424 11736 26430 12112
rect 26384 11724 26430 11736
rect 26502 12112 26548 12124
rect 26502 11736 26508 12112
rect 26542 11736 26548 12112
rect 26502 11724 26548 11736
rect 26620 12112 26666 12124
rect 26620 11736 26626 12112
rect 26660 11736 26666 12112
rect 26620 11724 26666 11736
rect 26739 12112 26785 12124
rect 26739 11736 26745 12112
rect 26779 11736 26785 12112
rect 26739 11724 26785 11736
rect 26857 12112 26903 12124
rect 26857 11736 26863 12112
rect 26897 11736 26903 12112
rect 26857 11724 26903 11736
rect 26975 12112 27021 12124
rect 26975 11736 26981 12112
rect 27015 11736 27021 12112
rect 26975 11724 27021 11736
rect 27093 12112 27139 12124
rect 27093 11736 27099 12112
rect 27133 11736 27139 12112
rect 27217 11924 27254 12211
rect 27093 11724 27139 11736
rect 27212 11912 27258 11924
rect 27212 11736 27218 11912
rect 27252 11736 27258 11912
rect 27212 11724 27258 11736
rect 27330 11912 27376 11924
rect 27330 11736 27336 11912
rect 27370 11736 27376 11912
rect 27330 11724 27376 11736
rect 27448 11912 27494 11924
rect 27448 11736 27454 11912
rect 27488 11736 27494 11912
rect 27448 11724 27494 11736
rect 27566 11912 27612 11924
rect 27566 11736 27572 11912
rect 27606 11736 27612 11912
rect 27566 11724 27612 11736
rect 25009 11538 25044 11724
rect 25918 11640 25952 11724
rect 27099 11640 27133 11724
rect 25918 11598 27133 11640
rect 27099 11578 27133 11598
rect 27099 11562 27456 11578
rect 25009 11521 26146 11538
rect 25009 11487 26096 11521
rect 26130 11487 26146 11521
rect 27099 11528 27406 11562
rect 27440 11528 27456 11562
rect 27099 11512 27456 11528
rect 25009 11471 26146 11487
rect 24750 11310 24926 11318
rect 24750 11242 24867 11310
rect 24924 11242 24934 11310
rect 24750 11234 24926 11242
rect 22922 11142 23014 11150
rect 22922 11077 22934 11142
rect 23002 11077 23014 11142
rect 22922 11065 23014 11077
rect 24428 10962 24463 11224
rect 21865 10914 23237 10961
rect 23559 10915 24463 10962
rect 24513 10930 24609 11224
rect 22699 10791 22733 10914
rect 23171 10901 23237 10914
rect 23171 10867 23187 10901
rect 23221 10867 23237 10901
rect 23171 10851 23237 10867
rect 23560 10791 23594 10915
rect 24513 10859 24525 10930
rect 24596 10859 24609 10930
rect 24513 10849 24609 10859
rect 24798 11142 24926 11150
rect 24798 11074 24867 11142
rect 24924 11074 24934 11142
rect 24798 11066 24926 11074
rect 22694 10779 22740 10791
rect 22694 10603 22700 10779
rect 22734 10603 22740 10779
rect 22694 10591 22740 10603
rect 22812 10779 22932 10791
rect 22812 10603 22818 10779
rect 22852 10603 22892 10779
rect 22812 10591 22892 10603
rect 22818 10224 22852 10591
rect 22886 10403 22892 10591
rect 22926 10403 22932 10779
rect 22886 10391 22932 10403
rect 23004 10779 23050 10791
rect 23004 10403 23010 10779
rect 23044 10403 23050 10779
rect 23004 10391 23050 10403
rect 23122 10779 23168 10791
rect 23122 10403 23128 10779
rect 23162 10403 23168 10779
rect 23122 10391 23168 10403
rect 23240 10779 23286 10791
rect 23240 10403 23246 10779
rect 23280 10403 23286 10779
rect 23240 10391 23286 10403
rect 23358 10779 23482 10791
rect 23358 10403 23364 10779
rect 23398 10603 23442 10779
rect 23476 10603 23482 10779
rect 23398 10591 23482 10603
rect 23554 10779 23600 10791
rect 23554 10603 23560 10779
rect 23594 10603 23600 10779
rect 23554 10591 23600 10603
rect 23398 10403 23404 10591
rect 23358 10391 23404 10403
rect 23128 10318 23162 10391
rect 23113 10302 23179 10318
rect 23113 10268 23129 10302
rect 23163 10268 23179 10302
rect 23113 10252 23179 10268
rect 23442 10224 23476 10591
rect 22818 10172 23476 10224
rect 23116 10150 23208 10172
rect 23116 10098 23128 10150
rect 23194 10098 23208 10150
rect 23116 10094 23208 10098
rect 24798 9875 24849 11066
rect 25009 10961 25044 11471
rect 25099 11425 25191 11438
rect 25099 11362 25111 11425
rect 25182 11362 25191 11425
rect 25099 11353 25191 11362
rect 26184 11425 26276 11435
rect 26184 11363 26196 11425
rect 26266 11363 26276 11425
rect 26184 11350 26276 11363
rect 27572 11370 27607 11724
rect 26431 11308 26496 11311
rect 26431 11305 26500 11308
rect 26431 11245 26437 11305
rect 26496 11245 26506 11305
rect 26431 11241 26500 11245
rect 26431 11239 26496 11241
rect 27572 11224 28052 11370
rect 26066 11142 26158 11150
rect 26066 11077 26078 11142
rect 26146 11077 26158 11142
rect 26066 11065 26158 11077
rect 27572 10962 27607 11224
rect 25009 10914 26381 10961
rect 26703 10915 27607 10962
rect 27948 10937 28052 10947
rect 25843 10791 25877 10914
rect 26315 10901 26381 10914
rect 26315 10867 26331 10901
rect 26365 10867 26381 10901
rect 26315 10851 26381 10867
rect 26704 10791 26738 10915
rect 27905 10867 27915 10937
rect 27974 10867 28052 10937
rect 27948 10859 28052 10867
rect 25838 10779 25884 10791
rect 25838 10603 25844 10779
rect 25878 10603 25884 10779
rect 25838 10591 25884 10603
rect 25956 10779 26076 10791
rect 25956 10603 25962 10779
rect 25996 10603 26036 10779
rect 25956 10591 26036 10603
rect 25962 10224 25996 10591
rect 26030 10403 26036 10591
rect 26070 10403 26076 10779
rect 26030 10391 26076 10403
rect 26148 10779 26194 10791
rect 26148 10403 26154 10779
rect 26188 10403 26194 10779
rect 26148 10391 26194 10403
rect 26266 10779 26312 10791
rect 26266 10403 26272 10779
rect 26306 10403 26312 10779
rect 26266 10391 26312 10403
rect 26384 10779 26430 10791
rect 26384 10403 26390 10779
rect 26424 10403 26430 10779
rect 26384 10391 26430 10403
rect 26502 10779 26626 10791
rect 26502 10403 26508 10779
rect 26542 10603 26586 10779
rect 26620 10603 26626 10779
rect 26542 10591 26626 10603
rect 26698 10779 26744 10791
rect 26698 10603 26704 10779
rect 26738 10603 26744 10779
rect 27903 10745 28052 10758
rect 27903 10682 27914 10745
rect 27975 10682 28052 10745
rect 27903 10672 28052 10682
rect 26698 10591 26744 10603
rect 26542 10403 26548 10591
rect 26502 10391 26548 10403
rect 26272 10318 26306 10391
rect 26257 10302 26323 10318
rect 26257 10268 26273 10302
rect 26307 10268 26323 10302
rect 26257 10252 26323 10268
rect 26586 10224 26620 10591
rect 27901 10525 28052 10542
rect 27901 10459 27913 10525
rect 27975 10459 28052 10525
rect 27901 10447 28052 10459
rect 27903 10329 28053 10346
rect 27903 10271 27913 10329
rect 27976 10271 28053 10329
rect 27903 10260 28053 10271
rect 25962 10172 26620 10224
rect 26260 10150 26352 10172
rect 26260 10098 26272 10150
rect 26338 10098 26352 10150
rect 26260 10094 26352 10098
rect 27901 9986 28054 10004
rect 27901 9925 27912 9986
rect 27976 9925 28054 9986
rect 27901 9914 28054 9925
rect 21614 9814 24599 9875
rect 23094 9576 23104 9636
rect 23184 9576 23194 9636
rect 23094 9536 23194 9576
rect 22297 9479 24100 9536
rect 22297 9392 22331 9479
rect 23472 9392 23506 9479
rect 22291 9380 22337 9392
rect 22291 9192 22297 9380
rect 21850 9180 21896 9192
rect 21850 9004 21856 9180
rect 21890 9004 21896 9180
rect 21850 8992 21896 9004
rect 21968 9180 22014 9192
rect 21968 9004 21974 9180
rect 22008 9004 22014 9180
rect 21968 8992 22014 9004
rect 22086 9180 22132 9192
rect 22086 9004 22092 9180
rect 22126 9004 22132 9180
rect 22086 8992 22132 9004
rect 22204 9180 22297 9192
rect 22204 9004 22210 9180
rect 22244 9004 22297 9180
rect 22331 9004 22337 9380
rect 22204 8992 22337 9004
rect 22409 9380 22455 9392
rect 22409 9004 22415 9380
rect 22449 9004 22455 9380
rect 22409 8992 22455 9004
rect 22527 9380 22573 9392
rect 22527 9004 22533 9380
rect 22567 9004 22573 9380
rect 22527 8992 22573 9004
rect 22645 9380 22691 9392
rect 22645 9004 22651 9380
rect 22685 9004 22691 9380
rect 22645 8992 22691 9004
rect 22758 9380 22804 9392
rect 22758 9004 22764 9380
rect 22798 9004 22804 9380
rect 22758 8992 22804 9004
rect 22876 9380 22922 9392
rect 22876 9004 22882 9380
rect 22916 9004 22922 9380
rect 22876 8992 22922 9004
rect 22994 9380 23040 9392
rect 22994 9004 23000 9380
rect 23034 9004 23040 9380
rect 22994 8992 23040 9004
rect 23112 9380 23158 9392
rect 23112 9004 23118 9380
rect 23152 9004 23158 9380
rect 23112 8992 23158 9004
rect 23230 9380 23276 9392
rect 23230 9004 23236 9380
rect 23270 9004 23276 9380
rect 23230 8992 23276 9004
rect 23348 9380 23394 9392
rect 23348 9004 23354 9380
rect 23388 9004 23394 9380
rect 23348 8992 23394 9004
rect 23466 9380 23512 9392
rect 23466 9004 23472 9380
rect 23506 9004 23512 9380
rect 23466 8992 23512 9004
rect 23585 9380 23631 9392
rect 23585 9004 23591 9380
rect 23625 9004 23631 9380
rect 23585 8992 23631 9004
rect 23703 9380 23749 9392
rect 23703 9004 23709 9380
rect 23743 9004 23749 9380
rect 23703 8992 23749 9004
rect 23821 9380 23867 9392
rect 23821 9004 23827 9380
rect 23861 9004 23867 9380
rect 23821 8992 23867 9004
rect 23939 9380 23985 9392
rect 23939 9004 23945 9380
rect 23979 9004 23985 9380
rect 24063 9192 24100 9479
rect 23939 8992 23985 9004
rect 24058 9180 24104 9192
rect 24058 9004 24064 9180
rect 24098 9004 24104 9180
rect 24058 8992 24104 9004
rect 24176 9180 24222 9192
rect 24176 9004 24182 9180
rect 24216 9004 24222 9180
rect 24176 8992 24222 9004
rect 24294 9180 24340 9192
rect 24294 9004 24300 9180
rect 24334 9004 24340 9180
rect 24294 8992 24340 9004
rect 24412 9180 24458 9192
rect 24412 9004 24418 9180
rect 24452 9004 24458 9180
rect 24412 8992 24458 9004
rect 21855 8806 21890 8992
rect 22764 8908 22798 8992
rect 23945 8908 23979 8992
rect 22764 8866 23979 8908
rect 23945 8846 23979 8866
rect 23945 8830 24302 8846
rect 21855 8789 22992 8806
rect 21855 8755 22942 8789
rect 22976 8755 22992 8789
rect 23945 8796 24252 8830
rect 24286 8796 24302 8830
rect 23945 8780 24302 8796
rect 21855 8739 22992 8755
rect 20145 8572 20210 8575
rect 20145 8569 20214 8572
rect 20145 8509 20151 8569
rect 20210 8509 20220 8569
rect 20145 8505 20214 8509
rect 20145 8503 20210 8505
rect 21286 8488 21467 8634
rect 21596 8694 21772 8702
rect 21596 8626 21713 8694
rect 21770 8626 21780 8694
rect 21596 8618 21772 8626
rect 21702 8578 21772 8586
rect 21702 8510 21713 8578
rect 21770 8510 21780 8578
rect 21702 8502 21772 8510
rect 19780 8406 19872 8414
rect 19780 8341 19792 8406
rect 19860 8341 19872 8406
rect 19780 8329 19872 8341
rect 21286 8226 21321 8488
rect 18723 8178 20095 8225
rect 20417 8179 21321 8226
rect 21653 8410 21772 8418
rect 21653 8342 21713 8410
rect 21770 8342 21780 8410
rect 21653 8334 21772 8342
rect 19557 8055 19591 8178
rect 20029 8165 20095 8178
rect 20029 8131 20045 8165
rect 20079 8131 20095 8165
rect 20029 8115 20095 8131
rect 20418 8055 20452 8179
rect 19552 8043 19598 8055
rect 19552 7867 19558 8043
rect 19592 7867 19598 8043
rect 19552 7855 19598 7867
rect 19670 8043 19790 8055
rect 19670 7867 19676 8043
rect 19710 7867 19750 8043
rect 19670 7855 19750 7867
rect 19676 7488 19710 7855
rect 19744 7667 19750 7855
rect 19784 7667 19790 8043
rect 19744 7655 19790 7667
rect 19862 8043 19908 8055
rect 19862 7667 19868 8043
rect 19902 7667 19908 8043
rect 19862 7655 19908 7667
rect 19980 8043 20026 8055
rect 19980 7667 19986 8043
rect 20020 7667 20026 8043
rect 19980 7655 20026 7667
rect 20098 8043 20144 8055
rect 20098 7667 20104 8043
rect 20138 7667 20144 8043
rect 20098 7655 20144 7667
rect 20216 8043 20340 8055
rect 20216 7667 20222 8043
rect 20256 7867 20300 8043
rect 20334 7867 20340 8043
rect 20256 7855 20340 7867
rect 20412 8043 20458 8055
rect 20412 7867 20418 8043
rect 20452 7867 20458 8043
rect 20412 7855 20458 7867
rect 20256 7667 20262 7855
rect 20216 7655 20262 7667
rect 19986 7582 20020 7655
rect 19971 7566 20037 7582
rect 19971 7532 19987 7566
rect 20021 7532 20037 7566
rect 19971 7516 20037 7532
rect 20300 7488 20334 7855
rect 19676 7436 20334 7488
rect 19974 7414 20066 7436
rect 19974 7362 19986 7414
rect 20052 7362 20066 7414
rect 19974 7358 20066 7362
rect 21653 7326 21701 8334
rect 21855 8229 21890 8739
rect 21945 8693 22037 8706
rect 21945 8630 21957 8693
rect 22028 8630 22037 8693
rect 21945 8621 22037 8630
rect 23030 8693 23122 8703
rect 23030 8631 23042 8693
rect 23112 8631 23122 8693
rect 23030 8618 23122 8631
rect 24418 8638 24453 8992
rect 24528 8638 24599 9814
rect 24798 9874 26152 9875
rect 24798 9813 27602 9874
rect 26238 9576 26248 9636
rect 26328 9576 26338 9636
rect 26238 9536 26338 9576
rect 25441 9479 27244 9536
rect 25441 9392 25475 9479
rect 26616 9392 26650 9479
rect 25435 9380 25481 9392
rect 25435 9192 25441 9380
rect 24994 9180 25040 9192
rect 24994 9004 25000 9180
rect 25034 9004 25040 9180
rect 24994 8992 25040 9004
rect 25112 9180 25158 9192
rect 25112 9004 25118 9180
rect 25152 9004 25158 9180
rect 25112 8992 25158 9004
rect 25230 9180 25276 9192
rect 25230 9004 25236 9180
rect 25270 9004 25276 9180
rect 25230 8992 25276 9004
rect 25348 9180 25441 9192
rect 25348 9004 25354 9180
rect 25388 9004 25441 9180
rect 25475 9004 25481 9380
rect 25348 8992 25481 9004
rect 25553 9380 25599 9392
rect 25553 9004 25559 9380
rect 25593 9004 25599 9380
rect 25553 8992 25599 9004
rect 25671 9380 25717 9392
rect 25671 9004 25677 9380
rect 25711 9004 25717 9380
rect 25671 8992 25717 9004
rect 25789 9380 25835 9392
rect 25789 9004 25795 9380
rect 25829 9004 25835 9380
rect 25789 8992 25835 9004
rect 25902 9380 25948 9392
rect 25902 9004 25908 9380
rect 25942 9004 25948 9380
rect 25902 8992 25948 9004
rect 26020 9380 26066 9392
rect 26020 9004 26026 9380
rect 26060 9004 26066 9380
rect 26020 8992 26066 9004
rect 26138 9380 26184 9392
rect 26138 9004 26144 9380
rect 26178 9004 26184 9380
rect 26138 8992 26184 9004
rect 26256 9380 26302 9392
rect 26256 9004 26262 9380
rect 26296 9004 26302 9380
rect 26256 8992 26302 9004
rect 26374 9380 26420 9392
rect 26374 9004 26380 9380
rect 26414 9004 26420 9380
rect 26374 8992 26420 9004
rect 26492 9380 26538 9392
rect 26492 9004 26498 9380
rect 26532 9004 26538 9380
rect 26492 8992 26538 9004
rect 26610 9380 26656 9392
rect 26610 9004 26616 9380
rect 26650 9004 26656 9380
rect 26610 8992 26656 9004
rect 26729 9380 26775 9392
rect 26729 9004 26735 9380
rect 26769 9004 26775 9380
rect 26729 8992 26775 9004
rect 26847 9380 26893 9392
rect 26847 9004 26853 9380
rect 26887 9004 26893 9380
rect 26847 8992 26893 9004
rect 26965 9380 27011 9392
rect 26965 9004 26971 9380
rect 27005 9004 27011 9380
rect 26965 8992 27011 9004
rect 27083 9380 27129 9392
rect 27083 9004 27089 9380
rect 27123 9004 27129 9380
rect 27207 9192 27244 9479
rect 27083 8992 27129 9004
rect 27202 9180 27248 9192
rect 27202 9004 27208 9180
rect 27242 9004 27248 9180
rect 27202 8992 27248 9004
rect 27320 9180 27366 9192
rect 27320 9004 27326 9180
rect 27360 9004 27366 9180
rect 27320 8992 27366 9004
rect 27438 9180 27484 9192
rect 27438 9004 27444 9180
rect 27478 9004 27484 9180
rect 27438 8992 27484 9004
rect 27556 9180 27602 9813
rect 27903 9814 28054 9831
rect 27903 9754 27914 9814
rect 27978 9754 28054 9814
rect 27903 9742 28054 9754
rect 27900 9460 28056 9480
rect 27900 9399 27913 9460
rect 27980 9399 28056 9460
rect 27900 9386 28056 9399
rect 27556 9004 27562 9180
rect 27596 9004 27602 9180
rect 27556 8992 27602 9004
rect 24999 8806 25034 8992
rect 25908 8908 25942 8992
rect 27089 8908 27123 8992
rect 25908 8866 27123 8908
rect 27089 8846 27123 8866
rect 27089 8830 27446 8846
rect 24999 8789 26136 8806
rect 24999 8755 26086 8789
rect 26120 8755 26136 8789
rect 27089 8796 27396 8830
rect 27430 8796 27446 8830
rect 27089 8780 27446 8796
rect 24999 8739 26136 8755
rect 23277 8576 23342 8579
rect 23277 8573 23346 8576
rect 23277 8513 23283 8573
rect 23342 8513 23352 8573
rect 23277 8509 23346 8513
rect 23277 8507 23342 8509
rect 24418 8492 24599 8638
rect 24740 8694 24916 8702
rect 24740 8626 24857 8694
rect 24914 8626 24924 8694
rect 24740 8618 24916 8626
rect 24846 8578 24916 8586
rect 24846 8510 24857 8578
rect 24914 8510 24924 8578
rect 24846 8502 24916 8510
rect 22912 8410 23004 8418
rect 22912 8345 22924 8410
rect 22992 8345 23004 8410
rect 22912 8333 23004 8345
rect 24418 8230 24453 8492
rect 21855 8182 23227 8229
rect 23549 8183 24453 8230
rect 24782 8418 24846 8419
rect 24782 8410 24916 8418
rect 24782 8342 24857 8410
rect 24914 8342 24924 8410
rect 24782 8334 24916 8342
rect 22689 8059 22723 8182
rect 23161 8169 23227 8182
rect 23161 8135 23177 8169
rect 23211 8135 23227 8169
rect 23161 8119 23227 8135
rect 23550 8059 23584 8183
rect 22684 8047 22730 8059
rect 22684 7871 22690 8047
rect 22724 7871 22730 8047
rect 22684 7859 22730 7871
rect 22802 8047 22922 8059
rect 22802 7871 22808 8047
rect 22842 7871 22882 8047
rect 22802 7859 22882 7871
rect 22808 7492 22842 7859
rect 22876 7671 22882 7859
rect 22916 7671 22922 8047
rect 22876 7659 22922 7671
rect 22994 8047 23040 8059
rect 22994 7671 23000 8047
rect 23034 7671 23040 8047
rect 22994 7659 23040 7671
rect 23112 8047 23158 8059
rect 23112 7671 23118 8047
rect 23152 7671 23158 8047
rect 23112 7659 23158 7671
rect 23230 8047 23276 8059
rect 23230 7671 23236 8047
rect 23270 7671 23276 8047
rect 23230 7659 23276 7671
rect 23348 8047 23472 8059
rect 23348 7671 23354 8047
rect 23388 7871 23432 8047
rect 23466 7871 23472 8047
rect 23388 7859 23472 7871
rect 23544 8047 23590 8059
rect 23544 7871 23550 8047
rect 23584 7871 23590 8047
rect 23544 7859 23590 7871
rect 23388 7671 23394 7859
rect 23348 7659 23394 7671
rect 23118 7586 23152 7659
rect 23103 7570 23169 7586
rect 23103 7536 23119 7570
rect 23153 7536 23169 7570
rect 23103 7520 23169 7536
rect 23432 7492 23466 7859
rect 22808 7440 23466 7492
rect 23106 7418 23198 7440
rect 23106 7366 23118 7418
rect 23184 7366 23198 7418
rect 23106 7362 23198 7366
rect 12176 7272 15348 7320
rect 15380 7274 18494 7323
rect 18522 7322 20129 7323
rect 18522 7274 21617 7322
rect 21653 7278 24373 7326
rect 15300 7246 15348 7272
rect 9016 7196 15272 7244
rect 15300 7198 18418 7246
rect 15224 7170 15272 7196
rect 15224 7122 18347 7170
rect 18299 7091 18347 7122
rect 18375 7168 18418 7198
rect 18446 7244 18494 7274
rect 21569 7250 21617 7274
rect 18446 7196 21497 7244
rect 21569 7202 23630 7250
rect 21449 7172 21497 7196
rect 18375 7120 21421 7168
rect 21449 7124 22897 7172
rect 21373 7096 21421 7120
rect 18299 7043 21345 7091
rect 21373 7048 22153 7096
rect 5884 6960 20659 7008
rect 2740 6851 19915 6899
rect 19575 6739 19585 6753
rect 19545 6733 19585 6739
rect 19661 6739 19671 6753
rect 19661 6733 19703 6739
rect 3512 6672 3522 6694
rect 3484 6640 3522 6672
rect 3576 6672 3586 6694
rect 5580 6674 5590 6696
rect 3576 6640 3618 6672
rect 3484 6589 3618 6640
rect 5552 6642 5590 6674
rect 5644 6674 5654 6696
rect 5644 6642 5686 6674
rect 7649 6672 7659 6694
rect 5552 6591 5686 6642
rect 7621 6640 7659 6672
rect 7713 6672 7723 6694
rect 9717 6674 9727 6696
rect 7713 6640 7755 6672
rect 2813 6546 4286 6589
rect 2813 6243 2847 6546
rect 3179 6443 3213 6546
rect 3415 6443 3449 6546
rect 3651 6443 3685 6546
rect 3887 6443 3921 6546
rect 3173 6431 3219 6443
rect 2689 6231 2735 6243
rect 2689 6055 2695 6231
rect 2729 6055 2735 6231
rect 2689 6043 2735 6055
rect 2807 6231 2853 6243
rect 2807 6055 2813 6231
rect 2847 6055 2853 6231
rect 2807 6043 2853 6055
rect 2925 6231 2971 6243
rect 2925 6055 2931 6231
rect 2965 6055 2971 6231
rect 2925 6043 2971 6055
rect 3043 6231 3089 6243
rect 3173 6231 3179 6431
rect 3043 6055 3049 6231
rect 3083 6055 3179 6231
rect 3213 6055 3219 6431
rect 3043 6043 3089 6055
rect 3173 6043 3219 6055
rect 3291 6431 3337 6443
rect 3291 6055 3297 6431
rect 3331 6055 3337 6431
rect 3291 6043 3337 6055
rect 3409 6431 3455 6443
rect 3409 6055 3415 6431
rect 3449 6055 3455 6431
rect 3409 6043 3455 6055
rect 3527 6431 3573 6443
rect 3527 6055 3533 6431
rect 3567 6055 3573 6431
rect 3527 6043 3573 6055
rect 3645 6431 3691 6443
rect 3645 6055 3651 6431
rect 3685 6055 3691 6431
rect 3645 6043 3691 6055
rect 3763 6431 3809 6443
rect 3763 6055 3769 6431
rect 3803 6055 3809 6431
rect 3763 6043 3809 6055
rect 3881 6431 3927 6443
rect 3881 6055 3887 6431
rect 3921 6231 3927 6431
rect 4252 6243 4286 6546
rect 4881 6548 6354 6591
rect 7621 6589 7755 6640
rect 9689 6642 9727 6674
rect 9781 6674 9791 6696
rect 11786 6674 11796 6696
rect 9781 6642 9823 6674
rect 9689 6591 9823 6642
rect 11758 6642 11796 6674
rect 11850 6674 11860 6696
rect 13854 6676 13864 6698
rect 11850 6642 11892 6674
rect 11758 6591 11892 6642
rect 13826 6644 13864 6676
rect 13918 6676 13928 6698
rect 13918 6644 13960 6676
rect 15923 6674 15933 6696
rect 13826 6593 13960 6644
rect 15895 6642 15933 6674
rect 15987 6674 15997 6696
rect 17991 6676 18001 6698
rect 15987 6642 16029 6674
rect 4881 6245 4915 6548
rect 5247 6445 5281 6548
rect 5483 6445 5517 6548
rect 5719 6445 5753 6548
rect 5955 6445 5989 6548
rect 5241 6433 5287 6445
rect 4010 6231 4056 6243
rect 3921 6055 4016 6231
rect 4050 6055 4056 6231
rect 3881 6043 3927 6055
rect 4010 6043 4056 6055
rect 4128 6231 4174 6243
rect 4128 6055 4134 6231
rect 4168 6055 4174 6231
rect 4128 6043 4174 6055
rect 4246 6231 4292 6243
rect 4246 6055 4252 6231
rect 4286 6055 4292 6231
rect 4246 6043 4292 6055
rect 4364 6231 4410 6243
rect 4364 6055 4370 6231
rect 4404 6055 4410 6231
rect 4364 6043 4410 6055
rect 4757 6233 4803 6245
rect 4757 6057 4763 6233
rect 4797 6057 4803 6233
rect 4757 6045 4803 6057
rect 4875 6233 4921 6245
rect 4875 6057 4881 6233
rect 4915 6057 4921 6233
rect 4875 6045 4921 6057
rect 4993 6233 5039 6245
rect 4993 6057 4999 6233
rect 5033 6057 5039 6233
rect 4993 6045 5039 6057
rect 5111 6233 5157 6245
rect 5241 6233 5247 6433
rect 5111 6057 5117 6233
rect 5151 6057 5247 6233
rect 5281 6057 5287 6433
rect 5111 6045 5157 6057
rect 5241 6045 5287 6057
rect 5359 6433 5405 6445
rect 5359 6057 5365 6433
rect 5399 6057 5405 6433
rect 5359 6045 5405 6057
rect 5477 6433 5523 6445
rect 5477 6057 5483 6433
rect 5517 6057 5523 6433
rect 5477 6045 5523 6057
rect 5595 6433 5641 6445
rect 5595 6057 5601 6433
rect 5635 6057 5641 6433
rect 5595 6045 5641 6057
rect 5713 6433 5759 6445
rect 5713 6057 5719 6433
rect 5753 6057 5759 6433
rect 5713 6045 5759 6057
rect 5831 6433 5877 6445
rect 5831 6057 5837 6433
rect 5871 6057 5877 6433
rect 5831 6045 5877 6057
rect 5949 6433 5995 6445
rect 5949 6057 5955 6433
rect 5989 6233 5995 6433
rect 6320 6245 6354 6548
rect 6950 6546 8423 6589
rect 6078 6233 6124 6245
rect 5989 6057 6084 6233
rect 6118 6057 6124 6233
rect 5949 6045 5995 6057
rect 6078 6045 6124 6057
rect 6196 6233 6242 6245
rect 6196 6057 6202 6233
rect 6236 6057 6242 6233
rect 6196 6045 6242 6057
rect 6314 6233 6360 6245
rect 6314 6057 6320 6233
rect 6354 6057 6360 6233
rect 6314 6045 6360 6057
rect 6432 6233 6478 6245
rect 6950 6243 6984 6546
rect 7316 6443 7350 6546
rect 7552 6443 7586 6546
rect 7788 6443 7822 6546
rect 8024 6443 8058 6546
rect 7310 6431 7356 6443
rect 6432 6057 6438 6233
rect 6472 6057 6478 6233
rect 6432 6045 6478 6057
rect 6826 6231 6872 6243
rect 6826 6055 6832 6231
rect 6866 6055 6872 6231
rect 2695 6009 2729 6043
rect 3297 6009 3331 6043
rect 3533 6009 3567 6043
rect 2695 5974 2854 6009
rect 3297 5974 3567 6009
rect 4134 6009 4168 6043
rect 4370 6009 4404 6043
rect 4134 5974 4404 6009
rect 4763 6011 4797 6045
rect 5365 6011 5399 6045
rect 5601 6011 5635 6045
rect 4763 5976 4922 6011
rect 5365 5976 5635 6011
rect 6202 6011 6236 6045
rect 6438 6011 6472 6045
rect 6826 6043 6872 6055
rect 6944 6231 6990 6243
rect 6944 6055 6950 6231
rect 6984 6055 6990 6231
rect 6944 6043 6990 6055
rect 7062 6231 7108 6243
rect 7062 6055 7068 6231
rect 7102 6055 7108 6231
rect 7062 6043 7108 6055
rect 7180 6231 7226 6243
rect 7310 6231 7316 6431
rect 7180 6055 7186 6231
rect 7220 6055 7316 6231
rect 7350 6055 7356 6431
rect 7180 6043 7226 6055
rect 7310 6043 7356 6055
rect 7428 6431 7474 6443
rect 7428 6055 7434 6431
rect 7468 6055 7474 6431
rect 7428 6043 7474 6055
rect 7546 6431 7592 6443
rect 7546 6055 7552 6431
rect 7586 6055 7592 6431
rect 7546 6043 7592 6055
rect 7664 6431 7710 6443
rect 7664 6055 7670 6431
rect 7704 6055 7710 6431
rect 7664 6043 7710 6055
rect 7782 6431 7828 6443
rect 7782 6055 7788 6431
rect 7822 6055 7828 6431
rect 7782 6043 7828 6055
rect 7900 6431 7946 6443
rect 7900 6055 7906 6431
rect 7940 6055 7946 6431
rect 7900 6043 7946 6055
rect 8018 6431 8064 6443
rect 8018 6055 8024 6431
rect 8058 6231 8064 6431
rect 8389 6243 8423 6546
rect 9018 6548 10491 6591
rect 9018 6245 9052 6548
rect 9384 6445 9418 6548
rect 9620 6445 9654 6548
rect 9856 6445 9890 6548
rect 10092 6445 10126 6548
rect 9378 6433 9424 6445
rect 8147 6231 8193 6243
rect 8058 6055 8153 6231
rect 8187 6055 8193 6231
rect 8018 6043 8064 6055
rect 8147 6043 8193 6055
rect 8265 6231 8311 6243
rect 8265 6055 8271 6231
rect 8305 6055 8311 6231
rect 8265 6043 8311 6055
rect 8383 6231 8429 6243
rect 8383 6055 8389 6231
rect 8423 6055 8429 6231
rect 8383 6043 8429 6055
rect 8501 6231 8547 6243
rect 8501 6055 8507 6231
rect 8541 6055 8547 6231
rect 8501 6043 8547 6055
rect 8894 6233 8940 6245
rect 8894 6057 8900 6233
rect 8934 6057 8940 6233
rect 8894 6045 8940 6057
rect 9012 6233 9058 6245
rect 9012 6057 9018 6233
rect 9052 6057 9058 6233
rect 9012 6045 9058 6057
rect 9130 6233 9176 6245
rect 9130 6057 9136 6233
rect 9170 6057 9176 6233
rect 9130 6045 9176 6057
rect 9248 6233 9294 6245
rect 9378 6233 9384 6433
rect 9248 6057 9254 6233
rect 9288 6057 9384 6233
rect 9418 6057 9424 6433
rect 9248 6045 9294 6057
rect 9378 6045 9424 6057
rect 9496 6433 9542 6445
rect 9496 6057 9502 6433
rect 9536 6057 9542 6433
rect 9496 6045 9542 6057
rect 9614 6433 9660 6445
rect 9614 6057 9620 6433
rect 9654 6057 9660 6433
rect 9614 6045 9660 6057
rect 9732 6433 9778 6445
rect 9732 6057 9738 6433
rect 9772 6057 9778 6433
rect 9732 6045 9778 6057
rect 9850 6433 9896 6445
rect 9850 6057 9856 6433
rect 9890 6057 9896 6433
rect 9850 6045 9896 6057
rect 9968 6433 10014 6445
rect 9968 6057 9974 6433
rect 10008 6057 10014 6433
rect 9968 6045 10014 6057
rect 10086 6433 10132 6445
rect 10086 6057 10092 6433
rect 10126 6233 10132 6433
rect 10457 6245 10491 6548
rect 11087 6548 12560 6591
rect 11087 6245 11121 6548
rect 11453 6445 11487 6548
rect 11689 6445 11723 6548
rect 11925 6445 11959 6548
rect 12161 6445 12195 6548
rect 11447 6433 11493 6445
rect 10215 6233 10261 6245
rect 10126 6057 10221 6233
rect 10255 6057 10261 6233
rect 10086 6045 10132 6057
rect 10215 6045 10261 6057
rect 10333 6233 10379 6245
rect 10333 6057 10339 6233
rect 10373 6057 10379 6233
rect 10333 6045 10379 6057
rect 10451 6233 10497 6245
rect 10451 6057 10457 6233
rect 10491 6057 10497 6233
rect 10451 6045 10497 6057
rect 10569 6233 10615 6245
rect 10569 6057 10575 6233
rect 10609 6057 10615 6233
rect 10569 6045 10615 6057
rect 10963 6233 11009 6245
rect 10963 6057 10969 6233
rect 11003 6057 11009 6233
rect 10963 6045 11009 6057
rect 11081 6233 11127 6245
rect 11081 6057 11087 6233
rect 11121 6057 11127 6233
rect 11081 6045 11127 6057
rect 11199 6233 11245 6245
rect 11199 6057 11205 6233
rect 11239 6057 11245 6233
rect 11199 6045 11245 6057
rect 11317 6233 11363 6245
rect 11447 6233 11453 6433
rect 11317 6057 11323 6233
rect 11357 6057 11453 6233
rect 11487 6057 11493 6433
rect 11317 6045 11363 6057
rect 11447 6045 11493 6057
rect 11565 6433 11611 6445
rect 11565 6057 11571 6433
rect 11605 6057 11611 6433
rect 11565 6045 11611 6057
rect 11683 6433 11729 6445
rect 11683 6057 11689 6433
rect 11723 6057 11729 6433
rect 11683 6045 11729 6057
rect 11801 6433 11847 6445
rect 11801 6057 11807 6433
rect 11841 6057 11847 6433
rect 11801 6045 11847 6057
rect 11919 6433 11965 6445
rect 11919 6057 11925 6433
rect 11959 6057 11965 6433
rect 11919 6045 11965 6057
rect 12037 6433 12083 6445
rect 12037 6057 12043 6433
rect 12077 6057 12083 6433
rect 12037 6045 12083 6057
rect 12155 6433 12201 6445
rect 12155 6057 12161 6433
rect 12195 6233 12201 6433
rect 12526 6245 12560 6548
rect 13155 6550 14628 6593
rect 15895 6591 16029 6642
rect 17963 6644 18001 6676
rect 18055 6676 18065 6698
rect 19545 6697 19571 6733
rect 19667 6697 19703 6733
rect 19545 6679 19585 6697
rect 19661 6679 19703 6697
rect 18055 6644 18097 6676
rect 17963 6593 18097 6644
rect 19545 6639 19703 6679
rect 19421 6593 19703 6639
rect 13155 6247 13189 6550
rect 13521 6447 13555 6550
rect 13757 6447 13791 6550
rect 13993 6447 14027 6550
rect 14229 6447 14263 6550
rect 13515 6435 13561 6447
rect 12284 6233 12330 6245
rect 12195 6057 12290 6233
rect 12324 6057 12330 6233
rect 12155 6045 12201 6057
rect 12284 6045 12330 6057
rect 12402 6233 12448 6245
rect 12402 6057 12408 6233
rect 12442 6057 12448 6233
rect 12402 6045 12448 6057
rect 12520 6233 12566 6245
rect 12520 6057 12526 6233
rect 12560 6057 12566 6233
rect 12520 6045 12566 6057
rect 12638 6233 12684 6245
rect 12638 6057 12644 6233
rect 12678 6057 12684 6233
rect 12638 6045 12684 6057
rect 13031 6235 13077 6247
rect 13031 6059 13037 6235
rect 13071 6059 13077 6235
rect 13031 6047 13077 6059
rect 13149 6235 13195 6247
rect 13149 6059 13155 6235
rect 13189 6059 13195 6235
rect 13149 6047 13195 6059
rect 13267 6235 13313 6247
rect 13267 6059 13273 6235
rect 13307 6059 13313 6235
rect 13267 6047 13313 6059
rect 13385 6235 13431 6247
rect 13515 6235 13521 6435
rect 13385 6059 13391 6235
rect 13425 6059 13521 6235
rect 13555 6059 13561 6435
rect 13385 6047 13431 6059
rect 13515 6047 13561 6059
rect 13633 6435 13679 6447
rect 13633 6059 13639 6435
rect 13673 6059 13679 6435
rect 13633 6047 13679 6059
rect 13751 6435 13797 6447
rect 13751 6059 13757 6435
rect 13791 6059 13797 6435
rect 13751 6047 13797 6059
rect 13869 6435 13915 6447
rect 13869 6059 13875 6435
rect 13909 6059 13915 6435
rect 13869 6047 13915 6059
rect 13987 6435 14033 6447
rect 13987 6059 13993 6435
rect 14027 6059 14033 6435
rect 13987 6047 14033 6059
rect 14105 6435 14151 6447
rect 14105 6059 14111 6435
rect 14145 6059 14151 6435
rect 14105 6047 14151 6059
rect 14223 6435 14269 6447
rect 14223 6059 14229 6435
rect 14263 6235 14269 6435
rect 14594 6247 14628 6550
rect 15224 6548 16697 6591
rect 14352 6235 14398 6247
rect 14263 6059 14358 6235
rect 14392 6059 14398 6235
rect 14223 6047 14269 6059
rect 14352 6047 14398 6059
rect 14470 6235 14516 6247
rect 14470 6059 14476 6235
rect 14510 6059 14516 6235
rect 14470 6047 14516 6059
rect 14588 6235 14634 6247
rect 14588 6059 14594 6235
rect 14628 6059 14634 6235
rect 14588 6047 14634 6059
rect 14706 6235 14752 6247
rect 15224 6245 15258 6548
rect 15590 6445 15624 6548
rect 15826 6445 15860 6548
rect 16062 6445 16096 6548
rect 16298 6445 16332 6548
rect 15584 6433 15630 6445
rect 14706 6059 14712 6235
rect 14746 6059 14752 6235
rect 14706 6047 14752 6059
rect 15100 6233 15146 6245
rect 15100 6057 15106 6233
rect 15140 6057 15146 6233
rect 6202 5976 6472 6011
rect 6832 6009 6866 6043
rect 7434 6009 7468 6043
rect 7670 6009 7704 6043
rect 1995 5841 2005 5901
rect 2069 5841 2079 5901
rect 2424 5885 2714 5892
rect 2005 4269 2069 5841
rect 2418 5832 2428 5885
rect 2488 5832 2714 5885
rect 2424 5826 2714 5832
rect 2780 5826 2790 5892
rect 2689 5702 2699 5704
rect 2424 5693 2699 5702
rect 2418 5635 2428 5693
rect 2480 5635 2699 5693
rect 2424 5630 2699 5635
rect 2689 5627 2699 5630
rect 2770 5627 2780 5704
rect 2820 5190 2854 5974
rect 3533 5912 3567 5974
rect 3122 5874 3864 5912
rect 3122 5750 3156 5874
rect 3358 5750 3392 5874
rect 3594 5750 3628 5874
rect 3830 5750 3864 5874
rect 4090 5886 4168 5892
rect 4090 5832 4102 5886
rect 4156 5832 4168 5886
rect 4090 5826 4168 5832
rect 3116 5738 3162 5750
rect 3116 5362 3122 5738
rect 3156 5362 3162 5738
rect 3116 5350 3162 5362
rect 3234 5738 3280 5750
rect 3234 5362 3240 5738
rect 3274 5362 3280 5738
rect 3234 5350 3280 5362
rect 3352 5738 3398 5750
rect 3352 5362 3358 5738
rect 3392 5362 3398 5738
rect 3352 5350 3398 5362
rect 3470 5738 3516 5750
rect 3470 5362 3476 5738
rect 3510 5362 3516 5738
rect 3470 5350 3516 5362
rect 3588 5738 3634 5750
rect 3588 5362 3594 5738
rect 3628 5362 3634 5738
rect 3588 5350 3634 5362
rect 3706 5738 3752 5750
rect 3706 5362 3712 5738
rect 3746 5362 3752 5738
rect 3706 5350 3752 5362
rect 3824 5738 3870 5750
rect 3824 5362 3830 5738
rect 3864 5362 3870 5738
rect 3824 5350 3870 5362
rect 4236 5191 4270 5974
rect 4708 5828 4782 5894
rect 4848 5828 4858 5894
rect 4708 5698 4848 5704
rect 4708 5638 4770 5698
rect 4836 5638 4848 5698
rect 4708 5632 4848 5638
rect 4322 5334 4448 5340
rect 4322 5232 4334 5334
rect 4436 5232 4448 5334
rect 4322 5226 4448 5232
rect 3963 5190 4270 5191
rect 2820 5185 3136 5190
rect 3850 5185 4270 5190
rect 2820 5174 3203 5185
rect 2820 5147 3152 5174
rect 2820 5018 2854 5147
rect 3136 5140 3152 5147
rect 3186 5140 3203 5174
rect 3136 5134 3203 5140
rect 3783 5174 4270 5185
rect 3783 5140 3800 5174
rect 3834 5147 4270 5174
rect 3834 5140 3850 5147
rect 3963 5146 4270 5147
rect 3783 5134 3850 5140
rect 2961 5107 3017 5119
rect 2961 5073 2967 5107
rect 3001 5106 3017 5107
rect 4074 5106 4130 5118
rect 3001 5090 3468 5106
rect 3001 5073 3418 5090
rect 2961 5057 3418 5073
rect 3402 5056 3418 5057
rect 3452 5056 3468 5090
rect 3402 5049 3468 5056
rect 3520 5091 4090 5106
rect 3520 5057 3536 5091
rect 3570 5072 4090 5091
rect 4124 5072 4130 5106
rect 3570 5057 4130 5072
rect 3520 5047 3587 5057
rect 4074 5056 4130 5057
rect 4236 5018 4270 5146
rect 2814 5006 2860 5018
rect 2814 4830 2820 5006
rect 2854 4830 2860 5006
rect 2814 4818 2860 4830
rect 2932 5006 2978 5018
rect 2932 4830 2938 5006
rect 2972 4830 2978 5006
rect 2932 4818 2978 4830
rect 3234 5006 3280 5018
rect 2937 4524 2971 4818
rect 3234 4630 3240 5006
rect 3274 4630 3280 5006
rect 3234 4618 3280 4630
rect 3352 5006 3398 5018
rect 3352 4630 3358 5006
rect 3392 4630 3398 5006
rect 3352 4618 3398 4630
rect 3470 5006 3516 5018
rect 3470 4630 3476 5006
rect 3510 4630 3516 5006
rect 3470 4618 3516 4630
rect 3588 5006 3634 5018
rect 3588 4630 3594 5006
rect 3628 4630 3634 5006
rect 3588 4618 3634 4630
rect 3706 5006 3752 5018
rect 3706 4630 3712 5006
rect 3746 4630 3752 5006
rect 4112 5006 4158 5018
rect 4112 4830 4118 5006
rect 4152 4830 4158 5006
rect 4112 4818 4158 4830
rect 4230 5006 4276 5018
rect 4230 4830 4236 5006
rect 4270 4830 4276 5006
rect 4230 4818 4276 4830
rect 3706 4618 3752 4630
rect 3594 4524 3628 4618
rect 4118 4524 4151 4818
rect 2937 4492 4151 4524
rect 3430 4470 3562 4492
rect 3430 4412 3464 4470
rect 3526 4412 3562 4470
rect 3430 4407 3562 4412
rect 4708 4269 4772 5632
rect 4888 5192 4922 5976
rect 5601 5914 5635 5976
rect 5190 5876 5932 5914
rect 5190 5752 5224 5876
rect 5426 5752 5460 5876
rect 5662 5752 5696 5876
rect 5898 5752 5932 5876
rect 6158 5888 6236 5894
rect 6158 5834 6170 5888
rect 6224 5834 6236 5888
rect 6158 5828 6236 5834
rect 5184 5740 5230 5752
rect 5184 5364 5190 5740
rect 5224 5364 5230 5740
rect 5184 5352 5230 5364
rect 5302 5740 5348 5752
rect 5302 5364 5308 5740
rect 5342 5364 5348 5740
rect 5302 5352 5348 5364
rect 5420 5740 5466 5752
rect 5420 5364 5426 5740
rect 5460 5364 5466 5740
rect 5420 5352 5466 5364
rect 5538 5740 5584 5752
rect 5538 5364 5544 5740
rect 5578 5364 5584 5740
rect 5538 5352 5584 5364
rect 5656 5740 5702 5752
rect 5656 5364 5662 5740
rect 5696 5364 5702 5740
rect 5656 5352 5702 5364
rect 5774 5740 5820 5752
rect 5774 5364 5780 5740
rect 5814 5364 5820 5740
rect 5774 5352 5820 5364
rect 5892 5740 5938 5752
rect 5892 5364 5898 5740
rect 5932 5364 5938 5740
rect 5892 5352 5938 5364
rect 6304 5193 6338 5976
rect 6832 5974 6991 6009
rect 7434 5974 7704 6009
rect 8271 6009 8305 6043
rect 8507 6009 8541 6043
rect 8271 5974 8541 6009
rect 8900 6011 8934 6045
rect 9502 6011 9536 6045
rect 9738 6011 9772 6045
rect 8900 5976 9059 6011
rect 9502 5976 9772 6011
rect 10339 6011 10373 6045
rect 10575 6011 10609 6045
rect 10339 5976 10609 6011
rect 10969 6011 11003 6045
rect 11571 6011 11605 6045
rect 11807 6011 11841 6045
rect 10969 5976 11128 6011
rect 11571 5976 11841 6011
rect 12408 6011 12442 6045
rect 12644 6011 12678 6045
rect 12408 5976 12678 6011
rect 13037 6013 13071 6047
rect 13639 6013 13673 6047
rect 13875 6013 13909 6047
rect 13037 5978 13196 6013
rect 13639 5978 13909 6013
rect 14476 6013 14510 6047
rect 14712 6013 14746 6047
rect 15100 6045 15146 6057
rect 15218 6233 15264 6245
rect 15218 6057 15224 6233
rect 15258 6057 15264 6233
rect 15218 6045 15264 6057
rect 15336 6233 15382 6245
rect 15336 6057 15342 6233
rect 15376 6057 15382 6233
rect 15336 6045 15382 6057
rect 15454 6233 15500 6245
rect 15584 6233 15590 6433
rect 15454 6057 15460 6233
rect 15494 6057 15590 6233
rect 15624 6057 15630 6433
rect 15454 6045 15500 6057
rect 15584 6045 15630 6057
rect 15702 6433 15748 6445
rect 15702 6057 15708 6433
rect 15742 6057 15748 6433
rect 15702 6045 15748 6057
rect 15820 6433 15866 6445
rect 15820 6057 15826 6433
rect 15860 6057 15866 6433
rect 15820 6045 15866 6057
rect 15938 6433 15984 6445
rect 15938 6057 15944 6433
rect 15978 6057 15984 6433
rect 15938 6045 15984 6057
rect 16056 6433 16102 6445
rect 16056 6057 16062 6433
rect 16096 6057 16102 6433
rect 16056 6045 16102 6057
rect 16174 6433 16220 6445
rect 16174 6057 16180 6433
rect 16214 6057 16220 6433
rect 16174 6045 16220 6057
rect 16292 6433 16338 6445
rect 16292 6057 16298 6433
rect 16332 6233 16338 6433
rect 16663 6245 16697 6548
rect 17292 6550 18765 6593
rect 17292 6247 17326 6550
rect 17658 6447 17692 6550
rect 17894 6447 17928 6550
rect 18130 6447 18164 6550
rect 18366 6447 18400 6550
rect 17652 6435 17698 6447
rect 16421 6233 16467 6245
rect 16332 6057 16427 6233
rect 16461 6057 16467 6233
rect 16292 6045 16338 6057
rect 16421 6045 16467 6057
rect 16539 6233 16585 6245
rect 16539 6057 16545 6233
rect 16579 6057 16585 6233
rect 16539 6045 16585 6057
rect 16657 6233 16703 6245
rect 16657 6057 16663 6233
rect 16697 6057 16703 6233
rect 16657 6045 16703 6057
rect 16775 6233 16821 6245
rect 16775 6057 16781 6233
rect 16815 6057 16821 6233
rect 16775 6045 16821 6057
rect 17168 6235 17214 6247
rect 17168 6059 17174 6235
rect 17208 6059 17214 6235
rect 17168 6047 17214 6059
rect 17286 6235 17332 6247
rect 17286 6059 17292 6235
rect 17326 6059 17332 6235
rect 17286 6047 17332 6059
rect 17404 6235 17450 6247
rect 17404 6059 17410 6235
rect 17444 6059 17450 6235
rect 17404 6047 17450 6059
rect 17522 6235 17568 6247
rect 17652 6235 17658 6435
rect 17522 6059 17528 6235
rect 17562 6059 17658 6235
rect 17692 6059 17698 6435
rect 17522 6047 17568 6059
rect 17652 6047 17698 6059
rect 17770 6435 17816 6447
rect 17770 6059 17776 6435
rect 17810 6059 17816 6435
rect 17770 6047 17816 6059
rect 17888 6435 17934 6447
rect 17888 6059 17894 6435
rect 17928 6059 17934 6435
rect 17888 6047 17934 6059
rect 18006 6435 18052 6447
rect 18006 6059 18012 6435
rect 18046 6059 18052 6435
rect 18006 6047 18052 6059
rect 18124 6435 18170 6447
rect 18124 6059 18130 6435
rect 18164 6059 18170 6435
rect 18124 6047 18170 6059
rect 18242 6435 18288 6447
rect 18242 6059 18248 6435
rect 18282 6059 18288 6435
rect 18242 6047 18288 6059
rect 18360 6435 18406 6447
rect 18360 6059 18366 6435
rect 18400 6235 18406 6435
rect 18731 6247 18765 6550
rect 19421 6547 19467 6593
rect 19421 6371 19427 6547
rect 19461 6371 19467 6547
rect 19421 6359 19467 6371
rect 19539 6547 19585 6559
rect 19539 6371 19545 6547
rect 19579 6371 19585 6547
rect 19539 6359 19585 6371
rect 19657 6547 19703 6593
rect 19657 6371 19663 6547
rect 19697 6371 19703 6547
rect 19657 6359 19703 6371
rect 19775 6547 19821 6559
rect 19775 6371 19781 6547
rect 19815 6371 19821 6547
rect 19775 6369 19821 6371
rect 19775 6282 19823 6369
rect 19851 6282 19915 6851
rect 20313 6737 20323 6751
rect 20283 6731 20323 6737
rect 20399 6737 20409 6751
rect 20399 6731 20441 6737
rect 20283 6695 20309 6731
rect 20405 6695 20441 6731
rect 20283 6677 20323 6695
rect 20399 6677 20441 6695
rect 20283 6637 20441 6677
rect 20159 6591 20441 6637
rect 20159 6551 20205 6591
rect 20159 6375 20165 6551
rect 20199 6375 20205 6551
rect 20159 6363 20205 6375
rect 20277 6551 20323 6563
rect 20277 6375 20283 6551
rect 20317 6375 20323 6551
rect 20277 6363 20323 6375
rect 20395 6551 20441 6591
rect 20395 6375 20401 6551
rect 20435 6375 20441 6551
rect 20395 6363 20441 6375
rect 20513 6551 20559 6563
rect 20513 6375 20519 6551
rect 20553 6375 20559 6551
rect 20513 6367 20559 6375
rect 20513 6284 20561 6367
rect 20595 6284 20659 6960
rect 21297 6987 21345 7043
rect 21297 6959 21384 6987
rect 21051 6737 21061 6751
rect 21021 6731 21061 6737
rect 21137 6737 21147 6751
rect 21137 6731 21179 6737
rect 21021 6695 21047 6731
rect 21143 6695 21179 6731
rect 21021 6677 21061 6695
rect 21137 6677 21179 6695
rect 21021 6637 21179 6677
rect 20897 6591 21179 6637
rect 20897 6547 20943 6591
rect 20897 6371 20903 6547
rect 20937 6371 20943 6547
rect 20897 6359 20943 6371
rect 21015 6547 21061 6559
rect 21015 6371 21021 6547
rect 21055 6371 21061 6547
rect 21015 6359 21061 6371
rect 21133 6547 21179 6591
rect 21133 6371 21139 6547
rect 21173 6371 21179 6547
rect 21133 6359 21179 6371
rect 21251 6547 21297 6559
rect 21251 6371 21257 6547
rect 21291 6371 21297 6547
rect 21251 6367 21297 6371
rect 21251 6286 21299 6367
rect 21336 6286 21384 6959
rect 21793 6737 21803 6751
rect 21763 6731 21803 6737
rect 21879 6737 21889 6751
rect 21879 6731 21921 6737
rect 21763 6695 21789 6731
rect 21885 6695 21921 6731
rect 21763 6677 21803 6695
rect 21879 6677 21921 6695
rect 21763 6637 21921 6677
rect 21639 6591 21921 6637
rect 21639 6545 21685 6591
rect 21639 6369 21645 6545
rect 21679 6369 21685 6545
rect 21639 6357 21685 6369
rect 21757 6545 21803 6557
rect 21757 6369 21763 6545
rect 21797 6369 21803 6545
rect 21757 6357 21803 6369
rect 21875 6545 21921 6591
rect 21875 6369 21881 6545
rect 21915 6369 21921 6545
rect 21875 6357 21921 6369
rect 21993 6545 22039 6557
rect 21993 6369 21999 6545
rect 22033 6369 22039 6545
rect 21993 6367 22039 6369
rect 19572 6265 19649 6271
rect 18489 6235 18535 6247
rect 18400 6059 18495 6235
rect 18529 6059 18535 6235
rect 18360 6047 18406 6059
rect 18489 6047 18535 6059
rect 18607 6235 18653 6247
rect 18607 6059 18613 6235
rect 18647 6059 18653 6235
rect 18607 6047 18653 6059
rect 18725 6235 18771 6247
rect 18725 6059 18731 6235
rect 18765 6059 18771 6235
rect 18725 6047 18771 6059
rect 18843 6235 18889 6247
rect 18843 6059 18849 6235
rect 18883 6059 18889 6235
rect 19572 6231 19603 6265
rect 19637 6231 19649 6265
rect 19572 6225 19649 6231
rect 19771 6221 19915 6282
rect 20301 6263 20387 6269
rect 20301 6229 20341 6263
rect 20375 6229 20387 6263
rect 20301 6223 20387 6229
rect 19775 6177 19823 6221
rect 20509 6220 20659 6284
rect 21046 6263 21125 6269
rect 21046 6229 21079 6263
rect 21113 6229 21125 6263
rect 21046 6223 21125 6229
rect 21247 6224 21384 6286
rect 21993 6285 22041 6367
rect 22089 6285 22153 7048
rect 22533 6737 22543 6751
rect 22503 6731 22543 6737
rect 22619 6737 22629 6751
rect 22619 6731 22661 6737
rect 22503 6695 22529 6731
rect 22625 6695 22661 6731
rect 22503 6677 22543 6695
rect 22619 6677 22661 6695
rect 22503 6637 22661 6677
rect 22379 6591 22661 6637
rect 22379 6545 22425 6591
rect 22379 6369 22385 6545
rect 22419 6369 22425 6545
rect 22379 6357 22425 6369
rect 22497 6545 22543 6557
rect 22497 6369 22503 6545
rect 22537 6369 22543 6545
rect 22497 6357 22543 6369
rect 22615 6545 22661 6591
rect 22615 6369 22621 6545
rect 22655 6369 22661 6545
rect 22615 6357 22661 6369
rect 22733 6545 22779 6557
rect 22733 6369 22739 6545
rect 22773 6369 22779 6545
rect 22733 6367 22779 6369
rect 22733 6285 22781 6367
rect 22833 6285 22897 7124
rect 23271 6737 23281 6751
rect 23241 6731 23281 6737
rect 23357 6737 23367 6751
rect 23357 6731 23399 6737
rect 23241 6695 23267 6731
rect 23363 6695 23399 6731
rect 23241 6677 23281 6695
rect 23357 6677 23399 6695
rect 23241 6637 23399 6677
rect 23117 6591 23399 6637
rect 23117 6545 23163 6591
rect 23117 6369 23123 6545
rect 23157 6369 23163 6545
rect 23117 6357 23163 6369
rect 23235 6545 23281 6557
rect 23235 6369 23241 6545
rect 23275 6369 23281 6545
rect 23235 6357 23281 6369
rect 23353 6545 23399 6591
rect 23353 6369 23359 6545
rect 23393 6369 23399 6545
rect 23353 6357 23399 6369
rect 23471 6545 23517 6557
rect 23471 6369 23477 6545
rect 23511 6369 23517 6545
rect 23471 6367 23517 6369
rect 23471 6285 23519 6367
rect 23566 6285 23630 7202
rect 24009 6737 24019 6751
rect 23979 6731 24019 6737
rect 24095 6737 24105 6751
rect 24095 6731 24137 6737
rect 23979 6695 24005 6731
rect 24101 6695 24137 6731
rect 23979 6677 24019 6695
rect 24095 6677 24137 6695
rect 23979 6637 24137 6677
rect 23855 6591 24137 6637
rect 23855 6545 23901 6591
rect 23855 6369 23861 6545
rect 23895 6369 23901 6545
rect 23855 6357 23901 6369
rect 23973 6545 24019 6557
rect 23973 6369 23979 6545
rect 24013 6369 24019 6545
rect 23973 6357 24019 6369
rect 24091 6545 24137 6591
rect 24091 6369 24097 6545
rect 24131 6369 24137 6545
rect 24091 6357 24137 6369
rect 24209 6545 24255 6557
rect 24209 6369 24215 6545
rect 24249 6369 24255 6545
rect 24209 6367 24255 6369
rect 21787 6263 21867 6269
rect 21787 6229 21821 6263
rect 21855 6229 21867 6263
rect 18843 6047 18889 6059
rect 19539 6161 19585 6173
rect 14476 5978 14746 6013
rect 15106 6011 15140 6045
rect 15708 6011 15742 6045
rect 15944 6011 15978 6045
rect 6777 5826 6851 5892
rect 6917 5826 6927 5892
rect 6742 5696 6917 5702
rect 6742 5636 6839 5696
rect 6905 5636 6917 5696
rect 6742 5630 6917 5636
rect 6390 5336 6516 5342
rect 6390 5234 6402 5336
rect 6504 5234 6516 5336
rect 6390 5228 6516 5234
rect 6031 5192 6338 5193
rect 4888 5187 5204 5192
rect 5918 5187 6338 5192
rect 4888 5176 5271 5187
rect 4888 5149 5220 5176
rect 4888 5020 4922 5149
rect 5204 5142 5220 5149
rect 5254 5142 5271 5176
rect 5204 5136 5271 5142
rect 5851 5176 6338 5187
rect 5851 5142 5868 5176
rect 5902 5149 6338 5176
rect 5902 5142 5918 5149
rect 6031 5148 6338 5149
rect 5851 5136 5918 5142
rect 5029 5109 5085 5121
rect 5029 5075 5035 5109
rect 5069 5108 5085 5109
rect 6142 5108 6198 5120
rect 5069 5092 5536 5108
rect 5069 5075 5486 5092
rect 5029 5059 5486 5075
rect 5470 5058 5486 5059
rect 5520 5058 5536 5092
rect 5470 5051 5536 5058
rect 5588 5093 6158 5108
rect 5588 5059 5604 5093
rect 5638 5074 6158 5093
rect 6192 5074 6198 5108
rect 5638 5059 6198 5074
rect 5588 5049 5655 5059
rect 6142 5058 6198 5059
rect 6304 5020 6338 5148
rect 4882 5008 4928 5020
rect 4882 4832 4888 5008
rect 4922 4832 4928 5008
rect 4882 4820 4928 4832
rect 5000 5008 5046 5020
rect 5000 4832 5006 5008
rect 5040 4832 5046 5008
rect 5000 4820 5046 4832
rect 5302 5008 5348 5020
rect 5005 4526 5039 4820
rect 5302 4632 5308 5008
rect 5342 4632 5348 5008
rect 5302 4620 5348 4632
rect 5420 5008 5466 5020
rect 5420 4632 5426 5008
rect 5460 4632 5466 5008
rect 5420 4620 5466 4632
rect 5538 5008 5584 5020
rect 5538 4632 5544 5008
rect 5578 4632 5584 5008
rect 5538 4620 5584 4632
rect 5656 5008 5702 5020
rect 5656 4632 5662 5008
rect 5696 4632 5702 5008
rect 5656 4620 5702 4632
rect 5774 5008 5820 5020
rect 5774 4632 5780 5008
rect 5814 4632 5820 5008
rect 6180 5008 6226 5020
rect 6180 4832 6186 5008
rect 6220 4832 6226 5008
rect 6180 4820 6226 4832
rect 6298 5008 6344 5020
rect 6298 4832 6304 5008
rect 6338 4832 6344 5008
rect 6298 4820 6344 4832
rect 5774 4620 5820 4632
rect 5662 4526 5696 4620
rect 6186 4526 6219 4820
rect 5005 4494 6219 4526
rect 5498 4472 5630 4494
rect 5498 4414 5532 4472
rect 5594 4414 5630 4472
rect 5498 4409 5630 4414
rect 2005 4205 4773 4269
rect 2005 4204 2310 4205
rect 4708 4061 4772 4205
rect 4703 4055 4778 4061
rect 4703 4004 4715 4055
rect 4766 4004 4778 4055
rect 4703 3998 4778 4004
rect 6742 3958 6806 5630
rect 6957 5190 6991 5974
rect 7670 5912 7704 5974
rect 7259 5874 8001 5912
rect 7259 5750 7293 5874
rect 7495 5750 7529 5874
rect 7731 5750 7765 5874
rect 7967 5750 8001 5874
rect 8227 5886 8305 5892
rect 8227 5832 8239 5886
rect 8293 5832 8305 5886
rect 8227 5826 8305 5832
rect 7253 5738 7299 5750
rect 7253 5362 7259 5738
rect 7293 5362 7299 5738
rect 7253 5350 7299 5362
rect 7371 5738 7417 5750
rect 7371 5362 7377 5738
rect 7411 5362 7417 5738
rect 7371 5350 7417 5362
rect 7489 5738 7535 5750
rect 7489 5362 7495 5738
rect 7529 5362 7535 5738
rect 7489 5350 7535 5362
rect 7607 5738 7653 5750
rect 7607 5362 7613 5738
rect 7647 5362 7653 5738
rect 7607 5350 7653 5362
rect 7725 5738 7771 5750
rect 7725 5362 7731 5738
rect 7765 5362 7771 5738
rect 7725 5350 7771 5362
rect 7843 5738 7889 5750
rect 7843 5362 7849 5738
rect 7883 5362 7889 5738
rect 7843 5350 7889 5362
rect 7961 5738 8007 5750
rect 7961 5362 7967 5738
rect 8001 5362 8007 5738
rect 7961 5350 8007 5362
rect 8373 5191 8407 5974
rect 8845 5828 8919 5894
rect 8985 5828 8995 5894
rect 8788 5698 8985 5704
rect 8788 5638 8907 5698
rect 8973 5638 8985 5698
rect 8788 5632 8985 5638
rect 8459 5334 8585 5340
rect 8459 5232 8471 5334
rect 8573 5232 8585 5334
rect 8459 5226 8585 5232
rect 8100 5190 8407 5191
rect 6957 5185 7273 5190
rect 7987 5185 8407 5190
rect 6957 5174 7340 5185
rect 6957 5147 7289 5174
rect 6957 5018 6991 5147
rect 7273 5140 7289 5147
rect 7323 5140 7340 5174
rect 7273 5134 7340 5140
rect 7920 5174 8407 5185
rect 7920 5140 7937 5174
rect 7971 5147 8407 5174
rect 7971 5140 7987 5147
rect 8100 5146 8407 5147
rect 7920 5134 7987 5140
rect 7098 5107 7154 5119
rect 7098 5073 7104 5107
rect 7138 5106 7154 5107
rect 8211 5106 8267 5118
rect 7138 5090 7605 5106
rect 7138 5073 7555 5090
rect 7098 5057 7555 5073
rect 7539 5056 7555 5057
rect 7589 5056 7605 5090
rect 7539 5049 7605 5056
rect 7657 5091 8227 5106
rect 7657 5057 7673 5091
rect 7707 5072 8227 5091
rect 8261 5072 8267 5106
rect 7707 5057 8267 5072
rect 7657 5047 7724 5057
rect 8211 5056 8267 5057
rect 8373 5018 8407 5146
rect 6951 5006 6997 5018
rect 6951 4830 6957 5006
rect 6991 4830 6997 5006
rect 6951 4818 6997 4830
rect 7069 5006 7115 5018
rect 7069 4830 7075 5006
rect 7109 4830 7115 5006
rect 7069 4818 7115 4830
rect 7371 5006 7417 5018
rect 7074 4524 7108 4818
rect 7371 4630 7377 5006
rect 7411 4630 7417 5006
rect 7371 4618 7417 4630
rect 7489 5006 7535 5018
rect 7489 4630 7495 5006
rect 7529 4630 7535 5006
rect 7489 4618 7535 4630
rect 7607 5006 7653 5018
rect 7607 4630 7613 5006
rect 7647 4630 7653 5006
rect 7607 4618 7653 4630
rect 7725 5006 7771 5018
rect 7725 4630 7731 5006
rect 7765 4630 7771 5006
rect 7725 4618 7771 4630
rect 7843 5006 7889 5018
rect 7843 4630 7849 5006
rect 7883 4630 7889 5006
rect 8249 5006 8295 5018
rect 8249 4830 8255 5006
rect 8289 4830 8295 5006
rect 8249 4818 8295 4830
rect 8367 5006 8413 5018
rect 8367 4830 8373 5006
rect 8407 4830 8413 5006
rect 8367 4818 8413 4830
rect 7843 4618 7889 4630
rect 7731 4524 7765 4618
rect 8255 4524 8288 4818
rect 7074 4492 8288 4524
rect 7567 4470 7699 4492
rect 7567 4412 7601 4470
rect 7663 4412 7699 4470
rect 7567 4407 7699 4412
rect 1775 3950 6806 3958
rect 1775 3896 6750 3950
rect 6797 3896 6806 3950
rect 1775 3877 6806 3896
rect 8788 3849 8852 5632
rect 9025 5192 9059 5976
rect 9738 5914 9772 5976
rect 9327 5876 10069 5914
rect 9327 5752 9361 5876
rect 9563 5752 9597 5876
rect 9799 5752 9833 5876
rect 10035 5752 10069 5876
rect 10295 5888 10373 5894
rect 10295 5834 10307 5888
rect 10361 5834 10373 5888
rect 10295 5828 10373 5834
rect 9321 5740 9367 5752
rect 9321 5364 9327 5740
rect 9361 5364 9367 5740
rect 9321 5352 9367 5364
rect 9439 5740 9485 5752
rect 9439 5364 9445 5740
rect 9479 5364 9485 5740
rect 9439 5352 9485 5364
rect 9557 5740 9603 5752
rect 9557 5364 9563 5740
rect 9597 5364 9603 5740
rect 9557 5352 9603 5364
rect 9675 5740 9721 5752
rect 9675 5364 9681 5740
rect 9715 5364 9721 5740
rect 9675 5352 9721 5364
rect 9793 5740 9839 5752
rect 9793 5364 9799 5740
rect 9833 5364 9839 5740
rect 9793 5352 9839 5364
rect 9911 5740 9957 5752
rect 9911 5364 9917 5740
rect 9951 5364 9957 5740
rect 9911 5352 9957 5364
rect 10029 5740 10075 5752
rect 10029 5364 10035 5740
rect 10069 5364 10075 5740
rect 10029 5352 10075 5364
rect 10441 5193 10475 5976
rect 10914 5828 10988 5894
rect 11054 5828 11064 5894
rect 10878 5698 11054 5704
rect 10878 5638 10976 5698
rect 11042 5638 11054 5698
rect 10878 5632 11054 5638
rect 10527 5336 10653 5342
rect 10527 5234 10539 5336
rect 10641 5234 10653 5336
rect 10527 5228 10653 5234
rect 10168 5192 10475 5193
rect 9025 5187 9341 5192
rect 10055 5187 10475 5192
rect 9025 5176 9408 5187
rect 9025 5149 9357 5176
rect 9025 5020 9059 5149
rect 9341 5142 9357 5149
rect 9391 5142 9408 5176
rect 9341 5136 9408 5142
rect 9988 5176 10475 5187
rect 9988 5142 10005 5176
rect 10039 5149 10475 5176
rect 10039 5142 10055 5149
rect 10168 5148 10475 5149
rect 9988 5136 10055 5142
rect 9166 5109 9222 5121
rect 9166 5075 9172 5109
rect 9206 5108 9222 5109
rect 10279 5108 10335 5120
rect 9206 5092 9673 5108
rect 9206 5075 9623 5092
rect 9166 5059 9623 5075
rect 9607 5058 9623 5059
rect 9657 5058 9673 5092
rect 9607 5051 9673 5058
rect 9725 5093 10295 5108
rect 9725 5059 9741 5093
rect 9775 5074 10295 5093
rect 10329 5074 10335 5108
rect 9775 5059 10335 5074
rect 9725 5049 9792 5059
rect 10279 5058 10335 5059
rect 10441 5020 10475 5148
rect 9019 5008 9065 5020
rect 9019 4832 9025 5008
rect 9059 4832 9065 5008
rect 9019 4820 9065 4832
rect 9137 5008 9183 5020
rect 9137 4832 9143 5008
rect 9177 4832 9183 5008
rect 9137 4820 9183 4832
rect 9439 5008 9485 5020
rect 9142 4526 9176 4820
rect 9439 4632 9445 5008
rect 9479 4632 9485 5008
rect 9439 4620 9485 4632
rect 9557 5008 9603 5020
rect 9557 4632 9563 5008
rect 9597 4632 9603 5008
rect 9557 4620 9603 4632
rect 9675 5008 9721 5020
rect 9675 4632 9681 5008
rect 9715 4632 9721 5008
rect 9675 4620 9721 4632
rect 9793 5008 9839 5020
rect 9793 4632 9799 5008
rect 9833 4632 9839 5008
rect 9793 4620 9839 4632
rect 9911 5008 9957 5020
rect 9911 4632 9917 5008
rect 9951 4632 9957 5008
rect 10317 5008 10363 5020
rect 10317 4832 10323 5008
rect 10357 4832 10363 5008
rect 10317 4820 10363 4832
rect 10435 5008 10481 5020
rect 10435 4832 10441 5008
rect 10475 4832 10481 5008
rect 10435 4820 10481 4832
rect 9911 4620 9957 4632
rect 9799 4526 9833 4620
rect 10323 4526 10356 4820
rect 9142 4494 10356 4526
rect 9635 4472 9767 4494
rect 9635 4414 9669 4472
rect 9731 4414 9767 4472
rect 9635 4409 9767 4414
rect 1578 3847 8852 3849
rect 1578 3793 8797 3847
rect 8844 3793 8852 3847
rect 1578 3757 8852 3793
rect 10878 3749 10942 5632
rect 11094 5192 11128 5976
rect 11807 5914 11841 5976
rect 11396 5876 12138 5914
rect 11396 5752 11430 5876
rect 11632 5752 11666 5876
rect 11868 5752 11902 5876
rect 12104 5752 12138 5876
rect 12364 5888 12442 5894
rect 12364 5834 12376 5888
rect 12430 5834 12442 5888
rect 12364 5828 12442 5834
rect 11390 5740 11436 5752
rect 11390 5364 11396 5740
rect 11430 5364 11436 5740
rect 11390 5352 11436 5364
rect 11508 5740 11554 5752
rect 11508 5364 11514 5740
rect 11548 5364 11554 5740
rect 11508 5352 11554 5364
rect 11626 5740 11672 5752
rect 11626 5364 11632 5740
rect 11666 5364 11672 5740
rect 11626 5352 11672 5364
rect 11744 5740 11790 5752
rect 11744 5364 11750 5740
rect 11784 5364 11790 5740
rect 11744 5352 11790 5364
rect 11862 5740 11908 5752
rect 11862 5364 11868 5740
rect 11902 5364 11908 5740
rect 11862 5352 11908 5364
rect 11980 5740 12026 5752
rect 11980 5364 11986 5740
rect 12020 5364 12026 5740
rect 11980 5352 12026 5364
rect 12098 5740 12144 5752
rect 12098 5364 12104 5740
rect 12138 5364 12144 5740
rect 12098 5352 12144 5364
rect 12510 5193 12544 5976
rect 12982 5830 13056 5896
rect 13122 5830 13132 5896
rect 12952 5700 13122 5706
rect 12952 5640 13044 5700
rect 13110 5640 13122 5700
rect 12952 5634 13122 5640
rect 12596 5336 12722 5342
rect 12596 5234 12608 5336
rect 12710 5234 12722 5336
rect 12596 5228 12722 5234
rect 12237 5192 12544 5193
rect 11094 5187 11410 5192
rect 12124 5187 12544 5192
rect 11094 5176 11477 5187
rect 11094 5149 11426 5176
rect 11094 5020 11128 5149
rect 11410 5142 11426 5149
rect 11460 5142 11477 5176
rect 11410 5136 11477 5142
rect 12057 5176 12544 5187
rect 12057 5142 12074 5176
rect 12108 5149 12544 5176
rect 12108 5142 12124 5149
rect 12237 5148 12544 5149
rect 12057 5136 12124 5142
rect 11235 5109 11291 5121
rect 11235 5075 11241 5109
rect 11275 5108 11291 5109
rect 12348 5108 12404 5120
rect 11275 5092 11742 5108
rect 11275 5075 11692 5092
rect 11235 5059 11692 5075
rect 11676 5058 11692 5059
rect 11726 5058 11742 5092
rect 11676 5051 11742 5058
rect 11794 5093 12364 5108
rect 11794 5059 11810 5093
rect 11844 5074 12364 5093
rect 12398 5074 12404 5108
rect 11844 5059 12404 5074
rect 11794 5049 11861 5059
rect 12348 5058 12404 5059
rect 12510 5020 12544 5148
rect 11088 5008 11134 5020
rect 11088 4832 11094 5008
rect 11128 4832 11134 5008
rect 11088 4820 11134 4832
rect 11206 5008 11252 5020
rect 11206 4832 11212 5008
rect 11246 4832 11252 5008
rect 11206 4820 11252 4832
rect 11508 5008 11554 5020
rect 11211 4526 11245 4820
rect 11508 4632 11514 5008
rect 11548 4632 11554 5008
rect 11508 4620 11554 4632
rect 11626 5008 11672 5020
rect 11626 4632 11632 5008
rect 11666 4632 11672 5008
rect 11626 4620 11672 4632
rect 11744 5008 11790 5020
rect 11744 4632 11750 5008
rect 11784 4632 11790 5008
rect 11744 4620 11790 4632
rect 11862 5008 11908 5020
rect 11862 4632 11868 5008
rect 11902 4632 11908 5008
rect 11862 4620 11908 4632
rect 11980 5008 12026 5020
rect 11980 4632 11986 5008
rect 12020 4632 12026 5008
rect 12386 5008 12432 5020
rect 12386 4832 12392 5008
rect 12426 4832 12432 5008
rect 12386 4820 12432 4832
rect 12504 5008 12550 5020
rect 12504 4832 12510 5008
rect 12544 4832 12550 5008
rect 12504 4820 12550 4832
rect 11980 4620 12026 4632
rect 11868 4526 11902 4620
rect 12392 4526 12425 4820
rect 11211 4494 12425 4526
rect 11704 4472 11836 4494
rect 11704 4414 11738 4472
rect 11800 4414 11836 4472
rect 11704 4409 11836 4414
rect 10878 3737 10943 3749
rect 1375 3729 1538 3730
rect 10878 3729 10887 3737
rect 1375 3686 10887 3729
rect 10937 3729 10943 3737
rect 10937 3686 10971 3729
rect 1375 3649 10971 3686
rect 1375 3648 1538 3649
rect 12952 3642 13016 5634
rect 13162 5194 13196 5978
rect 13875 5916 13909 5978
rect 13464 5878 14206 5916
rect 13464 5754 13498 5878
rect 13700 5754 13734 5878
rect 13936 5754 13970 5878
rect 14172 5754 14206 5878
rect 14432 5890 14510 5896
rect 14432 5836 14444 5890
rect 14498 5836 14510 5890
rect 14432 5830 14510 5836
rect 13458 5742 13504 5754
rect 13458 5366 13464 5742
rect 13498 5366 13504 5742
rect 13458 5354 13504 5366
rect 13576 5742 13622 5754
rect 13576 5366 13582 5742
rect 13616 5366 13622 5742
rect 13576 5354 13622 5366
rect 13694 5742 13740 5754
rect 13694 5366 13700 5742
rect 13734 5366 13740 5742
rect 13694 5354 13740 5366
rect 13812 5742 13858 5754
rect 13812 5366 13818 5742
rect 13852 5366 13858 5742
rect 13812 5354 13858 5366
rect 13930 5742 13976 5754
rect 13930 5366 13936 5742
rect 13970 5366 13976 5742
rect 13930 5354 13976 5366
rect 14048 5742 14094 5754
rect 14048 5366 14054 5742
rect 14088 5366 14094 5742
rect 14048 5354 14094 5366
rect 14166 5742 14212 5754
rect 14166 5366 14172 5742
rect 14206 5366 14212 5742
rect 14166 5354 14212 5366
rect 14578 5195 14612 5978
rect 15106 5976 15265 6011
rect 15708 5976 15978 6011
rect 16545 6011 16579 6045
rect 16781 6011 16815 6045
rect 16545 5976 16815 6011
rect 17174 6013 17208 6047
rect 17776 6013 17810 6047
rect 18012 6013 18046 6047
rect 17174 5978 17333 6013
rect 17776 5978 18046 6013
rect 18613 6013 18647 6047
rect 18849 6013 18883 6047
rect 18613 5978 18883 6013
rect 19539 5985 19545 6161
rect 19579 5985 19585 6161
rect 15051 5828 15125 5894
rect 15191 5828 15201 5894
rect 15051 5698 15191 5704
rect 15051 5638 15113 5698
rect 15179 5638 15191 5698
rect 15051 5632 15191 5638
rect 14664 5338 14790 5344
rect 14664 5236 14676 5338
rect 14778 5236 14790 5338
rect 14664 5230 14790 5236
rect 14305 5194 14612 5195
rect 13162 5189 13478 5194
rect 14192 5189 14612 5194
rect 13162 5178 13545 5189
rect 13162 5151 13494 5178
rect 13162 5022 13196 5151
rect 13478 5144 13494 5151
rect 13528 5144 13545 5178
rect 13478 5138 13545 5144
rect 14125 5178 14612 5189
rect 14125 5144 14142 5178
rect 14176 5151 14612 5178
rect 14176 5144 14192 5151
rect 14305 5150 14612 5151
rect 14125 5138 14192 5144
rect 13303 5111 13359 5123
rect 13303 5077 13309 5111
rect 13343 5110 13359 5111
rect 14416 5110 14472 5122
rect 13343 5094 13810 5110
rect 13343 5077 13760 5094
rect 13303 5061 13760 5077
rect 13744 5060 13760 5061
rect 13794 5060 13810 5094
rect 13744 5053 13810 5060
rect 13862 5095 14432 5110
rect 13862 5061 13878 5095
rect 13912 5076 14432 5095
rect 14466 5076 14472 5110
rect 13912 5061 14472 5076
rect 13862 5051 13929 5061
rect 14416 5060 14472 5061
rect 14578 5022 14612 5150
rect 13156 5010 13202 5022
rect 13156 4834 13162 5010
rect 13196 4834 13202 5010
rect 13156 4822 13202 4834
rect 13274 5010 13320 5022
rect 13274 4834 13280 5010
rect 13314 4834 13320 5010
rect 13274 4822 13320 4834
rect 13576 5010 13622 5022
rect 13279 4528 13313 4822
rect 13576 4634 13582 5010
rect 13616 4634 13622 5010
rect 13576 4622 13622 4634
rect 13694 5010 13740 5022
rect 13694 4634 13700 5010
rect 13734 4634 13740 5010
rect 13694 4622 13740 4634
rect 13812 5010 13858 5022
rect 13812 4634 13818 5010
rect 13852 4634 13858 5010
rect 13812 4622 13858 4634
rect 13930 5010 13976 5022
rect 13930 4634 13936 5010
rect 13970 4634 13976 5010
rect 13930 4622 13976 4634
rect 14048 5010 14094 5022
rect 14048 4634 14054 5010
rect 14088 4634 14094 5010
rect 14454 5010 14500 5022
rect 14454 4834 14460 5010
rect 14494 4834 14500 5010
rect 14454 4822 14500 4834
rect 14572 5010 14618 5022
rect 14572 4834 14578 5010
rect 14612 4834 14618 5010
rect 14572 4822 14618 4834
rect 14048 4622 14094 4634
rect 13936 4528 13970 4622
rect 14460 4528 14493 4822
rect 13279 4496 14493 4528
rect 13772 4474 13904 4496
rect 13772 4416 13806 4474
rect 13868 4416 13904 4474
rect 13772 4411 13904 4416
rect 12952 3602 12958 3642
rect 1203 3589 12958 3602
rect 13009 3602 13016 3642
rect 13009 3589 13017 3602
rect 1203 3534 13017 3589
rect 1203 3533 1267 3534
rect 15051 3503 15115 5632
rect 15231 5192 15265 5976
rect 15944 5914 15978 5976
rect 15533 5876 16275 5914
rect 15533 5752 15567 5876
rect 15769 5752 15803 5876
rect 16005 5752 16039 5876
rect 16241 5752 16275 5876
rect 16501 5888 16579 5894
rect 16501 5834 16513 5888
rect 16567 5834 16579 5888
rect 16501 5828 16579 5834
rect 15527 5740 15573 5752
rect 15527 5364 15533 5740
rect 15567 5364 15573 5740
rect 15527 5352 15573 5364
rect 15645 5740 15691 5752
rect 15645 5364 15651 5740
rect 15685 5364 15691 5740
rect 15645 5352 15691 5364
rect 15763 5740 15809 5752
rect 15763 5364 15769 5740
rect 15803 5364 15809 5740
rect 15763 5352 15809 5364
rect 15881 5740 15927 5752
rect 15881 5364 15887 5740
rect 15921 5364 15927 5740
rect 15881 5352 15927 5364
rect 15999 5740 16045 5752
rect 15999 5364 16005 5740
rect 16039 5364 16045 5740
rect 15999 5352 16045 5364
rect 16117 5740 16163 5752
rect 16117 5364 16123 5740
rect 16157 5364 16163 5740
rect 16117 5352 16163 5364
rect 16235 5740 16281 5752
rect 16235 5364 16241 5740
rect 16275 5364 16281 5740
rect 16235 5352 16281 5364
rect 16647 5193 16681 5976
rect 17119 5830 17193 5896
rect 17259 5830 17269 5896
rect 17122 5706 17186 5707
rect 17122 5700 17259 5706
rect 17122 5640 17181 5700
rect 17247 5640 17259 5700
rect 17122 5634 17259 5640
rect 16733 5336 16859 5342
rect 16733 5234 16745 5336
rect 16847 5234 16859 5336
rect 16733 5228 16859 5234
rect 16374 5192 16681 5193
rect 15231 5187 15547 5192
rect 16261 5187 16681 5192
rect 15231 5176 15614 5187
rect 15231 5149 15563 5176
rect 15231 5020 15265 5149
rect 15547 5142 15563 5149
rect 15597 5142 15614 5176
rect 15547 5136 15614 5142
rect 16194 5176 16681 5187
rect 16194 5142 16211 5176
rect 16245 5149 16681 5176
rect 16245 5142 16261 5149
rect 16374 5148 16681 5149
rect 16194 5136 16261 5142
rect 15372 5109 15428 5121
rect 15372 5075 15378 5109
rect 15412 5108 15428 5109
rect 16485 5108 16541 5120
rect 15412 5092 15879 5108
rect 15412 5075 15829 5092
rect 15372 5059 15829 5075
rect 15813 5058 15829 5059
rect 15863 5058 15879 5092
rect 15813 5051 15879 5058
rect 15931 5093 16501 5108
rect 15931 5059 15947 5093
rect 15981 5074 16501 5093
rect 16535 5074 16541 5108
rect 15981 5059 16541 5074
rect 15931 5049 15998 5059
rect 16485 5058 16541 5059
rect 16647 5020 16681 5148
rect 15225 5008 15271 5020
rect 15225 4832 15231 5008
rect 15265 4832 15271 5008
rect 15225 4820 15271 4832
rect 15343 5008 15389 5020
rect 15343 4832 15349 5008
rect 15383 4832 15389 5008
rect 15343 4820 15389 4832
rect 15645 5008 15691 5020
rect 15348 4526 15382 4820
rect 15645 4632 15651 5008
rect 15685 4632 15691 5008
rect 15645 4620 15691 4632
rect 15763 5008 15809 5020
rect 15763 4632 15769 5008
rect 15803 4632 15809 5008
rect 15763 4620 15809 4632
rect 15881 5008 15927 5020
rect 15881 4632 15887 5008
rect 15921 4632 15927 5008
rect 15881 4620 15927 4632
rect 15999 5008 16045 5020
rect 15999 4632 16005 5008
rect 16039 4632 16045 5008
rect 15999 4620 16045 4632
rect 16117 5008 16163 5020
rect 16117 4632 16123 5008
rect 16157 4632 16163 5008
rect 16523 5008 16569 5020
rect 16523 4832 16529 5008
rect 16563 4832 16569 5008
rect 16523 4820 16569 4832
rect 16641 5008 16687 5020
rect 16641 4832 16647 5008
rect 16681 4832 16687 5008
rect 16641 4820 16687 4832
rect 16117 4620 16163 4632
rect 16005 4526 16039 4620
rect 16529 4526 16562 4820
rect 15348 4494 16562 4526
rect 15841 4472 15973 4494
rect 15841 4414 15875 4472
rect 15937 4414 15973 4472
rect 15841 4409 15973 4414
rect 974 3498 15116 3503
rect 974 3447 15061 3498
rect 15105 3447 15116 3498
rect 974 3436 15116 3447
rect 974 3435 1054 3436
rect 15051 3435 15115 3436
rect 17122 3415 17186 5634
rect 17299 5194 17333 5978
rect 18012 5916 18046 5978
rect 17601 5878 18343 5916
rect 17601 5754 17635 5878
rect 17837 5754 17871 5878
rect 18073 5754 18107 5878
rect 18309 5754 18343 5878
rect 18569 5890 18647 5896
rect 18569 5836 18581 5890
rect 18635 5836 18647 5890
rect 18569 5830 18647 5836
rect 17595 5742 17641 5754
rect 17595 5366 17601 5742
rect 17635 5366 17641 5742
rect 17595 5354 17641 5366
rect 17713 5742 17759 5754
rect 17713 5366 17719 5742
rect 17753 5366 17759 5742
rect 17713 5354 17759 5366
rect 17831 5742 17877 5754
rect 17831 5366 17837 5742
rect 17871 5366 17877 5742
rect 17831 5354 17877 5366
rect 17949 5742 17995 5754
rect 17949 5366 17955 5742
rect 17989 5366 17995 5742
rect 17949 5354 17995 5366
rect 18067 5742 18113 5754
rect 18067 5366 18073 5742
rect 18107 5366 18113 5742
rect 18067 5354 18113 5366
rect 18185 5742 18231 5754
rect 18185 5366 18191 5742
rect 18225 5366 18231 5742
rect 18185 5354 18231 5366
rect 18303 5742 18349 5754
rect 18303 5366 18309 5742
rect 18343 5366 18349 5742
rect 18303 5354 18349 5366
rect 18715 5195 18749 5978
rect 19539 5871 19585 5985
rect 19657 6161 19823 6177
rect 20513 6175 20561 6220
rect 21251 6175 21299 6224
rect 21787 6223 21867 6229
rect 21989 6221 22153 6285
rect 22527 6263 22607 6269
rect 22527 6229 22561 6263
rect 22595 6229 22607 6263
rect 22527 6223 22607 6229
rect 22729 6221 22897 6285
rect 23263 6263 23345 6269
rect 23263 6229 23299 6263
rect 23333 6229 23345 6263
rect 23263 6223 23345 6229
rect 23467 6221 23630 6285
rect 24209 6282 24257 6367
rect 24309 6282 24373 7278
rect 24782 6954 24846 8334
rect 24999 8229 25034 8739
rect 25089 8693 25181 8706
rect 25089 8630 25101 8693
rect 25172 8630 25181 8693
rect 25089 8621 25181 8630
rect 26174 8693 26266 8703
rect 26174 8631 26186 8693
rect 26256 8631 26266 8693
rect 26174 8618 26266 8631
rect 27562 8638 27597 8992
rect 26421 8576 26486 8579
rect 26421 8573 26490 8576
rect 26421 8513 26427 8573
rect 26486 8513 26496 8573
rect 26421 8509 26490 8513
rect 26421 8507 26486 8509
rect 27562 8492 27598 8638
rect 26056 8410 26148 8418
rect 26056 8345 26068 8410
rect 26136 8345 26148 8410
rect 26056 8333 26148 8345
rect 27562 8230 27597 8492
rect 24999 8182 26371 8229
rect 26693 8183 27597 8230
rect 25833 8059 25867 8182
rect 26305 8169 26371 8182
rect 26305 8135 26321 8169
rect 26355 8135 26371 8169
rect 26305 8119 26371 8135
rect 26694 8059 26728 8183
rect 25828 8047 25874 8059
rect 25828 7871 25834 8047
rect 25868 7871 25874 8047
rect 25828 7859 25874 7871
rect 25946 8047 26066 8059
rect 25946 7871 25952 8047
rect 25986 7871 26026 8047
rect 25946 7859 26026 7871
rect 25952 7492 25986 7859
rect 26020 7671 26026 7859
rect 26060 7671 26066 8047
rect 26020 7659 26066 7671
rect 26138 8047 26184 8059
rect 26138 7671 26144 8047
rect 26178 7671 26184 8047
rect 26138 7659 26184 7671
rect 26256 8047 26302 8059
rect 26256 7671 26262 8047
rect 26296 7671 26302 8047
rect 26256 7659 26302 7671
rect 26374 8047 26420 8059
rect 26374 7671 26380 8047
rect 26414 7671 26420 8047
rect 26374 7659 26420 7671
rect 26492 8047 26616 8059
rect 26492 7671 26498 8047
rect 26532 7871 26576 8047
rect 26610 7871 26616 8047
rect 26532 7859 26616 7871
rect 26688 8047 26734 8059
rect 26688 7871 26694 8047
rect 26728 7871 26734 8047
rect 26688 7859 26734 7871
rect 26532 7671 26538 7859
rect 26492 7659 26538 7671
rect 26262 7586 26296 7659
rect 26247 7570 26313 7586
rect 26247 7536 26263 7570
rect 26297 7536 26313 7570
rect 26247 7520 26313 7536
rect 26576 7492 26610 7859
rect 25952 7440 26610 7492
rect 26250 7418 26342 7440
rect 26250 7366 26262 7418
rect 26328 7366 26342 7418
rect 26250 7362 26342 7366
rect 24782 6890 25113 6954
rect 24747 6737 24757 6751
rect 24717 6731 24757 6737
rect 24833 6737 24843 6751
rect 24833 6731 24875 6737
rect 24717 6695 24743 6731
rect 24839 6695 24875 6731
rect 24717 6677 24757 6695
rect 24833 6677 24875 6695
rect 24717 6637 24875 6677
rect 24593 6591 24875 6637
rect 24593 6545 24639 6591
rect 24593 6369 24599 6545
rect 24633 6369 24639 6545
rect 24593 6357 24639 6369
rect 24711 6545 24757 6557
rect 24711 6369 24717 6545
rect 24751 6369 24757 6545
rect 24711 6357 24757 6369
rect 24829 6545 24875 6591
rect 24829 6369 24835 6545
rect 24869 6369 24875 6545
rect 24829 6357 24875 6369
rect 24947 6545 24993 6557
rect 24947 6369 24953 6545
rect 24987 6369 24993 6545
rect 24947 6367 24993 6369
rect 24947 6285 24995 6367
rect 25049 6285 25113 6890
rect 23848 6269 23896 6281
rect 23848 6223 23854 6269
rect 23890 6263 24083 6269
rect 23890 6229 24037 6263
rect 24071 6229 24083 6263
rect 23890 6223 24083 6229
rect 21993 6175 22041 6221
rect 22733 6175 22781 6221
rect 23471 6175 23519 6221
rect 23848 6211 23896 6223
rect 24202 6218 24373 6282
rect 24585 6269 24635 6281
rect 24585 6223 24591 6269
rect 24629 6263 24821 6269
rect 24629 6229 24775 6263
rect 24809 6229 24821 6263
rect 24629 6223 24821 6229
rect 24209 6175 24257 6218
rect 24585 6211 24635 6223
rect 24943 6221 25113 6285
rect 24947 6175 24995 6221
rect 19657 5985 19663 6161
rect 19697 6147 19823 6161
rect 20277 6163 20323 6175
rect 19697 5985 19703 6147
rect 19657 5973 19703 5985
rect 20277 5987 20283 6163
rect 20317 5987 20323 6163
rect 19499 5805 19509 5871
rect 19611 5805 19621 5871
rect 20277 5869 20323 5987
rect 20395 6163 20561 6175
rect 20395 5987 20401 6163
rect 20435 6145 20561 6163
rect 21015 6159 21061 6171
rect 20435 5987 20441 6145
rect 20395 5975 20441 5987
rect 21015 5983 21021 6159
rect 21055 5983 21061 6159
rect 21015 5869 21061 5983
rect 21133 6159 21299 6175
rect 21133 5983 21139 6159
rect 21173 6145 21299 6159
rect 21757 6159 21803 6171
rect 21173 5983 21179 6145
rect 21133 5971 21179 5983
rect 21757 5983 21763 6159
rect 21797 5983 21803 6159
rect 21757 5869 21803 5983
rect 21875 6159 22041 6175
rect 21875 5983 21881 6159
rect 21915 6145 22041 6159
rect 22497 6159 22543 6171
rect 21915 5983 21921 6145
rect 21875 5971 21921 5983
rect 22497 5983 22503 6159
rect 22537 5983 22543 6159
rect 22497 5869 22543 5983
rect 22615 6159 22781 6175
rect 22615 5983 22621 6159
rect 22655 6145 22781 6159
rect 23235 6159 23281 6171
rect 22655 5983 22661 6145
rect 22615 5971 22661 5983
rect 23235 5983 23241 6159
rect 23275 5983 23281 6159
rect 23235 5869 23281 5983
rect 23353 6159 23519 6175
rect 23353 5983 23359 6159
rect 23393 6145 23519 6159
rect 23973 6163 24019 6175
rect 23393 5983 23399 6145
rect 23353 5971 23399 5983
rect 23973 5987 23979 6163
rect 24013 5987 24019 6163
rect 23973 5869 24019 5987
rect 24091 6163 24257 6175
rect 24091 5987 24097 6163
rect 24131 6145 24257 6163
rect 24711 6163 24757 6175
rect 24131 5987 24137 6145
rect 24091 5975 24137 5987
rect 24711 5987 24717 6163
rect 24751 5987 24757 6163
rect 24711 5869 24757 5987
rect 24829 6163 24995 6175
rect 24829 5987 24835 6163
rect 24869 6145 24995 6163
rect 24869 5987 24875 6145
rect 24829 5975 24875 5987
rect 20237 5803 20247 5869
rect 20349 5803 20359 5869
rect 20975 5803 20985 5869
rect 21087 5803 21097 5869
rect 21717 5803 21727 5869
rect 21829 5803 21839 5869
rect 22457 5803 22467 5869
rect 22569 5803 22579 5869
rect 23195 5803 23205 5869
rect 23307 5803 23317 5869
rect 23933 5803 23943 5869
rect 24045 5803 24055 5869
rect 24671 5803 24681 5869
rect 24783 5803 24793 5869
rect 18801 5338 18927 5344
rect 18801 5236 18813 5338
rect 18915 5236 18927 5338
rect 18801 5230 18927 5236
rect 18442 5194 18749 5195
rect 17299 5189 17615 5194
rect 18329 5189 18749 5194
rect 17299 5178 17682 5189
rect 17299 5151 17631 5178
rect 17299 5022 17333 5151
rect 17615 5144 17631 5151
rect 17665 5144 17682 5178
rect 17615 5138 17682 5144
rect 18262 5178 18749 5189
rect 18262 5144 18279 5178
rect 18313 5151 18749 5178
rect 18313 5144 18329 5151
rect 18442 5150 18749 5151
rect 18262 5138 18329 5144
rect 17440 5111 17496 5123
rect 17440 5077 17446 5111
rect 17480 5110 17496 5111
rect 18553 5110 18609 5122
rect 17480 5094 17947 5110
rect 17480 5077 17897 5094
rect 17440 5061 17897 5077
rect 17881 5060 17897 5061
rect 17931 5060 17947 5094
rect 17881 5053 17947 5060
rect 17999 5095 18569 5110
rect 17999 5061 18015 5095
rect 18049 5076 18569 5095
rect 18603 5076 18609 5110
rect 18049 5061 18609 5076
rect 17999 5051 18066 5061
rect 18553 5060 18609 5061
rect 18715 5022 18749 5150
rect 17293 5010 17339 5022
rect 17293 4834 17299 5010
rect 17333 4834 17339 5010
rect 17293 4822 17339 4834
rect 17411 5010 17457 5022
rect 17411 4834 17417 5010
rect 17451 4834 17457 5010
rect 17411 4822 17457 4834
rect 17713 5010 17759 5022
rect 17416 4528 17450 4822
rect 17713 4634 17719 5010
rect 17753 4634 17759 5010
rect 17713 4622 17759 4634
rect 17831 5010 17877 5022
rect 17831 4634 17837 5010
rect 17871 4634 17877 5010
rect 17831 4622 17877 4634
rect 17949 5010 17995 5022
rect 17949 4634 17955 5010
rect 17989 4634 17995 5010
rect 17949 4622 17995 4634
rect 18067 5010 18113 5022
rect 18067 4634 18073 5010
rect 18107 4634 18113 5010
rect 18067 4622 18113 4634
rect 18185 5010 18231 5022
rect 18185 4634 18191 5010
rect 18225 4634 18231 5010
rect 18591 5010 18637 5022
rect 18591 4834 18597 5010
rect 18631 4834 18637 5010
rect 18591 4822 18637 4834
rect 18709 5010 18755 5022
rect 18709 4834 18715 5010
rect 18749 4834 18755 5010
rect 18709 4822 18755 4834
rect 18185 4622 18231 4634
rect 18073 4528 18107 4622
rect 18597 4528 18630 4822
rect 17416 4496 18630 4528
rect 17909 4474 18041 4496
rect 17909 4416 17943 4474
rect 18005 4416 18041 4474
rect 17909 4411 18041 4416
rect 17122 3404 17188 3415
rect 721 3403 17188 3404
rect 721 3349 17129 3403
rect 17182 3349 17188 3403
rect 721 3326 17188 3349
rect 1498 2324 1508 2384
rect 1588 2324 1598 2384
rect 1498 2284 1598 2324
rect 4642 2324 4652 2384
rect 4732 2324 4742 2384
rect 4642 2284 4742 2324
rect 7774 2328 7784 2388
rect 7864 2328 7874 2388
rect 7774 2288 7874 2328
rect 10918 2328 10928 2388
rect 11008 2328 11018 2388
rect 10918 2288 11018 2328
rect 14120 2324 14130 2384
rect 14210 2324 14220 2384
rect 701 2227 2504 2284
rect 701 2140 735 2227
rect 1876 2140 1910 2227
rect 695 2128 741 2140
rect 695 1940 701 2128
rect 254 1928 300 1940
rect 254 1752 260 1928
rect 294 1752 300 1928
rect 254 1740 300 1752
rect 372 1928 418 1940
rect 372 1752 378 1928
rect 412 1752 418 1928
rect 372 1740 418 1752
rect 490 1928 536 1940
rect 490 1752 496 1928
rect 530 1752 536 1928
rect 490 1740 536 1752
rect 608 1928 701 1940
rect 608 1752 614 1928
rect 648 1752 701 1928
rect 735 1752 741 2128
rect 608 1740 741 1752
rect 813 2128 859 2140
rect 813 1752 819 2128
rect 853 1752 859 2128
rect 813 1740 859 1752
rect 931 2128 977 2140
rect 931 1752 937 2128
rect 971 1752 977 2128
rect 931 1740 977 1752
rect 1049 2128 1095 2140
rect 1049 1752 1055 2128
rect 1089 1752 1095 2128
rect 1049 1740 1095 1752
rect 1162 2128 1208 2140
rect 1162 1752 1168 2128
rect 1202 1752 1208 2128
rect 1162 1740 1208 1752
rect 1280 2128 1326 2140
rect 1280 1752 1286 2128
rect 1320 1752 1326 2128
rect 1280 1740 1326 1752
rect 1398 2128 1444 2140
rect 1398 1752 1404 2128
rect 1438 1752 1444 2128
rect 1398 1740 1444 1752
rect 1516 2128 1562 2140
rect 1516 1752 1522 2128
rect 1556 1752 1562 2128
rect 1516 1740 1562 1752
rect 1634 2128 1680 2140
rect 1634 1752 1640 2128
rect 1674 1752 1680 2128
rect 1634 1740 1680 1752
rect 1752 2128 1798 2140
rect 1752 1752 1758 2128
rect 1792 1752 1798 2128
rect 1752 1740 1798 1752
rect 1870 2128 1916 2140
rect 1870 1752 1876 2128
rect 1910 1752 1916 2128
rect 1870 1740 1916 1752
rect 1989 2128 2035 2140
rect 1989 1752 1995 2128
rect 2029 1752 2035 2128
rect 1989 1740 2035 1752
rect 2107 2128 2153 2140
rect 2107 1752 2113 2128
rect 2147 1752 2153 2128
rect 2107 1740 2153 1752
rect 2225 2128 2271 2140
rect 2225 1752 2231 2128
rect 2265 1752 2271 2128
rect 2225 1740 2271 1752
rect 2343 2128 2389 2140
rect 2343 1752 2349 2128
rect 2383 1752 2389 2128
rect 2467 1940 2504 2227
rect 3845 2227 5648 2284
rect 3845 2140 3879 2227
rect 5020 2140 5054 2227
rect 3839 2128 3885 2140
rect 3839 1940 3845 2128
rect 2343 1740 2389 1752
rect 2462 1928 2508 1940
rect 2462 1752 2468 1928
rect 2502 1752 2508 1928
rect 2462 1740 2508 1752
rect 2580 1928 2626 1940
rect 2580 1752 2586 1928
rect 2620 1752 2626 1928
rect 2580 1740 2626 1752
rect 2698 1928 2744 1940
rect 2698 1752 2704 1928
rect 2738 1752 2744 1928
rect 2698 1740 2744 1752
rect 2816 1928 2862 1940
rect 2816 1752 2822 1928
rect 2856 1752 2862 1928
rect 2816 1740 2862 1752
rect 3398 1928 3444 1940
rect 3398 1752 3404 1928
rect 3438 1752 3444 1928
rect 3398 1740 3444 1752
rect 3516 1928 3562 1940
rect 3516 1752 3522 1928
rect 3556 1752 3562 1928
rect 3516 1740 3562 1752
rect 3634 1928 3680 1940
rect 3634 1752 3640 1928
rect 3674 1752 3680 1928
rect 3634 1740 3680 1752
rect 3752 1928 3845 1940
rect 3752 1752 3758 1928
rect 3792 1752 3845 1928
rect 3879 1752 3885 2128
rect 3752 1740 3885 1752
rect 3957 2128 4003 2140
rect 3957 1752 3963 2128
rect 3997 1752 4003 2128
rect 3957 1740 4003 1752
rect 4075 2128 4121 2140
rect 4075 1752 4081 2128
rect 4115 1752 4121 2128
rect 4075 1740 4121 1752
rect 4193 2128 4239 2140
rect 4193 1752 4199 2128
rect 4233 1752 4239 2128
rect 4193 1740 4239 1752
rect 4306 2128 4352 2140
rect 4306 1752 4312 2128
rect 4346 1752 4352 2128
rect 4306 1740 4352 1752
rect 4424 2128 4470 2140
rect 4424 1752 4430 2128
rect 4464 1752 4470 2128
rect 4424 1740 4470 1752
rect 4542 2128 4588 2140
rect 4542 1752 4548 2128
rect 4582 1752 4588 2128
rect 4542 1740 4588 1752
rect 4660 2128 4706 2140
rect 4660 1752 4666 2128
rect 4700 1752 4706 2128
rect 4660 1740 4706 1752
rect 4778 2128 4824 2140
rect 4778 1752 4784 2128
rect 4818 1752 4824 2128
rect 4778 1740 4824 1752
rect 4896 2128 4942 2140
rect 4896 1752 4902 2128
rect 4936 1752 4942 2128
rect 4896 1740 4942 1752
rect 5014 2128 5060 2140
rect 5014 1752 5020 2128
rect 5054 1752 5060 2128
rect 5014 1740 5060 1752
rect 5133 2128 5179 2140
rect 5133 1752 5139 2128
rect 5173 1752 5179 2128
rect 5133 1740 5179 1752
rect 5251 2128 5297 2140
rect 5251 1752 5257 2128
rect 5291 1752 5297 2128
rect 5251 1740 5297 1752
rect 5369 2128 5415 2140
rect 5369 1752 5375 2128
rect 5409 1752 5415 2128
rect 5369 1740 5415 1752
rect 5487 2128 5533 2140
rect 5487 1752 5493 2128
rect 5527 1752 5533 2128
rect 5611 1940 5648 2227
rect 6977 2231 8780 2288
rect 6977 2144 7011 2231
rect 8152 2144 8186 2231
rect 6971 2132 7017 2144
rect 6971 1944 6977 2132
rect 5487 1740 5533 1752
rect 5606 1928 5652 1940
rect 5606 1752 5612 1928
rect 5646 1752 5652 1928
rect 5606 1740 5652 1752
rect 5724 1928 5770 1940
rect 5724 1752 5730 1928
rect 5764 1752 5770 1928
rect 5724 1740 5770 1752
rect 5842 1928 5888 1940
rect 5842 1752 5848 1928
rect 5882 1752 5888 1928
rect 5842 1740 5888 1752
rect 5960 1928 6006 1940
rect 5960 1752 5966 1928
rect 6000 1752 6006 1928
rect 5960 1740 6006 1752
rect 6530 1932 6576 1944
rect 6530 1756 6536 1932
rect 6570 1756 6576 1932
rect 6530 1744 6576 1756
rect 6648 1932 6694 1944
rect 6648 1756 6654 1932
rect 6688 1756 6694 1932
rect 6648 1744 6694 1756
rect 6766 1932 6812 1944
rect 6766 1756 6772 1932
rect 6806 1756 6812 1932
rect 6766 1744 6812 1756
rect 6884 1932 6977 1944
rect 6884 1756 6890 1932
rect 6924 1756 6977 1932
rect 7011 1756 7017 2132
rect 6884 1744 7017 1756
rect 7089 2132 7135 2144
rect 7089 1756 7095 2132
rect 7129 1756 7135 2132
rect 7089 1744 7135 1756
rect 7207 2132 7253 2144
rect 7207 1756 7213 2132
rect 7247 1756 7253 2132
rect 7207 1744 7253 1756
rect 7325 2132 7371 2144
rect 7325 1756 7331 2132
rect 7365 1756 7371 2132
rect 7325 1744 7371 1756
rect 7438 2132 7484 2144
rect 7438 1756 7444 2132
rect 7478 1756 7484 2132
rect 7438 1744 7484 1756
rect 7556 2132 7602 2144
rect 7556 1756 7562 2132
rect 7596 1756 7602 2132
rect 7556 1744 7602 1756
rect 7674 2132 7720 2144
rect 7674 1756 7680 2132
rect 7714 1756 7720 2132
rect 7674 1744 7720 1756
rect 7792 2132 7838 2144
rect 7792 1756 7798 2132
rect 7832 1756 7838 2132
rect 7792 1744 7838 1756
rect 7910 2132 7956 2144
rect 7910 1756 7916 2132
rect 7950 1756 7956 2132
rect 7910 1744 7956 1756
rect 8028 2132 8074 2144
rect 8028 1756 8034 2132
rect 8068 1756 8074 2132
rect 8028 1744 8074 1756
rect 8146 2132 8192 2144
rect 8146 1756 8152 2132
rect 8186 1756 8192 2132
rect 8146 1744 8192 1756
rect 8265 2132 8311 2144
rect 8265 1756 8271 2132
rect 8305 1756 8311 2132
rect 8265 1744 8311 1756
rect 8383 2132 8429 2144
rect 8383 1756 8389 2132
rect 8423 1756 8429 2132
rect 8383 1744 8429 1756
rect 8501 2132 8547 2144
rect 8501 1756 8507 2132
rect 8541 1756 8547 2132
rect 8501 1744 8547 1756
rect 8619 2132 8665 2144
rect 8619 1756 8625 2132
rect 8659 1756 8665 2132
rect 8743 1944 8780 2231
rect 10121 2231 11924 2288
rect 14120 2284 14220 2324
rect 17264 2324 17274 2384
rect 17354 2324 17364 2384
rect 17264 2284 17364 2324
rect 20396 2328 20406 2388
rect 20486 2328 20496 2388
rect 20396 2288 20496 2328
rect 23540 2328 23550 2388
rect 23630 2328 23640 2388
rect 23540 2288 23640 2328
rect 10121 2144 10155 2231
rect 11296 2144 11330 2231
rect 10115 2132 10161 2144
rect 10115 1944 10121 2132
rect 8619 1744 8665 1756
rect 8738 1932 8784 1944
rect 8738 1756 8744 1932
rect 8778 1756 8784 1932
rect 8738 1744 8784 1756
rect 8856 1932 8902 1944
rect 8856 1756 8862 1932
rect 8896 1756 8902 1932
rect 8856 1744 8902 1756
rect 8974 1932 9020 1944
rect 8974 1756 8980 1932
rect 9014 1756 9020 1932
rect 8974 1744 9020 1756
rect 9092 1932 9138 1944
rect 9092 1756 9098 1932
rect 9132 1756 9138 1932
rect 9092 1744 9138 1756
rect 9674 1932 9720 1944
rect 9674 1756 9680 1932
rect 9714 1756 9720 1932
rect 9674 1744 9720 1756
rect 9792 1932 9838 1944
rect 9792 1756 9798 1932
rect 9832 1756 9838 1932
rect 9792 1744 9838 1756
rect 9910 1932 9956 1944
rect 9910 1756 9916 1932
rect 9950 1756 9956 1932
rect 9910 1744 9956 1756
rect 10028 1932 10121 1944
rect 10028 1756 10034 1932
rect 10068 1756 10121 1932
rect 10155 1756 10161 2132
rect 10028 1744 10161 1756
rect 10233 2132 10279 2144
rect 10233 1756 10239 2132
rect 10273 1756 10279 2132
rect 10233 1744 10279 1756
rect 10351 2132 10397 2144
rect 10351 1756 10357 2132
rect 10391 1756 10397 2132
rect 10351 1744 10397 1756
rect 10469 2132 10515 2144
rect 10469 1756 10475 2132
rect 10509 1756 10515 2132
rect 10469 1744 10515 1756
rect 10582 2132 10628 2144
rect 10582 1756 10588 2132
rect 10622 1756 10628 2132
rect 10582 1744 10628 1756
rect 10700 2132 10746 2144
rect 10700 1756 10706 2132
rect 10740 1756 10746 2132
rect 10700 1744 10746 1756
rect 10818 2132 10864 2144
rect 10818 1756 10824 2132
rect 10858 1756 10864 2132
rect 10818 1744 10864 1756
rect 10936 2132 10982 2144
rect 10936 1756 10942 2132
rect 10976 1756 10982 2132
rect 10936 1744 10982 1756
rect 11054 2132 11100 2144
rect 11054 1756 11060 2132
rect 11094 1756 11100 2132
rect 11054 1744 11100 1756
rect 11172 2132 11218 2144
rect 11172 1756 11178 2132
rect 11212 1756 11218 2132
rect 11172 1744 11218 1756
rect 11290 2132 11336 2144
rect 11290 1756 11296 2132
rect 11330 1756 11336 2132
rect 11290 1744 11336 1756
rect 11409 2132 11455 2144
rect 11409 1756 11415 2132
rect 11449 1756 11455 2132
rect 11409 1744 11455 1756
rect 11527 2132 11573 2144
rect 11527 1756 11533 2132
rect 11567 1756 11573 2132
rect 11527 1744 11573 1756
rect 11645 2132 11691 2144
rect 11645 1756 11651 2132
rect 11685 1756 11691 2132
rect 11645 1744 11691 1756
rect 11763 2132 11809 2144
rect 11763 1756 11769 2132
rect 11803 1756 11809 2132
rect 11887 1944 11924 2231
rect 13323 2227 15126 2284
rect 13323 2140 13357 2227
rect 14498 2140 14532 2227
rect 13317 2128 13363 2140
rect 11763 1744 11809 1756
rect 11882 1932 11928 1944
rect 11882 1756 11888 1932
rect 11922 1756 11928 1932
rect 11882 1744 11928 1756
rect 12000 1932 12046 1944
rect 12000 1756 12006 1932
rect 12040 1756 12046 1932
rect 12000 1744 12046 1756
rect 12118 1932 12164 1944
rect 12118 1756 12124 1932
rect 12158 1756 12164 1932
rect 12118 1744 12164 1756
rect 12236 1932 12282 1944
rect 13317 1940 13323 2128
rect 12236 1756 12242 1932
rect 12276 1756 12282 1932
rect 12236 1744 12282 1756
rect 12876 1928 12922 1940
rect 12876 1752 12882 1928
rect 12916 1752 12922 1928
rect 259 1554 294 1740
rect 1168 1656 1202 1740
rect 2349 1656 2383 1740
rect 1168 1614 2383 1656
rect 2349 1594 2383 1614
rect 2349 1578 2706 1594
rect 259 1537 1396 1554
rect 259 1503 1346 1537
rect 1380 1503 1396 1537
rect 2349 1544 2656 1578
rect 2690 1544 2706 1578
rect 2349 1528 2706 1544
rect 259 1487 1396 1503
rect 0 1442 176 1450
rect 0 1374 117 1442
rect 174 1374 184 1442
rect 0 1366 176 1374
rect 0 1326 176 1334
rect 0 1258 117 1326
rect 174 1258 184 1326
rect 0 1250 176 1258
rect 0 1158 176 1166
rect 0 1090 117 1158
rect 174 1090 184 1158
rect 0 1082 176 1090
rect 259 977 294 1487
rect 349 1441 441 1454
rect 349 1378 361 1441
rect 432 1378 441 1441
rect 349 1369 441 1378
rect 1434 1441 1526 1451
rect 1434 1379 1446 1441
rect 1516 1379 1526 1441
rect 1434 1366 1526 1379
rect 2822 1386 2857 1740
rect 3403 1554 3438 1740
rect 4312 1656 4346 1740
rect 5493 1656 5527 1740
rect 4312 1614 5527 1656
rect 5493 1594 5527 1614
rect 5493 1578 5850 1594
rect 3403 1537 4540 1554
rect 3403 1503 4490 1537
rect 4524 1503 4540 1537
rect 5493 1544 5800 1578
rect 5834 1544 5850 1578
rect 5493 1528 5850 1544
rect 3403 1487 4540 1503
rect 3144 1442 3320 1450
rect 1681 1324 1746 1327
rect 1681 1321 1750 1324
rect 1681 1261 1687 1321
rect 1746 1261 1756 1321
rect 1681 1257 1750 1261
rect 1681 1255 1746 1257
rect 2822 1240 3003 1386
rect 3144 1374 3261 1442
rect 3318 1374 3328 1442
rect 3144 1366 3320 1374
rect 3144 1326 3320 1334
rect 3144 1258 3261 1326
rect 3318 1258 3328 1326
rect 3144 1250 3320 1258
rect 1316 1158 1408 1166
rect 1316 1093 1328 1158
rect 1396 1093 1408 1158
rect 1316 1081 1408 1093
rect 2822 978 2857 1240
rect 3144 1158 3320 1166
rect 3144 1090 3261 1158
rect 3318 1090 3328 1158
rect 3144 1082 3320 1090
rect 259 930 1631 977
rect 1953 931 2857 978
rect 3403 977 3438 1487
rect 3493 1441 3585 1454
rect 3493 1378 3505 1441
rect 3576 1378 3585 1441
rect 3493 1369 3585 1378
rect 4578 1441 4670 1451
rect 4578 1379 4590 1441
rect 4660 1379 4670 1441
rect 4578 1366 4670 1379
rect 5966 1386 6001 1740
rect 6535 1558 6570 1744
rect 7444 1660 7478 1744
rect 8625 1660 8659 1744
rect 7444 1618 8659 1660
rect 8625 1598 8659 1618
rect 8625 1582 8982 1598
rect 6535 1541 7672 1558
rect 6535 1507 7622 1541
rect 7656 1507 7672 1541
rect 8625 1548 8932 1582
rect 8966 1548 8982 1582
rect 8625 1532 8982 1548
rect 6535 1491 7672 1507
rect 6276 1446 6452 1454
rect 4825 1324 4890 1327
rect 4825 1321 4894 1324
rect 4825 1261 4831 1321
rect 4890 1261 4900 1321
rect 4825 1257 4894 1261
rect 4825 1255 4890 1257
rect 5966 1240 6147 1386
rect 6276 1378 6393 1446
rect 6450 1378 6460 1446
rect 6276 1370 6452 1378
rect 6276 1330 6452 1338
rect 6276 1262 6393 1330
rect 6450 1262 6460 1330
rect 6276 1254 6452 1262
rect 4460 1158 4552 1166
rect 4460 1093 4472 1158
rect 4540 1093 4552 1158
rect 4460 1081 4552 1093
rect 5966 978 6001 1240
rect 6276 1162 6452 1170
rect 6276 1094 6393 1162
rect 6450 1094 6460 1162
rect 6276 1086 6452 1094
rect 1093 807 1127 930
rect 1565 917 1631 930
rect 1565 883 1581 917
rect 1615 883 1631 917
rect 1565 867 1631 883
rect 1954 807 1988 931
rect 3403 930 4775 977
rect 5097 931 6001 978
rect 6535 981 6570 1491
rect 6625 1445 6717 1458
rect 6625 1382 6637 1445
rect 6708 1382 6717 1445
rect 6625 1373 6717 1382
rect 7710 1445 7802 1455
rect 7710 1383 7722 1445
rect 7792 1383 7802 1445
rect 7710 1370 7802 1383
rect 9098 1390 9133 1744
rect 9679 1558 9714 1744
rect 10588 1660 10622 1744
rect 11769 1660 11803 1744
rect 10588 1618 11803 1660
rect 11769 1598 11803 1618
rect 11769 1582 12126 1598
rect 9679 1541 10816 1558
rect 9679 1507 10766 1541
rect 10800 1507 10816 1541
rect 11769 1548 12076 1582
rect 12110 1548 12126 1582
rect 11769 1532 12126 1548
rect 9679 1491 10816 1507
rect 9420 1446 9596 1454
rect 7957 1328 8022 1331
rect 7957 1325 8026 1328
rect 7957 1265 7963 1325
rect 8022 1265 8032 1325
rect 7957 1261 8026 1265
rect 7957 1259 8022 1261
rect 9098 1244 9279 1390
rect 9420 1378 9537 1446
rect 9594 1378 9604 1446
rect 9420 1370 9596 1378
rect 9420 1330 9596 1338
rect 9420 1262 9537 1330
rect 9594 1262 9604 1330
rect 9420 1254 9596 1262
rect 7592 1162 7684 1170
rect 7592 1097 7604 1162
rect 7672 1097 7684 1162
rect 7592 1085 7684 1097
rect 9098 982 9133 1244
rect 9420 1162 9596 1170
rect 9420 1094 9537 1162
rect 9594 1094 9604 1162
rect 9420 1086 9596 1094
rect 6535 934 7907 981
rect 8229 935 9133 982
rect 9679 981 9714 1491
rect 9769 1445 9861 1458
rect 9769 1382 9781 1445
rect 9852 1382 9861 1445
rect 9769 1373 9861 1382
rect 10854 1445 10946 1455
rect 10854 1383 10866 1445
rect 10936 1383 10946 1445
rect 10854 1370 10946 1383
rect 12242 1390 12277 1744
rect 12876 1740 12922 1752
rect 12994 1928 13040 1940
rect 12994 1752 13000 1928
rect 13034 1752 13040 1928
rect 12994 1740 13040 1752
rect 13112 1928 13158 1940
rect 13112 1752 13118 1928
rect 13152 1752 13158 1928
rect 13112 1740 13158 1752
rect 13230 1928 13323 1940
rect 13230 1752 13236 1928
rect 13270 1752 13323 1928
rect 13357 1752 13363 2128
rect 13230 1740 13363 1752
rect 13435 2128 13481 2140
rect 13435 1752 13441 2128
rect 13475 1752 13481 2128
rect 13435 1740 13481 1752
rect 13553 2128 13599 2140
rect 13553 1752 13559 2128
rect 13593 1752 13599 2128
rect 13553 1740 13599 1752
rect 13671 2128 13717 2140
rect 13671 1752 13677 2128
rect 13711 1752 13717 2128
rect 13671 1740 13717 1752
rect 13784 2128 13830 2140
rect 13784 1752 13790 2128
rect 13824 1752 13830 2128
rect 13784 1740 13830 1752
rect 13902 2128 13948 2140
rect 13902 1752 13908 2128
rect 13942 1752 13948 2128
rect 13902 1740 13948 1752
rect 14020 2128 14066 2140
rect 14020 1752 14026 2128
rect 14060 1752 14066 2128
rect 14020 1740 14066 1752
rect 14138 2128 14184 2140
rect 14138 1752 14144 2128
rect 14178 1752 14184 2128
rect 14138 1740 14184 1752
rect 14256 2128 14302 2140
rect 14256 1752 14262 2128
rect 14296 1752 14302 2128
rect 14256 1740 14302 1752
rect 14374 2128 14420 2140
rect 14374 1752 14380 2128
rect 14414 1752 14420 2128
rect 14374 1740 14420 1752
rect 14492 2128 14538 2140
rect 14492 1752 14498 2128
rect 14532 1752 14538 2128
rect 14492 1740 14538 1752
rect 14611 2128 14657 2140
rect 14611 1752 14617 2128
rect 14651 1752 14657 2128
rect 14611 1740 14657 1752
rect 14729 2128 14775 2140
rect 14729 1752 14735 2128
rect 14769 1752 14775 2128
rect 14729 1740 14775 1752
rect 14847 2128 14893 2140
rect 14847 1752 14853 2128
rect 14887 1752 14893 2128
rect 14847 1740 14893 1752
rect 14965 2128 15011 2140
rect 14965 1752 14971 2128
rect 15005 1752 15011 2128
rect 15089 1940 15126 2227
rect 16467 2227 18270 2284
rect 16467 2140 16501 2227
rect 17642 2140 17676 2227
rect 16461 2128 16507 2140
rect 16461 1940 16467 2128
rect 14965 1740 15011 1752
rect 15084 1928 15130 1940
rect 15084 1752 15090 1928
rect 15124 1752 15130 1928
rect 15084 1740 15130 1752
rect 15202 1928 15248 1940
rect 15202 1752 15208 1928
rect 15242 1752 15248 1928
rect 15202 1740 15248 1752
rect 15320 1928 15366 1940
rect 15320 1752 15326 1928
rect 15360 1752 15366 1928
rect 15320 1740 15366 1752
rect 15438 1928 15484 1940
rect 15438 1752 15444 1928
rect 15478 1752 15484 1928
rect 15438 1740 15484 1752
rect 16020 1928 16066 1940
rect 16020 1752 16026 1928
rect 16060 1752 16066 1928
rect 16020 1740 16066 1752
rect 16138 1928 16184 1940
rect 16138 1752 16144 1928
rect 16178 1752 16184 1928
rect 16138 1740 16184 1752
rect 16256 1928 16302 1940
rect 16256 1752 16262 1928
rect 16296 1752 16302 1928
rect 16256 1740 16302 1752
rect 16374 1928 16467 1940
rect 16374 1752 16380 1928
rect 16414 1752 16467 1928
rect 16501 1752 16507 2128
rect 16374 1740 16507 1752
rect 16579 2128 16625 2140
rect 16579 1752 16585 2128
rect 16619 1752 16625 2128
rect 16579 1740 16625 1752
rect 16697 2128 16743 2140
rect 16697 1752 16703 2128
rect 16737 1752 16743 2128
rect 16697 1740 16743 1752
rect 16815 2128 16861 2140
rect 16815 1752 16821 2128
rect 16855 1752 16861 2128
rect 16815 1740 16861 1752
rect 16928 2128 16974 2140
rect 16928 1752 16934 2128
rect 16968 1752 16974 2128
rect 16928 1740 16974 1752
rect 17046 2128 17092 2140
rect 17046 1752 17052 2128
rect 17086 1752 17092 2128
rect 17046 1740 17092 1752
rect 17164 2128 17210 2140
rect 17164 1752 17170 2128
rect 17204 1752 17210 2128
rect 17164 1740 17210 1752
rect 17282 2128 17328 2140
rect 17282 1752 17288 2128
rect 17322 1752 17328 2128
rect 17282 1740 17328 1752
rect 17400 2128 17446 2140
rect 17400 1752 17406 2128
rect 17440 1752 17446 2128
rect 17400 1740 17446 1752
rect 17518 2128 17564 2140
rect 17518 1752 17524 2128
rect 17558 1752 17564 2128
rect 17518 1740 17564 1752
rect 17636 2128 17682 2140
rect 17636 1752 17642 2128
rect 17676 1752 17682 2128
rect 17636 1740 17682 1752
rect 17755 2128 17801 2140
rect 17755 1752 17761 2128
rect 17795 1752 17801 2128
rect 17755 1740 17801 1752
rect 17873 2128 17919 2140
rect 17873 1752 17879 2128
rect 17913 1752 17919 2128
rect 17873 1740 17919 1752
rect 17991 2128 18037 2140
rect 17991 1752 17997 2128
rect 18031 1752 18037 2128
rect 17991 1740 18037 1752
rect 18109 2128 18155 2140
rect 18109 1752 18115 2128
rect 18149 1752 18155 2128
rect 18233 1940 18270 2227
rect 19599 2231 21402 2288
rect 19599 2144 19633 2231
rect 20774 2144 20808 2231
rect 19593 2132 19639 2144
rect 19593 1944 19599 2132
rect 18109 1740 18155 1752
rect 18228 1928 18274 1940
rect 18228 1752 18234 1928
rect 18268 1752 18274 1928
rect 18228 1740 18274 1752
rect 18346 1928 18392 1940
rect 18346 1752 18352 1928
rect 18386 1752 18392 1928
rect 18346 1740 18392 1752
rect 18464 1928 18510 1940
rect 18464 1752 18470 1928
rect 18504 1752 18510 1928
rect 18464 1740 18510 1752
rect 18582 1928 18628 1940
rect 18582 1752 18588 1928
rect 18622 1752 18628 1928
rect 18582 1740 18628 1752
rect 19152 1932 19198 1944
rect 19152 1756 19158 1932
rect 19192 1756 19198 1932
rect 19152 1744 19198 1756
rect 19270 1932 19316 1944
rect 19270 1756 19276 1932
rect 19310 1756 19316 1932
rect 19270 1744 19316 1756
rect 19388 1932 19434 1944
rect 19388 1756 19394 1932
rect 19428 1756 19434 1932
rect 19388 1744 19434 1756
rect 19506 1932 19599 1944
rect 19506 1756 19512 1932
rect 19546 1756 19599 1932
rect 19633 1756 19639 2132
rect 19506 1744 19639 1756
rect 19711 2132 19757 2144
rect 19711 1756 19717 2132
rect 19751 1756 19757 2132
rect 19711 1744 19757 1756
rect 19829 2132 19875 2144
rect 19829 1756 19835 2132
rect 19869 1756 19875 2132
rect 19829 1744 19875 1756
rect 19947 2132 19993 2144
rect 19947 1756 19953 2132
rect 19987 1756 19993 2132
rect 19947 1744 19993 1756
rect 20060 2132 20106 2144
rect 20060 1756 20066 2132
rect 20100 1756 20106 2132
rect 20060 1744 20106 1756
rect 20178 2132 20224 2144
rect 20178 1756 20184 2132
rect 20218 1756 20224 2132
rect 20178 1744 20224 1756
rect 20296 2132 20342 2144
rect 20296 1756 20302 2132
rect 20336 1756 20342 2132
rect 20296 1744 20342 1756
rect 20414 2132 20460 2144
rect 20414 1756 20420 2132
rect 20454 1756 20460 2132
rect 20414 1744 20460 1756
rect 20532 2132 20578 2144
rect 20532 1756 20538 2132
rect 20572 1756 20578 2132
rect 20532 1744 20578 1756
rect 20650 2132 20696 2144
rect 20650 1756 20656 2132
rect 20690 1756 20696 2132
rect 20650 1744 20696 1756
rect 20768 2132 20814 2144
rect 20768 1756 20774 2132
rect 20808 1756 20814 2132
rect 20768 1744 20814 1756
rect 20887 2132 20933 2144
rect 20887 1756 20893 2132
rect 20927 1756 20933 2132
rect 20887 1744 20933 1756
rect 21005 2132 21051 2144
rect 21005 1756 21011 2132
rect 21045 1756 21051 2132
rect 21005 1744 21051 1756
rect 21123 2132 21169 2144
rect 21123 1756 21129 2132
rect 21163 1756 21169 2132
rect 21123 1744 21169 1756
rect 21241 2132 21287 2144
rect 21241 1756 21247 2132
rect 21281 1756 21287 2132
rect 21365 1944 21402 2231
rect 22743 2231 24546 2288
rect 22743 2144 22777 2231
rect 23918 2144 23952 2231
rect 22737 2132 22783 2144
rect 22737 1944 22743 2132
rect 21241 1744 21287 1756
rect 21360 1932 21406 1944
rect 21360 1756 21366 1932
rect 21400 1756 21406 1932
rect 21360 1744 21406 1756
rect 21478 1932 21524 1944
rect 21478 1756 21484 1932
rect 21518 1756 21524 1932
rect 21478 1744 21524 1756
rect 21596 1932 21642 1944
rect 21596 1756 21602 1932
rect 21636 1756 21642 1932
rect 21596 1744 21642 1756
rect 21714 1932 21760 1944
rect 21714 1756 21720 1932
rect 21754 1756 21760 1932
rect 21714 1744 21760 1756
rect 22296 1932 22342 1944
rect 22296 1756 22302 1932
rect 22336 1756 22342 1932
rect 22296 1744 22342 1756
rect 22414 1932 22460 1944
rect 22414 1756 22420 1932
rect 22454 1756 22460 1932
rect 22414 1744 22460 1756
rect 22532 1932 22578 1944
rect 22532 1756 22538 1932
rect 22572 1756 22578 1932
rect 22532 1744 22578 1756
rect 22650 1932 22743 1944
rect 22650 1756 22656 1932
rect 22690 1756 22743 1932
rect 22777 1756 22783 2132
rect 22650 1744 22783 1756
rect 22855 2132 22901 2144
rect 22855 1756 22861 2132
rect 22895 1756 22901 2132
rect 22855 1744 22901 1756
rect 22973 2132 23019 2144
rect 22973 1756 22979 2132
rect 23013 1756 23019 2132
rect 22973 1744 23019 1756
rect 23091 2132 23137 2144
rect 23091 1756 23097 2132
rect 23131 1756 23137 2132
rect 23091 1744 23137 1756
rect 23204 2132 23250 2144
rect 23204 1756 23210 2132
rect 23244 1756 23250 2132
rect 23204 1744 23250 1756
rect 23322 2132 23368 2144
rect 23322 1756 23328 2132
rect 23362 1756 23368 2132
rect 23322 1744 23368 1756
rect 23440 2132 23486 2144
rect 23440 1756 23446 2132
rect 23480 1756 23486 2132
rect 23440 1744 23486 1756
rect 23558 2132 23604 2144
rect 23558 1756 23564 2132
rect 23598 1756 23604 2132
rect 23558 1744 23604 1756
rect 23676 2132 23722 2144
rect 23676 1756 23682 2132
rect 23716 1756 23722 2132
rect 23676 1744 23722 1756
rect 23794 2132 23840 2144
rect 23794 1756 23800 2132
rect 23834 1756 23840 2132
rect 23794 1744 23840 1756
rect 23912 2132 23958 2144
rect 23912 1756 23918 2132
rect 23952 1756 23958 2132
rect 23912 1744 23958 1756
rect 24031 2132 24077 2144
rect 24031 1756 24037 2132
rect 24071 1756 24077 2132
rect 24031 1744 24077 1756
rect 24149 2132 24195 2144
rect 24149 1756 24155 2132
rect 24189 1756 24195 2132
rect 24149 1744 24195 1756
rect 24267 2132 24313 2144
rect 24267 1756 24273 2132
rect 24307 1756 24313 2132
rect 24267 1744 24313 1756
rect 24385 2132 24431 2144
rect 24385 1756 24391 2132
rect 24425 1756 24431 2132
rect 24509 1944 24546 2231
rect 24385 1744 24431 1756
rect 24504 1932 24550 1944
rect 24504 1756 24510 1932
rect 24544 1756 24550 1932
rect 24504 1744 24550 1756
rect 24622 1932 24668 1944
rect 24622 1756 24628 1932
rect 24662 1756 24668 1932
rect 24622 1744 24668 1756
rect 24740 1932 24786 1944
rect 24740 1756 24746 1932
rect 24780 1756 24786 1932
rect 24740 1744 24786 1756
rect 24858 1932 24904 1944
rect 24858 1756 24864 1932
rect 24898 1756 24904 1932
rect 24858 1744 24904 1756
rect 12881 1554 12916 1740
rect 13790 1656 13824 1740
rect 14971 1656 15005 1740
rect 13790 1614 15005 1656
rect 14971 1594 15005 1614
rect 14971 1578 15328 1594
rect 12881 1537 14018 1554
rect 12881 1503 13968 1537
rect 14002 1503 14018 1537
rect 14971 1544 15278 1578
rect 15312 1544 15328 1578
rect 14971 1528 15328 1544
rect 12881 1487 14018 1503
rect 12622 1442 12798 1450
rect 11101 1328 11166 1331
rect 11101 1325 11170 1328
rect 11101 1265 11107 1325
rect 11166 1265 11176 1325
rect 11101 1261 11170 1265
rect 11101 1259 11166 1261
rect 12242 1244 12423 1390
rect 12622 1374 12739 1442
rect 12796 1374 12806 1442
rect 12622 1366 12798 1374
rect 12622 1326 12798 1334
rect 12622 1258 12739 1326
rect 12796 1258 12806 1326
rect 12622 1250 12798 1258
rect 10736 1162 10828 1170
rect 10736 1097 10748 1162
rect 10816 1097 10828 1162
rect 10736 1085 10828 1097
rect 12242 982 12277 1244
rect 12622 1158 12798 1166
rect 12622 1090 12739 1158
rect 12796 1090 12806 1158
rect 12622 1082 12798 1090
rect 4237 807 4271 930
rect 4709 917 4775 930
rect 4709 883 4725 917
rect 4759 883 4775 917
rect 4709 867 4775 883
rect 5098 807 5132 931
rect 7369 811 7403 934
rect 7841 921 7907 934
rect 7841 887 7857 921
rect 7891 887 7907 921
rect 7841 871 7907 887
rect 8230 811 8264 935
rect 9679 934 11051 981
rect 11373 935 12277 982
rect 12881 977 12916 1487
rect 12971 1441 13063 1454
rect 12971 1378 12983 1441
rect 13054 1378 13063 1441
rect 12971 1369 13063 1378
rect 14056 1441 14148 1451
rect 14056 1379 14068 1441
rect 14138 1379 14148 1441
rect 14056 1366 14148 1379
rect 15444 1386 15479 1740
rect 16025 1554 16060 1740
rect 16934 1656 16968 1740
rect 18115 1656 18149 1740
rect 16934 1614 18149 1656
rect 18115 1594 18149 1614
rect 18115 1578 18472 1594
rect 16025 1537 17162 1554
rect 16025 1503 17112 1537
rect 17146 1503 17162 1537
rect 18115 1544 18422 1578
rect 18456 1544 18472 1578
rect 18115 1528 18472 1544
rect 16025 1487 17162 1503
rect 15766 1442 15942 1450
rect 14303 1324 14368 1327
rect 14303 1321 14372 1324
rect 14303 1261 14309 1321
rect 14368 1261 14378 1321
rect 14303 1257 14372 1261
rect 14303 1255 14368 1257
rect 15444 1240 15625 1386
rect 15766 1374 15883 1442
rect 15940 1374 15950 1442
rect 15766 1366 15942 1374
rect 15766 1326 15942 1334
rect 15766 1258 15883 1326
rect 15940 1258 15950 1326
rect 15766 1250 15942 1258
rect 13938 1158 14030 1166
rect 13938 1093 13950 1158
rect 14018 1093 14030 1158
rect 13938 1081 14030 1093
rect 15444 978 15479 1240
rect 15766 1158 15942 1166
rect 15766 1090 15883 1158
rect 15940 1090 15950 1158
rect 15766 1082 15942 1090
rect 10513 811 10547 934
rect 10985 921 11051 934
rect 10985 887 11001 921
rect 11035 887 11051 921
rect 10985 871 11051 887
rect 11374 811 11408 935
rect 12881 930 14253 977
rect 14575 931 15479 978
rect 16025 977 16060 1487
rect 16115 1441 16207 1454
rect 16115 1378 16127 1441
rect 16198 1378 16207 1441
rect 16115 1369 16207 1378
rect 17200 1441 17292 1451
rect 17200 1379 17212 1441
rect 17282 1379 17292 1441
rect 17200 1366 17292 1379
rect 18588 1386 18623 1740
rect 19157 1558 19192 1744
rect 20066 1660 20100 1744
rect 21247 1660 21281 1744
rect 20066 1618 21281 1660
rect 21247 1598 21281 1618
rect 21247 1582 21604 1598
rect 19157 1541 20294 1558
rect 19157 1507 20244 1541
rect 20278 1507 20294 1541
rect 21247 1548 21554 1582
rect 21588 1548 21604 1582
rect 21247 1532 21604 1548
rect 19157 1491 20294 1507
rect 18898 1446 19074 1454
rect 17447 1324 17512 1327
rect 17447 1321 17516 1324
rect 17447 1261 17453 1321
rect 17512 1261 17522 1321
rect 17447 1257 17516 1261
rect 17447 1255 17512 1257
rect 18588 1240 18769 1386
rect 18898 1378 19015 1446
rect 19072 1378 19082 1446
rect 18898 1370 19074 1378
rect 18898 1330 19074 1338
rect 18898 1262 19015 1330
rect 19072 1262 19082 1330
rect 18898 1254 19074 1262
rect 17082 1158 17174 1166
rect 17082 1093 17094 1158
rect 17162 1093 17174 1158
rect 17082 1081 17174 1093
rect 18588 978 18623 1240
rect 18898 1162 19074 1170
rect 18898 1094 19015 1162
rect 19072 1094 19082 1162
rect 18898 1086 19074 1094
rect 1088 795 1134 807
rect 1088 619 1094 795
rect 1128 619 1134 795
rect 1088 607 1134 619
rect 1206 795 1326 807
rect 1206 619 1212 795
rect 1246 619 1286 795
rect 1206 607 1286 619
rect 1212 240 1246 607
rect 1280 419 1286 607
rect 1320 419 1326 795
rect 1280 407 1326 419
rect 1398 795 1444 807
rect 1398 419 1404 795
rect 1438 419 1444 795
rect 1398 407 1444 419
rect 1516 795 1562 807
rect 1516 419 1522 795
rect 1556 419 1562 795
rect 1516 407 1562 419
rect 1634 795 1680 807
rect 1634 419 1640 795
rect 1674 419 1680 795
rect 1634 407 1680 419
rect 1752 795 1876 807
rect 1752 419 1758 795
rect 1792 619 1836 795
rect 1870 619 1876 795
rect 1792 607 1876 619
rect 1948 795 1994 807
rect 1948 619 1954 795
rect 1988 619 1994 795
rect 1948 607 1994 619
rect 4232 795 4278 807
rect 4232 619 4238 795
rect 4272 619 4278 795
rect 4232 607 4278 619
rect 4350 795 4470 807
rect 4350 619 4356 795
rect 4390 619 4430 795
rect 4350 607 4430 619
rect 1792 419 1798 607
rect 1752 407 1798 419
rect 1522 334 1556 407
rect 1507 318 1573 334
rect 1507 284 1523 318
rect 1557 284 1573 318
rect 1507 268 1573 284
rect 1836 240 1870 607
rect 1212 188 1870 240
rect 4356 240 4390 607
rect 4424 419 4430 607
rect 4464 419 4470 795
rect 4424 407 4470 419
rect 4542 795 4588 807
rect 4542 419 4548 795
rect 4582 419 4588 795
rect 4542 407 4588 419
rect 4660 795 4706 807
rect 4660 419 4666 795
rect 4700 419 4706 795
rect 4660 407 4706 419
rect 4778 795 4824 807
rect 4778 419 4784 795
rect 4818 419 4824 795
rect 4778 407 4824 419
rect 4896 795 5020 807
rect 4896 419 4902 795
rect 4936 619 4980 795
rect 5014 619 5020 795
rect 4936 607 5020 619
rect 5092 795 5138 807
rect 5092 619 5098 795
rect 5132 619 5138 795
rect 5092 607 5138 619
rect 7364 799 7410 811
rect 7364 623 7370 799
rect 7404 623 7410 799
rect 7364 611 7410 623
rect 7482 799 7602 811
rect 7482 623 7488 799
rect 7522 623 7562 799
rect 7482 611 7562 623
rect 4936 419 4942 607
rect 4896 407 4942 419
rect 4666 334 4700 407
rect 4651 318 4717 334
rect 4651 284 4667 318
rect 4701 284 4717 318
rect 4651 268 4717 284
rect 4980 240 5014 607
rect 4356 188 5014 240
rect 7488 244 7522 611
rect 7556 423 7562 611
rect 7596 423 7602 799
rect 7556 411 7602 423
rect 7674 799 7720 811
rect 7674 423 7680 799
rect 7714 423 7720 799
rect 7674 411 7720 423
rect 7792 799 7838 811
rect 7792 423 7798 799
rect 7832 423 7838 799
rect 7792 411 7838 423
rect 7910 799 7956 811
rect 7910 423 7916 799
rect 7950 423 7956 799
rect 7910 411 7956 423
rect 8028 799 8152 811
rect 8028 423 8034 799
rect 8068 623 8112 799
rect 8146 623 8152 799
rect 8068 611 8152 623
rect 8224 799 8270 811
rect 8224 623 8230 799
rect 8264 623 8270 799
rect 8224 611 8270 623
rect 10508 799 10554 811
rect 10508 623 10514 799
rect 10548 623 10554 799
rect 10508 611 10554 623
rect 10626 799 10746 811
rect 10626 623 10632 799
rect 10666 623 10706 799
rect 10626 611 10706 623
rect 8068 423 8074 611
rect 8028 411 8074 423
rect 7798 338 7832 411
rect 7783 322 7849 338
rect 7783 288 7799 322
rect 7833 288 7849 322
rect 7783 272 7849 288
rect 8112 244 8146 611
rect 7488 192 8146 244
rect 10632 244 10666 611
rect 10700 423 10706 611
rect 10740 423 10746 799
rect 10700 411 10746 423
rect 10818 799 10864 811
rect 10818 423 10824 799
rect 10858 423 10864 799
rect 10818 411 10864 423
rect 10936 799 10982 811
rect 10936 423 10942 799
rect 10976 423 10982 799
rect 10936 411 10982 423
rect 11054 799 11100 811
rect 11054 423 11060 799
rect 11094 423 11100 799
rect 11054 411 11100 423
rect 11172 799 11296 811
rect 11172 423 11178 799
rect 11212 623 11256 799
rect 11290 623 11296 799
rect 11212 611 11296 623
rect 11368 799 11414 811
rect 13715 807 13749 930
rect 14187 917 14253 930
rect 14187 883 14203 917
rect 14237 883 14253 917
rect 14187 867 14253 883
rect 14576 807 14610 931
rect 16025 930 17397 977
rect 17719 931 18623 978
rect 19157 981 19192 1491
rect 19247 1445 19339 1458
rect 19247 1382 19259 1445
rect 19330 1382 19339 1445
rect 19247 1373 19339 1382
rect 20332 1445 20424 1455
rect 20332 1383 20344 1445
rect 20414 1383 20424 1445
rect 20332 1370 20424 1383
rect 21720 1390 21755 1744
rect 22301 1558 22336 1744
rect 23210 1660 23244 1744
rect 24391 1660 24425 1744
rect 23210 1618 24425 1660
rect 24391 1598 24425 1618
rect 24391 1582 24748 1598
rect 22301 1541 23438 1558
rect 22301 1507 23388 1541
rect 23422 1507 23438 1541
rect 24391 1548 24698 1582
rect 24732 1548 24748 1582
rect 24391 1532 24748 1548
rect 22301 1491 23438 1507
rect 22042 1446 22218 1454
rect 20579 1328 20644 1331
rect 20579 1325 20648 1328
rect 20579 1265 20585 1325
rect 20644 1265 20654 1325
rect 20579 1261 20648 1265
rect 20579 1259 20644 1261
rect 21720 1244 21901 1390
rect 22042 1378 22159 1446
rect 22216 1378 22226 1446
rect 22042 1370 22218 1378
rect 22042 1330 22218 1338
rect 22042 1262 22159 1330
rect 22216 1262 22226 1330
rect 22042 1254 22218 1262
rect 20214 1162 20306 1170
rect 20214 1097 20226 1162
rect 20294 1097 20306 1162
rect 20214 1085 20306 1097
rect 21720 982 21755 1244
rect 22042 1162 22218 1170
rect 22042 1094 22159 1162
rect 22216 1094 22226 1162
rect 22042 1086 22218 1094
rect 19157 934 20529 981
rect 20851 935 21755 982
rect 22301 981 22336 1491
rect 22391 1445 22483 1458
rect 22391 1382 22403 1445
rect 22474 1382 22483 1445
rect 22391 1373 22483 1382
rect 23476 1445 23568 1455
rect 23476 1383 23488 1445
rect 23558 1383 23568 1445
rect 23476 1370 23568 1383
rect 24864 1390 24899 1744
rect 23723 1328 23788 1331
rect 23723 1325 23792 1328
rect 23723 1265 23729 1325
rect 23788 1265 23798 1325
rect 23723 1261 23792 1265
rect 23723 1259 23788 1261
rect 24864 1244 25045 1390
rect 23358 1162 23450 1170
rect 23358 1097 23370 1162
rect 23438 1097 23450 1162
rect 23358 1085 23450 1097
rect 24864 982 24899 1244
rect 16859 807 16893 930
rect 17331 917 17397 930
rect 17331 883 17347 917
rect 17381 883 17397 917
rect 17331 867 17397 883
rect 17720 807 17754 931
rect 19991 811 20025 934
rect 20463 921 20529 934
rect 20463 887 20479 921
rect 20513 887 20529 921
rect 20463 871 20529 887
rect 20852 811 20886 935
rect 22301 934 23673 981
rect 23995 935 24899 982
rect 23135 811 23169 934
rect 23607 921 23673 934
rect 23607 887 23623 921
rect 23657 887 23673 921
rect 23607 871 23673 887
rect 23996 811 24030 935
rect 11368 623 11374 799
rect 11408 623 11414 799
rect 11368 611 11414 623
rect 13710 795 13756 807
rect 13710 619 13716 795
rect 13750 619 13756 795
rect 11212 423 11218 611
rect 11172 411 11218 423
rect 10942 338 10976 411
rect 10927 322 10993 338
rect 10927 288 10943 322
rect 10977 288 10993 322
rect 10927 272 10993 288
rect 11256 244 11290 611
rect 13710 607 13756 619
rect 13828 795 13948 807
rect 13828 619 13834 795
rect 13868 619 13908 795
rect 13828 607 13908 619
rect 10632 192 11290 244
rect 13834 240 13868 607
rect 13902 419 13908 607
rect 13942 419 13948 795
rect 13902 407 13948 419
rect 14020 795 14066 807
rect 14020 419 14026 795
rect 14060 419 14066 795
rect 14020 407 14066 419
rect 14138 795 14184 807
rect 14138 419 14144 795
rect 14178 419 14184 795
rect 14138 407 14184 419
rect 14256 795 14302 807
rect 14256 419 14262 795
rect 14296 419 14302 795
rect 14256 407 14302 419
rect 14374 795 14498 807
rect 14374 419 14380 795
rect 14414 619 14458 795
rect 14492 619 14498 795
rect 14414 607 14498 619
rect 14570 795 14616 807
rect 14570 619 14576 795
rect 14610 619 14616 795
rect 14570 607 14616 619
rect 16854 795 16900 807
rect 16854 619 16860 795
rect 16894 619 16900 795
rect 16854 607 16900 619
rect 16972 795 17092 807
rect 16972 619 16978 795
rect 17012 619 17052 795
rect 16972 607 17052 619
rect 14414 419 14420 607
rect 14374 407 14420 419
rect 14144 334 14178 407
rect 14129 318 14195 334
rect 14129 284 14145 318
rect 14179 284 14195 318
rect 14129 268 14195 284
rect 14458 240 14492 607
rect 1510 166 1602 188
rect 1510 114 1522 166
rect 1588 114 1602 166
rect 1510 110 1602 114
rect 4654 166 4746 188
rect 4654 114 4666 166
rect 4732 114 4746 166
rect 7786 170 7878 192
rect 7786 118 7798 170
rect 7864 118 7878 170
rect 7786 114 7878 118
rect 10930 170 11022 192
rect 13834 188 14492 240
rect 16978 240 17012 607
rect 17046 419 17052 607
rect 17086 419 17092 795
rect 17046 407 17092 419
rect 17164 795 17210 807
rect 17164 419 17170 795
rect 17204 419 17210 795
rect 17164 407 17210 419
rect 17282 795 17328 807
rect 17282 419 17288 795
rect 17322 419 17328 795
rect 17282 407 17328 419
rect 17400 795 17446 807
rect 17400 419 17406 795
rect 17440 419 17446 795
rect 17400 407 17446 419
rect 17518 795 17642 807
rect 17518 419 17524 795
rect 17558 619 17602 795
rect 17636 619 17642 795
rect 17558 607 17642 619
rect 17714 795 17760 807
rect 17714 619 17720 795
rect 17754 619 17760 795
rect 17714 607 17760 619
rect 19986 799 20032 811
rect 19986 623 19992 799
rect 20026 623 20032 799
rect 19986 611 20032 623
rect 20104 799 20224 811
rect 20104 623 20110 799
rect 20144 623 20184 799
rect 20104 611 20184 623
rect 17558 419 17564 607
rect 17518 407 17564 419
rect 17288 334 17322 407
rect 17273 318 17339 334
rect 17273 284 17289 318
rect 17323 284 17339 318
rect 17273 268 17339 284
rect 17602 240 17636 607
rect 16978 188 17636 240
rect 20110 244 20144 611
rect 20178 423 20184 611
rect 20218 423 20224 799
rect 20178 411 20224 423
rect 20296 799 20342 811
rect 20296 423 20302 799
rect 20336 423 20342 799
rect 20296 411 20342 423
rect 20414 799 20460 811
rect 20414 423 20420 799
rect 20454 423 20460 799
rect 20414 411 20460 423
rect 20532 799 20578 811
rect 20532 423 20538 799
rect 20572 423 20578 799
rect 20532 411 20578 423
rect 20650 799 20774 811
rect 20650 423 20656 799
rect 20690 623 20734 799
rect 20768 623 20774 799
rect 20690 611 20774 623
rect 20846 799 20892 811
rect 20846 623 20852 799
rect 20886 623 20892 799
rect 20846 611 20892 623
rect 23130 799 23176 811
rect 23130 623 23136 799
rect 23170 623 23176 799
rect 23130 611 23176 623
rect 23248 799 23368 811
rect 23248 623 23254 799
rect 23288 623 23328 799
rect 23248 611 23328 623
rect 20690 423 20696 611
rect 20650 411 20696 423
rect 20420 338 20454 411
rect 20405 322 20471 338
rect 20405 288 20421 322
rect 20455 288 20471 322
rect 20405 272 20471 288
rect 20734 244 20768 611
rect 20110 192 20768 244
rect 23254 244 23288 611
rect 23322 423 23328 611
rect 23362 423 23368 799
rect 23322 411 23368 423
rect 23440 799 23486 811
rect 23440 423 23446 799
rect 23480 423 23486 799
rect 23440 411 23486 423
rect 23558 799 23604 811
rect 23558 423 23564 799
rect 23598 423 23604 799
rect 23558 411 23604 423
rect 23676 799 23722 811
rect 23676 423 23682 799
rect 23716 423 23722 799
rect 23676 411 23722 423
rect 23794 799 23918 811
rect 23794 423 23800 799
rect 23834 623 23878 799
rect 23912 623 23918 799
rect 23834 611 23918 623
rect 23990 799 24036 811
rect 23990 623 23996 799
rect 24030 623 24036 799
rect 23990 611 24036 623
rect 23834 423 23840 611
rect 23794 411 23840 423
rect 23564 338 23598 411
rect 23549 322 23615 338
rect 23549 288 23565 322
rect 23599 288 23615 322
rect 23549 272 23615 288
rect 23878 244 23912 611
rect 23254 192 23912 244
rect 10930 118 10942 170
rect 11008 118 11022 170
rect 10930 114 11022 118
rect 14132 166 14224 188
rect 14132 114 14144 166
rect 14210 114 14224 166
rect 4654 110 4746 114
rect 14132 110 14224 114
rect 17276 166 17368 188
rect 17276 114 17288 166
rect 17354 114 17368 166
rect 20408 170 20500 192
rect 20408 118 20420 170
rect 20486 118 20500 170
rect 20408 114 20500 118
rect 23552 170 23644 192
rect 23552 118 23564 170
rect 23630 118 23644 170
rect 23552 114 23644 118
rect 17276 110 17368 114
rect 1530 -1568 1540 -1508
rect 1620 -1568 1630 -1508
rect 1530 -1608 1630 -1568
rect 4674 -1568 4684 -1508
rect 4764 -1568 4774 -1508
rect 4674 -1608 4774 -1568
rect 7806 -1564 7816 -1504
rect 7896 -1564 7906 -1504
rect 7806 -1604 7906 -1564
rect 10950 -1564 10960 -1504
rect 11040 -1564 11050 -1504
rect 10950 -1604 11050 -1564
rect 14152 -1568 14162 -1508
rect 14242 -1568 14252 -1508
rect 733 -1665 2536 -1608
rect 733 -1752 767 -1665
rect 1908 -1752 1942 -1665
rect 727 -1764 773 -1752
rect 727 -1952 733 -1764
rect 286 -1964 332 -1952
rect 286 -2140 292 -1964
rect 326 -2140 332 -1964
rect 286 -2152 332 -2140
rect 404 -1964 450 -1952
rect 404 -2140 410 -1964
rect 444 -2140 450 -1964
rect 404 -2152 450 -2140
rect 522 -1964 568 -1952
rect 522 -2140 528 -1964
rect 562 -2140 568 -1964
rect 522 -2152 568 -2140
rect 640 -1964 733 -1952
rect 640 -2140 646 -1964
rect 680 -2140 733 -1964
rect 767 -2140 773 -1764
rect 640 -2152 773 -2140
rect 845 -1764 891 -1752
rect 845 -2140 851 -1764
rect 885 -2140 891 -1764
rect 845 -2152 891 -2140
rect 963 -1764 1009 -1752
rect 963 -2140 969 -1764
rect 1003 -2140 1009 -1764
rect 963 -2152 1009 -2140
rect 1081 -1764 1127 -1752
rect 1081 -2140 1087 -1764
rect 1121 -2140 1127 -1764
rect 1081 -2152 1127 -2140
rect 1194 -1764 1240 -1752
rect 1194 -2140 1200 -1764
rect 1234 -2140 1240 -1764
rect 1194 -2152 1240 -2140
rect 1312 -1764 1358 -1752
rect 1312 -2140 1318 -1764
rect 1352 -2140 1358 -1764
rect 1312 -2152 1358 -2140
rect 1430 -1764 1476 -1752
rect 1430 -2140 1436 -1764
rect 1470 -2140 1476 -1764
rect 1430 -2152 1476 -2140
rect 1548 -1764 1594 -1752
rect 1548 -2140 1554 -1764
rect 1588 -2140 1594 -1764
rect 1548 -2152 1594 -2140
rect 1666 -1764 1712 -1752
rect 1666 -2140 1672 -1764
rect 1706 -2140 1712 -1764
rect 1666 -2152 1712 -2140
rect 1784 -1764 1830 -1752
rect 1784 -2140 1790 -1764
rect 1824 -2140 1830 -1764
rect 1784 -2152 1830 -2140
rect 1902 -1764 1948 -1752
rect 1902 -2140 1908 -1764
rect 1942 -2140 1948 -1764
rect 1902 -2152 1948 -2140
rect 2021 -1764 2067 -1752
rect 2021 -2140 2027 -1764
rect 2061 -2140 2067 -1764
rect 2021 -2152 2067 -2140
rect 2139 -1764 2185 -1752
rect 2139 -2140 2145 -1764
rect 2179 -2140 2185 -1764
rect 2139 -2152 2185 -2140
rect 2257 -1764 2303 -1752
rect 2257 -2140 2263 -1764
rect 2297 -2140 2303 -1764
rect 2257 -2152 2303 -2140
rect 2375 -1764 2421 -1752
rect 2375 -2140 2381 -1764
rect 2415 -2140 2421 -1764
rect 2499 -1952 2536 -1665
rect 3877 -1665 5680 -1608
rect 3877 -1752 3911 -1665
rect 5052 -1752 5086 -1665
rect 3871 -1764 3917 -1752
rect 3871 -1952 3877 -1764
rect 2375 -2152 2421 -2140
rect 2494 -1964 2540 -1952
rect 2494 -2140 2500 -1964
rect 2534 -2140 2540 -1964
rect 2494 -2152 2540 -2140
rect 2612 -1964 2658 -1952
rect 2612 -2140 2618 -1964
rect 2652 -2140 2658 -1964
rect 2612 -2152 2658 -2140
rect 2730 -1964 2776 -1952
rect 2730 -2140 2736 -1964
rect 2770 -2140 2776 -1964
rect 2730 -2152 2776 -2140
rect 2848 -1964 2894 -1952
rect 2848 -2140 2854 -1964
rect 2888 -2140 2894 -1964
rect 2848 -2152 2894 -2140
rect 3430 -1964 3476 -1952
rect 3430 -2140 3436 -1964
rect 3470 -2140 3476 -1964
rect 3430 -2152 3476 -2140
rect 3548 -1964 3594 -1952
rect 3548 -2140 3554 -1964
rect 3588 -2140 3594 -1964
rect 3548 -2152 3594 -2140
rect 3666 -1964 3712 -1952
rect 3666 -2140 3672 -1964
rect 3706 -2140 3712 -1964
rect 3666 -2152 3712 -2140
rect 3784 -1964 3877 -1952
rect 3784 -2140 3790 -1964
rect 3824 -2140 3877 -1964
rect 3911 -2140 3917 -1764
rect 3784 -2152 3917 -2140
rect 3989 -1764 4035 -1752
rect 3989 -2140 3995 -1764
rect 4029 -2140 4035 -1764
rect 3989 -2152 4035 -2140
rect 4107 -1764 4153 -1752
rect 4107 -2140 4113 -1764
rect 4147 -2140 4153 -1764
rect 4107 -2152 4153 -2140
rect 4225 -1764 4271 -1752
rect 4225 -2140 4231 -1764
rect 4265 -2140 4271 -1764
rect 4225 -2152 4271 -2140
rect 4338 -1764 4384 -1752
rect 4338 -2140 4344 -1764
rect 4378 -2140 4384 -1764
rect 4338 -2152 4384 -2140
rect 4456 -1764 4502 -1752
rect 4456 -2140 4462 -1764
rect 4496 -2140 4502 -1764
rect 4456 -2152 4502 -2140
rect 4574 -1764 4620 -1752
rect 4574 -2140 4580 -1764
rect 4614 -2140 4620 -1764
rect 4574 -2152 4620 -2140
rect 4692 -1764 4738 -1752
rect 4692 -2140 4698 -1764
rect 4732 -2140 4738 -1764
rect 4692 -2152 4738 -2140
rect 4810 -1764 4856 -1752
rect 4810 -2140 4816 -1764
rect 4850 -2140 4856 -1764
rect 4810 -2152 4856 -2140
rect 4928 -1764 4974 -1752
rect 4928 -2140 4934 -1764
rect 4968 -2140 4974 -1764
rect 4928 -2152 4974 -2140
rect 5046 -1764 5092 -1752
rect 5046 -2140 5052 -1764
rect 5086 -2140 5092 -1764
rect 5046 -2152 5092 -2140
rect 5165 -1764 5211 -1752
rect 5165 -2140 5171 -1764
rect 5205 -2140 5211 -1764
rect 5165 -2152 5211 -2140
rect 5283 -1764 5329 -1752
rect 5283 -2140 5289 -1764
rect 5323 -2140 5329 -1764
rect 5283 -2152 5329 -2140
rect 5401 -1764 5447 -1752
rect 5401 -2140 5407 -1764
rect 5441 -2140 5447 -1764
rect 5401 -2152 5447 -2140
rect 5519 -1764 5565 -1752
rect 5519 -2140 5525 -1764
rect 5559 -2140 5565 -1764
rect 5643 -1952 5680 -1665
rect 7009 -1661 8812 -1604
rect 7009 -1748 7043 -1661
rect 8184 -1748 8218 -1661
rect 7003 -1760 7049 -1748
rect 7003 -1948 7009 -1760
rect 5519 -2152 5565 -2140
rect 5638 -1964 5684 -1952
rect 5638 -2140 5644 -1964
rect 5678 -2140 5684 -1964
rect 5638 -2152 5684 -2140
rect 5756 -1964 5802 -1952
rect 5756 -2140 5762 -1964
rect 5796 -2140 5802 -1964
rect 5756 -2152 5802 -2140
rect 5874 -1964 5920 -1952
rect 5874 -2140 5880 -1964
rect 5914 -2140 5920 -1964
rect 5874 -2152 5920 -2140
rect 5992 -1964 6038 -1952
rect 5992 -2140 5998 -1964
rect 6032 -2140 6038 -1964
rect 5992 -2152 6038 -2140
rect 6562 -1960 6608 -1948
rect 6562 -2136 6568 -1960
rect 6602 -2136 6608 -1960
rect 6562 -2148 6608 -2136
rect 6680 -1960 6726 -1948
rect 6680 -2136 6686 -1960
rect 6720 -2136 6726 -1960
rect 6680 -2148 6726 -2136
rect 6798 -1960 6844 -1948
rect 6798 -2136 6804 -1960
rect 6838 -2136 6844 -1960
rect 6798 -2148 6844 -2136
rect 6916 -1960 7009 -1948
rect 6916 -2136 6922 -1960
rect 6956 -2136 7009 -1960
rect 7043 -2136 7049 -1760
rect 6916 -2148 7049 -2136
rect 7121 -1760 7167 -1748
rect 7121 -2136 7127 -1760
rect 7161 -2136 7167 -1760
rect 7121 -2148 7167 -2136
rect 7239 -1760 7285 -1748
rect 7239 -2136 7245 -1760
rect 7279 -2136 7285 -1760
rect 7239 -2148 7285 -2136
rect 7357 -1760 7403 -1748
rect 7357 -2136 7363 -1760
rect 7397 -2136 7403 -1760
rect 7357 -2148 7403 -2136
rect 7470 -1760 7516 -1748
rect 7470 -2136 7476 -1760
rect 7510 -2136 7516 -1760
rect 7470 -2148 7516 -2136
rect 7588 -1760 7634 -1748
rect 7588 -2136 7594 -1760
rect 7628 -2136 7634 -1760
rect 7588 -2148 7634 -2136
rect 7706 -1760 7752 -1748
rect 7706 -2136 7712 -1760
rect 7746 -2136 7752 -1760
rect 7706 -2148 7752 -2136
rect 7824 -1760 7870 -1748
rect 7824 -2136 7830 -1760
rect 7864 -2136 7870 -1760
rect 7824 -2148 7870 -2136
rect 7942 -1760 7988 -1748
rect 7942 -2136 7948 -1760
rect 7982 -2136 7988 -1760
rect 7942 -2148 7988 -2136
rect 8060 -1760 8106 -1748
rect 8060 -2136 8066 -1760
rect 8100 -2136 8106 -1760
rect 8060 -2148 8106 -2136
rect 8178 -1760 8224 -1748
rect 8178 -2136 8184 -1760
rect 8218 -2136 8224 -1760
rect 8178 -2148 8224 -2136
rect 8297 -1760 8343 -1748
rect 8297 -2136 8303 -1760
rect 8337 -2136 8343 -1760
rect 8297 -2148 8343 -2136
rect 8415 -1760 8461 -1748
rect 8415 -2136 8421 -1760
rect 8455 -2136 8461 -1760
rect 8415 -2148 8461 -2136
rect 8533 -1760 8579 -1748
rect 8533 -2136 8539 -1760
rect 8573 -2136 8579 -1760
rect 8533 -2148 8579 -2136
rect 8651 -1760 8697 -1748
rect 8651 -2136 8657 -1760
rect 8691 -2136 8697 -1760
rect 8775 -1948 8812 -1661
rect 10153 -1661 11956 -1604
rect 14152 -1608 14252 -1568
rect 17296 -1568 17306 -1508
rect 17386 -1568 17396 -1508
rect 17296 -1608 17396 -1568
rect 20428 -1564 20438 -1504
rect 20518 -1564 20528 -1504
rect 20428 -1604 20528 -1564
rect 23572 -1564 23582 -1504
rect 23662 -1564 23672 -1504
rect 23572 -1604 23672 -1564
rect 10153 -1748 10187 -1661
rect 11328 -1748 11362 -1661
rect 10147 -1760 10193 -1748
rect 10147 -1948 10153 -1760
rect 8651 -2148 8697 -2136
rect 8770 -1960 8816 -1948
rect 8770 -2136 8776 -1960
rect 8810 -2136 8816 -1960
rect 8770 -2148 8816 -2136
rect 8888 -1960 8934 -1948
rect 8888 -2136 8894 -1960
rect 8928 -2136 8934 -1960
rect 8888 -2148 8934 -2136
rect 9006 -1960 9052 -1948
rect 9006 -2136 9012 -1960
rect 9046 -2136 9052 -1960
rect 9006 -2148 9052 -2136
rect 9124 -1960 9170 -1948
rect 9124 -2136 9130 -1960
rect 9164 -2136 9170 -1960
rect 9124 -2148 9170 -2136
rect 9706 -1960 9752 -1948
rect 9706 -2136 9712 -1960
rect 9746 -2136 9752 -1960
rect 9706 -2148 9752 -2136
rect 9824 -1960 9870 -1948
rect 9824 -2136 9830 -1960
rect 9864 -2136 9870 -1960
rect 9824 -2148 9870 -2136
rect 9942 -1960 9988 -1948
rect 9942 -2136 9948 -1960
rect 9982 -2136 9988 -1960
rect 9942 -2148 9988 -2136
rect 10060 -1960 10153 -1948
rect 10060 -2136 10066 -1960
rect 10100 -2136 10153 -1960
rect 10187 -2136 10193 -1760
rect 10060 -2148 10193 -2136
rect 10265 -1760 10311 -1748
rect 10265 -2136 10271 -1760
rect 10305 -2136 10311 -1760
rect 10265 -2148 10311 -2136
rect 10383 -1760 10429 -1748
rect 10383 -2136 10389 -1760
rect 10423 -2136 10429 -1760
rect 10383 -2148 10429 -2136
rect 10501 -1760 10547 -1748
rect 10501 -2136 10507 -1760
rect 10541 -2136 10547 -1760
rect 10501 -2148 10547 -2136
rect 10614 -1760 10660 -1748
rect 10614 -2136 10620 -1760
rect 10654 -2136 10660 -1760
rect 10614 -2148 10660 -2136
rect 10732 -1760 10778 -1748
rect 10732 -2136 10738 -1760
rect 10772 -2136 10778 -1760
rect 10732 -2148 10778 -2136
rect 10850 -1760 10896 -1748
rect 10850 -2136 10856 -1760
rect 10890 -2136 10896 -1760
rect 10850 -2148 10896 -2136
rect 10968 -1760 11014 -1748
rect 10968 -2136 10974 -1760
rect 11008 -2136 11014 -1760
rect 10968 -2148 11014 -2136
rect 11086 -1760 11132 -1748
rect 11086 -2136 11092 -1760
rect 11126 -2136 11132 -1760
rect 11086 -2148 11132 -2136
rect 11204 -1760 11250 -1748
rect 11204 -2136 11210 -1760
rect 11244 -2136 11250 -1760
rect 11204 -2148 11250 -2136
rect 11322 -1760 11368 -1748
rect 11322 -2136 11328 -1760
rect 11362 -2136 11368 -1760
rect 11322 -2148 11368 -2136
rect 11441 -1760 11487 -1748
rect 11441 -2136 11447 -1760
rect 11481 -2136 11487 -1760
rect 11441 -2148 11487 -2136
rect 11559 -1760 11605 -1748
rect 11559 -2136 11565 -1760
rect 11599 -2136 11605 -1760
rect 11559 -2148 11605 -2136
rect 11677 -1760 11723 -1748
rect 11677 -2136 11683 -1760
rect 11717 -2136 11723 -1760
rect 11677 -2148 11723 -2136
rect 11795 -1760 11841 -1748
rect 11795 -2136 11801 -1760
rect 11835 -2136 11841 -1760
rect 11919 -1948 11956 -1661
rect 13355 -1665 15158 -1608
rect 13355 -1752 13389 -1665
rect 14530 -1752 14564 -1665
rect 13349 -1764 13395 -1752
rect 11795 -2148 11841 -2136
rect 11914 -1960 11960 -1948
rect 11914 -2136 11920 -1960
rect 11954 -2136 11960 -1960
rect 11914 -2148 11960 -2136
rect 12032 -1960 12078 -1948
rect 12032 -2136 12038 -1960
rect 12072 -2136 12078 -1960
rect 12032 -2148 12078 -2136
rect 12150 -1960 12196 -1948
rect 12150 -2136 12156 -1960
rect 12190 -2136 12196 -1960
rect 12150 -2148 12196 -2136
rect 12268 -1960 12314 -1948
rect 13349 -1952 13355 -1764
rect 12268 -2136 12274 -1960
rect 12308 -2136 12314 -1960
rect 12268 -2148 12314 -2136
rect 12908 -1964 12954 -1952
rect 12908 -2140 12914 -1964
rect 12948 -2140 12954 -1964
rect 291 -2338 326 -2152
rect 1200 -2236 1234 -2152
rect 2381 -2236 2415 -2152
rect 1200 -2278 2415 -2236
rect 2381 -2298 2415 -2278
rect 2381 -2314 2738 -2298
rect 291 -2355 1428 -2338
rect 291 -2389 1378 -2355
rect 1412 -2389 1428 -2355
rect 2381 -2348 2688 -2314
rect 2722 -2348 2738 -2314
rect 2381 -2364 2738 -2348
rect 291 -2405 1428 -2389
rect 32 -2450 208 -2442
rect 32 -2518 149 -2450
rect 206 -2518 216 -2450
rect 32 -2526 208 -2518
rect 32 -2566 208 -2558
rect 32 -2634 149 -2566
rect 206 -2634 216 -2566
rect 32 -2642 208 -2634
rect 32 -2734 208 -2726
rect 32 -2802 149 -2734
rect 206 -2802 216 -2734
rect 32 -2810 208 -2802
rect 291 -2915 326 -2405
rect 381 -2451 473 -2438
rect 381 -2514 393 -2451
rect 464 -2514 473 -2451
rect 381 -2523 473 -2514
rect 1466 -2451 1558 -2441
rect 1466 -2513 1478 -2451
rect 1548 -2513 1558 -2451
rect 1466 -2526 1558 -2513
rect 2854 -2506 2889 -2152
rect 3435 -2338 3470 -2152
rect 4344 -2236 4378 -2152
rect 5525 -2236 5559 -2152
rect 4344 -2278 5559 -2236
rect 5525 -2298 5559 -2278
rect 5525 -2314 5882 -2298
rect 3435 -2355 4572 -2338
rect 3435 -2389 4522 -2355
rect 4556 -2389 4572 -2355
rect 5525 -2348 5832 -2314
rect 5866 -2348 5882 -2314
rect 5525 -2364 5882 -2348
rect 3435 -2405 4572 -2389
rect 3176 -2450 3352 -2442
rect 1713 -2568 1778 -2565
rect 1713 -2571 1782 -2568
rect 1713 -2631 1719 -2571
rect 1778 -2631 1788 -2571
rect 1713 -2635 1782 -2631
rect 1713 -2637 1778 -2635
rect 2854 -2652 3035 -2506
rect 3176 -2518 3293 -2450
rect 3350 -2518 3360 -2450
rect 3176 -2526 3352 -2518
rect 3176 -2566 3352 -2558
rect 3176 -2634 3293 -2566
rect 3350 -2634 3360 -2566
rect 3176 -2642 3352 -2634
rect 1348 -2734 1440 -2726
rect 1348 -2799 1360 -2734
rect 1428 -2799 1440 -2734
rect 1348 -2811 1440 -2799
rect 2854 -2914 2889 -2652
rect 3176 -2734 3352 -2726
rect 3176 -2802 3293 -2734
rect 3350 -2802 3360 -2734
rect 3176 -2810 3352 -2802
rect 291 -2962 1663 -2915
rect 1985 -2961 2889 -2914
rect 3435 -2915 3470 -2405
rect 3525 -2451 3617 -2438
rect 3525 -2514 3537 -2451
rect 3608 -2514 3617 -2451
rect 3525 -2523 3617 -2514
rect 4610 -2451 4702 -2441
rect 4610 -2513 4622 -2451
rect 4692 -2513 4702 -2451
rect 4610 -2526 4702 -2513
rect 5998 -2506 6033 -2152
rect 6567 -2334 6602 -2148
rect 7476 -2232 7510 -2148
rect 8657 -2232 8691 -2148
rect 7476 -2274 8691 -2232
rect 8657 -2294 8691 -2274
rect 8657 -2310 9014 -2294
rect 6567 -2351 7704 -2334
rect 6567 -2385 7654 -2351
rect 7688 -2385 7704 -2351
rect 8657 -2344 8964 -2310
rect 8998 -2344 9014 -2310
rect 8657 -2360 9014 -2344
rect 6567 -2401 7704 -2385
rect 6308 -2446 6484 -2438
rect 4857 -2568 4922 -2565
rect 4857 -2571 4926 -2568
rect 4857 -2631 4863 -2571
rect 4922 -2631 4932 -2571
rect 4857 -2635 4926 -2631
rect 4857 -2637 4922 -2635
rect 5998 -2652 6179 -2506
rect 6308 -2514 6425 -2446
rect 6482 -2514 6492 -2446
rect 6308 -2522 6484 -2514
rect 6308 -2562 6484 -2554
rect 6308 -2630 6425 -2562
rect 6482 -2630 6492 -2562
rect 6308 -2638 6484 -2630
rect 4492 -2734 4584 -2726
rect 4492 -2799 4504 -2734
rect 4572 -2799 4584 -2734
rect 4492 -2811 4584 -2799
rect 5998 -2914 6033 -2652
rect 6308 -2730 6484 -2722
rect 6308 -2798 6425 -2730
rect 6482 -2798 6492 -2730
rect 6308 -2806 6484 -2798
rect 1125 -3085 1159 -2962
rect 1597 -2975 1663 -2962
rect 1597 -3009 1613 -2975
rect 1647 -3009 1663 -2975
rect 1597 -3025 1663 -3009
rect 1986 -3085 2020 -2961
rect 3435 -2962 4807 -2915
rect 5129 -2961 6033 -2914
rect 6567 -2911 6602 -2401
rect 6657 -2447 6749 -2434
rect 6657 -2510 6669 -2447
rect 6740 -2510 6749 -2447
rect 6657 -2519 6749 -2510
rect 7742 -2447 7834 -2437
rect 7742 -2509 7754 -2447
rect 7824 -2509 7834 -2447
rect 7742 -2522 7834 -2509
rect 9130 -2502 9165 -2148
rect 9711 -2334 9746 -2148
rect 10620 -2232 10654 -2148
rect 11801 -2232 11835 -2148
rect 10620 -2274 11835 -2232
rect 11801 -2294 11835 -2274
rect 11801 -2310 12158 -2294
rect 9711 -2351 10848 -2334
rect 9711 -2385 10798 -2351
rect 10832 -2385 10848 -2351
rect 11801 -2344 12108 -2310
rect 12142 -2344 12158 -2310
rect 11801 -2360 12158 -2344
rect 9711 -2401 10848 -2385
rect 9452 -2446 9628 -2438
rect 7989 -2564 8054 -2561
rect 7989 -2567 8058 -2564
rect 7989 -2627 7995 -2567
rect 8054 -2627 8064 -2567
rect 7989 -2631 8058 -2627
rect 7989 -2633 8054 -2631
rect 9130 -2648 9311 -2502
rect 9452 -2514 9569 -2446
rect 9626 -2514 9636 -2446
rect 9452 -2522 9628 -2514
rect 9452 -2562 9628 -2554
rect 9452 -2630 9569 -2562
rect 9626 -2630 9636 -2562
rect 9452 -2638 9628 -2630
rect 7624 -2730 7716 -2722
rect 7624 -2795 7636 -2730
rect 7704 -2795 7716 -2730
rect 7624 -2807 7716 -2795
rect 9130 -2910 9165 -2648
rect 9452 -2730 9628 -2722
rect 9452 -2798 9569 -2730
rect 9626 -2798 9636 -2730
rect 9452 -2806 9628 -2798
rect 6567 -2958 7939 -2911
rect 8261 -2957 9165 -2910
rect 9711 -2911 9746 -2401
rect 9801 -2447 9893 -2434
rect 9801 -2510 9813 -2447
rect 9884 -2510 9893 -2447
rect 9801 -2519 9893 -2510
rect 10886 -2447 10978 -2437
rect 10886 -2509 10898 -2447
rect 10968 -2509 10978 -2447
rect 10886 -2522 10978 -2509
rect 12274 -2502 12309 -2148
rect 12908 -2152 12954 -2140
rect 13026 -1964 13072 -1952
rect 13026 -2140 13032 -1964
rect 13066 -2140 13072 -1964
rect 13026 -2152 13072 -2140
rect 13144 -1964 13190 -1952
rect 13144 -2140 13150 -1964
rect 13184 -2140 13190 -1964
rect 13144 -2152 13190 -2140
rect 13262 -1964 13355 -1952
rect 13262 -2140 13268 -1964
rect 13302 -2140 13355 -1964
rect 13389 -2140 13395 -1764
rect 13262 -2152 13395 -2140
rect 13467 -1764 13513 -1752
rect 13467 -2140 13473 -1764
rect 13507 -2140 13513 -1764
rect 13467 -2152 13513 -2140
rect 13585 -1764 13631 -1752
rect 13585 -2140 13591 -1764
rect 13625 -2140 13631 -1764
rect 13585 -2152 13631 -2140
rect 13703 -1764 13749 -1752
rect 13703 -2140 13709 -1764
rect 13743 -2140 13749 -1764
rect 13703 -2152 13749 -2140
rect 13816 -1764 13862 -1752
rect 13816 -2140 13822 -1764
rect 13856 -2140 13862 -1764
rect 13816 -2152 13862 -2140
rect 13934 -1764 13980 -1752
rect 13934 -2140 13940 -1764
rect 13974 -2140 13980 -1764
rect 13934 -2152 13980 -2140
rect 14052 -1764 14098 -1752
rect 14052 -2140 14058 -1764
rect 14092 -2140 14098 -1764
rect 14052 -2152 14098 -2140
rect 14170 -1764 14216 -1752
rect 14170 -2140 14176 -1764
rect 14210 -2140 14216 -1764
rect 14170 -2152 14216 -2140
rect 14288 -1764 14334 -1752
rect 14288 -2140 14294 -1764
rect 14328 -2140 14334 -1764
rect 14288 -2152 14334 -2140
rect 14406 -1764 14452 -1752
rect 14406 -2140 14412 -1764
rect 14446 -2140 14452 -1764
rect 14406 -2152 14452 -2140
rect 14524 -1764 14570 -1752
rect 14524 -2140 14530 -1764
rect 14564 -2140 14570 -1764
rect 14524 -2152 14570 -2140
rect 14643 -1764 14689 -1752
rect 14643 -2140 14649 -1764
rect 14683 -2140 14689 -1764
rect 14643 -2152 14689 -2140
rect 14761 -1764 14807 -1752
rect 14761 -2140 14767 -1764
rect 14801 -2140 14807 -1764
rect 14761 -2152 14807 -2140
rect 14879 -1764 14925 -1752
rect 14879 -2140 14885 -1764
rect 14919 -2140 14925 -1764
rect 14879 -2152 14925 -2140
rect 14997 -1764 15043 -1752
rect 14997 -2140 15003 -1764
rect 15037 -2140 15043 -1764
rect 15121 -1952 15158 -1665
rect 16499 -1665 18302 -1608
rect 16499 -1752 16533 -1665
rect 17674 -1752 17708 -1665
rect 16493 -1764 16539 -1752
rect 16493 -1952 16499 -1764
rect 14997 -2152 15043 -2140
rect 15116 -1964 15162 -1952
rect 15116 -2140 15122 -1964
rect 15156 -2140 15162 -1964
rect 15116 -2152 15162 -2140
rect 15234 -1964 15280 -1952
rect 15234 -2140 15240 -1964
rect 15274 -2140 15280 -1964
rect 15234 -2152 15280 -2140
rect 15352 -1964 15398 -1952
rect 15352 -2140 15358 -1964
rect 15392 -2140 15398 -1964
rect 15352 -2152 15398 -2140
rect 15470 -1964 15516 -1952
rect 15470 -2140 15476 -1964
rect 15510 -2140 15516 -1964
rect 15470 -2152 15516 -2140
rect 16052 -1964 16098 -1952
rect 16052 -2140 16058 -1964
rect 16092 -2140 16098 -1964
rect 16052 -2152 16098 -2140
rect 16170 -1964 16216 -1952
rect 16170 -2140 16176 -1964
rect 16210 -2140 16216 -1964
rect 16170 -2152 16216 -2140
rect 16288 -1964 16334 -1952
rect 16288 -2140 16294 -1964
rect 16328 -2140 16334 -1964
rect 16288 -2152 16334 -2140
rect 16406 -1964 16499 -1952
rect 16406 -2140 16412 -1964
rect 16446 -2140 16499 -1964
rect 16533 -2140 16539 -1764
rect 16406 -2152 16539 -2140
rect 16611 -1764 16657 -1752
rect 16611 -2140 16617 -1764
rect 16651 -2140 16657 -1764
rect 16611 -2152 16657 -2140
rect 16729 -1764 16775 -1752
rect 16729 -2140 16735 -1764
rect 16769 -2140 16775 -1764
rect 16729 -2152 16775 -2140
rect 16847 -1764 16893 -1752
rect 16847 -2140 16853 -1764
rect 16887 -2140 16893 -1764
rect 16847 -2152 16893 -2140
rect 16960 -1764 17006 -1752
rect 16960 -2140 16966 -1764
rect 17000 -2140 17006 -1764
rect 16960 -2152 17006 -2140
rect 17078 -1764 17124 -1752
rect 17078 -2140 17084 -1764
rect 17118 -2140 17124 -1764
rect 17078 -2152 17124 -2140
rect 17196 -1764 17242 -1752
rect 17196 -2140 17202 -1764
rect 17236 -2140 17242 -1764
rect 17196 -2152 17242 -2140
rect 17314 -1764 17360 -1752
rect 17314 -2140 17320 -1764
rect 17354 -2140 17360 -1764
rect 17314 -2152 17360 -2140
rect 17432 -1764 17478 -1752
rect 17432 -2140 17438 -1764
rect 17472 -2140 17478 -1764
rect 17432 -2152 17478 -2140
rect 17550 -1764 17596 -1752
rect 17550 -2140 17556 -1764
rect 17590 -2140 17596 -1764
rect 17550 -2152 17596 -2140
rect 17668 -1764 17714 -1752
rect 17668 -2140 17674 -1764
rect 17708 -2140 17714 -1764
rect 17668 -2152 17714 -2140
rect 17787 -1764 17833 -1752
rect 17787 -2140 17793 -1764
rect 17827 -2140 17833 -1764
rect 17787 -2152 17833 -2140
rect 17905 -1764 17951 -1752
rect 17905 -2140 17911 -1764
rect 17945 -2140 17951 -1764
rect 17905 -2152 17951 -2140
rect 18023 -1764 18069 -1752
rect 18023 -2140 18029 -1764
rect 18063 -2140 18069 -1764
rect 18023 -2152 18069 -2140
rect 18141 -1764 18187 -1752
rect 18141 -2140 18147 -1764
rect 18181 -2140 18187 -1764
rect 18265 -1952 18302 -1665
rect 19631 -1661 21434 -1604
rect 19631 -1748 19665 -1661
rect 20806 -1748 20840 -1661
rect 19625 -1760 19671 -1748
rect 19625 -1948 19631 -1760
rect 18141 -2152 18187 -2140
rect 18260 -1964 18306 -1952
rect 18260 -2140 18266 -1964
rect 18300 -2140 18306 -1964
rect 18260 -2152 18306 -2140
rect 18378 -1964 18424 -1952
rect 18378 -2140 18384 -1964
rect 18418 -2140 18424 -1964
rect 18378 -2152 18424 -2140
rect 18496 -1964 18542 -1952
rect 18496 -2140 18502 -1964
rect 18536 -2140 18542 -1964
rect 18496 -2152 18542 -2140
rect 18614 -1964 18660 -1952
rect 18614 -2140 18620 -1964
rect 18654 -2140 18660 -1964
rect 18614 -2152 18660 -2140
rect 19184 -1960 19230 -1948
rect 19184 -2136 19190 -1960
rect 19224 -2136 19230 -1960
rect 19184 -2148 19230 -2136
rect 19302 -1960 19348 -1948
rect 19302 -2136 19308 -1960
rect 19342 -2136 19348 -1960
rect 19302 -2148 19348 -2136
rect 19420 -1960 19466 -1948
rect 19420 -2136 19426 -1960
rect 19460 -2136 19466 -1960
rect 19420 -2148 19466 -2136
rect 19538 -1960 19631 -1948
rect 19538 -2136 19544 -1960
rect 19578 -2136 19631 -1960
rect 19665 -2136 19671 -1760
rect 19538 -2148 19671 -2136
rect 19743 -1760 19789 -1748
rect 19743 -2136 19749 -1760
rect 19783 -2136 19789 -1760
rect 19743 -2148 19789 -2136
rect 19861 -1760 19907 -1748
rect 19861 -2136 19867 -1760
rect 19901 -2136 19907 -1760
rect 19861 -2148 19907 -2136
rect 19979 -1760 20025 -1748
rect 19979 -2136 19985 -1760
rect 20019 -2136 20025 -1760
rect 19979 -2148 20025 -2136
rect 20092 -1760 20138 -1748
rect 20092 -2136 20098 -1760
rect 20132 -2136 20138 -1760
rect 20092 -2148 20138 -2136
rect 20210 -1760 20256 -1748
rect 20210 -2136 20216 -1760
rect 20250 -2136 20256 -1760
rect 20210 -2148 20256 -2136
rect 20328 -1760 20374 -1748
rect 20328 -2136 20334 -1760
rect 20368 -2136 20374 -1760
rect 20328 -2148 20374 -2136
rect 20446 -1760 20492 -1748
rect 20446 -2136 20452 -1760
rect 20486 -2136 20492 -1760
rect 20446 -2148 20492 -2136
rect 20564 -1760 20610 -1748
rect 20564 -2136 20570 -1760
rect 20604 -2136 20610 -1760
rect 20564 -2148 20610 -2136
rect 20682 -1760 20728 -1748
rect 20682 -2136 20688 -1760
rect 20722 -2136 20728 -1760
rect 20682 -2148 20728 -2136
rect 20800 -1760 20846 -1748
rect 20800 -2136 20806 -1760
rect 20840 -2136 20846 -1760
rect 20800 -2148 20846 -2136
rect 20919 -1760 20965 -1748
rect 20919 -2136 20925 -1760
rect 20959 -2136 20965 -1760
rect 20919 -2148 20965 -2136
rect 21037 -1760 21083 -1748
rect 21037 -2136 21043 -1760
rect 21077 -2136 21083 -1760
rect 21037 -2148 21083 -2136
rect 21155 -1760 21201 -1748
rect 21155 -2136 21161 -1760
rect 21195 -2136 21201 -1760
rect 21155 -2148 21201 -2136
rect 21273 -1760 21319 -1748
rect 21273 -2136 21279 -1760
rect 21313 -2136 21319 -1760
rect 21397 -1948 21434 -1661
rect 22775 -1661 24578 -1604
rect 22775 -1748 22809 -1661
rect 23950 -1748 23984 -1661
rect 22769 -1760 22815 -1748
rect 22769 -1948 22775 -1760
rect 21273 -2148 21319 -2136
rect 21392 -1960 21438 -1948
rect 21392 -2136 21398 -1960
rect 21432 -2136 21438 -1960
rect 21392 -2148 21438 -2136
rect 21510 -1960 21556 -1948
rect 21510 -2136 21516 -1960
rect 21550 -2136 21556 -1960
rect 21510 -2148 21556 -2136
rect 21628 -1960 21674 -1948
rect 21628 -2136 21634 -1960
rect 21668 -2136 21674 -1960
rect 21628 -2148 21674 -2136
rect 21746 -1960 21792 -1948
rect 21746 -2136 21752 -1960
rect 21786 -2136 21792 -1960
rect 21746 -2148 21792 -2136
rect 22328 -1960 22374 -1948
rect 22328 -2136 22334 -1960
rect 22368 -2136 22374 -1960
rect 22328 -2148 22374 -2136
rect 22446 -1960 22492 -1948
rect 22446 -2136 22452 -1960
rect 22486 -2136 22492 -1960
rect 22446 -2148 22492 -2136
rect 22564 -1960 22610 -1948
rect 22564 -2136 22570 -1960
rect 22604 -2136 22610 -1960
rect 22564 -2148 22610 -2136
rect 22682 -1960 22775 -1948
rect 22682 -2136 22688 -1960
rect 22722 -2136 22775 -1960
rect 22809 -2136 22815 -1760
rect 22682 -2148 22815 -2136
rect 22887 -1760 22933 -1748
rect 22887 -2136 22893 -1760
rect 22927 -2136 22933 -1760
rect 22887 -2148 22933 -2136
rect 23005 -1760 23051 -1748
rect 23005 -2136 23011 -1760
rect 23045 -2136 23051 -1760
rect 23005 -2148 23051 -2136
rect 23123 -1760 23169 -1748
rect 23123 -2136 23129 -1760
rect 23163 -2136 23169 -1760
rect 23123 -2148 23169 -2136
rect 23236 -1760 23282 -1748
rect 23236 -2136 23242 -1760
rect 23276 -2136 23282 -1760
rect 23236 -2148 23282 -2136
rect 23354 -1760 23400 -1748
rect 23354 -2136 23360 -1760
rect 23394 -2136 23400 -1760
rect 23354 -2148 23400 -2136
rect 23472 -1760 23518 -1748
rect 23472 -2136 23478 -1760
rect 23512 -2136 23518 -1760
rect 23472 -2148 23518 -2136
rect 23590 -1760 23636 -1748
rect 23590 -2136 23596 -1760
rect 23630 -2136 23636 -1760
rect 23590 -2148 23636 -2136
rect 23708 -1760 23754 -1748
rect 23708 -2136 23714 -1760
rect 23748 -2136 23754 -1760
rect 23708 -2148 23754 -2136
rect 23826 -1760 23872 -1748
rect 23826 -2136 23832 -1760
rect 23866 -2136 23872 -1760
rect 23826 -2148 23872 -2136
rect 23944 -1760 23990 -1748
rect 23944 -2136 23950 -1760
rect 23984 -2136 23990 -1760
rect 23944 -2148 23990 -2136
rect 24063 -1760 24109 -1748
rect 24063 -2136 24069 -1760
rect 24103 -2136 24109 -1760
rect 24063 -2148 24109 -2136
rect 24181 -1760 24227 -1748
rect 24181 -2136 24187 -1760
rect 24221 -2136 24227 -1760
rect 24181 -2148 24227 -2136
rect 24299 -1760 24345 -1748
rect 24299 -2136 24305 -1760
rect 24339 -2136 24345 -1760
rect 24299 -2148 24345 -2136
rect 24417 -1760 24463 -1748
rect 24417 -2136 24423 -1760
rect 24457 -2136 24463 -1760
rect 24541 -1948 24578 -1661
rect 24417 -2148 24463 -2136
rect 24536 -1960 24582 -1948
rect 24536 -2136 24542 -1960
rect 24576 -2136 24582 -1960
rect 24536 -2148 24582 -2136
rect 24654 -1960 24700 -1948
rect 24654 -2136 24660 -1960
rect 24694 -2136 24700 -1960
rect 24654 -2148 24700 -2136
rect 24772 -1960 24818 -1948
rect 24772 -2136 24778 -1960
rect 24812 -2136 24818 -1960
rect 24772 -2148 24818 -2136
rect 24890 -1960 24936 -1948
rect 24890 -2136 24896 -1960
rect 24930 -2136 24936 -1960
rect 24890 -2148 24936 -2136
rect 12913 -2338 12948 -2152
rect 13822 -2236 13856 -2152
rect 15003 -2236 15037 -2152
rect 13822 -2278 15037 -2236
rect 15003 -2298 15037 -2278
rect 15003 -2314 15360 -2298
rect 12913 -2355 14050 -2338
rect 12913 -2389 14000 -2355
rect 14034 -2389 14050 -2355
rect 15003 -2348 15310 -2314
rect 15344 -2348 15360 -2314
rect 15003 -2364 15360 -2348
rect 12913 -2405 14050 -2389
rect 12654 -2450 12830 -2442
rect 11133 -2564 11198 -2561
rect 11133 -2567 11202 -2564
rect 11133 -2627 11139 -2567
rect 11198 -2627 11208 -2567
rect 11133 -2631 11202 -2627
rect 11133 -2633 11198 -2631
rect 12274 -2648 12455 -2502
rect 12654 -2518 12771 -2450
rect 12828 -2518 12838 -2450
rect 12654 -2526 12830 -2518
rect 12654 -2566 12830 -2558
rect 12654 -2634 12771 -2566
rect 12828 -2634 12838 -2566
rect 12654 -2642 12830 -2634
rect 10768 -2730 10860 -2722
rect 10768 -2795 10780 -2730
rect 10848 -2795 10860 -2730
rect 10768 -2807 10860 -2795
rect 12274 -2910 12309 -2648
rect 12654 -2734 12830 -2726
rect 12654 -2802 12771 -2734
rect 12828 -2802 12838 -2734
rect 12654 -2810 12830 -2802
rect 4269 -3085 4303 -2962
rect 4741 -2975 4807 -2962
rect 4741 -3009 4757 -2975
rect 4791 -3009 4807 -2975
rect 4741 -3025 4807 -3009
rect 5130 -3085 5164 -2961
rect 7401 -3081 7435 -2958
rect 7873 -2971 7939 -2958
rect 7873 -3005 7889 -2971
rect 7923 -3005 7939 -2971
rect 7873 -3021 7939 -3005
rect 8262 -3081 8296 -2957
rect 9711 -2958 11083 -2911
rect 11405 -2957 12309 -2910
rect 12913 -2915 12948 -2405
rect 13003 -2451 13095 -2438
rect 13003 -2514 13015 -2451
rect 13086 -2514 13095 -2451
rect 13003 -2523 13095 -2514
rect 14088 -2451 14180 -2441
rect 14088 -2513 14100 -2451
rect 14170 -2513 14180 -2451
rect 14088 -2526 14180 -2513
rect 15476 -2506 15511 -2152
rect 16057 -2338 16092 -2152
rect 16966 -2236 17000 -2152
rect 18147 -2236 18181 -2152
rect 16966 -2278 18181 -2236
rect 18147 -2298 18181 -2278
rect 18147 -2314 18504 -2298
rect 16057 -2355 17194 -2338
rect 16057 -2389 17144 -2355
rect 17178 -2389 17194 -2355
rect 18147 -2348 18454 -2314
rect 18488 -2348 18504 -2314
rect 18147 -2364 18504 -2348
rect 16057 -2405 17194 -2389
rect 15798 -2450 15974 -2442
rect 14335 -2568 14400 -2565
rect 14335 -2571 14404 -2568
rect 14335 -2631 14341 -2571
rect 14400 -2631 14410 -2571
rect 14335 -2635 14404 -2631
rect 14335 -2637 14400 -2635
rect 15476 -2652 15657 -2506
rect 15798 -2518 15915 -2450
rect 15972 -2518 15982 -2450
rect 15798 -2526 15974 -2518
rect 15798 -2566 15974 -2558
rect 15798 -2634 15915 -2566
rect 15972 -2634 15982 -2566
rect 15798 -2642 15974 -2634
rect 13970 -2734 14062 -2726
rect 13970 -2799 13982 -2734
rect 14050 -2799 14062 -2734
rect 13970 -2811 14062 -2799
rect 15476 -2914 15511 -2652
rect 15798 -2734 15974 -2726
rect 15798 -2802 15915 -2734
rect 15972 -2802 15982 -2734
rect 15798 -2810 15974 -2802
rect 10545 -3081 10579 -2958
rect 11017 -2971 11083 -2958
rect 11017 -3005 11033 -2971
rect 11067 -3005 11083 -2971
rect 11017 -3021 11083 -3005
rect 11406 -3081 11440 -2957
rect 12913 -2962 14285 -2915
rect 14607 -2961 15511 -2914
rect 16057 -2915 16092 -2405
rect 16147 -2451 16239 -2438
rect 16147 -2514 16159 -2451
rect 16230 -2514 16239 -2451
rect 16147 -2523 16239 -2514
rect 17232 -2451 17324 -2441
rect 17232 -2513 17244 -2451
rect 17314 -2513 17324 -2451
rect 17232 -2526 17324 -2513
rect 18620 -2506 18655 -2152
rect 19189 -2334 19224 -2148
rect 20098 -2232 20132 -2148
rect 21279 -2232 21313 -2148
rect 20098 -2274 21313 -2232
rect 21279 -2294 21313 -2274
rect 21279 -2310 21636 -2294
rect 19189 -2351 20326 -2334
rect 19189 -2385 20276 -2351
rect 20310 -2385 20326 -2351
rect 21279 -2344 21586 -2310
rect 21620 -2344 21636 -2310
rect 21279 -2360 21636 -2344
rect 19189 -2401 20326 -2385
rect 18930 -2446 19106 -2438
rect 17479 -2568 17544 -2565
rect 17479 -2571 17548 -2568
rect 17479 -2631 17485 -2571
rect 17544 -2631 17554 -2571
rect 17479 -2635 17548 -2631
rect 17479 -2637 17544 -2635
rect 18620 -2652 18801 -2506
rect 18930 -2514 19047 -2446
rect 19104 -2514 19114 -2446
rect 18930 -2522 19106 -2514
rect 18930 -2562 19106 -2554
rect 18930 -2630 19047 -2562
rect 19104 -2630 19114 -2562
rect 18930 -2638 19106 -2630
rect 17114 -2734 17206 -2726
rect 17114 -2799 17126 -2734
rect 17194 -2799 17206 -2734
rect 17114 -2811 17206 -2799
rect 18620 -2914 18655 -2652
rect 18930 -2730 19106 -2722
rect 18930 -2798 19047 -2730
rect 19104 -2798 19114 -2730
rect 18930 -2806 19106 -2798
rect 1120 -3097 1166 -3085
rect 1120 -3273 1126 -3097
rect 1160 -3273 1166 -3097
rect 1120 -3285 1166 -3273
rect 1238 -3097 1358 -3085
rect 1238 -3273 1244 -3097
rect 1278 -3273 1318 -3097
rect 1238 -3285 1318 -3273
rect 1244 -3652 1278 -3285
rect 1312 -3473 1318 -3285
rect 1352 -3473 1358 -3097
rect 1312 -3485 1358 -3473
rect 1430 -3097 1476 -3085
rect 1430 -3473 1436 -3097
rect 1470 -3473 1476 -3097
rect 1430 -3485 1476 -3473
rect 1548 -3097 1594 -3085
rect 1548 -3473 1554 -3097
rect 1588 -3473 1594 -3097
rect 1548 -3485 1594 -3473
rect 1666 -3097 1712 -3085
rect 1666 -3473 1672 -3097
rect 1706 -3473 1712 -3097
rect 1666 -3485 1712 -3473
rect 1784 -3097 1908 -3085
rect 1784 -3473 1790 -3097
rect 1824 -3273 1868 -3097
rect 1902 -3273 1908 -3097
rect 1824 -3285 1908 -3273
rect 1980 -3097 2026 -3085
rect 1980 -3273 1986 -3097
rect 2020 -3273 2026 -3097
rect 1980 -3285 2026 -3273
rect 4264 -3097 4310 -3085
rect 4264 -3273 4270 -3097
rect 4304 -3273 4310 -3097
rect 4264 -3285 4310 -3273
rect 4382 -3097 4502 -3085
rect 4382 -3273 4388 -3097
rect 4422 -3273 4462 -3097
rect 4382 -3285 4462 -3273
rect 1824 -3473 1830 -3285
rect 1784 -3485 1830 -3473
rect 1554 -3558 1588 -3485
rect 1539 -3574 1605 -3558
rect 1539 -3608 1555 -3574
rect 1589 -3608 1605 -3574
rect 1539 -3624 1605 -3608
rect 1868 -3652 1902 -3285
rect 1244 -3704 1902 -3652
rect 4388 -3652 4422 -3285
rect 4456 -3473 4462 -3285
rect 4496 -3473 4502 -3097
rect 4456 -3485 4502 -3473
rect 4574 -3097 4620 -3085
rect 4574 -3473 4580 -3097
rect 4614 -3473 4620 -3097
rect 4574 -3485 4620 -3473
rect 4692 -3097 4738 -3085
rect 4692 -3473 4698 -3097
rect 4732 -3473 4738 -3097
rect 4692 -3485 4738 -3473
rect 4810 -3097 4856 -3085
rect 4810 -3473 4816 -3097
rect 4850 -3473 4856 -3097
rect 4810 -3485 4856 -3473
rect 4928 -3097 5052 -3085
rect 4928 -3473 4934 -3097
rect 4968 -3273 5012 -3097
rect 5046 -3273 5052 -3097
rect 4968 -3285 5052 -3273
rect 5124 -3097 5170 -3085
rect 5124 -3273 5130 -3097
rect 5164 -3273 5170 -3097
rect 5124 -3285 5170 -3273
rect 7396 -3093 7442 -3081
rect 7396 -3269 7402 -3093
rect 7436 -3269 7442 -3093
rect 7396 -3281 7442 -3269
rect 7514 -3093 7634 -3081
rect 7514 -3269 7520 -3093
rect 7554 -3269 7594 -3093
rect 7514 -3281 7594 -3269
rect 4968 -3473 4974 -3285
rect 4928 -3485 4974 -3473
rect 4698 -3558 4732 -3485
rect 4683 -3574 4749 -3558
rect 4683 -3608 4699 -3574
rect 4733 -3608 4749 -3574
rect 4683 -3624 4749 -3608
rect 5012 -3652 5046 -3285
rect 4388 -3704 5046 -3652
rect 7520 -3648 7554 -3281
rect 7588 -3469 7594 -3281
rect 7628 -3469 7634 -3093
rect 7588 -3481 7634 -3469
rect 7706 -3093 7752 -3081
rect 7706 -3469 7712 -3093
rect 7746 -3469 7752 -3093
rect 7706 -3481 7752 -3469
rect 7824 -3093 7870 -3081
rect 7824 -3469 7830 -3093
rect 7864 -3469 7870 -3093
rect 7824 -3481 7870 -3469
rect 7942 -3093 7988 -3081
rect 7942 -3469 7948 -3093
rect 7982 -3469 7988 -3093
rect 7942 -3481 7988 -3469
rect 8060 -3093 8184 -3081
rect 8060 -3469 8066 -3093
rect 8100 -3269 8144 -3093
rect 8178 -3269 8184 -3093
rect 8100 -3281 8184 -3269
rect 8256 -3093 8302 -3081
rect 8256 -3269 8262 -3093
rect 8296 -3269 8302 -3093
rect 8256 -3281 8302 -3269
rect 10540 -3093 10586 -3081
rect 10540 -3269 10546 -3093
rect 10580 -3269 10586 -3093
rect 10540 -3281 10586 -3269
rect 10658 -3093 10778 -3081
rect 10658 -3269 10664 -3093
rect 10698 -3269 10738 -3093
rect 10658 -3281 10738 -3269
rect 8100 -3469 8106 -3281
rect 8060 -3481 8106 -3469
rect 7830 -3554 7864 -3481
rect 7815 -3570 7881 -3554
rect 7815 -3604 7831 -3570
rect 7865 -3604 7881 -3570
rect 7815 -3620 7881 -3604
rect 8144 -3648 8178 -3281
rect 7520 -3700 8178 -3648
rect 10664 -3648 10698 -3281
rect 10732 -3469 10738 -3281
rect 10772 -3469 10778 -3093
rect 10732 -3481 10778 -3469
rect 10850 -3093 10896 -3081
rect 10850 -3469 10856 -3093
rect 10890 -3469 10896 -3093
rect 10850 -3481 10896 -3469
rect 10968 -3093 11014 -3081
rect 10968 -3469 10974 -3093
rect 11008 -3469 11014 -3093
rect 10968 -3481 11014 -3469
rect 11086 -3093 11132 -3081
rect 11086 -3469 11092 -3093
rect 11126 -3469 11132 -3093
rect 11086 -3481 11132 -3469
rect 11204 -3093 11328 -3081
rect 11204 -3469 11210 -3093
rect 11244 -3269 11288 -3093
rect 11322 -3269 11328 -3093
rect 11244 -3281 11328 -3269
rect 11400 -3093 11446 -3081
rect 13747 -3085 13781 -2962
rect 14219 -2975 14285 -2962
rect 14219 -3009 14235 -2975
rect 14269 -3009 14285 -2975
rect 14219 -3025 14285 -3009
rect 14608 -3085 14642 -2961
rect 16057 -2962 17429 -2915
rect 17751 -2961 18655 -2914
rect 19189 -2911 19224 -2401
rect 19279 -2447 19371 -2434
rect 19279 -2510 19291 -2447
rect 19362 -2510 19371 -2447
rect 19279 -2519 19371 -2510
rect 20364 -2447 20456 -2437
rect 20364 -2509 20376 -2447
rect 20446 -2509 20456 -2447
rect 20364 -2522 20456 -2509
rect 21752 -2502 21787 -2148
rect 22333 -2334 22368 -2148
rect 23242 -2232 23276 -2148
rect 24423 -2232 24457 -2148
rect 23242 -2274 24457 -2232
rect 24423 -2294 24457 -2274
rect 24423 -2310 24780 -2294
rect 22333 -2351 23470 -2334
rect 22333 -2385 23420 -2351
rect 23454 -2385 23470 -2351
rect 24423 -2344 24730 -2310
rect 24764 -2344 24780 -2310
rect 24423 -2360 24780 -2344
rect 22333 -2401 23470 -2385
rect 22074 -2446 22250 -2438
rect 20611 -2564 20676 -2561
rect 20611 -2567 20680 -2564
rect 20611 -2627 20617 -2567
rect 20676 -2627 20686 -2567
rect 20611 -2631 20680 -2627
rect 20611 -2633 20676 -2631
rect 21752 -2648 21933 -2502
rect 22074 -2514 22191 -2446
rect 22248 -2514 22258 -2446
rect 22074 -2522 22250 -2514
rect 22074 -2562 22250 -2554
rect 22074 -2630 22191 -2562
rect 22248 -2630 22258 -2562
rect 22074 -2638 22250 -2630
rect 20246 -2730 20338 -2722
rect 20246 -2795 20258 -2730
rect 20326 -2795 20338 -2730
rect 20246 -2807 20338 -2795
rect 21752 -2910 21787 -2648
rect 22074 -2730 22250 -2722
rect 22074 -2798 22191 -2730
rect 22248 -2798 22258 -2730
rect 22074 -2806 22250 -2798
rect 19189 -2958 20561 -2911
rect 20883 -2957 21787 -2910
rect 22333 -2911 22368 -2401
rect 22423 -2447 22515 -2434
rect 22423 -2510 22435 -2447
rect 22506 -2510 22515 -2447
rect 22423 -2519 22515 -2510
rect 23508 -2447 23600 -2437
rect 23508 -2509 23520 -2447
rect 23590 -2509 23600 -2447
rect 23508 -2522 23600 -2509
rect 24896 -2502 24931 -2148
rect 23755 -2564 23820 -2561
rect 23755 -2567 23824 -2564
rect 23755 -2627 23761 -2567
rect 23820 -2627 23830 -2567
rect 23755 -2631 23824 -2627
rect 23755 -2633 23820 -2631
rect 24896 -2648 25077 -2502
rect 23390 -2730 23482 -2722
rect 23390 -2795 23402 -2730
rect 23470 -2795 23482 -2730
rect 23390 -2807 23482 -2795
rect 24896 -2910 24931 -2648
rect 16891 -3085 16925 -2962
rect 17363 -2975 17429 -2962
rect 17363 -3009 17379 -2975
rect 17413 -3009 17429 -2975
rect 17363 -3025 17429 -3009
rect 17752 -3085 17786 -2961
rect 20023 -3081 20057 -2958
rect 20495 -2971 20561 -2958
rect 20495 -3005 20511 -2971
rect 20545 -3005 20561 -2971
rect 20495 -3021 20561 -3005
rect 20884 -3081 20918 -2957
rect 22333 -2958 23705 -2911
rect 24027 -2957 24931 -2910
rect 23167 -3081 23201 -2958
rect 23639 -2971 23705 -2958
rect 23639 -3005 23655 -2971
rect 23689 -3005 23705 -2971
rect 23639 -3021 23705 -3005
rect 24028 -3081 24062 -2957
rect 11400 -3269 11406 -3093
rect 11440 -3269 11446 -3093
rect 11400 -3281 11446 -3269
rect 13742 -3097 13788 -3085
rect 13742 -3273 13748 -3097
rect 13782 -3273 13788 -3097
rect 11244 -3469 11250 -3281
rect 11204 -3481 11250 -3469
rect 10974 -3554 11008 -3481
rect 10959 -3570 11025 -3554
rect 10959 -3604 10975 -3570
rect 11009 -3604 11025 -3570
rect 10959 -3620 11025 -3604
rect 11288 -3648 11322 -3281
rect 13742 -3285 13788 -3273
rect 13860 -3097 13980 -3085
rect 13860 -3273 13866 -3097
rect 13900 -3273 13940 -3097
rect 13860 -3285 13940 -3273
rect 10664 -3700 11322 -3648
rect 13866 -3652 13900 -3285
rect 13934 -3473 13940 -3285
rect 13974 -3473 13980 -3097
rect 13934 -3485 13980 -3473
rect 14052 -3097 14098 -3085
rect 14052 -3473 14058 -3097
rect 14092 -3473 14098 -3097
rect 14052 -3485 14098 -3473
rect 14170 -3097 14216 -3085
rect 14170 -3473 14176 -3097
rect 14210 -3473 14216 -3097
rect 14170 -3485 14216 -3473
rect 14288 -3097 14334 -3085
rect 14288 -3473 14294 -3097
rect 14328 -3473 14334 -3097
rect 14288 -3485 14334 -3473
rect 14406 -3097 14530 -3085
rect 14406 -3473 14412 -3097
rect 14446 -3273 14490 -3097
rect 14524 -3273 14530 -3097
rect 14446 -3285 14530 -3273
rect 14602 -3097 14648 -3085
rect 14602 -3273 14608 -3097
rect 14642 -3273 14648 -3097
rect 14602 -3285 14648 -3273
rect 16886 -3097 16932 -3085
rect 16886 -3273 16892 -3097
rect 16926 -3273 16932 -3097
rect 16886 -3285 16932 -3273
rect 17004 -3097 17124 -3085
rect 17004 -3273 17010 -3097
rect 17044 -3273 17084 -3097
rect 17004 -3285 17084 -3273
rect 14446 -3473 14452 -3285
rect 14406 -3485 14452 -3473
rect 14176 -3558 14210 -3485
rect 14161 -3574 14227 -3558
rect 14161 -3608 14177 -3574
rect 14211 -3608 14227 -3574
rect 14161 -3624 14227 -3608
rect 14490 -3652 14524 -3285
rect 1542 -3726 1634 -3704
rect 1542 -3778 1554 -3726
rect 1620 -3778 1634 -3726
rect 1542 -3782 1634 -3778
rect 4686 -3726 4778 -3704
rect 4686 -3778 4698 -3726
rect 4764 -3778 4778 -3726
rect 7818 -3722 7910 -3700
rect 7818 -3774 7830 -3722
rect 7896 -3774 7910 -3722
rect 7818 -3778 7910 -3774
rect 10962 -3722 11054 -3700
rect 13866 -3704 14524 -3652
rect 17010 -3652 17044 -3285
rect 17078 -3473 17084 -3285
rect 17118 -3473 17124 -3097
rect 17078 -3485 17124 -3473
rect 17196 -3097 17242 -3085
rect 17196 -3473 17202 -3097
rect 17236 -3473 17242 -3097
rect 17196 -3485 17242 -3473
rect 17314 -3097 17360 -3085
rect 17314 -3473 17320 -3097
rect 17354 -3473 17360 -3097
rect 17314 -3485 17360 -3473
rect 17432 -3097 17478 -3085
rect 17432 -3473 17438 -3097
rect 17472 -3473 17478 -3097
rect 17432 -3485 17478 -3473
rect 17550 -3097 17674 -3085
rect 17550 -3473 17556 -3097
rect 17590 -3273 17634 -3097
rect 17668 -3273 17674 -3097
rect 17590 -3285 17674 -3273
rect 17746 -3097 17792 -3085
rect 17746 -3273 17752 -3097
rect 17786 -3273 17792 -3097
rect 17746 -3285 17792 -3273
rect 20018 -3093 20064 -3081
rect 20018 -3269 20024 -3093
rect 20058 -3269 20064 -3093
rect 20018 -3281 20064 -3269
rect 20136 -3093 20256 -3081
rect 20136 -3269 20142 -3093
rect 20176 -3269 20216 -3093
rect 20136 -3281 20216 -3269
rect 17590 -3473 17596 -3285
rect 17550 -3485 17596 -3473
rect 17320 -3558 17354 -3485
rect 17305 -3574 17371 -3558
rect 17305 -3608 17321 -3574
rect 17355 -3608 17371 -3574
rect 17305 -3624 17371 -3608
rect 17634 -3652 17668 -3285
rect 17010 -3704 17668 -3652
rect 20142 -3648 20176 -3281
rect 20210 -3469 20216 -3281
rect 20250 -3469 20256 -3093
rect 20210 -3481 20256 -3469
rect 20328 -3093 20374 -3081
rect 20328 -3469 20334 -3093
rect 20368 -3469 20374 -3093
rect 20328 -3481 20374 -3469
rect 20446 -3093 20492 -3081
rect 20446 -3469 20452 -3093
rect 20486 -3469 20492 -3093
rect 20446 -3481 20492 -3469
rect 20564 -3093 20610 -3081
rect 20564 -3469 20570 -3093
rect 20604 -3469 20610 -3093
rect 20564 -3481 20610 -3469
rect 20682 -3093 20806 -3081
rect 20682 -3469 20688 -3093
rect 20722 -3269 20766 -3093
rect 20800 -3269 20806 -3093
rect 20722 -3281 20806 -3269
rect 20878 -3093 20924 -3081
rect 20878 -3269 20884 -3093
rect 20918 -3269 20924 -3093
rect 20878 -3281 20924 -3269
rect 23162 -3093 23208 -3081
rect 23162 -3269 23168 -3093
rect 23202 -3269 23208 -3093
rect 23162 -3281 23208 -3269
rect 23280 -3093 23400 -3081
rect 23280 -3269 23286 -3093
rect 23320 -3269 23360 -3093
rect 23280 -3281 23360 -3269
rect 20722 -3469 20728 -3281
rect 20682 -3481 20728 -3469
rect 20452 -3554 20486 -3481
rect 20437 -3570 20503 -3554
rect 20437 -3604 20453 -3570
rect 20487 -3604 20503 -3570
rect 20437 -3620 20503 -3604
rect 20766 -3648 20800 -3281
rect 20142 -3700 20800 -3648
rect 23286 -3648 23320 -3281
rect 23354 -3469 23360 -3281
rect 23394 -3469 23400 -3093
rect 23354 -3481 23400 -3469
rect 23472 -3093 23518 -3081
rect 23472 -3469 23478 -3093
rect 23512 -3469 23518 -3093
rect 23472 -3481 23518 -3469
rect 23590 -3093 23636 -3081
rect 23590 -3469 23596 -3093
rect 23630 -3469 23636 -3093
rect 23590 -3481 23636 -3469
rect 23708 -3093 23754 -3081
rect 23708 -3469 23714 -3093
rect 23748 -3469 23754 -3093
rect 23708 -3481 23754 -3469
rect 23826 -3093 23950 -3081
rect 23826 -3469 23832 -3093
rect 23866 -3269 23910 -3093
rect 23944 -3269 23950 -3093
rect 23866 -3281 23950 -3269
rect 24022 -3093 24068 -3081
rect 24022 -3269 24028 -3093
rect 24062 -3269 24068 -3093
rect 24022 -3281 24068 -3269
rect 23866 -3469 23872 -3281
rect 23826 -3481 23872 -3469
rect 23596 -3554 23630 -3481
rect 23581 -3570 23647 -3554
rect 23581 -3604 23597 -3570
rect 23631 -3604 23647 -3570
rect 23581 -3620 23647 -3604
rect 23910 -3648 23944 -3281
rect 23286 -3700 23944 -3648
rect 10962 -3774 10974 -3722
rect 11040 -3774 11054 -3722
rect 10962 -3778 11054 -3774
rect 14164 -3726 14256 -3704
rect 14164 -3778 14176 -3726
rect 14242 -3778 14256 -3726
rect 4686 -3782 4778 -3778
rect 14164 -3782 14256 -3778
rect 17308 -3726 17400 -3704
rect 17308 -3778 17320 -3726
rect 17386 -3778 17400 -3726
rect 20440 -3722 20532 -3700
rect 20440 -3774 20452 -3722
rect 20518 -3774 20532 -3722
rect 20440 -3778 20532 -3774
rect 23584 -3722 23676 -3700
rect 23584 -3774 23596 -3722
rect 23662 -3774 23676 -3722
rect 23584 -3778 23676 -3774
rect 17308 -3782 17400 -3778
<< via1 >>
rect 1714 22230 1794 22236
rect 1714 22176 1718 22230
rect 1718 22176 1790 22230
rect 1790 22176 1794 22230
rect 4858 22230 4938 22236
rect 4858 22176 4862 22230
rect 4862 22176 4934 22230
rect 4934 22176 4938 22230
rect 7990 22234 8070 22240
rect 7990 22180 7994 22234
rect 7994 22180 8066 22234
rect 8066 22180 8070 22234
rect 11134 22234 11214 22240
rect 11134 22180 11138 22234
rect 11138 22180 11210 22234
rect 11210 22180 11214 22234
rect 14336 22230 14416 22236
rect 14336 22176 14340 22230
rect 14340 22176 14412 22230
rect 14412 22176 14416 22230
rect 17480 22230 17560 22236
rect 17480 22176 17484 22230
rect 17484 22176 17556 22230
rect 17556 22176 17560 22230
rect 20612 22234 20692 22240
rect 20612 22180 20616 22234
rect 20616 22180 20688 22234
rect 20688 22180 20692 22234
rect 23756 22234 23836 22240
rect 23756 22180 23760 22234
rect 23760 22180 23832 22234
rect 23832 22180 23836 22234
rect 324 21381 378 21443
rect 323 21290 380 21294
rect 323 21230 327 21290
rect 327 21230 376 21290
rect 376 21230 380 21290
rect 323 21226 380 21230
rect 323 21006 380 21010
rect 323 20946 327 21006
rect 327 20946 376 21006
rect 376 20946 380 21006
rect 323 20942 380 20946
rect 567 21289 638 21293
rect 567 21234 571 21289
rect 571 21234 631 21289
rect 631 21234 638 21289
rect 567 21230 638 21234
rect 1652 21290 1722 21293
rect 1652 21235 1656 21290
rect 1656 21235 1716 21290
rect 1716 21235 1722 21290
rect 1652 21231 1722 21235
rect 3352 21343 3412 21396
rect 1893 21159 1952 21173
rect 1893 21125 1906 21159
rect 1906 21125 1940 21159
rect 1940 21125 1952 21159
rect 1893 21113 1952 21125
rect 3467 21174 3524 21178
rect 3467 21114 3471 21174
rect 3471 21114 3520 21174
rect 3520 21114 3524 21174
rect 3467 21110 3524 21114
rect 1534 21005 1602 21010
rect 1534 20950 1538 21005
rect 1538 20950 1598 21005
rect 1598 20950 1602 21005
rect 1534 20945 1602 20950
rect 323 20706 377 20768
rect 323 20571 377 20633
rect 325 20459 379 20521
rect 325 20334 379 20396
rect 330 20093 384 20155
rect 1728 19972 1732 20018
rect 1732 19972 1790 20018
rect 1790 19972 1794 20018
rect 1728 19966 1794 19972
rect 327 19871 381 19933
rect 3467 21006 3524 21010
rect 3467 20946 3471 21006
rect 3471 20946 3520 21006
rect 3520 20946 3524 21006
rect 3467 20942 3524 20946
rect 3711 21289 3782 21293
rect 3711 21234 3715 21289
rect 3715 21234 3775 21289
rect 3775 21234 3782 21289
rect 3711 21230 3782 21234
rect 4796 21290 4866 21293
rect 4796 21235 4800 21290
rect 4800 21235 4860 21290
rect 4860 21235 4866 21290
rect 4796 21231 4866 21235
rect 5037 21159 5096 21173
rect 5037 21125 5050 21159
rect 5050 21125 5084 21159
rect 5084 21125 5096 21159
rect 5037 21113 5096 21125
rect 4678 21005 4746 21010
rect 4678 20950 4682 21005
rect 4682 20950 4742 21005
rect 4742 20950 4746 21005
rect 4678 20945 4746 20950
rect 3362 20712 3432 20772
rect 6599 21010 6656 21014
rect 6599 20950 6603 21010
rect 6603 20950 6652 21010
rect 6652 20950 6656 21010
rect 6599 20946 6656 20950
rect 6843 21293 6914 21297
rect 6843 21238 6847 21293
rect 6847 21238 6907 21293
rect 6907 21238 6914 21293
rect 6843 21234 6914 21238
rect 7928 21294 7998 21297
rect 7928 21239 7932 21294
rect 7932 21239 7992 21294
rect 7992 21239 7998 21294
rect 7928 21235 7998 21239
rect 8169 21163 8228 21177
rect 8169 21129 8182 21163
rect 8182 21129 8216 21163
rect 8216 21129 8228 21163
rect 8169 21117 8228 21129
rect 9743 21178 9800 21182
rect 9743 21118 9747 21178
rect 9747 21118 9796 21178
rect 9796 21118 9800 21178
rect 9743 21114 9800 21118
rect 7810 21009 7878 21014
rect 7810 20954 7814 21009
rect 7814 20954 7874 21009
rect 7874 20954 7878 21009
rect 7810 20949 7878 20954
rect 6512 20574 6576 20631
rect 6244 20096 6303 20162
rect 9743 21010 9800 21014
rect 9743 20950 9747 21010
rect 9747 20950 9796 21010
rect 9796 20950 9800 21010
rect 9743 20946 9800 20950
rect 9987 21293 10058 21297
rect 9987 21238 9991 21293
rect 9991 21238 10051 21293
rect 10051 21238 10058 21293
rect 9987 21234 10058 21238
rect 11072 21294 11142 21297
rect 11072 21239 11076 21294
rect 11076 21239 11136 21294
rect 11136 21239 11142 21294
rect 11072 21235 11142 21239
rect 11313 21163 11372 21177
rect 11313 21129 11326 21163
rect 11326 21129 11360 21163
rect 11360 21129 11372 21163
rect 11313 21117 11372 21129
rect 10954 21009 11022 21014
rect 10954 20954 10958 21009
rect 10958 20954 11018 21009
rect 11018 20954 11022 21009
rect 10954 20949 11022 20954
rect 9654 20468 9708 20526
rect 9370 20222 9429 20279
rect 12545 20359 12607 20427
rect 12945 21006 13002 21010
rect 12945 20946 12949 21006
rect 12949 20946 12998 21006
rect 12998 20946 13002 21006
rect 12945 20942 13002 20946
rect 13189 21289 13260 21293
rect 13189 21234 13193 21289
rect 13193 21234 13253 21289
rect 13253 21234 13260 21289
rect 13189 21230 13260 21234
rect 14274 21290 14344 21293
rect 14274 21235 14278 21290
rect 14278 21235 14338 21290
rect 14338 21235 14344 21290
rect 14274 21231 14344 21235
rect 14515 21159 14574 21173
rect 14515 21125 14528 21159
rect 14528 21125 14562 21159
rect 14562 21125 14574 21159
rect 14515 21113 14574 21125
rect 16089 21174 16146 21178
rect 16089 21114 16093 21174
rect 16093 21114 16142 21174
rect 16142 21114 16146 21174
rect 16089 21110 16146 21114
rect 14156 21005 14224 21010
rect 14156 20950 14160 21005
rect 14160 20950 14220 21005
rect 14220 20950 14224 21005
rect 14156 20945 14224 20950
rect 12824 20241 12893 20302
rect 16089 21006 16146 21010
rect 16089 20946 16093 21006
rect 16093 20946 16142 21006
rect 16142 20946 16146 21006
rect 16089 20942 16146 20946
rect 15770 20509 15826 20578
rect 16333 21289 16404 21293
rect 16333 21234 16337 21289
rect 16337 21234 16397 21289
rect 16397 21234 16404 21289
rect 16333 21230 16404 21234
rect 17418 21290 17488 21293
rect 17418 21235 17422 21290
rect 17422 21235 17482 21290
rect 17482 21235 17488 21290
rect 17418 21231 17488 21235
rect 17659 21159 17718 21173
rect 17659 21125 17672 21159
rect 17672 21125 17706 21159
rect 17706 21125 17718 21159
rect 17659 21113 17718 21125
rect 19221 21178 19278 21182
rect 19221 21118 19225 21178
rect 19225 21118 19274 21178
rect 19274 21118 19278 21178
rect 19221 21114 19278 21118
rect 17300 21005 17368 21010
rect 17300 20950 17304 21005
rect 17304 20950 17364 21005
rect 17364 20950 17368 21005
rect 17300 20945 17368 20950
rect 19221 21010 19278 21014
rect 19221 20950 19225 21010
rect 19225 20950 19274 21010
rect 19274 20950 19278 21010
rect 19221 20946 19278 20950
rect 18906 20672 18970 20731
rect 15975 20100 16032 20167
rect 4872 19972 4876 20018
rect 4876 19972 4934 20018
rect 4934 19972 4938 20018
rect 4872 19966 4938 19972
rect 8004 19976 8008 20022
rect 8008 19976 8066 20022
rect 8066 19976 8070 20022
rect 8004 19970 8070 19976
rect 11148 19976 11152 20022
rect 11152 19976 11210 20022
rect 11210 19976 11214 20022
rect 11148 19970 11214 19976
rect 14350 19972 14354 20018
rect 14354 19972 14412 20018
rect 14412 19972 14416 20018
rect 14350 19966 14416 19972
rect 17494 19972 17498 20018
rect 17498 19972 17556 20018
rect 17556 19972 17560 20018
rect 17494 19966 17560 19972
rect 19465 21293 19536 21297
rect 19465 21238 19469 21293
rect 19469 21238 19529 21293
rect 19529 21238 19536 21293
rect 19465 21234 19536 21238
rect 20550 21294 20620 21297
rect 20550 21239 20554 21294
rect 20554 21239 20614 21294
rect 20614 21239 20620 21294
rect 20550 21235 20620 21239
rect 20791 21163 20850 21177
rect 20791 21129 20804 21163
rect 20804 21129 20838 21163
rect 20838 21129 20850 21163
rect 20791 21117 20850 21129
rect 22365 21178 22422 21182
rect 22365 21118 22369 21178
rect 22369 21118 22418 21178
rect 22418 21118 22422 21178
rect 22365 21114 22422 21118
rect 20432 21009 20500 21014
rect 20432 20954 20436 21009
rect 20436 20954 20496 21009
rect 20496 20954 20500 21009
rect 20432 20949 20500 20954
rect 22051 20801 22104 20858
rect 22609 21293 22680 21297
rect 22609 21238 22613 21293
rect 22613 21238 22673 21293
rect 22673 21238 22680 21293
rect 22609 21234 22680 21238
rect 23694 21294 23764 21297
rect 23694 21239 23698 21294
rect 23698 21239 23758 21294
rect 23758 21239 23764 21294
rect 23694 21235 23764 21239
rect 23935 21163 23994 21177
rect 23935 21129 23948 21163
rect 23948 21129 23982 21163
rect 23982 21129 23994 21163
rect 23935 21117 23994 21129
rect 23576 21009 23644 21014
rect 23576 20954 23580 21009
rect 23580 20954 23640 21009
rect 23640 20954 23644 21009
rect 23576 20949 23644 20954
rect 25549 20795 25620 20866
rect 25537 20670 25603 20730
rect 25527 20503 25591 20572
rect 25527 20357 25591 20426
rect 25527 20217 25591 20286
rect 25526 20078 25590 20147
rect 20626 19976 20630 20022
rect 20630 19976 20688 20022
rect 20688 19976 20692 20022
rect 20626 19970 20692 19976
rect 23770 19976 23774 20022
rect 23774 19976 23832 20022
rect 23832 19976 23836 20022
rect 23770 19970 23836 19976
rect 3111 19801 3184 19882
rect 19104 19875 19174 19951
rect 25526 19810 25590 19879
rect 230 18577 290 18636
rect 13012 18561 13066 18615
rect 13106 18468 13160 18522
rect 227 18374 287 18436
rect 220 18184 280 18246
rect 220 17995 280 18064
rect 207 17814 268 17877
rect 194 17614 265 17686
rect 211 15825 265 15880
rect 182 15451 238 15505
rect 201 11350 263 11425
rect 202 11023 264 11098
rect 11474 18376 11528 18430
rect 11649 18281 11703 18335
rect 471 7096 526 7157
rect 727 7099 795 7157
rect 471 6804 526 6865
rect 471 6499 526 6560
rect 471 6338 526 6399
rect 471 6187 527 6248
rect 471 6027 526 6088
rect 471 5840 526 5901
rect 471 5634 526 5695
rect 10013 18191 10067 18245
rect 986 6806 1042 6863
rect 10151 18097 10205 18151
rect 8511 18003 8565 18057
rect 8690 17909 8744 17963
rect 1204 6502 1265 6555
rect 7055 17819 7109 17873
rect 7183 17724 7237 17778
rect 1379 6340 1449 6398
rect 5602 17633 5656 17687
rect 1581 6190 1649 6248
rect 5733 17538 5787 17592
rect 4157 17447 4211 17501
rect 4267 17354 4321 17408
rect 1777 6031 1835 6085
rect 2415 16122 2486 16181
rect 3250 16775 3310 16837
rect 4698 16775 4758 16837
rect 6196 16777 6256 16839
rect 7644 16777 7704 16839
rect 9164 16775 9224 16837
rect 10612 16775 10672 16837
rect 12110 16777 12170 16839
rect 13558 16777 13618 16839
rect 15244 16973 15296 17025
rect 16412 16973 16464 17025
rect 2701 16021 2770 16085
rect 3472 15625 3534 15633
rect 3472 15579 3478 15625
rect 3478 15579 3530 15625
rect 3530 15579 3534 15625
rect 3472 15573 3534 15579
rect 4474 15958 4528 16012
rect 4359 15826 4413 15881
rect 4920 15625 4982 15633
rect 4920 15579 4926 15625
rect 4926 15579 4978 15625
rect 4978 15579 4982 15625
rect 4920 15573 4982 15579
rect 5968 15957 6022 16011
rect 5857 15825 5911 15879
rect 6418 15627 6480 15635
rect 6418 15581 6424 15627
rect 6424 15581 6476 15627
rect 6476 15581 6480 15627
rect 6418 15575 6480 15581
rect 2205 14070 2288 14158
rect 4216 15092 4296 15098
rect 4216 15038 4220 15092
rect 4220 15038 4292 15092
rect 4292 15038 4296 15092
rect 2825 14036 2882 14040
rect 2825 13976 2829 14036
rect 2829 13976 2878 14036
rect 2878 13976 2882 14036
rect 2825 13972 2882 13976
rect 2825 13868 2882 13872
rect 2825 13808 2829 13868
rect 2829 13808 2878 13868
rect 2878 13808 2882 13868
rect 2825 13804 2882 13808
rect 3069 14151 3140 14155
rect 3069 14096 3073 14151
rect 3073 14096 3133 14151
rect 3133 14096 3140 14151
rect 3069 14092 3140 14096
rect 4154 14152 4224 14155
rect 4154 14097 4158 14152
rect 4158 14097 4218 14152
rect 4218 14097 4224 14152
rect 4154 14093 4224 14097
rect 4395 14021 4454 14035
rect 4395 13987 4408 14021
rect 4408 13987 4442 14021
rect 4442 13987 4454 14021
rect 4395 13975 4454 13987
rect 7418 15960 7472 16014
rect 7305 15830 7359 15884
rect 17580 16973 17632 17025
rect 18748 16973 18800 17025
rect 7866 15627 7928 15635
rect 7866 15581 7872 15627
rect 7872 15581 7924 15627
rect 7924 15581 7928 15627
rect 7866 15575 7928 15581
rect 8937 15955 8991 16009
rect 8821 15830 8875 15884
rect 9386 15625 9448 15633
rect 9386 15579 9392 15625
rect 9392 15579 9444 15625
rect 9444 15579 9448 15625
rect 9386 15573 9448 15579
rect 10385 15962 10439 16016
rect 10273 15824 10327 15878
rect 10834 15625 10896 15633
rect 10834 15579 10840 15625
rect 10840 15579 10892 15625
rect 10892 15579 10896 15625
rect 10834 15573 10896 15579
rect 11882 15960 11936 16014
rect 11770 15830 11824 15884
rect 12332 15627 12394 15635
rect 12332 15581 12338 15627
rect 12338 15581 12390 15627
rect 12390 15581 12394 15627
rect 12332 15575 12394 15581
rect 13314 15942 13400 16030
rect 13200 15813 13286 15901
rect 13780 15627 13842 15635
rect 13780 15581 13786 15627
rect 13786 15581 13838 15627
rect 13838 15581 13842 15627
rect 13780 15575 13842 15581
rect 19922 16975 19974 17027
rect 21090 16975 21142 17027
rect 22258 16975 22310 17027
rect 23426 16975 23478 17027
rect 14773 15649 14825 15701
rect 15941 15649 15993 15701
rect 17109 15649 17161 15701
rect 18277 15649 18329 15701
rect 19451 15651 19503 15703
rect 20619 15651 20671 15703
rect 21787 15651 21839 15703
rect 22955 15651 23007 15703
rect 7360 15092 7440 15098
rect 7360 15038 7364 15092
rect 7364 15038 7436 15092
rect 7436 15038 7440 15092
rect 5969 14036 6026 14040
rect 5969 13976 5973 14036
rect 5973 13976 6022 14036
rect 6022 13976 6026 14036
rect 5969 13972 6026 13976
rect 4036 13867 4104 13872
rect 4036 13812 4040 13867
rect 4040 13812 4100 13867
rect 4100 13812 4104 13867
rect 4036 13807 4104 13812
rect 4230 12834 4234 12880
rect 4234 12834 4292 12880
rect 4292 12834 4296 12880
rect 4230 12828 4296 12834
rect 5969 13868 6026 13872
rect 5969 13808 5973 13868
rect 5973 13808 6022 13868
rect 6022 13808 6026 13868
rect 5969 13804 6026 13808
rect 6213 14151 6284 14155
rect 6213 14096 6217 14151
rect 6217 14096 6277 14151
rect 6277 14096 6284 14151
rect 6213 14092 6284 14096
rect 7298 14152 7368 14155
rect 7298 14097 7302 14152
rect 7302 14097 7362 14152
rect 7362 14097 7368 14152
rect 7298 14093 7368 14097
rect 7539 14021 7598 14035
rect 7539 13987 7552 14021
rect 7552 13987 7586 14021
rect 7586 13987 7598 14021
rect 7539 13975 7598 13987
rect 10492 15096 10572 15102
rect 10492 15042 10496 15096
rect 10496 15042 10568 15096
rect 10568 15042 10572 15096
rect 9101 14040 9158 14044
rect 9101 13980 9105 14040
rect 9105 13980 9154 14040
rect 9154 13980 9158 14040
rect 9101 13976 9158 13980
rect 7180 13867 7248 13872
rect 7180 13812 7184 13867
rect 7184 13812 7244 13867
rect 7244 13812 7248 13867
rect 7180 13807 7248 13812
rect 7374 12834 7378 12880
rect 7378 12834 7436 12880
rect 7436 12834 7440 12880
rect 7374 12828 7440 12834
rect 9101 13872 9158 13876
rect 9101 13812 9105 13872
rect 9105 13812 9154 13872
rect 9154 13812 9158 13872
rect 9101 13808 9158 13812
rect 9345 14155 9416 14159
rect 9345 14100 9349 14155
rect 9349 14100 9409 14155
rect 9409 14100 9416 14155
rect 9345 14096 9416 14100
rect 10430 14156 10500 14159
rect 10430 14101 10434 14156
rect 10434 14101 10494 14156
rect 10494 14101 10500 14156
rect 10430 14097 10500 14101
rect 10671 14025 10730 14039
rect 10671 13991 10684 14025
rect 10684 13991 10718 14025
rect 10718 13991 10730 14025
rect 10671 13979 10730 13991
rect 13636 15096 13716 15102
rect 13636 15042 13640 15096
rect 13640 15042 13712 15096
rect 13712 15042 13716 15096
rect 12245 14040 12302 14044
rect 12245 13980 12249 14040
rect 12249 13980 12298 14040
rect 12298 13980 12302 14040
rect 12245 13976 12302 13980
rect 10312 13871 10380 13876
rect 10312 13816 10316 13871
rect 10316 13816 10376 13871
rect 10376 13816 10380 13871
rect 10312 13811 10380 13816
rect 10506 12838 10510 12884
rect 10510 12838 10568 12884
rect 10568 12838 10572 12884
rect 10506 12832 10572 12838
rect 12489 14155 12560 14159
rect 12489 14100 12493 14155
rect 12493 14100 12553 14155
rect 12553 14100 12560 14155
rect 12489 14096 12560 14100
rect 13574 14156 13644 14159
rect 13574 14101 13578 14156
rect 13578 14101 13638 14156
rect 13638 14101 13644 14156
rect 13574 14097 13644 14101
rect 13815 14025 13874 14039
rect 13815 13991 13828 14025
rect 13828 13991 13862 14025
rect 13862 13991 13874 14025
rect 13815 13979 13874 13991
rect 16838 15092 16918 15098
rect 16838 15038 16842 15092
rect 16842 15038 16914 15092
rect 16914 15038 16918 15092
rect 15447 14036 15504 14040
rect 15447 13976 15451 14036
rect 15451 13976 15500 14036
rect 15500 13976 15504 14036
rect 15447 13972 15504 13976
rect 13650 12838 13654 12884
rect 13654 12838 13712 12884
rect 13712 12838 13716 12884
rect 13650 12832 13716 12838
rect 15691 14151 15762 14155
rect 15691 14096 15695 14151
rect 15695 14096 15755 14151
rect 15755 14096 15762 14151
rect 15691 14092 15762 14096
rect 16776 14152 16846 14155
rect 16776 14097 16780 14152
rect 16780 14097 16840 14152
rect 16840 14097 16846 14152
rect 16776 14093 16846 14097
rect 17017 14021 17076 14035
rect 17017 13987 17030 14021
rect 17030 13987 17064 14021
rect 17064 13987 17076 14021
rect 17017 13975 17076 13987
rect 19982 15092 20062 15098
rect 19982 15038 19986 15092
rect 19986 15038 20058 15092
rect 20058 15038 20062 15092
rect 18591 14036 18648 14040
rect 18591 13976 18595 14036
rect 18595 13976 18644 14036
rect 18644 13976 18648 14036
rect 18591 13972 18648 13976
rect 16852 12834 16856 12880
rect 16856 12834 16914 12880
rect 16914 12834 16918 12880
rect 16852 12828 16918 12834
rect 18591 13868 18648 13872
rect 18591 13808 18595 13868
rect 18595 13808 18644 13868
rect 18644 13808 18648 13868
rect 18591 13804 18648 13808
rect 18835 14151 18906 14155
rect 18835 14096 18839 14151
rect 18839 14096 18899 14151
rect 18899 14096 18906 14151
rect 18835 14092 18906 14096
rect 19920 14152 19990 14155
rect 19920 14097 19924 14152
rect 19924 14097 19984 14152
rect 19984 14097 19990 14152
rect 19920 14093 19990 14097
rect 20161 14021 20220 14035
rect 20161 13987 20174 14021
rect 20174 13987 20208 14021
rect 20208 13987 20220 14021
rect 20161 13975 20220 13987
rect 23114 15096 23194 15102
rect 23114 15042 23118 15096
rect 23118 15042 23190 15096
rect 23190 15042 23194 15096
rect 21723 14040 21780 14044
rect 21723 13980 21727 14040
rect 21727 13980 21776 14040
rect 21776 13980 21780 14040
rect 21723 13976 21780 13980
rect 19802 13867 19870 13872
rect 19802 13812 19806 13867
rect 19806 13812 19866 13867
rect 19866 13812 19870 13867
rect 19802 13807 19870 13812
rect 19996 12834 20000 12880
rect 20000 12834 20058 12880
rect 20058 12834 20062 12880
rect 19996 12828 20062 12834
rect 21723 13872 21780 13876
rect 21723 13812 21727 13872
rect 21727 13812 21776 13872
rect 21776 13812 21780 13872
rect 21723 13808 21780 13812
rect 21967 14155 22038 14159
rect 21967 14100 21971 14155
rect 21971 14100 22031 14155
rect 22031 14100 22038 14155
rect 21967 14096 22038 14100
rect 23052 14156 23122 14159
rect 23052 14101 23056 14156
rect 23056 14101 23116 14156
rect 23116 14101 23122 14156
rect 23052 14097 23122 14101
rect 23293 14025 23352 14039
rect 23293 13991 23306 14025
rect 23306 13991 23340 14025
rect 23340 13991 23352 14025
rect 23293 13979 23352 13991
rect 26258 15096 26338 15102
rect 26258 15042 26262 15096
rect 26262 15042 26334 15096
rect 26334 15042 26338 15096
rect 24867 14040 24924 14044
rect 24867 13980 24871 14040
rect 24871 13980 24920 14040
rect 24920 13980 24924 14040
rect 24867 13976 24924 13980
rect 22934 13871 23002 13876
rect 22934 13816 22938 13871
rect 22938 13816 22998 13871
rect 22998 13816 23002 13871
rect 22934 13811 23002 13816
rect 23128 12838 23132 12884
rect 23132 12838 23190 12884
rect 23190 12838 23194 12884
rect 23128 12832 23194 12838
rect 24867 13872 24924 13876
rect 24867 13812 24871 13872
rect 24871 13812 24920 13872
rect 24920 13812 24924 13872
rect 24867 13808 24924 13812
rect 25111 14155 25182 14159
rect 25111 14100 25115 14155
rect 25115 14100 25175 14155
rect 25175 14100 25182 14155
rect 25111 14096 25182 14100
rect 26196 14156 26266 14159
rect 26196 14101 26200 14156
rect 26200 14101 26260 14156
rect 26260 14101 26266 14156
rect 26196 14097 26266 14101
rect 26437 14025 26496 14039
rect 26437 13991 26450 14025
rect 26450 13991 26484 14025
rect 26484 13991 26496 14025
rect 26437 13979 26496 13991
rect 26078 13871 26146 13876
rect 26078 13816 26082 13871
rect 26082 13816 26142 13871
rect 26142 13816 26146 13871
rect 26078 13811 26146 13816
rect 26272 12838 26276 12884
rect 26276 12838 26334 12884
rect 26334 12838 26338 12884
rect 26272 12832 26338 12838
rect 4216 12358 4296 12364
rect 4216 12304 4220 12358
rect 4220 12304 4292 12358
rect 4292 12304 4296 12358
rect 2825 11302 2882 11306
rect 2825 11242 2829 11302
rect 2829 11242 2878 11302
rect 2878 11242 2882 11302
rect 2825 11238 2882 11242
rect 2212 11029 2279 11099
rect 2825 11134 2882 11138
rect 2825 11074 2829 11134
rect 2829 11074 2878 11134
rect 2878 11074 2882 11134
rect 2825 11070 2882 11074
rect 3069 11417 3140 11421
rect 3069 11362 3073 11417
rect 3073 11362 3133 11417
rect 3133 11362 3140 11417
rect 3069 11358 3140 11362
rect 4154 11418 4224 11421
rect 4154 11363 4158 11418
rect 4158 11363 4218 11418
rect 4218 11363 4224 11418
rect 4154 11359 4224 11363
rect 4395 11287 4454 11301
rect 4395 11253 4408 11287
rect 4408 11253 4442 11287
rect 4442 11253 4454 11287
rect 4395 11241 4454 11253
rect 7360 12358 7440 12364
rect 7360 12304 7364 12358
rect 7364 12304 7436 12358
rect 7436 12304 7440 12358
rect 5969 11302 6026 11306
rect 5969 11242 5973 11302
rect 5973 11242 6022 11302
rect 6022 11242 6026 11302
rect 5969 11238 6026 11242
rect 4036 11133 4104 11138
rect 4036 11078 4040 11133
rect 4040 11078 4100 11133
rect 4100 11078 4104 11133
rect 4036 11073 4104 11078
rect 5969 11134 6026 11138
rect 5969 11074 5973 11134
rect 5973 11074 6022 11134
rect 6022 11074 6026 11134
rect 5969 11070 6026 11074
rect 4230 10100 4234 10146
rect 4234 10100 4292 10146
rect 4292 10100 4296 10146
rect 4230 10094 4296 10100
rect 5644 10100 5708 10177
rect 6213 11417 6284 11421
rect 6213 11362 6217 11417
rect 6217 11362 6277 11417
rect 6277 11362 6284 11417
rect 6213 11358 6284 11362
rect 7298 11418 7368 11421
rect 7298 11363 7302 11418
rect 7302 11363 7362 11418
rect 7362 11363 7368 11418
rect 7298 11359 7368 11363
rect 7539 11287 7598 11301
rect 7539 11253 7552 11287
rect 7552 11253 7586 11287
rect 7586 11253 7598 11287
rect 7539 11241 7598 11253
rect 10492 12362 10572 12368
rect 10492 12308 10496 12362
rect 10496 12308 10568 12362
rect 10568 12308 10572 12362
rect 9101 11306 9158 11310
rect 9101 11246 9105 11306
rect 9105 11246 9154 11306
rect 9154 11246 9158 11306
rect 9101 11242 9158 11246
rect 7180 11133 7248 11138
rect 7180 11078 7184 11133
rect 7184 11078 7244 11133
rect 7244 11078 7248 11133
rect 7180 11073 7248 11078
rect 7374 10100 7378 10146
rect 7378 10100 7436 10146
rect 7436 10100 7440 10146
rect 7374 10094 7440 10100
rect 8754 10046 8822 10118
rect 9101 11138 9158 11142
rect 9101 11078 9105 11138
rect 9105 11078 9154 11138
rect 9154 11078 9158 11138
rect 9101 11074 9158 11078
rect 9345 11421 9416 11425
rect 9345 11366 9349 11421
rect 9349 11366 9409 11421
rect 9409 11366 9416 11421
rect 9345 11362 9416 11366
rect 10430 11422 10500 11425
rect 10430 11367 10434 11422
rect 10434 11367 10494 11422
rect 10494 11367 10500 11422
rect 10430 11363 10500 11367
rect 10671 11291 10730 11305
rect 10671 11257 10684 11291
rect 10684 11257 10718 11291
rect 10718 11257 10730 11291
rect 10671 11245 10730 11257
rect 13636 12362 13716 12368
rect 13636 12308 13640 12362
rect 13640 12308 13712 12362
rect 13712 12308 13716 12362
rect 12245 11306 12302 11310
rect 12245 11246 12249 11306
rect 12249 11246 12298 11306
rect 12298 11246 12302 11306
rect 12245 11242 12302 11246
rect 10312 11137 10380 11142
rect 10312 11082 10316 11137
rect 10316 11082 10376 11137
rect 10376 11082 10380 11137
rect 10312 11077 10380 11082
rect 10506 10104 10510 10150
rect 10510 10104 10568 10150
rect 10568 10104 10572 10150
rect 10506 10098 10572 10104
rect 11890 9924 11957 9992
rect 12245 11138 12302 11142
rect 12245 11078 12249 11138
rect 12249 11078 12298 11138
rect 12298 11078 12302 11138
rect 12245 11074 12302 11078
rect 12489 11421 12560 11425
rect 12489 11366 12493 11421
rect 12493 11366 12553 11421
rect 12553 11366 12560 11421
rect 12489 11362 12560 11366
rect 13574 11422 13644 11425
rect 13574 11367 13578 11422
rect 13578 11367 13638 11422
rect 13638 11367 13644 11422
rect 13574 11363 13644 11367
rect 13815 11291 13874 11305
rect 13815 11257 13828 11291
rect 13828 11257 13862 11291
rect 13862 11257 13874 11291
rect 13815 11245 13874 11257
rect 16838 12358 16918 12364
rect 16838 12304 16842 12358
rect 16842 12304 16914 12358
rect 16914 12304 16918 12358
rect 15447 11302 15504 11306
rect 15447 11242 15451 11302
rect 15451 11242 15500 11302
rect 15500 11242 15504 11302
rect 15447 11238 15504 11242
rect 13456 11137 13524 11142
rect 13456 11082 13460 11137
rect 13460 11082 13520 11137
rect 13520 11082 13524 11137
rect 13456 11077 13524 11082
rect 15037 10267 15115 10336
rect 15447 11134 15504 11138
rect 15447 11074 15451 11134
rect 15451 11074 15500 11134
rect 15500 11074 15504 11134
rect 15447 11070 15504 11074
rect 13650 10104 13654 10150
rect 13654 10104 13712 10150
rect 13712 10104 13716 10150
rect 13650 10098 13716 10104
rect 15691 11417 15762 11421
rect 15691 11362 15695 11417
rect 15695 11362 15755 11417
rect 15755 11362 15762 11417
rect 15691 11358 15762 11362
rect 16776 11418 16846 11421
rect 16776 11363 16780 11418
rect 16780 11363 16840 11418
rect 16840 11363 16846 11418
rect 16776 11359 16846 11363
rect 17017 11287 17076 11301
rect 17017 11253 17030 11287
rect 17030 11253 17064 11287
rect 17064 11253 17076 11287
rect 17017 11241 17076 11253
rect 19982 12358 20062 12364
rect 19982 12304 19986 12358
rect 19986 12304 20058 12358
rect 20058 12304 20062 12358
rect 18591 11418 18648 11422
rect 18591 11358 18595 11418
rect 18595 11358 18644 11418
rect 18644 11358 18648 11418
rect 18591 11354 18648 11358
rect 18591 11302 18648 11306
rect 18591 11242 18595 11302
rect 18595 11242 18644 11302
rect 18644 11242 18648 11302
rect 18591 11238 18648 11242
rect 16658 11133 16726 11138
rect 16658 11078 16662 11133
rect 16662 11078 16722 11133
rect 16722 11078 16726 11133
rect 16658 11073 16726 11078
rect 18591 11134 18648 11138
rect 18591 11074 18595 11134
rect 18595 11074 18644 11134
rect 18644 11074 18648 11134
rect 18591 11070 18648 11074
rect 18237 10445 18333 10540
rect 16852 10100 16856 10146
rect 16856 10100 16914 10146
rect 16914 10100 16918 10146
rect 16852 10094 16918 10100
rect 18835 11417 18906 11421
rect 18835 11362 18839 11417
rect 18839 11362 18899 11417
rect 18899 11362 18906 11417
rect 18835 11358 18906 11362
rect 19920 11418 19990 11421
rect 19920 11363 19924 11418
rect 19924 11363 19984 11418
rect 19984 11363 19990 11418
rect 19920 11359 19990 11363
rect 20161 11287 20220 11301
rect 20161 11253 20174 11287
rect 20174 11253 20208 11287
rect 20208 11253 20220 11287
rect 20161 11241 20220 11253
rect 23114 12362 23194 12368
rect 23114 12308 23118 12362
rect 23118 12308 23190 12362
rect 23190 12308 23194 12362
rect 21723 11306 21780 11310
rect 21723 11246 21727 11306
rect 21727 11246 21776 11306
rect 21776 11246 21780 11306
rect 21723 11242 21780 11246
rect 19802 11133 19870 11138
rect 19802 11078 19806 11133
rect 19806 11078 19866 11133
rect 19866 11078 19870 11133
rect 19802 11073 19870 11078
rect 21396 10678 21466 10771
rect 21723 11138 21780 11142
rect 21723 11078 21727 11138
rect 21727 11078 21776 11138
rect 21776 11078 21780 11138
rect 21723 11074 21780 11078
rect 19996 10100 20000 10146
rect 20000 10100 20058 10146
rect 20058 10100 20062 10146
rect 19996 10094 20062 10100
rect 4206 9626 4286 9632
rect 4206 9572 4210 9626
rect 4210 9572 4282 9626
rect 4282 9572 4286 9626
rect 2815 8686 2872 8690
rect 2815 8626 2819 8686
rect 2819 8626 2868 8686
rect 2868 8626 2872 8686
rect 2815 8622 2872 8626
rect 2815 8570 2872 8574
rect 2815 8510 2819 8570
rect 2819 8510 2868 8570
rect 2868 8510 2872 8570
rect 2815 8506 2872 8510
rect 2815 8402 2872 8406
rect 2815 8342 2819 8402
rect 2819 8342 2868 8402
rect 2868 8342 2872 8402
rect 2815 8338 2872 8342
rect 3059 8685 3130 8689
rect 3059 8630 3063 8685
rect 3063 8630 3123 8685
rect 3123 8630 3130 8685
rect 3059 8626 3130 8630
rect 4144 8686 4214 8689
rect 4144 8631 4148 8686
rect 4148 8631 4208 8686
rect 4208 8631 4214 8686
rect 4144 8627 4214 8631
rect 7350 9626 7430 9632
rect 7350 9572 7354 9626
rect 7354 9572 7426 9626
rect 7426 9572 7430 9626
rect 4385 8555 4444 8569
rect 4385 8521 4398 8555
rect 4398 8521 4432 8555
rect 4432 8521 4444 8555
rect 4385 8509 4444 8521
rect 5959 8686 6016 8690
rect 5959 8626 5963 8686
rect 5963 8626 6012 8686
rect 6012 8626 6016 8686
rect 5959 8622 6016 8626
rect 5959 8570 6016 8574
rect 5959 8510 5963 8570
rect 5963 8510 6012 8570
rect 6012 8510 6016 8570
rect 5959 8506 6016 8510
rect 4026 8401 4094 8406
rect 4026 8346 4030 8401
rect 4030 8346 4090 8401
rect 4090 8346 4094 8401
rect 4026 8341 4094 8346
rect 5959 8402 6016 8406
rect 5959 8342 5963 8402
rect 5963 8342 6012 8402
rect 6012 8342 6016 8402
rect 5959 8338 6016 8342
rect 4220 7368 4224 7414
rect 4224 7368 4282 7414
rect 4282 7368 4286 7414
rect 4220 7362 4286 7368
rect 6203 8685 6274 8689
rect 6203 8630 6207 8685
rect 6207 8630 6267 8685
rect 6267 8630 6274 8685
rect 6203 8626 6274 8630
rect 7288 8686 7358 8689
rect 7288 8631 7292 8686
rect 7292 8631 7352 8686
rect 7352 8631 7358 8686
rect 7288 8627 7358 8631
rect 10482 9630 10562 9636
rect 10482 9576 10486 9630
rect 10486 9576 10558 9630
rect 10558 9576 10562 9630
rect 7529 8555 7588 8569
rect 7529 8521 7542 8555
rect 7542 8521 7576 8555
rect 7576 8521 7588 8555
rect 7529 8509 7588 8521
rect 9091 8690 9148 8694
rect 9091 8630 9095 8690
rect 9095 8630 9144 8690
rect 9144 8630 9148 8690
rect 9091 8626 9148 8630
rect 9091 8574 9148 8578
rect 9091 8514 9095 8574
rect 9095 8514 9144 8574
rect 9144 8514 9148 8574
rect 9091 8510 9148 8514
rect 7170 8401 7238 8406
rect 7170 8346 7174 8401
rect 7174 8346 7234 8401
rect 7234 8346 7238 8401
rect 7170 8341 7238 8346
rect 9091 8406 9148 8410
rect 9091 8346 9095 8406
rect 9095 8346 9144 8406
rect 9144 8346 9148 8406
rect 9091 8342 9148 8346
rect 7364 7368 7368 7414
rect 7368 7368 7426 7414
rect 7426 7368 7430 7414
rect 7364 7362 7430 7368
rect 9335 8689 9406 8693
rect 9335 8634 9339 8689
rect 9339 8634 9399 8689
rect 9399 8634 9406 8689
rect 9335 8630 9406 8634
rect 10420 8690 10490 8693
rect 10420 8635 10424 8690
rect 10424 8635 10484 8690
rect 10484 8635 10490 8690
rect 10420 8631 10490 8635
rect 13626 9630 13706 9636
rect 13626 9576 13630 9630
rect 13630 9576 13702 9630
rect 13702 9576 13706 9630
rect 10661 8559 10720 8573
rect 10661 8525 10674 8559
rect 10674 8525 10708 8559
rect 10708 8525 10720 8559
rect 10661 8513 10720 8525
rect 12235 8690 12292 8694
rect 12235 8630 12239 8690
rect 12239 8630 12288 8690
rect 12288 8630 12292 8690
rect 12235 8626 12292 8630
rect 12235 8574 12292 8578
rect 12235 8514 12239 8574
rect 12239 8514 12288 8574
rect 12288 8514 12292 8574
rect 12235 8510 12292 8514
rect 10302 8405 10370 8410
rect 10302 8350 10306 8405
rect 10306 8350 10366 8405
rect 10366 8350 10370 8405
rect 10302 8345 10370 8350
rect 12235 8406 12292 8410
rect 12235 8346 12239 8406
rect 12239 8346 12288 8406
rect 12288 8346 12292 8406
rect 12235 8342 12292 8346
rect 10496 7372 10500 7418
rect 10500 7372 10558 7418
rect 10558 7372 10562 7418
rect 10496 7366 10562 7372
rect 12479 8689 12550 8693
rect 12479 8634 12483 8689
rect 12483 8634 12543 8689
rect 12543 8634 12550 8689
rect 12479 8630 12550 8634
rect 13564 8690 13634 8693
rect 13564 8635 13568 8690
rect 13568 8635 13628 8690
rect 13628 8635 13634 8690
rect 13564 8631 13634 8635
rect 16828 9626 16908 9632
rect 16828 9572 16832 9626
rect 16832 9572 16904 9626
rect 16904 9572 16908 9626
rect 19972 9626 20052 9632
rect 19972 9572 19976 9626
rect 19976 9572 20048 9626
rect 20048 9572 20052 9626
rect 13805 8559 13864 8573
rect 13805 8525 13818 8559
rect 13818 8525 13852 8559
rect 13852 8525 13864 8559
rect 13805 8513 13864 8525
rect 15437 8686 15494 8690
rect 15437 8626 15441 8686
rect 15441 8626 15490 8686
rect 15490 8626 15494 8686
rect 15437 8622 15494 8626
rect 15437 8570 15494 8574
rect 15437 8510 15441 8570
rect 15441 8510 15490 8570
rect 15490 8510 15494 8570
rect 15437 8506 15494 8510
rect 13446 8405 13514 8410
rect 13446 8350 13450 8405
rect 13450 8350 13510 8405
rect 13510 8350 13514 8405
rect 13446 8345 13514 8350
rect 15437 8402 15494 8406
rect 15437 8342 15441 8402
rect 15441 8342 15490 8402
rect 15490 8342 15494 8402
rect 15437 8338 15494 8342
rect 13640 7372 13644 7418
rect 13644 7372 13702 7418
rect 13702 7372 13706 7418
rect 13640 7366 13706 7372
rect 15681 8685 15752 8689
rect 15681 8630 15685 8685
rect 15685 8630 15745 8685
rect 15745 8630 15752 8685
rect 15681 8626 15752 8630
rect 16766 8686 16836 8689
rect 16766 8631 16770 8686
rect 16770 8631 16830 8686
rect 16830 8631 16836 8686
rect 16766 8627 16836 8631
rect 17007 8555 17066 8569
rect 17007 8521 17020 8555
rect 17020 8521 17054 8555
rect 17054 8521 17066 8555
rect 17007 8509 17066 8521
rect 16648 8401 16716 8406
rect 16648 8346 16652 8401
rect 16652 8346 16712 8401
rect 16712 8346 16716 8401
rect 16648 8341 16716 8346
rect 18581 8686 18638 8690
rect 18581 8626 18585 8686
rect 18585 8626 18634 8686
rect 18634 8626 18638 8686
rect 18581 8622 18638 8626
rect 18581 8570 18638 8574
rect 18581 8510 18585 8570
rect 18585 8510 18634 8570
rect 18634 8510 18638 8570
rect 18581 8506 18638 8510
rect 18581 8402 18638 8406
rect 18581 8342 18585 8402
rect 18585 8342 18634 8402
rect 18634 8342 18638 8402
rect 18581 8338 18638 8342
rect 16842 7368 16846 7414
rect 16846 7368 16904 7414
rect 16904 7368 16908 7414
rect 16842 7362 16908 7368
rect 18825 8685 18896 8689
rect 18825 8630 18829 8685
rect 18829 8630 18889 8685
rect 18889 8630 18896 8685
rect 18825 8626 18896 8630
rect 19910 8686 19980 8689
rect 19910 8631 19914 8686
rect 19914 8631 19974 8686
rect 19974 8631 19980 8686
rect 19910 8627 19980 8631
rect 21967 11421 22038 11425
rect 21967 11366 21971 11421
rect 21971 11366 22031 11421
rect 22031 11366 22038 11421
rect 21967 11362 22038 11366
rect 23052 11422 23122 11425
rect 23052 11367 23056 11422
rect 23056 11367 23116 11422
rect 23116 11367 23122 11422
rect 23052 11363 23122 11367
rect 23293 11291 23352 11305
rect 23293 11257 23306 11291
rect 23306 11257 23340 11291
rect 23340 11257 23352 11291
rect 23293 11245 23352 11257
rect 26258 12362 26338 12368
rect 26258 12308 26262 12362
rect 26262 12308 26334 12362
rect 26334 12308 26338 12362
rect 24867 11306 24924 11310
rect 24867 11246 24871 11306
rect 24871 11246 24920 11306
rect 24920 11246 24924 11306
rect 24867 11242 24924 11246
rect 22934 11137 23002 11142
rect 22934 11082 22938 11137
rect 22938 11082 22998 11137
rect 22998 11082 23002 11137
rect 22934 11077 23002 11082
rect 24525 10859 24596 10930
rect 24867 11138 24924 11142
rect 24867 11078 24871 11138
rect 24871 11078 24920 11138
rect 24920 11078 24924 11138
rect 24867 11074 24924 11078
rect 23128 10104 23132 10150
rect 23132 10104 23190 10150
rect 23190 10104 23194 10150
rect 23128 10098 23194 10104
rect 25111 11421 25182 11425
rect 25111 11366 25115 11421
rect 25115 11366 25175 11421
rect 25175 11366 25182 11421
rect 25111 11362 25182 11366
rect 26196 11422 26266 11425
rect 26196 11367 26200 11422
rect 26200 11367 26260 11422
rect 26260 11367 26266 11422
rect 26196 11363 26266 11367
rect 26437 11291 26496 11305
rect 26437 11257 26450 11291
rect 26450 11257 26484 11291
rect 26484 11257 26496 11291
rect 26437 11245 26496 11257
rect 26078 11137 26146 11142
rect 26078 11082 26082 11137
rect 26082 11082 26142 11137
rect 26142 11082 26146 11137
rect 26078 11077 26146 11082
rect 27915 10867 27974 10937
rect 27914 10682 27975 10745
rect 27913 10459 27975 10525
rect 27913 10271 27976 10329
rect 26272 10104 26276 10150
rect 26276 10104 26334 10150
rect 26334 10104 26338 10150
rect 26272 10098 26338 10104
rect 27912 9925 27976 9986
rect 23104 9630 23184 9636
rect 23104 9576 23108 9630
rect 23108 9576 23180 9630
rect 23180 9576 23184 9630
rect 20151 8555 20210 8569
rect 20151 8521 20164 8555
rect 20164 8521 20198 8555
rect 20198 8521 20210 8555
rect 20151 8509 20210 8521
rect 21713 8690 21770 8694
rect 21713 8630 21717 8690
rect 21717 8630 21766 8690
rect 21766 8630 21770 8690
rect 21713 8626 21770 8630
rect 21713 8574 21770 8578
rect 21713 8514 21717 8574
rect 21717 8514 21766 8574
rect 21766 8514 21770 8574
rect 21713 8510 21770 8514
rect 19792 8401 19860 8406
rect 19792 8346 19796 8401
rect 19796 8346 19856 8401
rect 19856 8346 19860 8401
rect 19792 8341 19860 8346
rect 21713 8406 21770 8410
rect 21713 8346 21717 8406
rect 21717 8346 21766 8406
rect 21766 8346 21770 8406
rect 21713 8342 21770 8346
rect 19986 7368 19990 7414
rect 19990 7368 20048 7414
rect 20048 7368 20052 7414
rect 19986 7362 20052 7368
rect 21957 8689 22028 8693
rect 21957 8634 21961 8689
rect 21961 8634 22021 8689
rect 22021 8634 22028 8689
rect 21957 8630 22028 8634
rect 23042 8690 23112 8693
rect 23042 8635 23046 8690
rect 23046 8635 23106 8690
rect 23106 8635 23112 8690
rect 23042 8631 23112 8635
rect 26248 9630 26328 9636
rect 26248 9576 26252 9630
rect 26252 9576 26324 9630
rect 26324 9576 26328 9630
rect 27914 9754 27978 9814
rect 27913 9399 27980 9460
rect 23283 8559 23342 8573
rect 23283 8525 23296 8559
rect 23296 8525 23330 8559
rect 23330 8525 23342 8559
rect 23283 8513 23342 8525
rect 24857 8690 24914 8694
rect 24857 8630 24861 8690
rect 24861 8630 24910 8690
rect 24910 8630 24914 8690
rect 24857 8626 24914 8630
rect 24857 8574 24914 8578
rect 24857 8514 24861 8574
rect 24861 8514 24910 8574
rect 24910 8514 24914 8574
rect 24857 8510 24914 8514
rect 22924 8405 22992 8410
rect 22924 8350 22928 8405
rect 22928 8350 22988 8405
rect 22988 8350 22992 8405
rect 22924 8345 22992 8350
rect 24857 8406 24914 8410
rect 24857 8346 24861 8406
rect 24861 8346 24910 8406
rect 24910 8346 24914 8406
rect 24857 8342 24914 8346
rect 23118 7372 23122 7418
rect 23122 7372 23180 7418
rect 23180 7372 23184 7418
rect 23118 7366 23184 7372
rect 19585 6733 19661 6753
rect 3522 6686 3576 6694
rect 3522 6648 3532 6686
rect 3532 6648 3570 6686
rect 3570 6648 3576 6686
rect 5590 6688 5644 6696
rect 3522 6640 3576 6648
rect 5590 6650 5600 6688
rect 5600 6650 5638 6688
rect 5638 6650 5644 6688
rect 5590 6642 5644 6650
rect 7659 6686 7713 6694
rect 7659 6648 7669 6686
rect 7669 6648 7707 6686
rect 7707 6648 7713 6686
rect 9727 6688 9781 6696
rect 7659 6640 7713 6648
rect 9727 6650 9737 6688
rect 9737 6650 9775 6688
rect 9775 6650 9781 6688
rect 11796 6688 11850 6696
rect 9727 6642 9781 6650
rect 11796 6650 11806 6688
rect 11806 6650 11844 6688
rect 11844 6650 11850 6688
rect 13864 6690 13918 6698
rect 11796 6642 11850 6650
rect 13864 6652 13874 6690
rect 13874 6652 13912 6690
rect 13912 6652 13918 6690
rect 13864 6644 13918 6652
rect 15933 6688 15987 6696
rect 15933 6650 15943 6688
rect 15943 6650 15981 6688
rect 15981 6650 15987 6688
rect 18001 6690 18055 6698
rect 15933 6642 15987 6650
rect 18001 6652 18011 6690
rect 18011 6652 18049 6690
rect 18049 6652 18055 6690
rect 19585 6697 19661 6733
rect 19585 6679 19661 6697
rect 18001 6644 18055 6652
rect 2005 5841 2069 5901
rect 2428 5832 2488 5885
rect 2714 5826 2780 5892
rect 2699 5696 2770 5704
rect 2428 5635 2480 5693
rect 2699 5636 2702 5696
rect 2702 5636 2768 5696
rect 2768 5636 2770 5696
rect 2699 5627 2770 5636
rect 4102 5832 4156 5886
rect 4782 5828 4848 5894
rect 3464 4464 3526 4470
rect 3464 4422 3470 4464
rect 3470 4422 3520 4464
rect 3520 4422 3526 4464
rect 3464 4412 3526 4422
rect 6170 5834 6224 5888
rect 20323 6731 20399 6751
rect 20323 6695 20399 6731
rect 20323 6677 20399 6695
rect 21061 6731 21137 6751
rect 21061 6695 21137 6731
rect 21061 6677 21137 6695
rect 21803 6731 21879 6751
rect 21803 6695 21879 6731
rect 21803 6677 21879 6695
rect 22543 6731 22619 6751
rect 22543 6695 22619 6731
rect 22543 6677 22619 6695
rect 23281 6731 23357 6751
rect 23281 6695 23357 6731
rect 23281 6677 23357 6695
rect 24019 6731 24095 6751
rect 24019 6695 24095 6731
rect 24019 6677 24095 6695
rect 6851 5826 6917 5892
rect 5532 4466 5594 4472
rect 5532 4424 5538 4466
rect 5538 4424 5588 4466
rect 5588 4424 5594 4466
rect 5532 4414 5594 4424
rect 8239 5832 8293 5886
rect 8919 5828 8985 5894
rect 7601 4464 7663 4470
rect 7601 4422 7607 4464
rect 7607 4422 7657 4464
rect 7657 4422 7663 4464
rect 7601 4412 7663 4422
rect 10307 5834 10361 5888
rect 10988 5828 11054 5894
rect 9669 4466 9731 4472
rect 9669 4424 9675 4466
rect 9675 4424 9725 4466
rect 9725 4424 9731 4466
rect 9669 4414 9731 4424
rect 12376 5834 12430 5888
rect 13056 5830 13122 5896
rect 11738 4466 11800 4472
rect 11738 4424 11744 4466
rect 11744 4424 11794 4466
rect 11794 4424 11800 4466
rect 11738 4414 11800 4424
rect 14444 5836 14498 5890
rect 15125 5828 15191 5894
rect 13806 4468 13868 4474
rect 13806 4426 13812 4468
rect 13812 4426 13862 4468
rect 13862 4426 13868 4468
rect 13806 4416 13868 4426
rect 16513 5834 16567 5888
rect 17193 5830 17259 5896
rect 15875 4466 15937 4472
rect 15875 4424 15881 4466
rect 15881 4424 15931 4466
rect 15931 4424 15937 4466
rect 15875 4414 15937 4424
rect 18581 5836 18635 5890
rect 25101 8689 25172 8693
rect 25101 8634 25105 8689
rect 25105 8634 25165 8689
rect 25165 8634 25172 8689
rect 25101 8630 25172 8634
rect 26186 8690 26256 8693
rect 26186 8635 26190 8690
rect 26190 8635 26250 8690
rect 26250 8635 26256 8690
rect 26186 8631 26256 8635
rect 26427 8559 26486 8573
rect 26427 8525 26440 8559
rect 26440 8525 26474 8559
rect 26474 8525 26486 8559
rect 26427 8513 26486 8525
rect 26068 8405 26136 8410
rect 26068 8350 26072 8405
rect 26072 8350 26132 8405
rect 26132 8350 26136 8405
rect 26068 8345 26136 8350
rect 26262 7372 26266 7418
rect 26266 7372 26324 7418
rect 26324 7372 26328 7418
rect 26262 7366 26328 7372
rect 24757 6731 24833 6751
rect 24757 6695 24833 6731
rect 24757 6677 24833 6695
rect 19509 5865 19611 5871
rect 19509 5811 19521 5865
rect 19521 5811 19599 5865
rect 19599 5811 19611 5865
rect 19509 5805 19611 5811
rect 20247 5863 20349 5869
rect 20247 5809 20259 5863
rect 20259 5809 20337 5863
rect 20337 5809 20349 5863
rect 20247 5803 20349 5809
rect 20985 5863 21087 5869
rect 20985 5809 20997 5863
rect 20997 5809 21075 5863
rect 21075 5809 21087 5863
rect 20985 5803 21087 5809
rect 21727 5863 21829 5869
rect 21727 5809 21739 5863
rect 21739 5809 21817 5863
rect 21817 5809 21829 5863
rect 21727 5803 21829 5809
rect 22467 5863 22569 5869
rect 22467 5809 22479 5863
rect 22479 5809 22557 5863
rect 22557 5809 22569 5863
rect 22467 5803 22569 5809
rect 23205 5863 23307 5869
rect 23205 5809 23217 5863
rect 23217 5809 23295 5863
rect 23295 5809 23307 5863
rect 23205 5803 23307 5809
rect 23943 5863 24045 5869
rect 23943 5809 23955 5863
rect 23955 5809 24033 5863
rect 24033 5809 24045 5863
rect 23943 5803 24045 5809
rect 24681 5863 24783 5869
rect 24681 5809 24693 5863
rect 24693 5809 24771 5863
rect 24771 5809 24783 5863
rect 24681 5803 24783 5809
rect 17943 4468 18005 4474
rect 17943 4426 17949 4468
rect 17949 4426 17999 4468
rect 17999 4426 18005 4468
rect 17943 4416 18005 4426
rect 1508 2378 1588 2384
rect 1508 2324 1512 2378
rect 1512 2324 1584 2378
rect 1584 2324 1588 2378
rect 4652 2378 4732 2384
rect 4652 2324 4656 2378
rect 4656 2324 4728 2378
rect 4728 2324 4732 2378
rect 7784 2382 7864 2388
rect 7784 2328 7788 2382
rect 7788 2328 7860 2382
rect 7860 2328 7864 2382
rect 10928 2382 11008 2388
rect 10928 2328 10932 2382
rect 10932 2328 11004 2382
rect 11004 2328 11008 2382
rect 14130 2378 14210 2384
rect 14130 2324 14134 2378
rect 14134 2324 14206 2378
rect 14206 2324 14210 2378
rect 17274 2378 17354 2384
rect 17274 2324 17278 2378
rect 17278 2324 17350 2378
rect 17350 2324 17354 2378
rect 20406 2382 20486 2388
rect 20406 2328 20410 2382
rect 20410 2328 20482 2382
rect 20482 2328 20486 2382
rect 23550 2382 23630 2388
rect 23550 2328 23554 2382
rect 23554 2328 23626 2382
rect 23626 2328 23630 2382
rect 117 1438 174 1442
rect 117 1378 121 1438
rect 121 1378 170 1438
rect 170 1378 174 1438
rect 117 1374 174 1378
rect 117 1322 174 1326
rect 117 1262 121 1322
rect 121 1262 170 1322
rect 170 1262 174 1322
rect 117 1258 174 1262
rect 117 1154 174 1158
rect 117 1094 121 1154
rect 121 1094 170 1154
rect 170 1094 174 1154
rect 117 1090 174 1094
rect 361 1437 432 1441
rect 361 1382 365 1437
rect 365 1382 425 1437
rect 425 1382 432 1437
rect 361 1378 432 1382
rect 1446 1438 1516 1441
rect 1446 1383 1450 1438
rect 1450 1383 1510 1438
rect 1510 1383 1516 1438
rect 1446 1379 1516 1383
rect 1687 1307 1746 1321
rect 1687 1273 1700 1307
rect 1700 1273 1734 1307
rect 1734 1273 1746 1307
rect 1687 1261 1746 1273
rect 3261 1438 3318 1442
rect 3261 1378 3265 1438
rect 3265 1378 3314 1438
rect 3314 1378 3318 1438
rect 3261 1374 3318 1378
rect 3261 1322 3318 1326
rect 3261 1262 3265 1322
rect 3265 1262 3314 1322
rect 3314 1262 3318 1322
rect 3261 1258 3318 1262
rect 1328 1153 1396 1158
rect 1328 1098 1332 1153
rect 1332 1098 1392 1153
rect 1392 1098 1396 1153
rect 1328 1093 1396 1098
rect 3261 1154 3318 1158
rect 3261 1094 3265 1154
rect 3265 1094 3314 1154
rect 3314 1094 3318 1154
rect 3261 1090 3318 1094
rect 3505 1437 3576 1441
rect 3505 1382 3509 1437
rect 3509 1382 3569 1437
rect 3569 1382 3576 1437
rect 3505 1378 3576 1382
rect 4590 1438 4660 1441
rect 4590 1383 4594 1438
rect 4594 1383 4654 1438
rect 4654 1383 4660 1438
rect 4590 1379 4660 1383
rect 4831 1307 4890 1321
rect 4831 1273 4844 1307
rect 4844 1273 4878 1307
rect 4878 1273 4890 1307
rect 4831 1261 4890 1273
rect 6393 1442 6450 1446
rect 6393 1382 6397 1442
rect 6397 1382 6446 1442
rect 6446 1382 6450 1442
rect 6393 1378 6450 1382
rect 6393 1326 6450 1330
rect 6393 1266 6397 1326
rect 6397 1266 6446 1326
rect 6446 1266 6450 1326
rect 6393 1262 6450 1266
rect 4472 1153 4540 1158
rect 4472 1098 4476 1153
rect 4476 1098 4536 1153
rect 4536 1098 4540 1153
rect 4472 1093 4540 1098
rect 6393 1158 6450 1162
rect 6393 1098 6397 1158
rect 6397 1098 6446 1158
rect 6446 1098 6450 1158
rect 6393 1094 6450 1098
rect 6637 1441 6708 1445
rect 6637 1386 6641 1441
rect 6641 1386 6701 1441
rect 6701 1386 6708 1441
rect 6637 1382 6708 1386
rect 7722 1442 7792 1445
rect 7722 1387 7726 1442
rect 7726 1387 7786 1442
rect 7786 1387 7792 1442
rect 7722 1383 7792 1387
rect 7963 1311 8022 1325
rect 7963 1277 7976 1311
rect 7976 1277 8010 1311
rect 8010 1277 8022 1311
rect 7963 1265 8022 1277
rect 9537 1442 9594 1446
rect 9537 1382 9541 1442
rect 9541 1382 9590 1442
rect 9590 1382 9594 1442
rect 9537 1378 9594 1382
rect 9537 1326 9594 1330
rect 9537 1266 9541 1326
rect 9541 1266 9590 1326
rect 9590 1266 9594 1326
rect 9537 1262 9594 1266
rect 7604 1157 7672 1162
rect 7604 1102 7608 1157
rect 7608 1102 7668 1157
rect 7668 1102 7672 1157
rect 7604 1097 7672 1102
rect 9537 1158 9594 1162
rect 9537 1098 9541 1158
rect 9541 1098 9590 1158
rect 9590 1098 9594 1158
rect 9537 1094 9594 1098
rect 9781 1441 9852 1445
rect 9781 1386 9785 1441
rect 9785 1386 9845 1441
rect 9845 1386 9852 1441
rect 9781 1382 9852 1386
rect 10866 1442 10936 1445
rect 10866 1387 10870 1442
rect 10870 1387 10930 1442
rect 10930 1387 10936 1442
rect 10866 1383 10936 1387
rect 11107 1311 11166 1325
rect 11107 1277 11120 1311
rect 11120 1277 11154 1311
rect 11154 1277 11166 1311
rect 11107 1265 11166 1277
rect 12739 1438 12796 1442
rect 12739 1378 12743 1438
rect 12743 1378 12792 1438
rect 12792 1378 12796 1438
rect 12739 1374 12796 1378
rect 12739 1322 12796 1326
rect 12739 1262 12743 1322
rect 12743 1262 12792 1322
rect 12792 1262 12796 1322
rect 12739 1258 12796 1262
rect 10748 1157 10816 1162
rect 10748 1102 10752 1157
rect 10752 1102 10812 1157
rect 10812 1102 10816 1157
rect 10748 1097 10816 1102
rect 12739 1154 12796 1158
rect 12739 1094 12743 1154
rect 12743 1094 12792 1154
rect 12792 1094 12796 1154
rect 12739 1090 12796 1094
rect 12983 1437 13054 1441
rect 12983 1382 12987 1437
rect 12987 1382 13047 1437
rect 13047 1382 13054 1437
rect 12983 1378 13054 1382
rect 14068 1438 14138 1441
rect 14068 1383 14072 1438
rect 14072 1383 14132 1438
rect 14132 1383 14138 1438
rect 14068 1379 14138 1383
rect 14309 1307 14368 1321
rect 14309 1273 14322 1307
rect 14322 1273 14356 1307
rect 14356 1273 14368 1307
rect 14309 1261 14368 1273
rect 15883 1438 15940 1442
rect 15883 1378 15887 1438
rect 15887 1378 15936 1438
rect 15936 1378 15940 1438
rect 15883 1374 15940 1378
rect 15883 1322 15940 1326
rect 15883 1262 15887 1322
rect 15887 1262 15936 1322
rect 15936 1262 15940 1322
rect 15883 1258 15940 1262
rect 13950 1153 14018 1158
rect 13950 1098 13954 1153
rect 13954 1098 14014 1153
rect 14014 1098 14018 1153
rect 13950 1093 14018 1098
rect 15883 1154 15940 1158
rect 15883 1094 15887 1154
rect 15887 1094 15936 1154
rect 15936 1094 15940 1154
rect 15883 1090 15940 1094
rect 16127 1437 16198 1441
rect 16127 1382 16131 1437
rect 16131 1382 16191 1437
rect 16191 1382 16198 1437
rect 16127 1378 16198 1382
rect 17212 1438 17282 1441
rect 17212 1383 17216 1438
rect 17216 1383 17276 1438
rect 17276 1383 17282 1438
rect 17212 1379 17282 1383
rect 17453 1307 17512 1321
rect 17453 1273 17466 1307
rect 17466 1273 17500 1307
rect 17500 1273 17512 1307
rect 17453 1261 17512 1273
rect 19015 1442 19072 1446
rect 19015 1382 19019 1442
rect 19019 1382 19068 1442
rect 19068 1382 19072 1442
rect 19015 1378 19072 1382
rect 19015 1326 19072 1330
rect 19015 1266 19019 1326
rect 19019 1266 19068 1326
rect 19068 1266 19072 1326
rect 19015 1262 19072 1266
rect 17094 1153 17162 1158
rect 17094 1098 17098 1153
rect 17098 1098 17158 1153
rect 17158 1098 17162 1153
rect 17094 1093 17162 1098
rect 19015 1158 19072 1162
rect 19015 1098 19019 1158
rect 19019 1098 19068 1158
rect 19068 1098 19072 1158
rect 19015 1094 19072 1098
rect 19259 1441 19330 1445
rect 19259 1386 19263 1441
rect 19263 1386 19323 1441
rect 19323 1386 19330 1441
rect 19259 1382 19330 1386
rect 20344 1442 20414 1445
rect 20344 1387 20348 1442
rect 20348 1387 20408 1442
rect 20408 1387 20414 1442
rect 20344 1383 20414 1387
rect 20585 1311 20644 1325
rect 20585 1277 20598 1311
rect 20598 1277 20632 1311
rect 20632 1277 20644 1311
rect 20585 1265 20644 1277
rect 22159 1442 22216 1446
rect 22159 1382 22163 1442
rect 22163 1382 22212 1442
rect 22212 1382 22216 1442
rect 22159 1378 22216 1382
rect 22159 1326 22216 1330
rect 22159 1266 22163 1326
rect 22163 1266 22212 1326
rect 22212 1266 22216 1326
rect 22159 1262 22216 1266
rect 20226 1157 20294 1162
rect 20226 1102 20230 1157
rect 20230 1102 20290 1157
rect 20290 1102 20294 1157
rect 20226 1097 20294 1102
rect 22159 1158 22216 1162
rect 22159 1098 22163 1158
rect 22163 1098 22212 1158
rect 22212 1098 22216 1158
rect 22159 1094 22216 1098
rect 22403 1441 22474 1445
rect 22403 1386 22407 1441
rect 22407 1386 22467 1441
rect 22467 1386 22474 1441
rect 22403 1382 22474 1386
rect 23488 1442 23558 1445
rect 23488 1387 23492 1442
rect 23492 1387 23552 1442
rect 23552 1387 23558 1442
rect 23488 1383 23558 1387
rect 23729 1311 23788 1325
rect 23729 1277 23742 1311
rect 23742 1277 23776 1311
rect 23776 1277 23788 1311
rect 23729 1265 23788 1277
rect 23370 1157 23438 1162
rect 23370 1102 23374 1157
rect 23374 1102 23434 1157
rect 23434 1102 23438 1157
rect 23370 1097 23438 1102
rect 1522 120 1526 166
rect 1526 120 1584 166
rect 1584 120 1588 166
rect 1522 114 1588 120
rect 4666 120 4670 166
rect 4670 120 4728 166
rect 4728 120 4732 166
rect 4666 114 4732 120
rect 7798 124 7802 170
rect 7802 124 7860 170
rect 7860 124 7864 170
rect 7798 118 7864 124
rect 10942 124 10946 170
rect 10946 124 11004 170
rect 11004 124 11008 170
rect 10942 118 11008 124
rect 14144 120 14148 166
rect 14148 120 14206 166
rect 14206 120 14210 166
rect 14144 114 14210 120
rect 17288 120 17292 166
rect 17292 120 17350 166
rect 17350 120 17354 166
rect 17288 114 17354 120
rect 20420 124 20424 170
rect 20424 124 20482 170
rect 20482 124 20486 170
rect 20420 118 20486 124
rect 23564 124 23568 170
rect 23568 124 23626 170
rect 23626 124 23630 170
rect 23564 118 23630 124
rect 1540 -1514 1620 -1508
rect 1540 -1568 1544 -1514
rect 1544 -1568 1616 -1514
rect 1616 -1568 1620 -1514
rect 4684 -1514 4764 -1508
rect 4684 -1568 4688 -1514
rect 4688 -1568 4760 -1514
rect 4760 -1568 4764 -1514
rect 7816 -1510 7896 -1504
rect 7816 -1564 7820 -1510
rect 7820 -1564 7892 -1510
rect 7892 -1564 7896 -1510
rect 10960 -1510 11040 -1504
rect 10960 -1564 10964 -1510
rect 10964 -1564 11036 -1510
rect 11036 -1564 11040 -1510
rect 14162 -1514 14242 -1508
rect 14162 -1568 14166 -1514
rect 14166 -1568 14238 -1514
rect 14238 -1568 14242 -1514
rect 17306 -1514 17386 -1508
rect 17306 -1568 17310 -1514
rect 17310 -1568 17382 -1514
rect 17382 -1568 17386 -1514
rect 20438 -1510 20518 -1504
rect 20438 -1564 20442 -1510
rect 20442 -1564 20514 -1510
rect 20514 -1564 20518 -1510
rect 23582 -1510 23662 -1504
rect 23582 -1564 23586 -1510
rect 23586 -1564 23658 -1510
rect 23658 -1564 23662 -1510
rect 149 -2454 206 -2450
rect 149 -2514 153 -2454
rect 153 -2514 202 -2454
rect 202 -2514 206 -2454
rect 149 -2518 206 -2514
rect 149 -2570 206 -2566
rect 149 -2630 153 -2570
rect 153 -2630 202 -2570
rect 202 -2630 206 -2570
rect 149 -2634 206 -2630
rect 149 -2738 206 -2734
rect 149 -2798 153 -2738
rect 153 -2798 202 -2738
rect 202 -2798 206 -2738
rect 149 -2802 206 -2798
rect 393 -2455 464 -2451
rect 393 -2510 397 -2455
rect 397 -2510 457 -2455
rect 457 -2510 464 -2455
rect 393 -2514 464 -2510
rect 1478 -2454 1548 -2451
rect 1478 -2509 1482 -2454
rect 1482 -2509 1542 -2454
rect 1542 -2509 1548 -2454
rect 1478 -2513 1548 -2509
rect 1719 -2585 1778 -2571
rect 1719 -2619 1732 -2585
rect 1732 -2619 1766 -2585
rect 1766 -2619 1778 -2585
rect 1719 -2631 1778 -2619
rect 3293 -2454 3350 -2450
rect 3293 -2514 3297 -2454
rect 3297 -2514 3346 -2454
rect 3346 -2514 3350 -2454
rect 3293 -2518 3350 -2514
rect 3293 -2570 3350 -2566
rect 3293 -2630 3297 -2570
rect 3297 -2630 3346 -2570
rect 3346 -2630 3350 -2570
rect 3293 -2634 3350 -2630
rect 1360 -2739 1428 -2734
rect 1360 -2794 1364 -2739
rect 1364 -2794 1424 -2739
rect 1424 -2794 1428 -2739
rect 1360 -2799 1428 -2794
rect 3293 -2738 3350 -2734
rect 3293 -2798 3297 -2738
rect 3297 -2798 3346 -2738
rect 3346 -2798 3350 -2738
rect 3293 -2802 3350 -2798
rect 3537 -2455 3608 -2451
rect 3537 -2510 3541 -2455
rect 3541 -2510 3601 -2455
rect 3601 -2510 3608 -2455
rect 3537 -2514 3608 -2510
rect 4622 -2454 4692 -2451
rect 4622 -2509 4626 -2454
rect 4626 -2509 4686 -2454
rect 4686 -2509 4692 -2454
rect 4622 -2513 4692 -2509
rect 4863 -2585 4922 -2571
rect 4863 -2619 4876 -2585
rect 4876 -2619 4910 -2585
rect 4910 -2619 4922 -2585
rect 4863 -2631 4922 -2619
rect 6425 -2450 6482 -2446
rect 6425 -2510 6429 -2450
rect 6429 -2510 6478 -2450
rect 6478 -2510 6482 -2450
rect 6425 -2514 6482 -2510
rect 6425 -2566 6482 -2562
rect 6425 -2626 6429 -2566
rect 6429 -2626 6478 -2566
rect 6478 -2626 6482 -2566
rect 6425 -2630 6482 -2626
rect 4504 -2739 4572 -2734
rect 4504 -2794 4508 -2739
rect 4508 -2794 4568 -2739
rect 4568 -2794 4572 -2739
rect 4504 -2799 4572 -2794
rect 6425 -2734 6482 -2730
rect 6425 -2794 6429 -2734
rect 6429 -2794 6478 -2734
rect 6478 -2794 6482 -2734
rect 6425 -2798 6482 -2794
rect 6669 -2451 6740 -2447
rect 6669 -2506 6673 -2451
rect 6673 -2506 6733 -2451
rect 6733 -2506 6740 -2451
rect 6669 -2510 6740 -2506
rect 7754 -2450 7824 -2447
rect 7754 -2505 7758 -2450
rect 7758 -2505 7818 -2450
rect 7818 -2505 7824 -2450
rect 7754 -2509 7824 -2505
rect 7995 -2581 8054 -2567
rect 7995 -2615 8008 -2581
rect 8008 -2615 8042 -2581
rect 8042 -2615 8054 -2581
rect 7995 -2627 8054 -2615
rect 9569 -2450 9626 -2446
rect 9569 -2510 9573 -2450
rect 9573 -2510 9622 -2450
rect 9622 -2510 9626 -2450
rect 9569 -2514 9626 -2510
rect 9569 -2566 9626 -2562
rect 9569 -2626 9573 -2566
rect 9573 -2626 9622 -2566
rect 9622 -2626 9626 -2566
rect 9569 -2630 9626 -2626
rect 7636 -2735 7704 -2730
rect 7636 -2790 7640 -2735
rect 7640 -2790 7700 -2735
rect 7700 -2790 7704 -2735
rect 7636 -2795 7704 -2790
rect 9569 -2734 9626 -2730
rect 9569 -2794 9573 -2734
rect 9573 -2794 9622 -2734
rect 9622 -2794 9626 -2734
rect 9569 -2798 9626 -2794
rect 9813 -2451 9884 -2447
rect 9813 -2506 9817 -2451
rect 9817 -2506 9877 -2451
rect 9877 -2506 9884 -2451
rect 9813 -2510 9884 -2506
rect 10898 -2450 10968 -2447
rect 10898 -2505 10902 -2450
rect 10902 -2505 10962 -2450
rect 10962 -2505 10968 -2450
rect 10898 -2509 10968 -2505
rect 11139 -2581 11198 -2567
rect 11139 -2615 11152 -2581
rect 11152 -2615 11186 -2581
rect 11186 -2615 11198 -2581
rect 11139 -2627 11198 -2615
rect 12771 -2454 12828 -2450
rect 12771 -2514 12775 -2454
rect 12775 -2514 12824 -2454
rect 12824 -2514 12828 -2454
rect 12771 -2518 12828 -2514
rect 12771 -2570 12828 -2566
rect 12771 -2630 12775 -2570
rect 12775 -2630 12824 -2570
rect 12824 -2630 12828 -2570
rect 12771 -2634 12828 -2630
rect 10780 -2735 10848 -2730
rect 10780 -2790 10784 -2735
rect 10784 -2790 10844 -2735
rect 10844 -2790 10848 -2735
rect 10780 -2795 10848 -2790
rect 12771 -2738 12828 -2734
rect 12771 -2798 12775 -2738
rect 12775 -2798 12824 -2738
rect 12824 -2798 12828 -2738
rect 12771 -2802 12828 -2798
rect 13015 -2455 13086 -2451
rect 13015 -2510 13019 -2455
rect 13019 -2510 13079 -2455
rect 13079 -2510 13086 -2455
rect 13015 -2514 13086 -2510
rect 14100 -2454 14170 -2451
rect 14100 -2509 14104 -2454
rect 14104 -2509 14164 -2454
rect 14164 -2509 14170 -2454
rect 14100 -2513 14170 -2509
rect 14341 -2585 14400 -2571
rect 14341 -2619 14354 -2585
rect 14354 -2619 14388 -2585
rect 14388 -2619 14400 -2585
rect 14341 -2631 14400 -2619
rect 15915 -2454 15972 -2450
rect 15915 -2514 15919 -2454
rect 15919 -2514 15968 -2454
rect 15968 -2514 15972 -2454
rect 15915 -2518 15972 -2514
rect 15915 -2570 15972 -2566
rect 15915 -2630 15919 -2570
rect 15919 -2630 15968 -2570
rect 15968 -2630 15972 -2570
rect 15915 -2634 15972 -2630
rect 13982 -2739 14050 -2734
rect 13982 -2794 13986 -2739
rect 13986 -2794 14046 -2739
rect 14046 -2794 14050 -2739
rect 13982 -2799 14050 -2794
rect 15915 -2738 15972 -2734
rect 15915 -2798 15919 -2738
rect 15919 -2798 15968 -2738
rect 15968 -2798 15972 -2738
rect 15915 -2802 15972 -2798
rect 16159 -2455 16230 -2451
rect 16159 -2510 16163 -2455
rect 16163 -2510 16223 -2455
rect 16223 -2510 16230 -2455
rect 16159 -2514 16230 -2510
rect 17244 -2454 17314 -2451
rect 17244 -2509 17248 -2454
rect 17248 -2509 17308 -2454
rect 17308 -2509 17314 -2454
rect 17244 -2513 17314 -2509
rect 17485 -2585 17544 -2571
rect 17485 -2619 17498 -2585
rect 17498 -2619 17532 -2585
rect 17532 -2619 17544 -2585
rect 17485 -2631 17544 -2619
rect 19047 -2450 19104 -2446
rect 19047 -2510 19051 -2450
rect 19051 -2510 19100 -2450
rect 19100 -2510 19104 -2450
rect 19047 -2514 19104 -2510
rect 19047 -2566 19104 -2562
rect 19047 -2626 19051 -2566
rect 19051 -2626 19100 -2566
rect 19100 -2626 19104 -2566
rect 19047 -2630 19104 -2626
rect 17126 -2739 17194 -2734
rect 17126 -2794 17130 -2739
rect 17130 -2794 17190 -2739
rect 17190 -2794 17194 -2739
rect 17126 -2799 17194 -2794
rect 19047 -2734 19104 -2730
rect 19047 -2794 19051 -2734
rect 19051 -2794 19100 -2734
rect 19100 -2794 19104 -2734
rect 19047 -2798 19104 -2794
rect 19291 -2451 19362 -2447
rect 19291 -2506 19295 -2451
rect 19295 -2506 19355 -2451
rect 19355 -2506 19362 -2451
rect 19291 -2510 19362 -2506
rect 20376 -2450 20446 -2447
rect 20376 -2505 20380 -2450
rect 20380 -2505 20440 -2450
rect 20440 -2505 20446 -2450
rect 20376 -2509 20446 -2505
rect 20617 -2581 20676 -2567
rect 20617 -2615 20630 -2581
rect 20630 -2615 20664 -2581
rect 20664 -2615 20676 -2581
rect 20617 -2627 20676 -2615
rect 22191 -2450 22248 -2446
rect 22191 -2510 22195 -2450
rect 22195 -2510 22244 -2450
rect 22244 -2510 22248 -2450
rect 22191 -2514 22248 -2510
rect 22191 -2566 22248 -2562
rect 22191 -2626 22195 -2566
rect 22195 -2626 22244 -2566
rect 22244 -2626 22248 -2566
rect 22191 -2630 22248 -2626
rect 20258 -2735 20326 -2730
rect 20258 -2790 20262 -2735
rect 20262 -2790 20322 -2735
rect 20322 -2790 20326 -2735
rect 20258 -2795 20326 -2790
rect 22191 -2734 22248 -2730
rect 22191 -2794 22195 -2734
rect 22195 -2794 22244 -2734
rect 22244 -2794 22248 -2734
rect 22191 -2798 22248 -2794
rect 22435 -2451 22506 -2447
rect 22435 -2506 22439 -2451
rect 22439 -2506 22499 -2451
rect 22499 -2506 22506 -2451
rect 22435 -2510 22506 -2506
rect 23520 -2450 23590 -2447
rect 23520 -2505 23524 -2450
rect 23524 -2505 23584 -2450
rect 23584 -2505 23590 -2450
rect 23520 -2509 23590 -2505
rect 23761 -2581 23820 -2567
rect 23761 -2615 23774 -2581
rect 23774 -2615 23808 -2581
rect 23808 -2615 23820 -2581
rect 23761 -2627 23820 -2615
rect 23402 -2735 23470 -2730
rect 23402 -2790 23406 -2735
rect 23406 -2790 23466 -2735
rect 23466 -2790 23470 -2735
rect 23402 -2795 23470 -2790
rect 1554 -3772 1558 -3726
rect 1558 -3772 1616 -3726
rect 1616 -3772 1620 -3726
rect 1554 -3778 1620 -3772
rect 4698 -3772 4702 -3726
rect 4702 -3772 4760 -3726
rect 4760 -3772 4764 -3726
rect 4698 -3778 4764 -3772
rect 7830 -3768 7834 -3722
rect 7834 -3768 7892 -3722
rect 7892 -3768 7896 -3722
rect 7830 -3774 7896 -3768
rect 10974 -3768 10978 -3722
rect 10978 -3768 11036 -3722
rect 11036 -3768 11040 -3722
rect 10974 -3774 11040 -3768
rect 14176 -3772 14180 -3726
rect 14180 -3772 14238 -3726
rect 14238 -3772 14242 -3726
rect 14176 -3778 14242 -3772
rect 17320 -3772 17324 -3726
rect 17324 -3772 17382 -3726
rect 17382 -3772 17386 -3726
rect 17320 -3778 17386 -3772
rect 20452 -3768 20456 -3722
rect 20456 -3768 20514 -3722
rect 20514 -3768 20518 -3722
rect 20452 -3774 20518 -3768
rect 23596 -3768 23600 -3722
rect 23600 -3768 23658 -3722
rect 23658 -3768 23662 -3722
rect 23596 -3774 23662 -3768
<< metal2 >>
rect 1702 22264 1802 22274
rect 1702 22162 1802 22172
rect 4846 22264 4946 22274
rect 4846 22162 4946 22172
rect 7978 22268 8078 22278
rect 7978 22166 8078 22176
rect 11122 22268 11222 22278
rect 11122 22166 11222 22176
rect 14324 22264 14424 22274
rect 14324 22162 14424 22172
rect 17468 22264 17568 22274
rect 17468 22162 17568 22172
rect 20600 22268 20700 22278
rect 20600 22166 20700 22176
rect 23744 22268 23844 22278
rect 23744 22166 23844 22176
rect 324 21445 378 21453
rect 313 21443 3412 21445
rect 313 21381 324 21443
rect 378 21396 3412 21443
rect 378 21381 3352 21396
rect 313 21380 392 21381
rect 324 21371 378 21380
rect 3352 21333 3412 21343
rect 6832 21307 6925 21309
rect 9976 21307 10069 21309
rect 19454 21307 19547 21309
rect 22598 21307 22691 21309
rect 323 21303 380 21304
rect 556 21303 649 21305
rect 3700 21303 3793 21305
rect 4743 21303 11151 21307
rect 13178 21303 13271 21305
rect 16322 21303 16415 21305
rect 17406 21303 23773 21307
rect 315 21302 1731 21303
rect 3526 21302 23773 21303
rect 312 21297 23773 21302
rect 312 21294 6843 21297
rect 312 21226 323 21294
rect 380 21293 6843 21294
rect 380 21230 567 21293
rect 638 21231 1652 21293
rect 1722 21231 3711 21293
rect 638 21230 3711 21231
rect 3782 21231 4796 21293
rect 4866 21234 6843 21293
rect 6914 21235 7928 21297
rect 7998 21235 9987 21297
rect 6914 21234 9987 21235
rect 10058 21235 11072 21297
rect 11142 21293 19465 21297
rect 11142 21235 13189 21293
rect 10058 21234 13189 21235
rect 4866 21231 13189 21234
rect 3782 21230 13189 21231
rect 13260 21231 14274 21293
rect 14344 21231 16333 21293
rect 13260 21230 16333 21231
rect 16404 21231 17418 21293
rect 17488 21234 19465 21293
rect 19536 21235 20550 21297
rect 20620 21235 22609 21297
rect 19536 21234 22609 21235
rect 22680 21235 23694 21297
rect 23764 21235 23773 21297
rect 22680 21234 23773 21235
rect 17488 21231 23773 21234
rect 16404 21230 23773 21231
rect 380 21226 23773 21230
rect 312 21223 23773 21226
rect 312 21222 6666 21223
rect 312 21219 6556 21222
rect 12934 21219 19285 21223
rect 312 21218 390 21219
rect 1688 21218 3534 21219
rect 14262 21218 16156 21219
rect 323 21216 380 21218
rect 9743 21190 9800 21192
rect 3467 21186 3524 21188
rect 9732 21187 9828 21190
rect 3456 21183 3552 21186
rect 312 21173 1952 21183
rect 312 21169 1893 21173
rect 312 21113 322 21169
rect 378 21113 1893 21169
rect 312 21104 1952 21113
rect 322 21103 378 21104
rect 1893 21103 1952 21104
rect 3456 21178 5096 21183
rect 3456 21110 3467 21178
rect 3524 21173 5096 21178
rect 3524 21113 5037 21173
rect 3524 21110 5096 21113
rect 3456 21104 5096 21110
rect 3456 21101 3552 21104
rect 5037 21103 5096 21104
rect 6410 21177 8228 21187
rect 6410 21117 8169 21177
rect 6410 21108 8228 21117
rect 3467 21100 3524 21101
rect 6410 21064 6467 21108
rect 8169 21107 8228 21108
rect 9732 21182 11372 21187
rect 9732 21114 9743 21182
rect 9800 21177 11372 21182
rect 9800 21117 11313 21177
rect 9800 21114 11372 21117
rect 9732 21108 11372 21114
rect 9732 21105 9828 21108
rect 11313 21107 11372 21108
rect 12667 21173 14574 21183
rect 12667 21113 14515 21173
rect 9743 21104 9800 21105
rect 12667 21104 14574 21113
rect 16078 21178 17718 21183
rect 16078 21110 16089 21178
rect 16146 21173 17718 21178
rect 16146 21113 17659 21173
rect 16146 21110 17718 21113
rect 16078 21104 17718 21110
rect 323 21019 380 21020
rect 3467 21019 3524 21020
rect 6252 21019 6467 21064
rect 6599 21023 6656 21024
rect 9743 21023 9800 21024
rect 6588 21022 6684 21023
rect 9732 21022 9828 21023
rect 312 21018 408 21019
rect 3456 21018 3552 21019
rect 312 21010 3145 21018
rect 312 20942 323 21010
rect 380 20945 1534 21010
rect 1602 20945 3145 21010
rect 380 20942 3145 20945
rect 312 20934 3145 20942
rect 3456 21010 4757 21018
rect 3456 20942 3467 21010
rect 3524 20945 4678 21010
rect 4746 20945 4757 21010
rect 3524 20942 4757 20945
rect 3456 20934 4757 20942
rect 323 20932 380 20934
rect 3070 20893 3145 20934
rect 3467 20932 3524 20934
rect 6252 20893 6324 21019
rect 6588 21014 9366 21022
rect 6588 20946 6599 21014
rect 6656 20949 7810 21014
rect 7878 20949 9366 21014
rect 6656 20946 9366 20949
rect 6588 20938 9366 20946
rect 9732 21014 11033 21022
rect 9732 20946 9743 21014
rect 9800 20949 10954 21014
rect 11022 20949 11033 21014
rect 9800 20946 11033 20949
rect 9732 20938 11033 20946
rect 6599 20936 6656 20938
rect 3070 20828 6324 20893
rect 9287 20855 9366 20938
rect 9743 20936 9800 20938
rect 12667 20855 12757 21104
rect 14515 21103 14574 21104
rect 17659 21103 17718 21104
rect 18988 21182 20850 21187
rect 18988 21114 19221 21182
rect 19278 21177 20850 21182
rect 19278 21117 20791 21177
rect 19278 21114 20850 21117
rect 18988 21108 20850 21114
rect 22354 21182 23994 21187
rect 22354 21114 22365 21182
rect 22422 21177 23994 21182
rect 22422 21117 23935 21177
rect 22422 21114 23994 21117
rect 22354 21108 23994 21114
rect 12945 21019 13002 21020
rect 16089 21019 16146 21020
rect 12934 21018 13030 21019
rect 16078 21018 16174 21019
rect 12934 21010 14236 21018
rect 12934 20942 12945 21010
rect 13002 20945 14156 21010
rect 14224 20945 14236 21010
rect 13002 20942 14236 20945
rect 12934 20934 14236 20942
rect 16078 21010 17379 21018
rect 16078 20942 16089 21010
rect 16146 20945 17300 21010
rect 17368 20945 17379 21010
rect 16146 20942 17379 20945
rect 16078 20934 17379 20942
rect 12945 20932 13002 20934
rect 9287 20787 12757 20855
rect 14155 20877 14236 20934
rect 16089 20932 16146 20934
rect 18988 20877 19069 21108
rect 20791 21107 20850 21108
rect 23935 21107 23994 21108
rect 22354 21024 22433 21034
rect 19221 21023 19278 21024
rect 19210 21022 19306 21023
rect 19210 21014 20511 21022
rect 19210 20946 19221 21014
rect 19278 20949 20432 21014
rect 20500 20949 20511 21014
rect 19278 20946 20511 20949
rect 19210 20938 20511 20946
rect 19221 20936 19278 20938
rect 22433 21022 22450 21023
rect 22433 21014 23655 21022
rect 22433 20949 23576 21014
rect 23644 20949 23655 21014
rect 22433 20938 23655 20949
rect 22354 20925 22433 20935
rect 14155 20798 19069 20877
rect 22051 20876 25585 20877
rect 22051 20866 25620 20876
rect 22051 20858 25549 20866
rect 22104 20801 25549 20858
rect 22051 20795 25549 20801
rect 22051 20787 25620 20795
rect 25549 20785 25620 20787
rect 323 20769 377 20778
rect 3362 20772 3432 20782
rect 312 20768 3362 20769
rect 312 20706 323 20768
rect 377 20712 3362 20768
rect 3432 20712 3439 20769
rect 377 20706 3439 20712
rect 312 20705 3439 20706
rect 18906 20731 18970 20741
rect 323 20696 377 20705
rect 3362 20702 3432 20705
rect 18906 20662 18970 20672
rect 25537 20730 25603 20740
rect 25537 20660 25603 20670
rect 323 20634 377 20643
rect 6512 20634 6576 20641
rect 312 20633 6576 20634
rect 312 20571 323 20633
rect 377 20631 6576 20633
rect 377 20574 6512 20631
rect 377 20571 6576 20574
rect 312 20570 6576 20571
rect 323 20561 377 20570
rect 6512 20564 6576 20570
rect 15770 20578 15826 20588
rect 325 20522 379 20531
rect 9654 20526 9708 20536
rect 314 20521 9654 20522
rect 314 20459 325 20521
rect 379 20468 9654 20521
rect 15770 20499 15826 20509
rect 25527 20572 25591 20582
rect 25527 20493 25591 20503
rect 379 20459 9708 20468
rect 314 20458 9708 20459
rect 325 20449 379 20458
rect 12545 20427 12607 20437
rect 325 20397 379 20406
rect 314 20396 541 20397
rect 314 20334 325 20396
rect 379 20334 12421 20396
rect 12545 20349 12607 20359
rect 25527 20426 25591 20436
rect 25527 20347 25591 20357
rect 314 20333 12421 20334
rect 325 20324 379 20333
rect 12353 20298 12421 20333
rect 12824 20302 12893 20312
rect 9370 20279 9429 20289
rect 6018 20203 6465 20267
rect 12353 20241 12824 20298
rect 12353 20234 12893 20241
rect 12824 20231 12893 20234
rect 25527 20286 25591 20296
rect 9370 20212 9429 20222
rect 25527 20207 25591 20217
rect 330 20163 384 20165
rect 6018 20163 6082 20203
rect 313 20155 6082 20163
rect 313 20098 330 20155
rect 319 20093 330 20098
rect 384 20098 6082 20155
rect 6244 20162 6303 20172
rect 384 20093 395 20098
rect 319 20092 395 20093
rect 6401 20162 6465 20203
rect 15975 20167 16032 20177
rect 6401 20100 15975 20162
rect 6401 20098 16032 20100
rect 330 20083 384 20092
rect 6244 20086 6303 20096
rect 15975 20090 16032 20098
rect 25526 20147 25590 20157
rect 25526 20068 25590 20078
rect 1722 20020 1798 20030
rect 1722 19952 1798 19962
rect 4866 20020 4942 20030
rect 4866 19952 4942 19962
rect 7998 20024 8074 20034
rect 7998 19956 8074 19966
rect 11142 20024 11218 20034
rect 11142 19956 11218 19966
rect 14344 20020 14420 20030
rect 14344 19952 14420 19962
rect 17488 20020 17564 20030
rect 17488 19952 17564 19962
rect 20620 20024 20696 20034
rect 19104 19951 19174 19961
rect 20620 19956 20696 19966
rect 23764 20024 23840 20034
rect 23764 19956 23840 19966
rect 327 19934 381 19941
rect 316 19933 434 19934
rect 316 19871 327 19933
rect 381 19923 434 19933
rect 381 19871 2972 19923
rect 316 19870 2972 19871
rect 327 19861 381 19870
rect 2908 19762 2972 19870
rect 3111 19882 3184 19892
rect 3243 19875 19104 19924
rect 3243 19870 19174 19875
rect 3243 19865 3306 19870
rect 19104 19865 19174 19870
rect 25526 19879 25590 19889
rect 3111 19791 3184 19801
rect 3242 19762 3306 19865
rect 25526 19800 25590 19810
rect 2908 19734 3306 19762
rect 230 18636 290 18646
rect 290 18615 13066 18625
rect 290 18577 13012 18615
rect 230 18567 290 18577
rect 13012 18551 13066 18561
rect 227 18439 287 18446
rect 11474 18439 11528 18440
rect 227 18436 11531 18439
rect 287 18430 11531 18436
rect 287 18376 11474 18430
rect 11528 18376 11531 18430
rect 287 18374 11531 18376
rect 227 18364 287 18374
rect 220 18250 280 18256
rect 10013 18250 10067 18255
rect 220 18246 10068 18250
rect 280 18245 10068 18246
rect 280 18191 10013 18245
rect 10067 18191 10068 18245
rect 280 18184 10068 18191
rect 220 18174 280 18184
rect 220 18064 280 18074
rect 8511 18064 8565 18067
rect 280 18057 8565 18064
rect 280 18003 8511 18057
rect 280 17995 8565 18003
rect 220 17985 280 17995
rect 8510 17993 8565 17995
rect 207 17877 268 17887
rect 7055 17877 7109 17883
rect 268 17873 7109 17877
rect 268 17819 7055 17873
rect 268 17814 7109 17819
rect 207 17804 268 17814
rect 194 17686 265 17696
rect 5602 17687 5656 17697
rect 265 17633 5602 17686
rect 265 17614 5656 17633
rect 194 17604 265 17614
rect 4157 17501 4211 17511
rect 3250 16837 3310 16847
rect 3250 16765 3310 16775
rect 2415 16181 2486 16191
rect 2415 16112 2486 16122
rect 2701 16085 2770 16095
rect 2701 16011 2770 16021
rect 211 15880 265 15890
rect 4157 15882 4211 17447
rect 4267 17416 4321 17418
rect 4266 17408 4321 17416
rect 4266 17354 4267 17408
rect 4266 16012 4321 17354
rect 4698 16837 4758 16847
rect 4698 16765 4758 16775
rect 4474 16012 4528 16022
rect 4266 15958 4474 16012
rect 4474 15948 4528 15958
rect 4348 15899 4424 15909
rect 686 15881 4218 15882
rect 469 15880 4348 15881
rect 265 15826 4348 15880
rect 265 15825 4218 15826
rect 211 15815 265 15825
rect 5602 15879 5656 17614
rect 5733 17592 5787 17602
rect 5733 16011 5787 17538
rect 6196 16839 6256 16849
rect 6196 16767 6256 16777
rect 5968 16011 6022 16021
rect 5733 15957 5968 16011
rect 5968 15947 6022 15957
rect 5850 15891 5914 15901
rect 5602 15825 5850 15879
rect 7055 15884 7109 17814
rect 7183 17778 7237 17788
rect 7183 16014 7237 17724
rect 7644 16839 7704 16849
rect 7644 16767 7704 16777
rect 7394 16014 7472 16024
rect 7183 15960 7418 16014
rect 7183 15959 7472 15960
rect 7394 15950 7472 15959
rect 7299 15897 7366 15907
rect 7055 15830 7299 15884
rect 8510 15884 8564 17993
rect 8690 17963 8744 17973
rect 8690 16009 8744 17909
rect 9164 16837 9224 16847
rect 9164 16765 9224 16775
rect 8937 16009 8991 16019
rect 8690 15955 8937 16009
rect 8937 15945 8991 15955
rect 8818 15895 8878 15905
rect 8510 15830 8818 15884
rect 4348 15802 4424 15812
rect 5850 15807 5914 15817
rect 7299 15809 7366 15819
rect 10013 15878 10067 18184
rect 10151 18151 10205 18161
rect 10151 16017 10205 18097
rect 10612 16837 10672 16847
rect 10612 16765 10672 16775
rect 10385 16017 10439 16026
rect 10151 16016 10439 16017
rect 10151 15962 10385 16016
rect 10385 15952 10439 15962
rect 10268 15888 10328 15898
rect 10013 15824 10268 15878
rect 11474 15884 11528 18374
rect 11649 18335 11703 18345
rect 11649 16104 11703 18281
rect 12110 16839 12170 16849
rect 12110 16767 12170 16777
rect 11649 16050 11936 16104
rect 11882 16014 11936 16050
rect 11882 15950 11936 15960
rect 11767 15897 11828 15907
rect 11474 15830 11767 15884
rect 8818 15810 8878 15820
rect 10268 15810 10328 15820
rect 11767 15808 11828 15818
rect 13015 15901 13065 18551
rect 13106 18522 13160 18532
rect 13106 18458 13160 18468
rect 13108 16121 13158 18458
rect 15222 17046 15312 17056
rect 15222 16945 15312 16955
rect 16390 17046 16480 17056
rect 16390 16945 16480 16955
rect 17558 17046 17648 17056
rect 17558 16945 17648 16955
rect 18726 17046 18816 17056
rect 18726 16945 18816 16955
rect 19900 17048 19990 17058
rect 19900 16947 19990 16957
rect 21068 17048 21158 17058
rect 21068 16947 21158 16957
rect 22236 17048 22326 17058
rect 22236 16947 22326 16957
rect 23404 17048 23494 17058
rect 23404 16947 23494 16957
rect 13558 16839 13618 16849
rect 13558 16767 13618 16777
rect 13108 16071 13386 16121
rect 13335 16040 13385 16071
rect 13314 16030 13400 16040
rect 13314 15932 13400 15942
rect 13201 15911 13286 15912
rect 13200 15902 13286 15911
rect 13200 15901 13201 15902
rect 13015 15813 13200 15901
rect 13200 15812 13201 15813
rect 13200 15803 13286 15812
rect 13201 15802 13286 15803
rect 14757 15719 14847 15729
rect 6418 15643 6480 15645
rect 7866 15643 7928 15645
rect 12332 15643 12394 15645
rect 13780 15643 13842 15645
rect 3472 15641 3534 15643
rect 4920 15641 4982 15643
rect 3472 15633 3536 15641
rect 3534 15631 3536 15633
rect 3472 15559 3536 15569
rect 4920 15633 4984 15641
rect 4982 15631 4984 15633
rect 4920 15559 4984 15569
rect 6418 15635 6482 15643
rect 6480 15633 6482 15635
rect 6418 15561 6482 15571
rect 7866 15635 7930 15643
rect 7928 15633 7930 15635
rect 7866 15561 7930 15571
rect 9386 15641 9448 15643
rect 10834 15641 10896 15643
rect 9386 15633 9450 15641
rect 9448 15631 9450 15633
rect 9386 15559 9450 15569
rect 10834 15633 10898 15641
rect 10896 15631 10898 15633
rect 10834 15559 10898 15569
rect 12332 15635 12396 15643
rect 12394 15633 12396 15635
rect 12332 15561 12396 15571
rect 13780 15635 13844 15643
rect 13842 15633 13844 15635
rect 14757 15618 14847 15628
rect 15925 15719 16015 15729
rect 15925 15618 16015 15628
rect 17093 15719 17183 15729
rect 17093 15618 17183 15628
rect 18261 15719 18351 15729
rect 18261 15618 18351 15628
rect 19435 15721 19525 15731
rect 19435 15620 19525 15630
rect 20603 15721 20693 15731
rect 20603 15620 20693 15630
rect 21771 15721 21861 15731
rect 21771 15620 21861 15630
rect 22939 15721 23029 15731
rect 22939 15620 23029 15630
rect 13780 15561 13844 15571
rect 181 15506 239 15516
rect 181 15440 239 15450
rect 4204 15126 4304 15136
rect 4204 15024 4304 15034
rect 7348 15126 7448 15136
rect 7348 15024 7448 15034
rect 10480 15130 10580 15140
rect 10480 15028 10580 15038
rect 13624 15130 13724 15140
rect 13624 15028 13724 15038
rect 16826 15126 16926 15136
rect 16826 15024 16926 15034
rect 19970 15126 20070 15136
rect 19970 15024 20070 15034
rect 23102 15130 23202 15140
rect 23102 15028 23202 15038
rect 26246 15130 26346 15140
rect 26246 15028 26346 15038
rect 9334 14169 9427 14171
rect 12478 14169 12571 14171
rect 21956 14169 22049 14171
rect 25100 14169 25193 14171
rect 3058 14165 3151 14167
rect 6202 14165 6295 14167
rect 9090 14165 10509 14169
rect 12234 14165 13653 14169
rect 15680 14165 15773 14167
rect 18824 14165 18917 14167
rect 21712 14165 23131 14169
rect 24856 14165 26275 14169
rect 2189 14159 26275 14165
rect 2189 14158 9345 14159
rect 2189 14081 2205 14158
rect 2288 14155 9345 14158
rect 2288 14092 3069 14155
rect 3140 14093 4154 14155
rect 4224 14093 6213 14155
rect 3140 14092 6213 14093
rect 6284 14093 7298 14155
rect 7368 14096 9345 14155
rect 9416 14097 10430 14159
rect 10500 14097 12489 14159
rect 9416 14096 12489 14097
rect 12560 14097 13574 14159
rect 13644 14155 21967 14159
rect 13644 14097 15691 14155
rect 12560 14096 15691 14097
rect 7368 14093 15691 14096
rect 6284 14092 15691 14093
rect 15762 14093 16776 14155
rect 16846 14093 18835 14155
rect 15762 14092 18835 14093
rect 18906 14093 19920 14155
rect 19990 14096 21967 14155
rect 22038 14097 23052 14159
rect 23122 14097 25111 14159
rect 22038 14096 25111 14097
rect 25182 14097 26196 14159
rect 26266 14097 26275 14159
rect 25182 14096 26275 14097
rect 19990 14093 26275 14096
rect 18906 14092 26275 14093
rect 2288 14081 26275 14092
rect 2205 14060 2288 14070
rect 5969 14048 6026 14050
rect 2814 14045 2910 14048
rect 5958 14045 6054 14048
rect 2814 14040 4454 14045
rect 2814 13972 2825 14040
rect 2882 14035 4454 14040
rect 2882 13975 4395 14035
rect 2882 13972 4454 13975
rect 2814 13966 4454 13972
rect 2814 13963 2910 13966
rect 4395 13965 4454 13966
rect 5958 14040 7598 14045
rect 5958 13972 5969 14040
rect 6026 14035 7598 14040
rect 6026 13975 7539 14035
rect 6026 13972 7598 13975
rect 5958 13966 7598 13972
rect 9090 14044 10730 14049
rect 9090 13976 9101 14044
rect 9158 14039 10730 14044
rect 9158 13979 10671 14039
rect 9158 13976 10730 13979
rect 9090 13970 10730 13976
rect 10671 13969 10730 13970
rect 12234 14044 13874 14049
rect 12234 13976 12245 14044
rect 12302 14039 13874 14044
rect 12302 13979 13815 14039
rect 12302 13976 13874 13979
rect 12234 13970 13874 13976
rect 12234 13967 12330 13970
rect 13815 13969 13874 13970
rect 15436 14045 15532 14048
rect 18580 14045 18676 14048
rect 15436 14040 17076 14045
rect 15436 13972 15447 14040
rect 15504 14035 17076 14040
rect 15504 13975 17017 14035
rect 15504 13972 17076 13975
rect 12245 13966 12302 13967
rect 15436 13966 17076 13972
rect 5958 13963 6054 13966
rect 7539 13965 7598 13966
rect 15436 13963 15532 13966
rect 17017 13965 17076 13966
rect 18580 14040 20220 14045
rect 18580 13972 18591 14040
rect 18648 14035 20220 14040
rect 18648 13975 20161 14035
rect 18648 13972 20220 13975
rect 18580 13966 20220 13972
rect 21712 14044 23352 14049
rect 21712 13976 21723 14044
rect 21780 14039 23352 14044
rect 21780 13979 23293 14039
rect 21780 13976 23352 13979
rect 21712 13970 23352 13976
rect 21712 13967 21808 13970
rect 23293 13969 23352 13970
rect 24856 14044 26496 14049
rect 24856 13976 24867 14044
rect 24924 14039 26496 14044
rect 24924 13979 26437 14039
rect 24924 13976 26496 13979
rect 24856 13970 26496 13976
rect 24856 13967 24952 13970
rect 26437 13969 26496 13970
rect 21723 13966 21780 13967
rect 24867 13966 24924 13967
rect 18580 13963 18676 13966
rect 20161 13965 20220 13966
rect 2825 13962 2882 13963
rect 5969 13962 6026 13963
rect 15447 13962 15504 13963
rect 18591 13962 18648 13963
rect 9101 13885 9158 13886
rect 21723 13885 21780 13886
rect 24867 13885 24924 13886
rect 9090 13884 9186 13885
rect 21712 13884 21808 13885
rect 24856 13884 24952 13885
rect 2825 13881 2882 13882
rect 5969 13881 6026 13882
rect 2814 13880 2910 13881
rect 5958 13880 6054 13881
rect 2814 13872 4115 13880
rect 2814 13804 2825 13872
rect 2882 13807 4036 13872
rect 4104 13807 4115 13872
rect 2882 13804 4115 13807
rect 2814 13796 4115 13804
rect 5958 13872 7259 13880
rect 5958 13804 5969 13872
rect 6026 13807 7180 13872
rect 7248 13807 7259 13872
rect 6026 13804 7259 13807
rect 5958 13796 7259 13804
rect 9090 13876 10391 13884
rect 18591 13881 18648 13882
rect 9090 13808 9101 13876
rect 9158 13811 10312 13876
rect 10380 13811 10391 13876
rect 9158 13808 10391 13811
rect 9090 13800 10391 13808
rect 18580 13880 18676 13881
rect 18580 13872 19881 13880
rect 18580 13804 18591 13872
rect 18648 13807 19802 13872
rect 19870 13807 19881 13872
rect 18648 13804 19881 13807
rect 9101 13798 9158 13800
rect 18580 13796 19881 13804
rect 21712 13876 23013 13884
rect 21712 13808 21723 13876
rect 21780 13811 22934 13876
rect 23002 13811 23013 13876
rect 21780 13808 23013 13811
rect 21712 13800 23013 13808
rect 24856 13876 26157 13884
rect 24856 13808 24867 13876
rect 24924 13811 26078 13876
rect 26146 13811 26157 13876
rect 24924 13808 26157 13811
rect 24856 13800 26157 13808
rect 21723 13798 21780 13800
rect 24867 13798 24924 13800
rect 2825 13794 2882 13796
rect 5969 13794 6026 13796
rect 18591 13794 18648 13796
rect 4224 12882 4300 12892
rect 4224 12814 4300 12824
rect 7368 12882 7444 12892
rect 7368 12814 7444 12824
rect 10500 12886 10576 12896
rect 10500 12818 10576 12828
rect 13644 12886 13720 12896
rect 13644 12818 13720 12828
rect 16846 12882 16922 12892
rect 16846 12814 16922 12824
rect 19990 12882 20066 12892
rect 19990 12814 20066 12824
rect 23122 12886 23198 12896
rect 23122 12818 23198 12828
rect 26266 12886 26342 12896
rect 26266 12818 26342 12828
rect 4204 12392 4304 12402
rect 4204 12290 4304 12300
rect 7348 12392 7448 12402
rect 7348 12290 7448 12300
rect 10480 12396 10580 12406
rect 10480 12294 10580 12304
rect 13624 12396 13724 12406
rect 13624 12294 13724 12304
rect 16826 12392 16926 12402
rect 16826 12290 16926 12300
rect 19970 12392 20070 12402
rect 19970 12290 20070 12300
rect 23102 12396 23202 12406
rect 23102 12294 23202 12304
rect 26246 12396 26346 12406
rect 26246 12294 26346 12304
rect 12478 11435 12571 11437
rect 21956 11435 22049 11437
rect 25100 11435 25193 11437
rect 201 11431 263 11435
rect 9093 11434 13653 11435
rect 21715 11434 23131 11435
rect 24859 11434 26275 11435
rect 3058 11431 3151 11433
rect 6202 11431 6295 11433
rect 9090 11431 13653 11434
rect 15680 11431 15773 11433
rect 18824 11431 18917 11433
rect 19937 11431 26275 11434
rect 196 11430 13653 11431
rect 15439 11430 16855 11431
rect 18583 11430 26275 11431
rect 196 11429 16855 11430
rect 18580 11429 26275 11430
rect 196 11425 26275 11429
rect 196 11350 201 11425
rect 263 11421 9345 11425
rect 263 11358 3069 11421
rect 3140 11359 4154 11421
rect 4224 11359 6213 11421
rect 3140 11358 6213 11359
rect 6284 11359 7298 11421
rect 7368 11362 9345 11421
rect 9416 11363 10430 11425
rect 10500 11363 12489 11425
rect 9416 11362 12489 11363
rect 12560 11363 13574 11425
rect 13644 11422 21967 11425
rect 13644 11421 18591 11422
rect 13644 11363 15691 11421
rect 12560 11362 15691 11363
rect 7368 11359 15691 11362
rect 6284 11358 15691 11359
rect 15762 11359 16776 11421
rect 16846 11359 18591 11421
rect 15762 11358 18591 11359
rect 263 11354 18591 11358
rect 18648 11421 21967 11422
rect 18648 11358 18835 11421
rect 18906 11359 19920 11421
rect 19990 11362 21967 11421
rect 22038 11363 23052 11425
rect 23122 11363 25111 11425
rect 22038 11362 25111 11363
rect 25182 11363 26196 11425
rect 26266 11363 26275 11425
rect 25182 11362 26275 11363
rect 19990 11359 26275 11362
rect 18906 11358 26275 11359
rect 18648 11354 26275 11358
rect 263 11351 26275 11354
rect 263 11350 9168 11351
rect 196 11348 9158 11350
rect 196 11347 9121 11348
rect 15436 11347 21744 11351
rect 196 11346 2724 11347
rect 201 11340 263 11346
rect 12245 11318 12302 11320
rect 24867 11318 24924 11320
rect 2825 11314 2882 11316
rect 5969 11314 6026 11316
rect 12234 11315 12330 11318
rect 2814 11311 2910 11314
rect 5958 11311 6054 11314
rect 2814 11306 4454 11311
rect 2814 11238 2825 11306
rect 2882 11301 4454 11306
rect 2882 11241 4395 11301
rect 2882 11238 4454 11241
rect 2814 11232 4454 11238
rect 2814 11229 2910 11232
rect 4395 11231 4454 11232
rect 5958 11306 7598 11311
rect 5958 11238 5969 11306
rect 6026 11301 7598 11306
rect 6026 11241 7539 11301
rect 6026 11238 7598 11241
rect 5958 11232 7598 11238
rect 9090 11310 10730 11315
rect 9090 11242 9101 11310
rect 9158 11305 10730 11310
rect 9158 11245 10671 11305
rect 9158 11242 10730 11245
rect 9090 11236 10730 11242
rect 9090 11233 9186 11236
rect 10671 11235 10730 11236
rect 12234 11310 13874 11315
rect 18591 11314 18648 11316
rect 24856 11315 24952 11318
rect 12234 11242 12245 11310
rect 12302 11305 13874 11310
rect 12302 11245 13815 11305
rect 12302 11242 13874 11245
rect 12234 11236 13874 11242
rect 12234 11233 12330 11236
rect 13815 11235 13874 11236
rect 15436 11311 15532 11314
rect 18580 11311 18676 11314
rect 15436 11306 17076 11311
rect 15436 11238 15447 11306
rect 15504 11301 17076 11306
rect 15504 11241 17017 11301
rect 15504 11238 17076 11241
rect 9101 11232 9158 11233
rect 12245 11232 12302 11233
rect 15436 11232 17076 11238
rect 5958 11229 6054 11232
rect 7539 11231 7598 11232
rect 15436 11229 15532 11232
rect 17017 11231 17076 11232
rect 18580 11306 20220 11311
rect 18580 11238 18591 11306
rect 18648 11301 20220 11306
rect 18648 11241 20161 11301
rect 18648 11238 20220 11241
rect 18580 11232 20220 11238
rect 21712 11310 23352 11315
rect 21712 11242 21723 11310
rect 21780 11305 23352 11310
rect 21780 11245 23293 11305
rect 21780 11242 23352 11245
rect 21712 11236 23352 11242
rect 21712 11233 21808 11236
rect 23293 11235 23352 11236
rect 24856 11310 26496 11315
rect 24856 11242 24867 11310
rect 24924 11305 26496 11310
rect 24924 11245 26437 11305
rect 24924 11242 26496 11245
rect 24856 11236 26496 11242
rect 24856 11233 24952 11236
rect 26437 11235 26496 11236
rect 21723 11232 21780 11233
rect 24867 11232 24924 11233
rect 18580 11229 18676 11232
rect 20161 11231 20220 11232
rect 2825 11228 2882 11229
rect 5969 11228 6026 11229
rect 15447 11228 15504 11229
rect 18591 11228 18648 11229
rect 9101 11151 9158 11152
rect 12245 11151 12302 11152
rect 21723 11151 21780 11152
rect 24867 11151 24924 11152
rect 9090 11150 9186 11151
rect 12234 11150 12330 11151
rect 21712 11150 21808 11151
rect 24856 11150 24952 11151
rect 2825 11147 2882 11148
rect 5969 11147 6026 11148
rect 2814 11146 2910 11147
rect 5958 11146 6054 11147
rect 2814 11138 4115 11146
rect 202 11106 264 11108
rect 2212 11106 2279 11109
rect 202 11104 2299 11106
rect 197 11099 2299 11104
rect 197 11098 2212 11099
rect 197 11023 202 11098
rect 264 11029 2212 11098
rect 2279 11029 2299 11099
rect 2814 11070 2825 11138
rect 2882 11073 4036 11138
rect 4104 11073 4115 11138
rect 2882 11070 4115 11073
rect 2814 11062 4115 11070
rect 5958 11138 7259 11146
rect 5958 11070 5969 11138
rect 6026 11073 7180 11138
rect 7248 11073 7259 11138
rect 6026 11070 7259 11073
rect 5958 11062 7259 11070
rect 9090 11142 10391 11150
rect 9090 11074 9101 11142
rect 9158 11077 10312 11142
rect 10380 11077 10391 11142
rect 9158 11074 10391 11077
rect 9090 11066 10391 11074
rect 12234 11142 13535 11150
rect 15447 11147 15504 11148
rect 18591 11147 18648 11148
rect 12234 11074 12245 11142
rect 12302 11077 13456 11142
rect 13524 11077 13535 11142
rect 12302 11074 13535 11077
rect 12234 11066 13535 11074
rect 15436 11146 15532 11147
rect 18580 11146 18676 11147
rect 15436 11138 16737 11146
rect 15436 11070 15447 11138
rect 15504 11073 16658 11138
rect 16726 11073 16737 11138
rect 15504 11070 16737 11073
rect 9101 11064 9158 11066
rect 12245 11064 12302 11066
rect 15436 11062 16737 11070
rect 18580 11138 19881 11146
rect 18580 11070 18591 11138
rect 18648 11073 19802 11138
rect 19870 11073 19881 11138
rect 18648 11070 19881 11073
rect 18580 11062 19881 11070
rect 21712 11142 23013 11150
rect 21712 11074 21723 11142
rect 21780 11077 22934 11142
rect 23002 11077 23013 11142
rect 21780 11074 23013 11077
rect 21712 11066 23013 11074
rect 24856 11142 26157 11150
rect 24856 11074 24867 11142
rect 24924 11077 26078 11142
rect 26146 11077 26157 11142
rect 24924 11074 26157 11077
rect 24856 11066 26157 11074
rect 21723 11064 21780 11066
rect 24867 11064 24924 11066
rect 2825 11060 2882 11062
rect 5969 11060 6026 11062
rect 15447 11060 15504 11062
rect 18591 11060 18648 11062
rect 264 11023 2299 11029
rect 197 11020 2299 11023
rect 197 11019 288 11020
rect 2212 11019 2279 11020
rect 202 11013 264 11019
rect 24525 10937 27974 10947
rect 24525 10930 27915 10937
rect 24596 10867 27915 10930
rect 24596 10859 27974 10867
rect 24525 10849 24596 10859
rect 27915 10857 27974 10859
rect 21396 10771 21466 10781
rect 21466 10745 27976 10758
rect 21466 10682 27914 10745
rect 27975 10682 27976 10745
rect 21466 10678 27976 10682
rect 21396 10672 27976 10678
rect 21396 10668 21466 10672
rect 18237 10542 18333 10550
rect 18237 10540 27976 10542
rect 18333 10525 27976 10540
rect 18333 10459 27913 10525
rect 27975 10459 27976 10525
rect 18333 10448 27976 10459
rect 18237 10435 18333 10445
rect 15037 10336 27977 10346
rect 15115 10329 27977 10336
rect 15115 10271 27913 10329
rect 27976 10271 27977 10329
rect 15115 10267 27977 10271
rect 15037 10260 27977 10267
rect 15037 10257 15115 10260
rect 5644 10184 5708 10187
rect 5634 10177 5719 10184
rect 4224 10148 4300 10158
rect 4224 10080 4300 10090
rect 5634 10100 5644 10177
rect 5708 10100 5719 10177
rect 4194 9660 4294 9670
rect 4194 9558 4294 9568
rect 5634 9479 5719 10100
rect 7368 10148 7444 10158
rect 10500 10152 10576 10162
rect 8754 10118 8822 10128
rect 7368 10080 7444 10090
rect 8745 10046 8754 10106
rect 8822 10046 8832 10106
rect 10500 10084 10576 10094
rect 13644 10152 13720 10162
rect 13644 10084 13720 10094
rect 16846 10148 16922 10158
rect 16846 10080 16922 10090
rect 19990 10148 20066 10158
rect 19990 10080 20066 10090
rect 23122 10152 23198 10162
rect 23122 10084 23198 10094
rect 26266 10152 26342 10162
rect 26266 10084 26342 10094
rect 8745 9830 8832 10046
rect 11892 10002 27977 10003
rect 11890 9992 27977 10002
rect 11957 9986 27977 9992
rect 11957 9925 27912 9986
rect 27976 9925 27977 9986
rect 11957 9924 27977 9925
rect 11890 9914 27977 9924
rect 8745 9814 27980 9830
rect 8745 9754 27914 9814
rect 27978 9754 27980 9814
rect 8745 9743 27980 9754
rect 7338 9660 7438 9670
rect 7338 9558 7438 9568
rect 10470 9664 10570 9674
rect 10470 9562 10570 9572
rect 13614 9664 13714 9674
rect 13614 9562 13714 9572
rect 16816 9660 16916 9670
rect 16816 9558 16916 9568
rect 19960 9660 20060 9670
rect 19960 9558 20060 9568
rect 23092 9664 23192 9674
rect 23092 9562 23192 9572
rect 26236 9664 26336 9674
rect 26236 9562 26336 9572
rect 5634 9460 27980 9479
rect 5634 9399 27913 9460
rect 5634 9387 27980 9399
rect 5634 9386 5719 9387
rect 9091 8703 9148 8704
rect 9324 8703 9417 8705
rect 12235 8703 12292 8704
rect 12468 8703 12561 8705
rect 21713 8703 21770 8704
rect 21946 8703 22039 8705
rect 24857 8703 24914 8704
rect 25090 8703 25183 8705
rect 9083 8702 10499 8703
rect 12227 8702 13643 8703
rect 21705 8702 23121 8703
rect 24849 8702 26265 8703
rect 2815 8699 2872 8700
rect 3048 8699 3141 8701
rect 5959 8699 6016 8700
rect 6192 8699 6285 8701
rect 9080 8699 10499 8702
rect 12224 8699 13643 8702
rect 15437 8699 15494 8700
rect 15670 8699 15763 8701
rect 18581 8699 18638 8700
rect 18814 8699 18907 8701
rect 21702 8699 23121 8702
rect 24846 8699 26265 8702
rect 2804 8694 26265 8699
rect 2804 8690 9091 8694
rect 2804 8622 2815 8690
rect 2872 8689 5959 8690
rect 2872 8626 3059 8689
rect 3130 8627 4144 8689
rect 4214 8627 5959 8689
rect 3130 8626 5959 8627
rect 2872 8622 5959 8626
rect 6016 8689 9091 8690
rect 6016 8626 6203 8689
rect 6274 8627 7288 8689
rect 7358 8627 9091 8689
rect 6274 8626 9091 8627
rect 9148 8693 12235 8694
rect 9148 8630 9335 8693
rect 9406 8631 10420 8693
rect 10490 8631 12235 8693
rect 9406 8630 12235 8631
rect 9148 8626 12235 8630
rect 12292 8693 21713 8694
rect 12292 8630 12479 8693
rect 12550 8631 13564 8693
rect 13634 8690 21713 8693
rect 13634 8631 15437 8690
rect 12550 8630 15437 8631
rect 12292 8626 15437 8630
rect 6016 8622 15437 8626
rect 15494 8689 18581 8690
rect 15494 8626 15681 8689
rect 15752 8627 16766 8689
rect 16836 8627 18581 8689
rect 15752 8626 18581 8627
rect 15494 8622 18581 8626
rect 18638 8689 21713 8690
rect 18638 8626 18825 8689
rect 18896 8627 19910 8689
rect 19980 8627 21713 8689
rect 18896 8626 21713 8627
rect 21770 8693 24857 8694
rect 21770 8630 21957 8693
rect 22028 8631 23042 8693
rect 23112 8631 24857 8693
rect 22028 8630 24857 8631
rect 21770 8626 24857 8630
rect 24914 8693 26265 8694
rect 24914 8630 25101 8693
rect 25172 8631 26186 8693
rect 26256 8631 26265 8693
rect 25172 8630 26265 8631
rect 24914 8626 26265 8630
rect 18638 8622 26265 8626
rect 2804 8614 26265 8622
rect 2815 8612 2872 8614
rect 5959 8612 6016 8614
rect 15437 8612 15494 8614
rect 18581 8612 18638 8614
rect 2815 8582 2872 8584
rect 5959 8582 6016 8584
rect 2804 8579 2900 8582
rect 5948 8579 6044 8582
rect 2804 8574 4444 8579
rect 2804 8506 2815 8574
rect 2872 8569 4444 8574
rect 2872 8509 4385 8569
rect 2872 8506 4444 8509
rect 2804 8500 4444 8506
rect 2804 8497 2900 8500
rect 4385 8499 4444 8500
rect 5948 8574 7588 8579
rect 5948 8506 5959 8574
rect 6016 8569 7588 8574
rect 6016 8509 7529 8569
rect 6016 8506 7588 8509
rect 5948 8500 7588 8506
rect 9080 8578 10720 8583
rect 9080 8510 9091 8578
rect 9148 8573 10720 8578
rect 9148 8513 10661 8573
rect 9148 8510 10720 8513
rect 9080 8504 10720 8510
rect 9080 8501 9176 8504
rect 10661 8503 10720 8504
rect 12224 8578 13864 8583
rect 15437 8582 15494 8584
rect 18581 8582 18638 8584
rect 12224 8510 12235 8578
rect 12292 8573 13864 8578
rect 12292 8513 13805 8573
rect 12292 8510 13864 8513
rect 12224 8504 13864 8510
rect 12224 8501 12320 8504
rect 13805 8503 13864 8504
rect 15426 8579 15522 8582
rect 18570 8579 18666 8582
rect 15426 8574 17066 8579
rect 15426 8506 15437 8574
rect 15494 8569 17066 8574
rect 15494 8509 17007 8569
rect 15494 8506 17066 8509
rect 9091 8500 9148 8501
rect 12235 8500 12292 8501
rect 15426 8500 17066 8506
rect 5948 8497 6044 8500
rect 7529 8499 7588 8500
rect 15426 8497 15522 8500
rect 17007 8499 17066 8500
rect 18570 8574 20210 8579
rect 18570 8506 18581 8574
rect 18638 8569 20210 8574
rect 18638 8509 20151 8569
rect 18638 8506 20210 8509
rect 18570 8500 20210 8506
rect 21702 8578 23342 8583
rect 21702 8510 21713 8578
rect 21770 8573 23342 8578
rect 21770 8513 23283 8573
rect 21770 8510 23342 8513
rect 21702 8504 23342 8510
rect 21702 8501 21798 8504
rect 23283 8503 23342 8504
rect 24846 8578 26486 8583
rect 24846 8510 24857 8578
rect 24914 8573 26486 8578
rect 24914 8513 26427 8573
rect 24914 8510 26486 8513
rect 24846 8504 26486 8510
rect 24846 8501 24942 8504
rect 26427 8503 26486 8504
rect 21713 8500 21770 8501
rect 24857 8500 24914 8501
rect 18570 8497 18666 8500
rect 20151 8499 20210 8500
rect 2815 8496 2872 8497
rect 5959 8496 6016 8497
rect 15437 8496 15494 8497
rect 18581 8496 18638 8497
rect 9091 8419 9148 8420
rect 12235 8419 12292 8420
rect 21713 8419 21770 8420
rect 24857 8419 24914 8420
rect 9080 8418 9176 8419
rect 12224 8418 12320 8419
rect 21702 8418 21798 8419
rect 24846 8418 24942 8419
rect 2815 8415 2872 8416
rect 5959 8415 6016 8416
rect 2804 8414 2900 8415
rect 5948 8414 6044 8415
rect 2804 8406 4105 8414
rect 2804 8338 2815 8406
rect 2872 8341 4026 8406
rect 4094 8341 4105 8406
rect 2872 8338 4105 8341
rect 2804 8330 4105 8338
rect 5948 8406 7249 8414
rect 5948 8338 5959 8406
rect 6016 8341 7170 8406
rect 7238 8341 7249 8406
rect 6016 8338 7249 8341
rect 5948 8330 7249 8338
rect 9080 8410 10381 8418
rect 9080 8342 9091 8410
rect 9148 8345 10302 8410
rect 10370 8345 10381 8410
rect 9148 8342 10381 8345
rect 9080 8334 10381 8342
rect 12224 8410 13525 8418
rect 15437 8415 15494 8416
rect 18581 8415 18638 8416
rect 12224 8342 12235 8410
rect 12292 8345 13446 8410
rect 13514 8345 13525 8410
rect 12292 8342 13525 8345
rect 12224 8334 13525 8342
rect 15426 8414 15522 8415
rect 18570 8414 18666 8415
rect 15426 8406 16727 8414
rect 15426 8338 15437 8406
rect 15494 8341 16648 8406
rect 16716 8341 16727 8406
rect 15494 8338 16727 8341
rect 9091 8332 9148 8334
rect 12235 8332 12292 8334
rect 15426 8330 16727 8338
rect 18570 8406 19871 8414
rect 18570 8338 18581 8406
rect 18638 8341 19792 8406
rect 19860 8341 19871 8406
rect 18638 8338 19871 8341
rect 18570 8330 19871 8338
rect 21702 8410 23003 8418
rect 21702 8342 21713 8410
rect 21770 8345 22924 8410
rect 22992 8345 23003 8410
rect 21770 8342 23003 8345
rect 21702 8334 23003 8342
rect 24846 8410 26147 8418
rect 24846 8342 24857 8410
rect 24914 8345 26068 8410
rect 26136 8345 26147 8410
rect 24914 8342 26147 8345
rect 24846 8334 26147 8342
rect 21713 8332 21770 8334
rect 24857 8332 24914 8334
rect 2815 8328 2872 8330
rect 5959 8328 6016 8330
rect 15437 8328 15494 8330
rect 18581 8328 18638 8330
rect 4214 7416 4290 7426
rect 4214 7348 4290 7358
rect 7358 7416 7434 7426
rect 7358 7348 7434 7358
rect 10490 7420 10566 7430
rect 10490 7352 10566 7362
rect 13634 7420 13710 7430
rect 13634 7352 13710 7362
rect 16836 7416 16912 7426
rect 16836 7348 16912 7358
rect 19980 7416 20056 7426
rect 19980 7348 20056 7358
rect 23112 7420 23188 7430
rect 23112 7352 23188 7362
rect 26256 7420 26332 7430
rect 26256 7352 26332 7362
rect 471 7158 526 7167
rect 727 7158 795 7167
rect 471 7157 799 7158
rect 526 7099 727 7157
rect 795 7099 799 7157
rect 526 7096 799 7099
rect 471 7086 526 7096
rect 727 7089 795 7096
rect 471 6866 526 6875
rect 471 6865 541 6866
rect 986 6865 1042 6873
rect 526 6863 1053 6865
rect 526 6806 986 6863
rect 1042 6806 1053 6863
rect 526 6804 1053 6806
rect 471 6794 526 6804
rect 986 6796 1042 6804
rect 19577 6763 19671 6773
rect 3510 6702 3588 6712
rect 3510 6622 3588 6632
rect 5578 6704 5656 6714
rect 5578 6624 5656 6634
rect 7647 6702 7725 6712
rect 7647 6622 7725 6632
rect 9715 6704 9793 6714
rect 9715 6624 9793 6634
rect 11784 6704 11862 6714
rect 11784 6624 11862 6634
rect 13852 6706 13930 6716
rect 13852 6626 13930 6636
rect 15921 6704 15999 6714
rect 15921 6624 15999 6634
rect 17989 6706 18067 6716
rect 19577 6669 19671 6679
rect 20315 6761 20409 6771
rect 20315 6667 20409 6677
rect 21053 6761 21147 6771
rect 21053 6667 21147 6677
rect 21795 6761 21889 6771
rect 21795 6667 21889 6677
rect 22535 6761 22629 6771
rect 22535 6667 22629 6677
rect 23273 6761 23367 6771
rect 23273 6667 23367 6677
rect 24011 6761 24105 6771
rect 24011 6667 24105 6677
rect 24749 6761 24843 6771
rect 24749 6667 24843 6677
rect 17989 6626 18067 6636
rect 471 6561 526 6570
rect 471 6560 541 6561
rect 1204 6560 1265 6565
rect 526 6555 1267 6560
rect 526 6502 1204 6555
rect 1265 6502 1267 6555
rect 526 6499 1267 6502
rect 471 6489 526 6499
rect 1204 6492 1265 6499
rect 471 6400 526 6409
rect 471 6399 541 6400
rect 1379 6399 1449 6408
rect 526 6398 1454 6399
rect 526 6340 1379 6398
rect 1449 6340 1454 6398
rect 526 6338 1454 6340
rect 471 6328 526 6338
rect 1379 6330 1449 6338
rect 471 6249 527 6258
rect 471 6248 528 6249
rect 1581 6248 1649 6258
rect 527 6190 1581 6248
rect 1649 6190 1652 6248
rect 527 6187 1652 6190
rect 471 6177 527 6187
rect 1581 6180 1649 6187
rect 471 6089 526 6098
rect 471 6088 541 6089
rect 1777 6088 1835 6095
rect 526 6085 1839 6088
rect 526 6031 1777 6085
rect 1835 6031 1839 6085
rect 526 6027 1839 6031
rect 471 6017 526 6027
rect 1777 6021 1835 6027
rect 471 5902 526 5911
rect 2005 5902 2069 5911
rect 4777 5910 4852 5920
rect 471 5901 2070 5902
rect 526 5841 2005 5901
rect 2069 5841 2070 5901
rect 526 5840 2070 5841
rect 2426 5886 2492 5896
rect 471 5830 526 5840
rect 2005 5831 2069 5840
rect 2426 5819 2492 5829
rect 2708 5826 2714 5892
rect 2780 5886 4156 5892
rect 2780 5832 4102 5886
rect 2780 5826 4156 5832
rect 4776 5828 4777 5894
rect 4852 5888 6224 5894
rect 6848 5892 6917 5902
rect 8920 5894 8984 5903
rect 10988 5896 11055 5906
rect 13051 5896 13116 5906
rect 17186 5905 17269 5915
rect 4852 5834 6170 5888
rect 4852 5828 6224 5834
rect 6845 5826 6848 5892
rect 6917 5886 8293 5892
rect 6917 5832 8239 5886
rect 6917 5826 8293 5832
rect 8913 5828 8919 5894
rect 8985 5888 10361 5894
rect 8985 5834 10307 5888
rect 8985 5828 10361 5834
rect 10982 5828 10988 5894
rect 11055 5888 12430 5894
rect 11055 5834 12376 5888
rect 11055 5828 12430 5834
rect 13050 5830 13051 5896
rect 13122 5890 14498 5896
rect 15122 5894 15189 5903
rect 13122 5836 14444 5890
rect 13122 5830 14498 5836
rect 15119 5893 15125 5894
rect 15119 5829 15122 5893
rect 15191 5888 16567 5894
rect 15191 5834 16513 5888
rect 15119 5828 15125 5829
rect 15191 5828 16567 5834
rect 17269 5890 18635 5896
rect 17269 5836 18581 5890
rect 17269 5830 18635 5836
rect 19509 5875 19611 5881
rect 19509 5871 19613 5875
rect 4777 5814 4852 5824
rect 6848 5816 6917 5826
rect 8920 5818 8984 5828
rect 10988 5817 11055 5827
rect 13051 5818 13116 5828
rect 15122 5819 15189 5828
rect 17186 5815 17269 5825
rect 19611 5805 19613 5871
rect 19509 5797 19613 5805
rect 20247 5873 20349 5879
rect 20985 5873 21087 5879
rect 21727 5873 21829 5879
rect 22467 5873 22569 5879
rect 23205 5873 23307 5879
rect 23943 5873 24045 5879
rect 24681 5873 24783 5879
rect 20247 5869 20351 5873
rect 20349 5803 20351 5869
rect 19509 5795 19611 5797
rect 20247 5795 20351 5803
rect 20985 5869 21089 5873
rect 21087 5803 21089 5869
rect 20985 5795 21089 5803
rect 21727 5869 21831 5873
rect 21829 5803 21831 5869
rect 21727 5795 21831 5803
rect 22467 5869 22571 5873
rect 22569 5803 22571 5869
rect 22467 5795 22571 5803
rect 23205 5869 23309 5873
rect 23307 5803 23309 5869
rect 23205 5795 23309 5803
rect 23943 5869 24047 5873
rect 24045 5803 24047 5869
rect 23943 5795 24047 5803
rect 24681 5869 24785 5873
rect 24783 5803 24785 5869
rect 24681 5795 24785 5803
rect 20247 5793 20349 5795
rect 20985 5793 21087 5795
rect 21727 5793 21829 5795
rect 22467 5793 22569 5795
rect 23205 5793 23307 5795
rect 23943 5793 24045 5795
rect 24681 5793 24783 5795
rect 471 5695 526 5705
rect 2699 5704 2770 5714
rect 2428 5694 2480 5703
rect 526 5693 2480 5694
rect 526 5635 2428 5693
rect 471 5624 526 5634
rect 2428 5625 2480 5635
rect 2699 5617 2770 5627
rect 3458 4472 3530 4482
rect 3458 4392 3530 4402
rect 5526 4474 5598 4484
rect 5526 4394 5598 4404
rect 7595 4472 7667 4482
rect 7595 4392 7667 4402
rect 9663 4474 9735 4484
rect 9663 4394 9735 4404
rect 11732 4474 11804 4484
rect 11732 4394 11804 4404
rect 13800 4476 13872 4486
rect 13800 4396 13872 4406
rect 15869 4474 15941 4484
rect 15869 4394 15941 4404
rect 17937 4476 18009 4486
rect 17937 4396 18009 4406
rect 1496 2412 1596 2422
rect 1496 2310 1596 2320
rect 4640 2412 4740 2422
rect 4640 2310 4740 2320
rect 7772 2416 7872 2426
rect 7772 2314 7872 2324
rect 10916 2416 11016 2426
rect 10916 2314 11016 2324
rect 14118 2412 14218 2422
rect 14118 2310 14218 2320
rect 17262 2412 17362 2422
rect 17262 2310 17362 2320
rect 20394 2416 20494 2426
rect 20394 2314 20494 2324
rect 23538 2416 23638 2426
rect 23538 2314 23638 2324
rect 6393 1455 6450 1456
rect 6626 1455 6719 1457
rect 9537 1455 9594 1456
rect 9770 1455 9863 1457
rect 19015 1455 19072 1456
rect 19248 1455 19341 1457
rect 22159 1455 22216 1456
rect 22392 1455 22485 1457
rect 6385 1454 7801 1455
rect 9529 1454 10945 1455
rect 19007 1454 20423 1455
rect 22151 1454 23567 1455
rect 117 1451 174 1452
rect 350 1451 443 1453
rect 3261 1451 3318 1452
rect 3494 1451 3587 1453
rect 109 1450 1525 1451
rect 3253 1450 4669 1451
rect 106 1442 1525 1450
rect 106 1374 117 1442
rect 174 1441 1525 1442
rect 174 1378 361 1441
rect 432 1379 1446 1441
rect 1516 1379 1525 1441
rect 432 1378 1525 1379
rect 174 1374 1525 1378
rect 106 1367 1525 1374
rect 3250 1442 4669 1450
rect 3250 1374 3261 1442
rect 3318 1441 4669 1442
rect 3318 1378 3505 1441
rect 3576 1379 4590 1441
rect 4660 1379 4669 1441
rect 3576 1378 4669 1379
rect 3318 1374 4669 1378
rect 3250 1367 4669 1374
rect 6382 1446 7801 1454
rect 6382 1378 6393 1446
rect 6450 1445 7801 1446
rect 6450 1382 6637 1445
rect 6708 1383 7722 1445
rect 7792 1383 7801 1445
rect 6708 1382 7801 1383
rect 6450 1378 7801 1382
rect 6382 1371 7801 1378
rect 9526 1446 10945 1454
rect 12739 1451 12796 1452
rect 12972 1451 13065 1453
rect 15883 1451 15940 1452
rect 16116 1451 16209 1453
rect 12731 1450 14147 1451
rect 15875 1450 17291 1451
rect 9526 1378 9537 1446
rect 9594 1445 10945 1446
rect 9594 1382 9781 1445
rect 9852 1383 10866 1445
rect 10936 1383 10945 1445
rect 9852 1382 10945 1383
rect 9594 1378 10945 1382
rect 9526 1371 10945 1378
rect 12728 1442 14147 1450
rect 12728 1374 12739 1442
rect 12796 1441 14147 1442
rect 12796 1378 12983 1441
rect 13054 1379 14068 1441
rect 14138 1379 14147 1441
rect 13054 1378 14147 1379
rect 12796 1374 14147 1378
rect 6382 1370 6460 1371
rect 9526 1370 9604 1371
rect 6393 1368 6450 1370
rect 9537 1368 9594 1370
rect 12728 1367 14147 1374
rect 15872 1442 17291 1450
rect 15872 1374 15883 1442
rect 15940 1441 17291 1442
rect 15940 1378 16127 1441
rect 16198 1379 17212 1441
rect 17282 1379 17291 1441
rect 16198 1378 17291 1379
rect 15940 1374 17291 1378
rect 15872 1367 17291 1374
rect 19004 1446 20423 1454
rect 19004 1378 19015 1446
rect 19072 1445 20423 1446
rect 19072 1382 19259 1445
rect 19330 1383 20344 1445
rect 20414 1383 20423 1445
rect 19330 1382 20423 1383
rect 19072 1378 20423 1382
rect 19004 1371 20423 1378
rect 22148 1446 23567 1454
rect 22148 1378 22159 1446
rect 22216 1445 23567 1446
rect 22216 1382 22403 1445
rect 22474 1383 23488 1445
rect 23558 1383 23567 1445
rect 22474 1382 23567 1383
rect 22216 1378 23567 1382
rect 22148 1371 23567 1378
rect 19004 1370 19082 1371
rect 22148 1370 22226 1371
rect 19015 1368 19072 1370
rect 22159 1368 22216 1370
rect 106 1366 184 1367
rect 3250 1366 3328 1367
rect 12728 1366 12806 1367
rect 15872 1366 15950 1367
rect 117 1364 174 1366
rect 3261 1364 3318 1366
rect 12739 1364 12796 1366
rect 15883 1364 15940 1366
rect 6393 1338 6450 1340
rect 9537 1338 9594 1340
rect 19015 1338 19072 1340
rect 22159 1338 22216 1340
rect 117 1334 174 1336
rect 3261 1334 3318 1336
rect 6382 1335 6478 1338
rect 9526 1335 9622 1338
rect 106 1331 202 1334
rect 3250 1331 3346 1334
rect 106 1326 1746 1331
rect 106 1258 117 1326
rect 174 1321 1746 1326
rect 174 1261 1687 1321
rect 174 1258 1746 1261
rect 106 1252 1746 1258
rect 106 1249 202 1252
rect 1687 1251 1746 1252
rect 3250 1326 4890 1331
rect 3250 1258 3261 1326
rect 3318 1321 4890 1326
rect 3318 1261 4831 1321
rect 3318 1258 4890 1261
rect 3250 1252 4890 1258
rect 6382 1330 8022 1335
rect 6382 1262 6393 1330
rect 6450 1325 8022 1330
rect 6450 1265 7963 1325
rect 6450 1262 8022 1265
rect 6382 1256 8022 1262
rect 6382 1253 6478 1256
rect 7963 1255 8022 1256
rect 9526 1330 11166 1335
rect 12739 1334 12796 1336
rect 15883 1334 15940 1336
rect 19004 1335 19100 1338
rect 22148 1335 22244 1338
rect 9526 1262 9537 1330
rect 9594 1325 11166 1330
rect 9594 1265 11107 1325
rect 9594 1262 11166 1265
rect 9526 1256 11166 1262
rect 9526 1253 9622 1256
rect 11107 1255 11166 1256
rect 12728 1331 12824 1334
rect 15872 1331 15968 1334
rect 12728 1326 14368 1331
rect 12728 1258 12739 1326
rect 12796 1321 14368 1326
rect 12796 1261 14309 1321
rect 12796 1258 14368 1261
rect 6393 1252 6450 1253
rect 9537 1252 9594 1253
rect 12728 1252 14368 1258
rect 3250 1249 3346 1252
rect 4831 1251 4890 1252
rect 12728 1249 12824 1252
rect 14309 1251 14368 1252
rect 15872 1326 17512 1331
rect 15872 1258 15883 1326
rect 15940 1321 17512 1326
rect 15940 1261 17453 1321
rect 15940 1258 17512 1261
rect 15872 1252 17512 1258
rect 19004 1330 20644 1335
rect 19004 1262 19015 1330
rect 19072 1325 20644 1330
rect 19072 1265 20585 1325
rect 19072 1262 20644 1265
rect 19004 1256 20644 1262
rect 19004 1253 19100 1256
rect 20585 1255 20644 1256
rect 22148 1330 23788 1335
rect 22148 1262 22159 1330
rect 22216 1325 23788 1330
rect 22216 1265 23729 1325
rect 22216 1262 23788 1265
rect 22148 1256 23788 1262
rect 22148 1253 22244 1256
rect 23729 1255 23788 1256
rect 19015 1252 19072 1253
rect 22159 1252 22216 1253
rect 15872 1249 15968 1252
rect 17453 1251 17512 1252
rect 117 1248 174 1249
rect 3261 1248 3318 1249
rect 12739 1248 12796 1249
rect 15883 1248 15940 1249
rect 6393 1171 6450 1172
rect 9537 1171 9594 1172
rect 19015 1171 19072 1172
rect 22159 1171 22216 1172
rect 6382 1170 6478 1171
rect 9526 1170 9622 1171
rect 19004 1170 19100 1171
rect 22148 1170 22244 1171
rect 117 1167 174 1168
rect 3261 1167 3318 1168
rect 106 1166 202 1167
rect 3250 1166 3346 1167
rect 106 1158 1407 1166
rect 106 1090 117 1158
rect 174 1093 1328 1158
rect 1396 1093 1407 1158
rect 174 1090 1407 1093
rect 106 1082 1407 1090
rect 3250 1158 4551 1166
rect 3250 1090 3261 1158
rect 3318 1093 4472 1158
rect 4540 1093 4551 1158
rect 3318 1090 4551 1093
rect 3250 1082 4551 1090
rect 6382 1162 7683 1170
rect 6382 1094 6393 1162
rect 6450 1097 7604 1162
rect 7672 1097 7683 1162
rect 6450 1094 7683 1097
rect 6382 1086 7683 1094
rect 9526 1162 10827 1170
rect 12739 1167 12796 1168
rect 15883 1167 15940 1168
rect 9526 1094 9537 1162
rect 9594 1097 10748 1162
rect 10816 1097 10827 1162
rect 9594 1094 10827 1097
rect 9526 1086 10827 1094
rect 12728 1166 12824 1167
rect 15872 1166 15968 1167
rect 12728 1158 14029 1166
rect 12728 1090 12739 1158
rect 12796 1093 13950 1158
rect 14018 1093 14029 1158
rect 12796 1090 14029 1093
rect 6393 1084 6450 1086
rect 9537 1084 9594 1086
rect 12728 1082 14029 1090
rect 15872 1158 17173 1166
rect 15872 1090 15883 1158
rect 15940 1093 17094 1158
rect 17162 1093 17173 1158
rect 15940 1090 17173 1093
rect 15872 1082 17173 1090
rect 19004 1162 20305 1170
rect 19004 1094 19015 1162
rect 19072 1097 20226 1162
rect 20294 1097 20305 1162
rect 19072 1094 20305 1097
rect 19004 1086 20305 1094
rect 22148 1162 23449 1170
rect 22148 1094 22159 1162
rect 22216 1097 23370 1162
rect 23438 1097 23449 1162
rect 22216 1094 23449 1097
rect 22148 1086 23449 1094
rect 19015 1084 19072 1086
rect 22159 1084 22216 1086
rect 117 1080 174 1082
rect 3261 1080 3318 1082
rect 12739 1080 12796 1082
rect 15883 1080 15940 1082
rect 1516 168 1592 178
rect 1516 100 1592 110
rect 4660 168 4736 178
rect 4660 100 4736 110
rect 7792 172 7868 182
rect 7792 104 7868 114
rect 10936 172 11012 182
rect 10936 104 11012 114
rect 14138 168 14214 178
rect 14138 100 14214 110
rect 17282 168 17358 178
rect 17282 100 17358 110
rect 20414 172 20490 182
rect 20414 104 20490 114
rect 23558 172 23634 182
rect 23558 104 23634 114
rect 1528 -1480 1628 -1470
rect 1528 -1582 1628 -1572
rect 4672 -1480 4772 -1470
rect 4672 -1582 4772 -1572
rect 7804 -1476 7904 -1466
rect 7804 -1578 7904 -1568
rect 10948 -1476 11048 -1466
rect 10948 -1578 11048 -1568
rect 14150 -1480 14250 -1470
rect 14150 -1582 14250 -1572
rect 17294 -1480 17394 -1470
rect 17294 -1582 17394 -1572
rect 20426 -1476 20526 -1466
rect 20426 -1578 20526 -1568
rect 23570 -1476 23670 -1466
rect 23570 -1578 23670 -1568
rect 6425 -2437 6482 -2436
rect 6658 -2437 6751 -2435
rect 9569 -2437 9626 -2436
rect 9802 -2437 9895 -2435
rect 19047 -2437 19104 -2436
rect 19280 -2437 19373 -2435
rect 22191 -2437 22248 -2436
rect 22424 -2437 22517 -2435
rect 6417 -2438 7833 -2437
rect 9561 -2438 10977 -2437
rect 19039 -2438 20455 -2437
rect 22183 -2438 23599 -2437
rect 149 -2441 206 -2440
rect 382 -2441 475 -2439
rect 3293 -2441 3350 -2440
rect 3526 -2441 3619 -2439
rect 141 -2442 1557 -2441
rect 3285 -2442 4701 -2441
rect 138 -2450 1557 -2442
rect 138 -2518 149 -2450
rect 206 -2451 1557 -2450
rect 206 -2514 393 -2451
rect 464 -2513 1478 -2451
rect 1548 -2513 1557 -2451
rect 464 -2514 1557 -2513
rect 206 -2518 1557 -2514
rect 138 -2525 1557 -2518
rect 3282 -2450 4701 -2442
rect 3282 -2518 3293 -2450
rect 3350 -2451 4701 -2450
rect 3350 -2514 3537 -2451
rect 3608 -2513 4622 -2451
rect 4692 -2513 4701 -2451
rect 3608 -2514 4701 -2513
rect 3350 -2518 4701 -2514
rect 3282 -2525 4701 -2518
rect 6414 -2446 7833 -2438
rect 6414 -2514 6425 -2446
rect 6482 -2447 7833 -2446
rect 6482 -2510 6669 -2447
rect 6740 -2509 7754 -2447
rect 7824 -2509 7833 -2447
rect 6740 -2510 7833 -2509
rect 6482 -2514 7833 -2510
rect 6414 -2521 7833 -2514
rect 9558 -2446 10977 -2438
rect 12771 -2441 12828 -2440
rect 13004 -2441 13097 -2439
rect 15915 -2441 15972 -2440
rect 16148 -2441 16241 -2439
rect 12763 -2442 14179 -2441
rect 15907 -2442 17323 -2441
rect 9558 -2514 9569 -2446
rect 9626 -2447 10977 -2446
rect 9626 -2510 9813 -2447
rect 9884 -2509 10898 -2447
rect 10968 -2509 10977 -2447
rect 9884 -2510 10977 -2509
rect 9626 -2514 10977 -2510
rect 9558 -2521 10977 -2514
rect 12760 -2450 14179 -2442
rect 12760 -2518 12771 -2450
rect 12828 -2451 14179 -2450
rect 12828 -2514 13015 -2451
rect 13086 -2513 14100 -2451
rect 14170 -2513 14179 -2451
rect 13086 -2514 14179 -2513
rect 12828 -2518 14179 -2514
rect 6414 -2522 6492 -2521
rect 9558 -2522 9636 -2521
rect 6425 -2524 6482 -2522
rect 9569 -2524 9626 -2522
rect 12760 -2525 14179 -2518
rect 15904 -2450 17323 -2442
rect 15904 -2518 15915 -2450
rect 15972 -2451 17323 -2450
rect 15972 -2514 16159 -2451
rect 16230 -2513 17244 -2451
rect 17314 -2513 17323 -2451
rect 16230 -2514 17323 -2513
rect 15972 -2518 17323 -2514
rect 15904 -2525 17323 -2518
rect 19036 -2446 20455 -2438
rect 19036 -2514 19047 -2446
rect 19104 -2447 20455 -2446
rect 19104 -2510 19291 -2447
rect 19362 -2509 20376 -2447
rect 20446 -2509 20455 -2447
rect 19362 -2510 20455 -2509
rect 19104 -2514 20455 -2510
rect 19036 -2521 20455 -2514
rect 22180 -2446 23599 -2438
rect 22180 -2514 22191 -2446
rect 22248 -2447 23599 -2446
rect 22248 -2510 22435 -2447
rect 22506 -2509 23520 -2447
rect 23590 -2509 23599 -2447
rect 22506 -2510 23599 -2509
rect 22248 -2514 23599 -2510
rect 22180 -2521 23599 -2514
rect 19036 -2522 19114 -2521
rect 22180 -2522 22258 -2521
rect 19047 -2524 19104 -2522
rect 22191 -2524 22248 -2522
rect 138 -2526 216 -2525
rect 3282 -2526 3360 -2525
rect 12760 -2526 12838 -2525
rect 15904 -2526 15982 -2525
rect 149 -2528 206 -2526
rect 3293 -2528 3350 -2526
rect 12771 -2528 12828 -2526
rect 15915 -2528 15972 -2526
rect 6425 -2554 6482 -2552
rect 9569 -2554 9626 -2552
rect 19047 -2554 19104 -2552
rect 22191 -2554 22248 -2552
rect 149 -2558 206 -2556
rect 3293 -2558 3350 -2556
rect 6414 -2557 6510 -2554
rect 9558 -2557 9654 -2554
rect 138 -2561 234 -2558
rect 3282 -2561 3378 -2558
rect 138 -2566 1778 -2561
rect 138 -2634 149 -2566
rect 206 -2571 1778 -2566
rect 206 -2631 1719 -2571
rect 206 -2634 1778 -2631
rect 138 -2640 1778 -2634
rect 138 -2643 234 -2640
rect 1719 -2641 1778 -2640
rect 3282 -2566 4922 -2561
rect 3282 -2634 3293 -2566
rect 3350 -2571 4922 -2566
rect 3350 -2631 4863 -2571
rect 3350 -2634 4922 -2631
rect 3282 -2640 4922 -2634
rect 6414 -2562 8054 -2557
rect 6414 -2630 6425 -2562
rect 6482 -2567 8054 -2562
rect 6482 -2627 7995 -2567
rect 6482 -2630 8054 -2627
rect 6414 -2636 8054 -2630
rect 6414 -2639 6510 -2636
rect 7995 -2637 8054 -2636
rect 9558 -2562 11198 -2557
rect 12771 -2558 12828 -2556
rect 15915 -2558 15972 -2556
rect 19036 -2557 19132 -2554
rect 22180 -2557 22276 -2554
rect 9558 -2630 9569 -2562
rect 9626 -2567 11198 -2562
rect 9626 -2627 11139 -2567
rect 9626 -2630 11198 -2627
rect 9558 -2636 11198 -2630
rect 9558 -2639 9654 -2636
rect 11139 -2637 11198 -2636
rect 12760 -2561 12856 -2558
rect 15904 -2561 16000 -2558
rect 12760 -2566 14400 -2561
rect 12760 -2634 12771 -2566
rect 12828 -2571 14400 -2566
rect 12828 -2631 14341 -2571
rect 12828 -2634 14400 -2631
rect 6425 -2640 6482 -2639
rect 9569 -2640 9626 -2639
rect 12760 -2640 14400 -2634
rect 3282 -2643 3378 -2640
rect 4863 -2641 4922 -2640
rect 12760 -2643 12856 -2640
rect 14341 -2641 14400 -2640
rect 15904 -2566 17544 -2561
rect 15904 -2634 15915 -2566
rect 15972 -2571 17544 -2566
rect 15972 -2631 17485 -2571
rect 15972 -2634 17544 -2631
rect 15904 -2640 17544 -2634
rect 19036 -2562 20676 -2557
rect 19036 -2630 19047 -2562
rect 19104 -2567 20676 -2562
rect 19104 -2627 20617 -2567
rect 19104 -2630 20676 -2627
rect 19036 -2636 20676 -2630
rect 19036 -2639 19132 -2636
rect 20617 -2637 20676 -2636
rect 22180 -2562 23820 -2557
rect 22180 -2630 22191 -2562
rect 22248 -2567 23820 -2562
rect 22248 -2627 23761 -2567
rect 22248 -2630 23820 -2627
rect 22180 -2636 23820 -2630
rect 22180 -2639 22276 -2636
rect 23761 -2637 23820 -2636
rect 19047 -2640 19104 -2639
rect 22191 -2640 22248 -2639
rect 15904 -2643 16000 -2640
rect 17485 -2641 17544 -2640
rect 149 -2644 206 -2643
rect 3293 -2644 3350 -2643
rect 12771 -2644 12828 -2643
rect 15915 -2644 15972 -2643
rect 6425 -2721 6482 -2720
rect 9569 -2721 9626 -2720
rect 19047 -2721 19104 -2720
rect 22191 -2721 22248 -2720
rect 6414 -2722 6510 -2721
rect 9558 -2722 9654 -2721
rect 19036 -2722 19132 -2721
rect 22180 -2722 22276 -2721
rect 149 -2725 206 -2724
rect 3293 -2725 3350 -2724
rect 138 -2726 234 -2725
rect 3282 -2726 3378 -2725
rect 138 -2734 1439 -2726
rect 138 -2802 149 -2734
rect 206 -2799 1360 -2734
rect 1428 -2799 1439 -2734
rect 206 -2802 1439 -2799
rect 138 -2810 1439 -2802
rect 3282 -2734 4583 -2726
rect 3282 -2802 3293 -2734
rect 3350 -2799 4504 -2734
rect 4572 -2799 4583 -2734
rect 3350 -2802 4583 -2799
rect 3282 -2810 4583 -2802
rect 6414 -2730 7715 -2722
rect 6414 -2798 6425 -2730
rect 6482 -2795 7636 -2730
rect 7704 -2795 7715 -2730
rect 6482 -2798 7715 -2795
rect 6414 -2806 7715 -2798
rect 9558 -2730 10859 -2722
rect 12771 -2725 12828 -2724
rect 15915 -2725 15972 -2724
rect 9558 -2798 9569 -2730
rect 9626 -2795 10780 -2730
rect 10848 -2795 10859 -2730
rect 9626 -2798 10859 -2795
rect 9558 -2806 10859 -2798
rect 12760 -2726 12856 -2725
rect 15904 -2726 16000 -2725
rect 12760 -2734 14061 -2726
rect 12760 -2802 12771 -2734
rect 12828 -2799 13982 -2734
rect 14050 -2799 14061 -2734
rect 12828 -2802 14061 -2799
rect 6425 -2808 6482 -2806
rect 9569 -2808 9626 -2806
rect 12760 -2810 14061 -2802
rect 15904 -2734 17205 -2726
rect 15904 -2802 15915 -2734
rect 15972 -2799 17126 -2734
rect 17194 -2799 17205 -2734
rect 15972 -2802 17205 -2799
rect 15904 -2810 17205 -2802
rect 19036 -2730 20337 -2722
rect 19036 -2798 19047 -2730
rect 19104 -2795 20258 -2730
rect 20326 -2795 20337 -2730
rect 19104 -2798 20337 -2795
rect 19036 -2806 20337 -2798
rect 22180 -2730 23481 -2722
rect 22180 -2798 22191 -2730
rect 22248 -2795 23402 -2730
rect 23470 -2795 23481 -2730
rect 22248 -2798 23481 -2795
rect 22180 -2806 23481 -2798
rect 19047 -2808 19104 -2806
rect 22191 -2808 22248 -2806
rect 149 -2812 206 -2810
rect 3293 -2812 3350 -2810
rect 12771 -2812 12828 -2810
rect 15915 -2812 15972 -2810
rect 1548 -3724 1624 -3714
rect 1548 -3792 1624 -3782
rect 4692 -3724 4768 -3714
rect 4692 -3792 4768 -3782
rect 7824 -3720 7900 -3710
rect 7824 -3788 7900 -3778
rect 10968 -3720 11044 -3710
rect 10968 -3788 11044 -3778
rect 14170 -3724 14246 -3714
rect 14170 -3792 14246 -3782
rect 17314 -3724 17390 -3714
rect 17314 -3792 17390 -3782
rect 20446 -3720 20522 -3710
rect 20446 -3788 20522 -3778
rect 23590 -3720 23666 -3710
rect 23590 -3788 23666 -3778
<< via2 >>
rect 1702 22236 1802 22264
rect 1702 22176 1714 22236
rect 1714 22176 1794 22236
rect 1794 22176 1802 22236
rect 1702 22172 1802 22176
rect 4846 22236 4946 22264
rect 4846 22176 4858 22236
rect 4858 22176 4938 22236
rect 4938 22176 4946 22236
rect 4846 22172 4946 22176
rect 7978 22240 8078 22268
rect 7978 22180 7990 22240
rect 7990 22180 8070 22240
rect 8070 22180 8078 22240
rect 7978 22176 8078 22180
rect 11122 22240 11222 22268
rect 11122 22180 11134 22240
rect 11134 22180 11214 22240
rect 11214 22180 11222 22240
rect 11122 22176 11222 22180
rect 14324 22236 14424 22264
rect 14324 22176 14336 22236
rect 14336 22176 14416 22236
rect 14416 22176 14424 22236
rect 14324 22172 14424 22176
rect 17468 22236 17568 22264
rect 17468 22176 17480 22236
rect 17480 22176 17560 22236
rect 17560 22176 17568 22236
rect 17468 22172 17568 22176
rect 20600 22240 20700 22268
rect 20600 22180 20612 22240
rect 20612 22180 20692 22240
rect 20692 22180 20700 22240
rect 20600 22176 20700 22180
rect 23744 22240 23844 22268
rect 23744 22180 23756 22240
rect 23756 22180 23836 22240
rect 23836 22180 23844 22240
rect 23744 22176 23844 22180
rect 322 21113 378 21169
rect 22354 20935 22433 21024
rect 18906 20672 18970 20731
rect 25537 20670 25603 20730
rect 15770 20509 15826 20578
rect 25527 20503 25591 20572
rect 12545 20359 12607 20427
rect 25527 20357 25591 20426
rect 9370 20222 9429 20279
rect 25527 20217 25591 20286
rect 6244 20096 6303 20162
rect 25526 20078 25590 20147
rect 1722 20018 1798 20020
rect 1722 19966 1728 20018
rect 1728 19966 1794 20018
rect 1794 19966 1798 20018
rect 1722 19962 1798 19966
rect 4866 20018 4942 20020
rect 4866 19966 4872 20018
rect 4872 19966 4938 20018
rect 4938 19966 4942 20018
rect 4866 19962 4942 19966
rect 7998 20022 8074 20024
rect 7998 19970 8004 20022
rect 8004 19970 8070 20022
rect 8070 19970 8074 20022
rect 7998 19966 8074 19970
rect 11142 20022 11218 20024
rect 11142 19970 11148 20022
rect 11148 19970 11214 20022
rect 11214 19970 11218 20022
rect 11142 19966 11218 19970
rect 14344 20018 14420 20020
rect 14344 19966 14350 20018
rect 14350 19966 14416 20018
rect 14416 19966 14420 20018
rect 14344 19962 14420 19966
rect 17488 20018 17564 20020
rect 17488 19966 17494 20018
rect 17494 19966 17560 20018
rect 17560 19966 17564 20018
rect 17488 19962 17564 19966
rect 20620 20022 20696 20024
rect 20620 19970 20626 20022
rect 20626 19970 20692 20022
rect 20692 19970 20696 20022
rect 20620 19966 20696 19970
rect 23764 20022 23840 20024
rect 23764 19970 23770 20022
rect 23770 19970 23836 20022
rect 23836 19970 23840 20022
rect 23764 19966 23840 19970
rect 3111 19801 3184 19882
rect 25526 19810 25590 19879
rect 3250 16775 3310 16837
rect 2415 16122 2486 16181
rect 2701 16021 2770 16085
rect 4698 16775 4758 16837
rect 4348 15881 4424 15899
rect 4348 15826 4359 15881
rect 4359 15826 4413 15881
rect 4413 15826 4424 15881
rect 4348 15812 4424 15826
rect 6196 16777 6256 16839
rect 5850 15879 5914 15891
rect 5850 15825 5857 15879
rect 5857 15825 5911 15879
rect 5911 15825 5914 15879
rect 7644 16777 7704 16839
rect 7299 15884 7366 15897
rect 7299 15830 7305 15884
rect 7305 15830 7359 15884
rect 7359 15830 7366 15884
rect 9164 16775 9224 16837
rect 8818 15884 8878 15895
rect 8818 15830 8821 15884
rect 8821 15830 8875 15884
rect 8875 15830 8878 15884
rect 5850 15817 5914 15825
rect 7299 15819 7366 15830
rect 8818 15820 8878 15830
rect 10612 16775 10672 16837
rect 10268 15878 10328 15888
rect 10268 15824 10273 15878
rect 10273 15824 10327 15878
rect 10327 15824 10328 15878
rect 12110 16777 12170 16839
rect 11767 15884 11828 15897
rect 11767 15830 11770 15884
rect 11770 15830 11824 15884
rect 11824 15830 11828 15884
rect 10268 15820 10328 15824
rect 11767 15818 11828 15830
rect 15222 17025 15312 17046
rect 15222 16973 15244 17025
rect 15244 16973 15296 17025
rect 15296 16973 15312 17025
rect 15222 16955 15312 16973
rect 16390 17025 16480 17046
rect 16390 16973 16412 17025
rect 16412 16973 16464 17025
rect 16464 16973 16480 17025
rect 16390 16955 16480 16973
rect 17558 17025 17648 17046
rect 17558 16973 17580 17025
rect 17580 16973 17632 17025
rect 17632 16973 17648 17025
rect 17558 16955 17648 16973
rect 18726 17025 18816 17046
rect 18726 16973 18748 17025
rect 18748 16973 18800 17025
rect 18800 16973 18816 17025
rect 18726 16955 18816 16973
rect 19900 17027 19990 17048
rect 19900 16975 19922 17027
rect 19922 16975 19974 17027
rect 19974 16975 19990 17027
rect 19900 16957 19990 16975
rect 21068 17027 21158 17048
rect 21068 16975 21090 17027
rect 21090 16975 21142 17027
rect 21142 16975 21158 17027
rect 21068 16957 21158 16975
rect 22236 17027 22326 17048
rect 22236 16975 22258 17027
rect 22258 16975 22310 17027
rect 22310 16975 22326 17027
rect 22236 16957 22326 16975
rect 23404 17027 23494 17048
rect 23404 16975 23426 17027
rect 23426 16975 23478 17027
rect 23478 16975 23494 17027
rect 23404 16957 23494 16975
rect 13558 16777 13618 16839
rect 13201 15901 13286 15902
rect 13201 15813 13286 15901
rect 13201 15812 13286 15813
rect 14757 15701 14847 15719
rect 14757 15649 14773 15701
rect 14773 15649 14825 15701
rect 14825 15649 14847 15701
rect 3472 15573 3534 15631
rect 3534 15573 3536 15631
rect 3472 15569 3536 15573
rect 4920 15573 4982 15631
rect 4982 15573 4984 15631
rect 4920 15569 4984 15573
rect 6418 15575 6480 15633
rect 6480 15575 6482 15633
rect 6418 15571 6482 15575
rect 7866 15575 7928 15633
rect 7928 15575 7930 15633
rect 7866 15571 7930 15575
rect 9386 15573 9448 15631
rect 9448 15573 9450 15631
rect 9386 15569 9450 15573
rect 10834 15573 10896 15631
rect 10896 15573 10898 15631
rect 10834 15569 10898 15573
rect 12332 15575 12394 15633
rect 12394 15575 12396 15633
rect 12332 15571 12396 15575
rect 13780 15575 13842 15633
rect 13842 15575 13844 15633
rect 14757 15628 14847 15649
rect 15925 15701 16015 15719
rect 15925 15649 15941 15701
rect 15941 15649 15993 15701
rect 15993 15649 16015 15701
rect 15925 15628 16015 15649
rect 17093 15701 17183 15719
rect 17093 15649 17109 15701
rect 17109 15649 17161 15701
rect 17161 15649 17183 15701
rect 17093 15628 17183 15649
rect 18261 15701 18351 15719
rect 18261 15649 18277 15701
rect 18277 15649 18329 15701
rect 18329 15649 18351 15701
rect 18261 15628 18351 15649
rect 19435 15703 19525 15721
rect 19435 15651 19451 15703
rect 19451 15651 19503 15703
rect 19503 15651 19525 15703
rect 19435 15630 19525 15651
rect 20603 15703 20693 15721
rect 20603 15651 20619 15703
rect 20619 15651 20671 15703
rect 20671 15651 20693 15703
rect 20603 15630 20693 15651
rect 21771 15703 21861 15721
rect 21771 15651 21787 15703
rect 21787 15651 21839 15703
rect 21839 15651 21861 15703
rect 21771 15630 21861 15651
rect 22939 15703 23029 15721
rect 22939 15651 22955 15703
rect 22955 15651 23007 15703
rect 23007 15651 23029 15703
rect 22939 15630 23029 15651
rect 13780 15571 13844 15575
rect 181 15505 239 15506
rect 181 15451 182 15505
rect 182 15451 238 15505
rect 238 15451 239 15505
rect 181 15450 239 15451
rect 4204 15098 4304 15126
rect 4204 15038 4216 15098
rect 4216 15038 4296 15098
rect 4296 15038 4304 15098
rect 4204 15034 4304 15038
rect 7348 15098 7448 15126
rect 7348 15038 7360 15098
rect 7360 15038 7440 15098
rect 7440 15038 7448 15098
rect 7348 15034 7448 15038
rect 10480 15102 10580 15130
rect 10480 15042 10492 15102
rect 10492 15042 10572 15102
rect 10572 15042 10580 15102
rect 10480 15038 10580 15042
rect 13624 15102 13724 15130
rect 13624 15042 13636 15102
rect 13636 15042 13716 15102
rect 13716 15042 13724 15102
rect 13624 15038 13724 15042
rect 16826 15098 16926 15126
rect 16826 15038 16838 15098
rect 16838 15038 16918 15098
rect 16918 15038 16926 15098
rect 16826 15034 16926 15038
rect 19970 15098 20070 15126
rect 19970 15038 19982 15098
rect 19982 15038 20062 15098
rect 20062 15038 20070 15098
rect 19970 15034 20070 15038
rect 23102 15102 23202 15130
rect 23102 15042 23114 15102
rect 23114 15042 23194 15102
rect 23194 15042 23202 15102
rect 23102 15038 23202 15042
rect 26246 15102 26346 15130
rect 26246 15042 26258 15102
rect 26258 15042 26338 15102
rect 26338 15042 26346 15102
rect 26246 15038 26346 15042
rect 4224 12880 4300 12882
rect 4224 12828 4230 12880
rect 4230 12828 4296 12880
rect 4296 12828 4300 12880
rect 4224 12824 4300 12828
rect 7368 12880 7444 12882
rect 7368 12828 7374 12880
rect 7374 12828 7440 12880
rect 7440 12828 7444 12880
rect 7368 12824 7444 12828
rect 10500 12884 10576 12886
rect 10500 12832 10506 12884
rect 10506 12832 10572 12884
rect 10572 12832 10576 12884
rect 10500 12828 10576 12832
rect 13644 12884 13720 12886
rect 13644 12832 13650 12884
rect 13650 12832 13716 12884
rect 13716 12832 13720 12884
rect 13644 12828 13720 12832
rect 16846 12880 16922 12882
rect 16846 12828 16852 12880
rect 16852 12828 16918 12880
rect 16918 12828 16922 12880
rect 16846 12824 16922 12828
rect 19990 12880 20066 12882
rect 19990 12828 19996 12880
rect 19996 12828 20062 12880
rect 20062 12828 20066 12880
rect 19990 12824 20066 12828
rect 23122 12884 23198 12886
rect 23122 12832 23128 12884
rect 23128 12832 23194 12884
rect 23194 12832 23198 12884
rect 23122 12828 23198 12832
rect 26266 12884 26342 12886
rect 26266 12832 26272 12884
rect 26272 12832 26338 12884
rect 26338 12832 26342 12884
rect 26266 12828 26342 12832
rect 4204 12364 4304 12392
rect 4204 12304 4216 12364
rect 4216 12304 4296 12364
rect 4296 12304 4304 12364
rect 4204 12300 4304 12304
rect 7348 12364 7448 12392
rect 7348 12304 7360 12364
rect 7360 12304 7440 12364
rect 7440 12304 7448 12364
rect 7348 12300 7448 12304
rect 10480 12368 10580 12396
rect 10480 12308 10492 12368
rect 10492 12308 10572 12368
rect 10572 12308 10580 12368
rect 10480 12304 10580 12308
rect 13624 12368 13724 12396
rect 13624 12308 13636 12368
rect 13636 12308 13716 12368
rect 13716 12308 13724 12368
rect 13624 12304 13724 12308
rect 16826 12364 16926 12392
rect 16826 12304 16838 12364
rect 16838 12304 16918 12364
rect 16918 12304 16926 12364
rect 16826 12300 16926 12304
rect 19970 12364 20070 12392
rect 19970 12304 19982 12364
rect 19982 12304 20062 12364
rect 20062 12304 20070 12364
rect 19970 12300 20070 12304
rect 23102 12368 23202 12396
rect 23102 12308 23114 12368
rect 23114 12308 23194 12368
rect 23194 12308 23202 12368
rect 23102 12304 23202 12308
rect 26246 12368 26346 12396
rect 26246 12308 26258 12368
rect 26258 12308 26338 12368
rect 26338 12308 26346 12368
rect 26246 12304 26346 12308
rect 4224 10146 4300 10148
rect 4224 10094 4230 10146
rect 4230 10094 4296 10146
rect 4296 10094 4300 10146
rect 4224 10090 4300 10094
rect 4194 9632 4294 9660
rect 4194 9572 4206 9632
rect 4206 9572 4286 9632
rect 4286 9572 4294 9632
rect 4194 9568 4294 9572
rect 7368 10146 7444 10148
rect 7368 10094 7374 10146
rect 7374 10094 7440 10146
rect 7440 10094 7444 10146
rect 10500 10150 10576 10152
rect 7368 10090 7444 10094
rect 10500 10098 10506 10150
rect 10506 10098 10572 10150
rect 10572 10098 10576 10150
rect 10500 10094 10576 10098
rect 13644 10150 13720 10152
rect 13644 10098 13650 10150
rect 13650 10098 13716 10150
rect 13716 10098 13720 10150
rect 13644 10094 13720 10098
rect 16846 10146 16922 10148
rect 16846 10094 16852 10146
rect 16852 10094 16918 10146
rect 16918 10094 16922 10146
rect 16846 10090 16922 10094
rect 19990 10146 20066 10148
rect 19990 10094 19996 10146
rect 19996 10094 20062 10146
rect 20062 10094 20066 10146
rect 19990 10090 20066 10094
rect 23122 10150 23198 10152
rect 23122 10098 23128 10150
rect 23128 10098 23194 10150
rect 23194 10098 23198 10150
rect 23122 10094 23198 10098
rect 26266 10150 26342 10152
rect 26266 10098 26272 10150
rect 26272 10098 26338 10150
rect 26338 10098 26342 10150
rect 26266 10094 26342 10098
rect 7338 9632 7438 9660
rect 7338 9572 7350 9632
rect 7350 9572 7430 9632
rect 7430 9572 7438 9632
rect 7338 9568 7438 9572
rect 10470 9636 10570 9664
rect 10470 9576 10482 9636
rect 10482 9576 10562 9636
rect 10562 9576 10570 9636
rect 10470 9572 10570 9576
rect 13614 9636 13714 9664
rect 13614 9576 13626 9636
rect 13626 9576 13706 9636
rect 13706 9576 13714 9636
rect 13614 9572 13714 9576
rect 16816 9632 16916 9660
rect 16816 9572 16828 9632
rect 16828 9572 16908 9632
rect 16908 9572 16916 9632
rect 16816 9568 16916 9572
rect 19960 9632 20060 9660
rect 19960 9572 19972 9632
rect 19972 9572 20052 9632
rect 20052 9572 20060 9632
rect 19960 9568 20060 9572
rect 23092 9636 23192 9664
rect 23092 9576 23104 9636
rect 23104 9576 23184 9636
rect 23184 9576 23192 9636
rect 23092 9572 23192 9576
rect 26236 9636 26336 9664
rect 26236 9576 26248 9636
rect 26248 9576 26328 9636
rect 26328 9576 26336 9636
rect 26236 9572 26336 9576
rect 4214 7414 4290 7416
rect 4214 7362 4220 7414
rect 4220 7362 4286 7414
rect 4286 7362 4290 7414
rect 4214 7358 4290 7362
rect 7358 7414 7434 7416
rect 7358 7362 7364 7414
rect 7364 7362 7430 7414
rect 7430 7362 7434 7414
rect 7358 7358 7434 7362
rect 10490 7418 10566 7420
rect 10490 7366 10496 7418
rect 10496 7366 10562 7418
rect 10562 7366 10566 7418
rect 10490 7362 10566 7366
rect 13634 7418 13710 7420
rect 13634 7366 13640 7418
rect 13640 7366 13706 7418
rect 13706 7366 13710 7418
rect 13634 7362 13710 7366
rect 16836 7414 16912 7416
rect 16836 7362 16842 7414
rect 16842 7362 16908 7414
rect 16908 7362 16912 7414
rect 16836 7358 16912 7362
rect 19980 7414 20056 7416
rect 19980 7362 19986 7414
rect 19986 7362 20052 7414
rect 20052 7362 20056 7414
rect 19980 7358 20056 7362
rect 23112 7418 23188 7420
rect 23112 7366 23118 7418
rect 23118 7366 23184 7418
rect 23184 7366 23188 7418
rect 23112 7362 23188 7366
rect 26256 7418 26332 7420
rect 26256 7366 26262 7418
rect 26262 7366 26328 7418
rect 26328 7366 26332 7418
rect 26256 7362 26332 7366
rect 19577 6753 19671 6763
rect 3510 6694 3588 6702
rect 3510 6640 3522 6694
rect 3522 6640 3576 6694
rect 3576 6640 3588 6694
rect 3510 6632 3588 6640
rect 5578 6696 5656 6704
rect 5578 6642 5590 6696
rect 5590 6642 5644 6696
rect 5644 6642 5656 6696
rect 5578 6634 5656 6642
rect 7647 6694 7725 6702
rect 7647 6640 7659 6694
rect 7659 6640 7713 6694
rect 7713 6640 7725 6694
rect 7647 6632 7725 6640
rect 9715 6696 9793 6704
rect 9715 6642 9727 6696
rect 9727 6642 9781 6696
rect 9781 6642 9793 6696
rect 9715 6634 9793 6642
rect 11784 6696 11862 6704
rect 11784 6642 11796 6696
rect 11796 6642 11850 6696
rect 11850 6642 11862 6696
rect 11784 6634 11862 6642
rect 13852 6698 13930 6706
rect 13852 6644 13864 6698
rect 13864 6644 13918 6698
rect 13918 6644 13930 6698
rect 13852 6636 13930 6644
rect 15921 6696 15999 6704
rect 15921 6642 15933 6696
rect 15933 6642 15987 6696
rect 15987 6642 15999 6696
rect 15921 6634 15999 6642
rect 17989 6698 18067 6706
rect 17989 6644 18001 6698
rect 18001 6644 18055 6698
rect 18055 6644 18067 6698
rect 19577 6679 19585 6753
rect 19585 6679 19661 6753
rect 19661 6679 19671 6753
rect 20315 6751 20409 6761
rect 20315 6677 20323 6751
rect 20323 6677 20399 6751
rect 20399 6677 20409 6751
rect 21053 6751 21147 6761
rect 21053 6677 21061 6751
rect 21061 6677 21137 6751
rect 21137 6677 21147 6751
rect 21795 6751 21889 6761
rect 21795 6677 21803 6751
rect 21803 6677 21879 6751
rect 21879 6677 21889 6751
rect 22535 6751 22629 6761
rect 22535 6677 22543 6751
rect 22543 6677 22619 6751
rect 22619 6677 22629 6751
rect 23273 6751 23367 6761
rect 23273 6677 23281 6751
rect 23281 6677 23357 6751
rect 23357 6677 23367 6751
rect 24011 6751 24105 6761
rect 24011 6677 24019 6751
rect 24019 6677 24095 6751
rect 24095 6677 24105 6751
rect 24749 6751 24843 6761
rect 24749 6677 24757 6751
rect 24757 6677 24833 6751
rect 24833 6677 24843 6751
rect 17989 6636 18067 6644
rect 4777 5894 4852 5910
rect 2426 5885 2492 5886
rect 2426 5832 2428 5885
rect 2428 5832 2488 5885
rect 2488 5832 2492 5885
rect 2426 5829 2492 5832
rect 4777 5828 4782 5894
rect 4782 5828 4848 5894
rect 4848 5828 4852 5894
rect 10988 5894 11055 5896
rect 4777 5824 4852 5828
rect 6848 5826 6851 5892
rect 6851 5826 6917 5892
rect 8920 5828 8984 5893
rect 10988 5828 11054 5894
rect 11054 5828 11055 5894
rect 13051 5830 13056 5896
rect 13056 5830 13116 5896
rect 17186 5896 17269 5905
rect 13051 5828 13116 5830
rect 15122 5829 15125 5893
rect 15125 5829 15189 5893
rect 17186 5830 17193 5896
rect 17193 5830 17259 5896
rect 17259 5830 17269 5896
rect 10988 5827 11055 5828
rect 17186 5825 17269 5830
rect 19525 5807 19591 5865
rect 20263 5805 20329 5863
rect 21001 5805 21067 5863
rect 21743 5805 21809 5863
rect 22483 5805 22549 5863
rect 23221 5805 23287 5863
rect 23959 5805 24025 5863
rect 24697 5805 24763 5863
rect 2699 5627 2770 5704
rect 3458 4470 3530 4472
rect 3458 4412 3464 4470
rect 3464 4412 3526 4470
rect 3526 4412 3530 4470
rect 3458 4402 3530 4412
rect 5526 4472 5598 4474
rect 5526 4414 5532 4472
rect 5532 4414 5594 4472
rect 5594 4414 5598 4472
rect 5526 4404 5598 4414
rect 7595 4470 7667 4472
rect 7595 4412 7601 4470
rect 7601 4412 7663 4470
rect 7663 4412 7667 4470
rect 7595 4402 7667 4412
rect 9663 4472 9735 4474
rect 9663 4414 9669 4472
rect 9669 4414 9731 4472
rect 9731 4414 9735 4472
rect 9663 4404 9735 4414
rect 11732 4472 11804 4474
rect 11732 4414 11738 4472
rect 11738 4414 11800 4472
rect 11800 4414 11804 4472
rect 11732 4404 11804 4414
rect 13800 4474 13872 4476
rect 13800 4416 13806 4474
rect 13806 4416 13868 4474
rect 13868 4416 13872 4474
rect 13800 4406 13872 4416
rect 15869 4472 15941 4474
rect 15869 4414 15875 4472
rect 15875 4414 15937 4472
rect 15937 4414 15941 4472
rect 15869 4404 15941 4414
rect 17937 4474 18009 4476
rect 17937 4416 17943 4474
rect 17943 4416 18005 4474
rect 18005 4416 18009 4474
rect 17937 4406 18009 4416
rect 1496 2384 1596 2412
rect 1496 2324 1508 2384
rect 1508 2324 1588 2384
rect 1588 2324 1596 2384
rect 1496 2320 1596 2324
rect 4640 2384 4740 2412
rect 4640 2324 4652 2384
rect 4652 2324 4732 2384
rect 4732 2324 4740 2384
rect 4640 2320 4740 2324
rect 7772 2388 7872 2416
rect 7772 2328 7784 2388
rect 7784 2328 7864 2388
rect 7864 2328 7872 2388
rect 7772 2324 7872 2328
rect 10916 2388 11016 2416
rect 10916 2328 10928 2388
rect 10928 2328 11008 2388
rect 11008 2328 11016 2388
rect 10916 2324 11016 2328
rect 14118 2384 14218 2412
rect 14118 2324 14130 2384
rect 14130 2324 14210 2384
rect 14210 2324 14218 2384
rect 14118 2320 14218 2324
rect 17262 2384 17362 2412
rect 17262 2324 17274 2384
rect 17274 2324 17354 2384
rect 17354 2324 17362 2384
rect 17262 2320 17362 2324
rect 20394 2388 20494 2416
rect 20394 2328 20406 2388
rect 20406 2328 20486 2388
rect 20486 2328 20494 2388
rect 20394 2324 20494 2328
rect 23538 2388 23638 2416
rect 23538 2328 23550 2388
rect 23550 2328 23630 2388
rect 23630 2328 23638 2388
rect 23538 2324 23638 2328
rect 1516 166 1592 168
rect 1516 114 1522 166
rect 1522 114 1588 166
rect 1588 114 1592 166
rect 1516 110 1592 114
rect 4660 166 4736 168
rect 4660 114 4666 166
rect 4666 114 4732 166
rect 4732 114 4736 166
rect 4660 110 4736 114
rect 7792 170 7868 172
rect 7792 118 7798 170
rect 7798 118 7864 170
rect 7864 118 7868 170
rect 7792 114 7868 118
rect 10936 170 11012 172
rect 10936 118 10942 170
rect 10942 118 11008 170
rect 11008 118 11012 170
rect 10936 114 11012 118
rect 14138 166 14214 168
rect 14138 114 14144 166
rect 14144 114 14210 166
rect 14210 114 14214 166
rect 14138 110 14214 114
rect 17282 166 17358 168
rect 17282 114 17288 166
rect 17288 114 17354 166
rect 17354 114 17358 166
rect 17282 110 17358 114
rect 20414 170 20490 172
rect 20414 118 20420 170
rect 20420 118 20486 170
rect 20486 118 20490 170
rect 20414 114 20490 118
rect 23558 170 23634 172
rect 23558 118 23564 170
rect 23564 118 23630 170
rect 23630 118 23634 170
rect 23558 114 23634 118
rect 1528 -1508 1628 -1480
rect 1528 -1568 1540 -1508
rect 1540 -1568 1620 -1508
rect 1620 -1568 1628 -1508
rect 1528 -1572 1628 -1568
rect 4672 -1508 4772 -1480
rect 4672 -1568 4684 -1508
rect 4684 -1568 4764 -1508
rect 4764 -1568 4772 -1508
rect 4672 -1572 4772 -1568
rect 7804 -1504 7904 -1476
rect 7804 -1564 7816 -1504
rect 7816 -1564 7896 -1504
rect 7896 -1564 7904 -1504
rect 7804 -1568 7904 -1564
rect 10948 -1504 11048 -1476
rect 10948 -1564 10960 -1504
rect 10960 -1564 11040 -1504
rect 11040 -1564 11048 -1504
rect 10948 -1568 11048 -1564
rect 14150 -1508 14250 -1480
rect 14150 -1568 14162 -1508
rect 14162 -1568 14242 -1508
rect 14242 -1568 14250 -1508
rect 14150 -1572 14250 -1568
rect 17294 -1508 17394 -1480
rect 17294 -1568 17306 -1508
rect 17306 -1568 17386 -1508
rect 17386 -1568 17394 -1508
rect 17294 -1572 17394 -1568
rect 20426 -1504 20526 -1476
rect 20426 -1564 20438 -1504
rect 20438 -1564 20518 -1504
rect 20518 -1564 20526 -1504
rect 20426 -1568 20526 -1564
rect 23570 -1504 23670 -1476
rect 23570 -1564 23582 -1504
rect 23582 -1564 23662 -1504
rect 23662 -1564 23670 -1504
rect 23570 -1568 23670 -1564
rect 1548 -3726 1624 -3724
rect 1548 -3778 1554 -3726
rect 1554 -3778 1620 -3726
rect 1620 -3778 1624 -3726
rect 1548 -3782 1624 -3778
rect 4692 -3726 4768 -3724
rect 4692 -3778 4698 -3726
rect 4698 -3778 4764 -3726
rect 4764 -3778 4768 -3726
rect 4692 -3782 4768 -3778
rect 7824 -3722 7900 -3720
rect 7824 -3774 7830 -3722
rect 7830 -3774 7896 -3722
rect 7896 -3774 7900 -3722
rect 7824 -3778 7900 -3774
rect 10968 -3722 11044 -3720
rect 10968 -3774 10974 -3722
rect 10974 -3774 11040 -3722
rect 11040 -3774 11044 -3722
rect 10968 -3778 11044 -3774
rect 14170 -3726 14246 -3724
rect 14170 -3778 14176 -3726
rect 14176 -3778 14242 -3726
rect 14242 -3778 14246 -3726
rect 14170 -3782 14246 -3778
rect 17314 -3726 17390 -3724
rect 17314 -3778 17320 -3726
rect 17320 -3778 17386 -3726
rect 17386 -3778 17390 -3726
rect 17314 -3782 17390 -3778
rect 20446 -3722 20522 -3720
rect 20446 -3774 20452 -3722
rect 20452 -3774 20518 -3722
rect 20518 -3774 20522 -3722
rect 20446 -3778 20522 -3774
rect 23590 -3722 23666 -3720
rect 23590 -3774 23596 -3722
rect 23596 -3774 23662 -3722
rect 23662 -3774 23666 -3722
rect 23590 -3778 23666 -3774
<< metal3 >>
rect 1692 22264 1812 22269
rect 1692 22170 1702 22264
rect 1802 22170 1812 22264
rect 1692 22167 1812 22170
rect 4836 22264 4956 22269
rect 4836 22170 4846 22264
rect 4946 22170 4956 22264
rect 7968 22268 8088 22273
rect 7968 22174 7978 22268
rect 8078 22174 8088 22268
rect 7968 22171 8088 22174
rect 11112 22268 11232 22273
rect 11112 22174 11122 22268
rect 11222 22174 11232 22268
rect 11112 22171 11232 22174
rect 14314 22264 14434 22269
rect 4836 22167 4956 22170
rect 14314 22170 14324 22264
rect 14424 22170 14434 22264
rect 14314 22167 14434 22170
rect 17458 22264 17578 22269
rect 17458 22170 17468 22264
rect 17568 22170 17578 22264
rect 20590 22268 20710 22273
rect 20590 22174 20600 22268
rect 20700 22174 20710 22268
rect 20590 22171 20710 22174
rect 23734 22268 23854 22273
rect 23734 22174 23744 22268
rect 23844 22174 23854 22268
rect 23734 22171 23854 22174
rect 17458 22167 17578 22170
rect 302 21183 399 21184
rect 302 21100 312 21183
rect 389 21100 399 21183
rect 302 21081 399 21100
rect 22333 20925 22343 21034
rect 22443 20925 22453 21034
rect 18896 20735 25609 20736
rect 18896 20731 25613 20735
rect 18896 20672 18906 20731
rect 18970 20730 25613 20731
rect 18970 20672 25537 20730
rect 18896 20670 25537 20672
rect 25603 20670 25613 20730
rect 18896 20667 25613 20670
rect 25527 20665 25613 20667
rect 15760 20578 15836 20583
rect 15760 20509 15770 20578
rect 15826 20572 15836 20578
rect 25517 20572 25601 20577
rect 15826 20509 25527 20572
rect 15760 20504 25527 20509
rect 25517 20503 25527 20504
rect 25591 20503 25601 20572
rect 25517 20498 25601 20503
rect 12535 20427 12617 20432
rect 12535 20359 12545 20427
rect 12607 20426 12617 20427
rect 25517 20426 25601 20431
rect 12607 20359 25527 20426
rect 12535 20358 25527 20359
rect 12535 20354 12617 20358
rect 25517 20357 25527 20358
rect 25591 20357 25601 20426
rect 25517 20352 25601 20357
rect 25517 20286 25601 20291
rect 9415 20284 25527 20286
rect 9360 20279 25527 20284
rect 9360 20222 9370 20279
rect 9429 20222 25527 20279
rect 9360 20218 25527 20222
rect 9360 20217 9439 20218
rect 25517 20217 25527 20218
rect 25591 20217 25601 20286
rect 25517 20212 25601 20217
rect 6234 20162 6313 20167
rect 6234 20096 6244 20162
rect 6303 20153 6313 20162
rect 23980 20153 25389 20158
rect 6303 20148 25389 20153
rect 25456 20148 25600 20152
rect 6303 20147 25600 20148
rect 6303 20096 25526 20147
rect 6234 20092 25526 20096
rect 6234 20091 6313 20092
rect 23980 20084 25526 20092
rect 25424 20079 25526 20084
rect 25516 20078 25526 20079
rect 25590 20078 25600 20147
rect 25516 20073 25600 20078
rect 1682 20020 1848 20028
rect 1682 19952 1716 20020
rect 1800 19952 1848 20020
rect 1682 19948 1848 19952
rect 4826 20020 4992 20028
rect 4826 19952 4860 20020
rect 4944 19952 4992 20020
rect 7958 20024 8124 20032
rect 7958 19956 7992 20024
rect 8076 19956 8124 20024
rect 7958 19952 8124 19956
rect 11102 20024 11268 20032
rect 11102 19956 11136 20024
rect 11220 19956 11268 20024
rect 11102 19952 11268 19956
rect 14304 20020 14470 20028
rect 14304 19952 14338 20020
rect 14422 19952 14470 20020
rect 4826 19948 4992 19952
rect 14304 19948 14470 19952
rect 17448 20020 17614 20028
rect 17448 19952 17482 20020
rect 17566 19952 17614 20020
rect 20580 20024 20746 20032
rect 20580 19956 20614 20024
rect 20698 19956 20746 20024
rect 20580 19952 20746 19956
rect 23724 20024 23890 20032
rect 23724 19956 23758 20024
rect 23842 19956 23890 20024
rect 23724 19952 23890 19956
rect 17448 19948 17614 19952
rect 3101 19882 3194 19887
rect 25433 19882 25600 19884
rect 3101 19801 3111 19882
rect 3184 19879 25600 19882
rect 3184 19810 25526 19879
rect 25590 19810 25600 19879
rect 3184 19805 25600 19810
rect 3184 19802 25540 19805
rect 3184 19801 3194 19802
rect 3101 19796 3194 19801
rect 15194 16940 15204 17060
rect 15326 16940 15336 17060
rect 16362 17046 16504 17060
rect 16362 16955 16390 17046
rect 16480 16955 16504 17046
rect 16362 16940 16504 16955
rect 17530 17046 17672 17060
rect 17530 16955 17558 17046
rect 17648 16955 17672 17046
rect 17530 16940 17672 16955
rect 18698 17046 18840 17060
rect 18698 16955 18726 17046
rect 18816 16955 18840 17046
rect 18698 16940 18840 16955
rect 19872 17048 20014 17062
rect 19872 16957 19900 17048
rect 19990 16957 20014 17048
rect 19872 16942 20014 16957
rect 21040 17048 21182 17062
rect 21040 16957 21068 17048
rect 21158 16957 21182 17048
rect 21040 16942 21182 16957
rect 22208 17048 22350 17062
rect 22208 16957 22236 17048
rect 22326 16957 22350 17048
rect 22208 16942 22350 16957
rect 23376 17048 23518 17062
rect 23376 16957 23404 17048
rect 23494 16957 23518 17048
rect 23376 16942 23518 16957
rect 3234 16841 3332 16859
rect 3234 16769 3244 16841
rect 3314 16769 3332 16841
rect 3234 16761 3332 16769
rect 4682 16841 4780 16859
rect 4682 16769 4692 16841
rect 4762 16769 4780 16841
rect 4682 16761 4780 16769
rect 6180 16843 6278 16861
rect 6180 16771 6190 16843
rect 6260 16771 6278 16843
rect 6180 16763 6278 16771
rect 7628 16843 7726 16861
rect 7628 16771 7638 16843
rect 7708 16771 7726 16843
rect 7628 16763 7726 16771
rect 9148 16841 9246 16859
rect 9148 16769 9158 16841
rect 9228 16769 9246 16841
rect 9148 16761 9246 16769
rect 10596 16841 10694 16859
rect 10596 16769 10606 16841
rect 10676 16769 10694 16841
rect 10596 16761 10694 16769
rect 12094 16843 12192 16861
rect 12094 16771 12104 16843
rect 12174 16771 12192 16843
rect 12094 16763 12192 16771
rect 13542 16843 13640 16861
rect 13542 16771 13552 16843
rect 13622 16771 13640 16843
rect 13542 16763 13640 16771
rect 2415 16186 2487 16191
rect 2405 16181 2496 16186
rect 2405 16122 2415 16181
rect 2486 16122 2496 16181
rect 2405 16117 2496 16122
rect 171 15509 249 15511
rect 2415 15509 2487 16117
rect 2691 16085 2780 16090
rect 2691 16021 2701 16085
rect 2770 16021 2780 16085
rect 2691 16016 2780 16021
rect 171 15506 2487 15509
rect 171 15450 181 15506
rect 239 15450 2487 15506
rect 171 15447 2487 15450
rect 171 15445 249 15447
rect 2415 5891 2487 15447
rect 2415 5886 2502 5891
rect 2415 5829 2426 5886
rect 2492 5829 2502 5886
rect 2415 5824 2502 5829
rect 2415 5815 2487 5824
rect 2699 5749 2771 16016
rect 4338 15899 4824 15911
rect 11757 15903 12618 15905
rect 4338 15812 4348 15899
rect 4424 15812 4824 15899
rect 4338 15806 4824 15812
rect 5837 15891 6902 15902
rect 5837 15817 5850 15891
rect 5914 15817 6902 15891
rect 5837 15811 6902 15817
rect 3452 15637 3554 15653
rect 3452 15569 3466 15637
rect 3540 15569 3554 15637
rect 3452 15555 3554 15569
rect 4194 15126 4314 15131
rect 4194 15032 4204 15126
rect 4304 15032 4314 15126
rect 4194 15029 4314 15032
rect 4184 12882 4350 12890
rect 4184 12814 4218 12882
rect 4302 12814 4350 12882
rect 4184 12810 4350 12814
rect 4194 12392 4314 12397
rect 4194 12298 4204 12392
rect 4304 12298 4314 12392
rect 4194 12295 4314 12298
rect 4184 10148 4350 10156
rect 4184 10080 4218 10148
rect 4302 10080 4350 10148
rect 4184 10076 4350 10080
rect 4184 9660 4304 9665
rect 4184 9566 4194 9660
rect 4294 9566 4304 9660
rect 4184 9563 4304 9566
rect 4174 7416 4340 7424
rect 4174 7348 4208 7416
rect 4292 7348 4340 7416
rect 4174 7344 4340 7348
rect 3440 6704 3654 6708
rect 3440 6632 3510 6704
rect 3586 6702 3654 6704
rect 3588 6632 3654 6702
rect 3440 6630 3654 6632
rect 3500 6627 3598 6630
rect 4759 5915 4824 15806
rect 4900 15637 5002 15653
rect 4900 15569 4914 15637
rect 4988 15569 5002 15637
rect 4900 15555 5002 15569
rect 6398 15639 6500 15655
rect 6398 15571 6412 15639
rect 6486 15571 6500 15639
rect 6398 15557 6500 15571
rect 5508 6706 5722 6710
rect 5508 6634 5578 6706
rect 5654 6704 5722 6706
rect 5656 6634 5722 6704
rect 5508 6632 5722 6634
rect 5568 6629 5666 6632
rect 4759 5910 4862 5915
rect 4759 5824 4777 5910
rect 4852 5824 4862 5910
rect 4759 5819 4862 5824
rect 6838 5897 6902 15811
rect 7289 15897 7376 15902
rect 9058 15900 9124 15901
rect 7289 15819 7299 15897
rect 7366 15819 7376 15897
rect 7289 15682 7376 15819
rect 8808 15895 9124 15900
rect 8808 15820 8818 15895
rect 8878 15820 9124 15895
rect 11757 15897 12673 15903
rect 10335 15893 11353 15894
rect 8808 15816 9124 15820
rect 8808 15815 8888 15816
rect 7290 15481 7376 15682
rect 7846 15639 7948 15655
rect 7846 15571 7860 15639
rect 7934 15571 7948 15639
rect 7846 15557 7948 15571
rect 7290 15409 8976 15481
rect 7338 15126 7458 15131
rect 7338 15032 7348 15126
rect 7448 15032 7458 15126
rect 7338 15029 7458 15032
rect 7328 12882 7494 12890
rect 7328 12814 7362 12882
rect 7446 12814 7494 12882
rect 7328 12810 7494 12814
rect 7338 12392 7458 12397
rect 7338 12298 7348 12392
rect 7448 12298 7458 12392
rect 7338 12295 7458 12298
rect 7328 10148 7494 10156
rect 7328 10080 7362 10148
rect 7446 10080 7494 10148
rect 7328 10076 7494 10080
rect 7328 9660 7448 9665
rect 7328 9566 7338 9660
rect 7438 9566 7448 9660
rect 7328 9563 7448 9566
rect 7318 7416 7484 7424
rect 7318 7348 7352 7416
rect 7436 7348 7484 7416
rect 7318 7344 7484 7348
rect 7577 6704 7791 6708
rect 7577 6632 7647 6704
rect 7723 6702 7791 6704
rect 7725 6632 7791 6702
rect 7577 6630 7791 6632
rect 7637 6627 7735 6630
rect 8909 5898 8976 15409
rect 9058 15451 9124 15816
rect 10258 15888 11353 15893
rect 10258 15820 10268 15888
rect 10328 15820 11353 15888
rect 10258 15816 11353 15820
rect 10258 15815 10338 15816
rect 9366 15637 9468 15653
rect 9366 15569 9380 15637
rect 9454 15569 9468 15637
rect 9366 15555 9468 15569
rect 10814 15637 10916 15653
rect 10814 15569 10828 15637
rect 10902 15569 10916 15637
rect 10814 15555 10916 15569
rect 11271 15460 11353 15816
rect 11757 15818 11767 15897
rect 11828 15818 12673 15897
rect 11757 15813 12673 15818
rect 12610 15667 12673 15813
rect 13191 15902 13296 15907
rect 13191 15812 13201 15902
rect 13286 15894 13296 15902
rect 16559 15894 16644 15895
rect 13286 15817 16644 15894
rect 13286 15812 13296 15817
rect 13191 15807 13296 15812
rect 13106 15667 13542 15668
rect 12312 15639 12414 15655
rect 12312 15571 12326 15639
rect 12400 15571 12414 15639
rect 12610 15582 13542 15667
rect 12312 15557 12414 15571
rect 13481 15476 13542 15582
rect 13760 15639 13862 15655
rect 13760 15571 13774 15639
rect 13848 15571 13862 15639
rect 14737 15618 14747 15729
rect 14857 15618 14867 15729
rect 15905 15618 15915 15729
rect 16025 15618 16035 15729
rect 13760 15557 13862 15571
rect 13040 15460 13106 15462
rect 10979 15451 11053 15452
rect 9058 15376 11053 15451
rect 9058 15375 9124 15376
rect 10470 15130 10590 15135
rect 10470 15036 10480 15130
rect 10580 15036 10590 15130
rect 10470 15033 10590 15036
rect 10460 12886 10626 12894
rect 10460 12818 10494 12886
rect 10578 12818 10626 12886
rect 10460 12814 10626 12818
rect 10470 12396 10590 12401
rect 10470 12302 10480 12396
rect 10580 12302 10590 12396
rect 10470 12299 10590 12302
rect 10460 10152 10626 10160
rect 10460 10084 10494 10152
rect 10578 10084 10626 10152
rect 10460 10080 10626 10084
rect 10460 9664 10580 9669
rect 10460 9570 10470 9664
rect 10570 9570 10580 9664
rect 10460 9567 10580 9570
rect 10450 7420 10616 7428
rect 10450 7352 10484 7420
rect 10568 7352 10616 7420
rect 10450 7348 10616 7352
rect 9645 6706 9859 6710
rect 9645 6634 9715 6706
rect 9791 6704 9859 6706
rect 9793 6634 9859 6704
rect 9645 6632 9859 6634
rect 9705 6629 9803 6632
rect 10979 5901 11053 15376
rect 11271 15371 13110 15460
rect 13481 15416 14792 15476
rect 11271 15369 11353 15371
rect 11714 6706 11928 6710
rect 11714 6634 11784 6706
rect 11860 6704 11928 6706
rect 11862 6634 11928 6704
rect 11714 6632 11928 6634
rect 11774 6629 11872 6632
rect 13040 5901 13106 15371
rect 13614 15130 13734 15135
rect 13614 15036 13624 15130
rect 13724 15036 13734 15130
rect 13614 15033 13734 15036
rect 13604 12886 13770 12894
rect 13604 12818 13638 12886
rect 13722 12818 13770 12886
rect 13604 12814 13770 12818
rect 13614 12396 13734 12401
rect 13614 12302 13624 12396
rect 13724 12302 13734 12396
rect 13614 12299 13734 12302
rect 13604 10152 13770 10160
rect 13604 10084 13638 10152
rect 13722 10084 13770 10152
rect 13604 10080 13770 10084
rect 13604 9664 13724 9669
rect 13604 9570 13614 9664
rect 13714 9570 13724 9664
rect 13604 9567 13724 9570
rect 13594 7420 13760 7428
rect 13594 7352 13628 7420
rect 13712 7352 13760 7420
rect 13594 7348 13760 7352
rect 13782 6708 13996 6712
rect 13782 6636 13852 6708
rect 13928 6706 13996 6708
rect 13930 6636 13996 6706
rect 13782 6634 13996 6636
rect 13842 6631 13940 6634
rect 6838 5892 6927 5897
rect 6838 5826 6848 5892
rect 6917 5826 6927 5892
rect 6838 5821 6927 5826
rect 8909 5893 8994 5898
rect 8909 5828 8920 5893
rect 8984 5828 8994 5893
rect 8909 5823 8994 5828
rect 10978 5896 11065 5901
rect 10978 5827 10988 5896
rect 11055 5827 11065 5896
rect 4759 5805 4824 5819
rect 6838 5814 6902 5821
rect 8909 5815 8976 5823
rect 10978 5822 11065 5827
rect 13040 5896 13126 5901
rect 13040 5828 13051 5896
rect 13116 5828 13126 5896
rect 13040 5823 13126 5828
rect 14727 5899 14792 15416
rect 16559 15385 16644 15817
rect 17073 15618 17083 15729
rect 17193 15618 17203 15729
rect 18241 15618 18251 15729
rect 18361 15618 18371 15729
rect 19415 15620 19425 15731
rect 19535 15620 19545 15731
rect 20583 15620 20593 15731
rect 20703 15620 20713 15731
rect 21751 15620 21761 15731
rect 21871 15620 21881 15731
rect 22919 15620 22929 15731
rect 23039 15620 23049 15731
rect 16559 15380 17148 15385
rect 16560 15315 17148 15380
rect 16816 15126 16936 15131
rect 16816 15032 16826 15126
rect 16926 15032 16936 15126
rect 16816 15029 16936 15032
rect 16806 12882 16972 12890
rect 16806 12814 16840 12882
rect 16924 12814 16972 12882
rect 16806 12810 16972 12814
rect 16816 12392 16936 12397
rect 16816 12298 16826 12392
rect 16926 12298 16936 12392
rect 16816 12295 16936 12298
rect 16806 10148 16972 10156
rect 16806 10080 16840 10148
rect 16924 10080 16972 10148
rect 16806 10076 16972 10080
rect 16806 9660 16926 9665
rect 16806 9566 16816 9660
rect 16916 9566 16926 9660
rect 16806 9563 16926 9566
rect 16796 7416 16962 7424
rect 16796 7348 16830 7416
rect 16914 7348 16962 7416
rect 16796 7344 16962 7348
rect 15851 6706 16065 6710
rect 15851 6634 15921 6706
rect 15997 6704 16065 6706
rect 15999 6634 16065 6704
rect 15851 6632 16065 6634
rect 15911 6629 16009 6632
rect 17075 5910 17146 15315
rect 19960 15126 20080 15131
rect 19960 15032 19970 15126
rect 20070 15032 20080 15126
rect 23092 15130 23212 15135
rect 23092 15036 23102 15130
rect 23202 15036 23212 15130
rect 23092 15033 23212 15036
rect 26236 15130 26356 15135
rect 26236 15036 26246 15130
rect 26346 15036 26356 15130
rect 26236 15033 26356 15036
rect 19960 15029 20080 15032
rect 19950 12882 20116 12890
rect 19950 12814 19984 12882
rect 20068 12814 20116 12882
rect 23082 12886 23248 12894
rect 23082 12818 23116 12886
rect 23200 12818 23248 12886
rect 23082 12814 23248 12818
rect 26226 12886 26392 12894
rect 26226 12818 26260 12886
rect 26344 12818 26392 12886
rect 26226 12814 26392 12818
rect 19950 12810 20116 12814
rect 19960 12392 20080 12397
rect 19960 12298 19970 12392
rect 20070 12298 20080 12392
rect 23092 12396 23212 12401
rect 23092 12302 23102 12396
rect 23202 12302 23212 12396
rect 23092 12299 23212 12302
rect 26236 12396 26356 12401
rect 26236 12302 26246 12396
rect 26346 12302 26356 12396
rect 26236 12299 26356 12302
rect 19960 12295 20080 12298
rect 19950 10148 20116 10156
rect 19950 10080 19984 10148
rect 20068 10080 20116 10148
rect 23082 10152 23248 10160
rect 23082 10084 23116 10152
rect 23200 10084 23248 10152
rect 23082 10080 23248 10084
rect 26226 10152 26392 10160
rect 26226 10084 26260 10152
rect 26344 10084 26392 10152
rect 26226 10080 26392 10084
rect 19950 10076 20116 10080
rect 19950 9660 20070 9665
rect 19950 9566 19960 9660
rect 20060 9566 20070 9660
rect 23082 9664 23202 9669
rect 23082 9570 23092 9664
rect 23192 9570 23202 9664
rect 23082 9567 23202 9570
rect 26226 9664 26346 9669
rect 26226 9570 26236 9664
rect 26336 9570 26346 9664
rect 26226 9567 26346 9570
rect 19950 9563 20070 9566
rect 19940 7416 20106 7424
rect 19940 7348 19974 7416
rect 20058 7348 20106 7416
rect 23072 7420 23238 7428
rect 23072 7352 23106 7420
rect 23190 7352 23238 7420
rect 23072 7348 23238 7352
rect 26216 7420 26382 7428
rect 26216 7352 26250 7420
rect 26334 7352 26382 7420
rect 26216 7348 26382 7352
rect 19940 7344 20106 7348
rect 19421 6777 19815 6783
rect 17919 6708 18133 6712
rect 17919 6636 17989 6708
rect 18065 6706 18133 6708
rect 18067 6636 18133 6706
rect 17919 6634 18133 6636
rect 19421 6669 19569 6777
rect 19679 6669 19815 6777
rect 17979 6631 18077 6634
rect 19421 6633 19815 6669
rect 20159 6775 20553 6781
rect 20159 6667 20307 6775
rect 20417 6667 20553 6775
rect 20159 6631 20553 6667
rect 20897 6775 21291 6781
rect 20897 6667 21045 6775
rect 21155 6667 21291 6775
rect 20897 6631 21291 6667
rect 21639 6775 22033 6781
rect 21639 6667 21787 6775
rect 21897 6667 22033 6775
rect 21639 6631 22033 6667
rect 22379 6775 22773 6781
rect 22379 6667 22527 6775
rect 22637 6667 22773 6775
rect 22379 6631 22773 6667
rect 23117 6775 23511 6781
rect 23117 6667 23265 6775
rect 23375 6667 23511 6775
rect 23117 6631 23511 6667
rect 23855 6775 24249 6781
rect 23855 6667 24003 6775
rect 24113 6667 24249 6775
rect 23855 6631 24249 6667
rect 24593 6775 24987 6781
rect 24593 6667 24741 6775
rect 24851 6667 24987 6775
rect 24593 6631 24987 6667
rect 17075 5905 17279 5910
rect 14727 5898 15147 5899
rect 14727 5893 15199 5898
rect 14727 5829 15122 5893
rect 15189 5829 15199 5893
rect 14727 5825 15199 5829
rect 14727 5824 14792 5825
rect 15012 5824 15199 5825
rect 17075 5825 17186 5905
rect 17269 5825 17279 5905
rect 19479 5885 19639 5887
rect 19479 5875 19509 5885
rect 10979 5810 11053 5822
rect 13040 5814 13106 5823
rect 17075 5812 17279 5825
rect 19477 5793 19509 5875
rect 19479 5785 19509 5793
rect 19611 5785 19639 5885
rect 20217 5883 20377 5885
rect 20217 5873 20247 5883
rect 20215 5791 20247 5873
rect 19479 5779 19639 5785
rect 20217 5783 20247 5791
rect 20349 5783 20377 5883
rect 20955 5883 21115 5885
rect 20955 5873 20985 5883
rect 20953 5791 20985 5873
rect 20217 5777 20377 5783
rect 20955 5783 20985 5791
rect 21087 5783 21115 5883
rect 21697 5883 21857 5885
rect 21697 5873 21727 5883
rect 21695 5791 21727 5873
rect 20955 5777 21115 5783
rect 21697 5783 21727 5791
rect 21829 5783 21857 5883
rect 22437 5883 22597 5885
rect 22437 5873 22467 5883
rect 22435 5791 22467 5873
rect 21697 5777 21857 5783
rect 22437 5783 22467 5791
rect 22569 5783 22597 5883
rect 23175 5883 23335 5885
rect 23175 5873 23205 5883
rect 23173 5791 23205 5873
rect 22437 5777 22597 5783
rect 23175 5783 23205 5791
rect 23307 5783 23335 5883
rect 23913 5883 24073 5885
rect 23913 5873 23943 5883
rect 23911 5791 23943 5873
rect 23175 5777 23335 5783
rect 23913 5783 23943 5791
rect 24045 5783 24073 5883
rect 24651 5883 24811 5885
rect 24651 5873 24681 5883
rect 24649 5791 24681 5873
rect 23913 5777 24073 5783
rect 24651 5783 24681 5791
rect 24783 5783 24811 5883
rect 24651 5777 24811 5783
rect 2679 5704 2789 5749
rect 2679 5627 2699 5704
rect 2770 5627 2789 5704
rect 2679 5607 2789 5627
rect 13762 4490 13914 4492
rect 17899 4490 18051 4492
rect 5488 4488 5640 4490
rect 9625 4488 9777 4490
rect 11694 4488 11846 4490
rect 3420 4486 3572 4488
rect 3418 4482 3572 4486
rect 3418 4394 3448 4482
rect 3542 4394 3572 4482
rect 3418 4388 3572 4394
rect 5486 4484 5640 4488
rect 7557 4486 7709 4488
rect 5486 4396 5516 4484
rect 5610 4396 5640 4484
rect 5486 4390 5640 4396
rect 3420 4378 3572 4388
rect 5488 4380 5640 4390
rect 7555 4482 7709 4486
rect 7555 4394 7585 4482
rect 7679 4394 7709 4482
rect 7555 4388 7709 4394
rect 9623 4484 9777 4488
rect 9623 4396 9653 4484
rect 9747 4396 9777 4484
rect 9623 4390 9777 4396
rect 11692 4484 11846 4488
rect 11692 4396 11722 4484
rect 11816 4396 11846 4484
rect 11692 4390 11846 4396
rect 13760 4486 13914 4490
rect 15831 4488 15983 4490
rect 13760 4398 13790 4486
rect 13884 4398 13914 4486
rect 13760 4392 13914 4398
rect 7557 4378 7709 4388
rect 9625 4380 9777 4390
rect 11694 4380 11846 4390
rect 13762 4382 13914 4392
rect 15829 4484 15983 4488
rect 15829 4396 15859 4484
rect 15953 4396 15983 4484
rect 15829 4390 15983 4396
rect 17897 4486 18051 4490
rect 17897 4398 17927 4486
rect 18021 4398 18051 4486
rect 17897 4392 18051 4398
rect 15831 4380 15983 4390
rect 17899 4382 18051 4392
rect 1486 2412 1606 2417
rect 1486 2318 1496 2412
rect 1596 2318 1606 2412
rect 1486 2315 1606 2318
rect 4630 2412 4750 2417
rect 4630 2318 4640 2412
rect 4740 2318 4750 2412
rect 7762 2416 7882 2421
rect 7762 2322 7772 2416
rect 7872 2322 7882 2416
rect 7762 2319 7882 2322
rect 10906 2416 11026 2421
rect 10906 2322 10916 2416
rect 11016 2322 11026 2416
rect 10906 2319 11026 2322
rect 14108 2412 14228 2417
rect 4630 2315 4750 2318
rect 14108 2318 14118 2412
rect 14218 2318 14228 2412
rect 14108 2315 14228 2318
rect 17252 2412 17372 2417
rect 17252 2318 17262 2412
rect 17362 2318 17372 2412
rect 20384 2416 20504 2421
rect 20384 2322 20394 2416
rect 20494 2322 20504 2416
rect 20384 2319 20504 2322
rect 23528 2416 23648 2421
rect 23528 2322 23538 2416
rect 23638 2322 23648 2416
rect 23528 2319 23648 2322
rect 17252 2315 17372 2318
rect 1476 168 1642 176
rect 1476 100 1510 168
rect 1594 100 1642 168
rect 1476 96 1642 100
rect 4620 168 4786 176
rect 4620 100 4654 168
rect 4738 100 4786 168
rect 7752 172 7918 180
rect 7752 104 7786 172
rect 7870 104 7918 172
rect 7752 100 7918 104
rect 10896 172 11062 180
rect 10896 104 10930 172
rect 11014 104 11062 172
rect 10896 100 11062 104
rect 14098 168 14264 176
rect 14098 100 14132 168
rect 14216 100 14264 168
rect 4620 96 4786 100
rect 14098 96 14264 100
rect 17242 168 17408 176
rect 17242 100 17276 168
rect 17360 100 17408 168
rect 20374 172 20540 180
rect 20374 104 20408 172
rect 20492 104 20540 172
rect 20374 100 20540 104
rect 23518 172 23684 180
rect 23518 104 23552 172
rect 23636 104 23684 172
rect 23518 100 23684 104
rect 17242 96 17408 100
rect 1518 -1480 1638 -1475
rect 1518 -1574 1528 -1480
rect 1628 -1574 1638 -1480
rect 1518 -1577 1638 -1574
rect 4662 -1480 4782 -1475
rect 4662 -1574 4672 -1480
rect 4772 -1574 4782 -1480
rect 7794 -1476 7914 -1471
rect 7794 -1570 7804 -1476
rect 7904 -1570 7914 -1476
rect 7794 -1573 7914 -1570
rect 10938 -1476 11058 -1471
rect 10938 -1570 10948 -1476
rect 11048 -1570 11058 -1476
rect 10938 -1573 11058 -1570
rect 14140 -1480 14260 -1475
rect 4662 -1577 4782 -1574
rect 14140 -1574 14150 -1480
rect 14250 -1574 14260 -1480
rect 14140 -1577 14260 -1574
rect 17284 -1480 17404 -1475
rect 17284 -1574 17294 -1480
rect 17394 -1574 17404 -1480
rect 20416 -1476 20536 -1471
rect 20416 -1570 20426 -1476
rect 20526 -1570 20536 -1476
rect 20416 -1573 20536 -1570
rect 23560 -1476 23680 -1471
rect 23560 -1570 23570 -1476
rect 23670 -1570 23680 -1476
rect 23560 -1573 23680 -1570
rect 17284 -1577 17404 -1574
rect 1508 -3724 1674 -3716
rect 1508 -3792 1542 -3724
rect 1626 -3792 1674 -3724
rect 1508 -3796 1674 -3792
rect 4652 -3724 4818 -3716
rect 4652 -3792 4686 -3724
rect 4770 -3792 4818 -3724
rect 7784 -3720 7950 -3712
rect 7784 -3788 7818 -3720
rect 7902 -3788 7950 -3720
rect 7784 -3792 7950 -3788
rect 10928 -3720 11094 -3712
rect 10928 -3788 10962 -3720
rect 11046 -3788 11094 -3720
rect 10928 -3792 11094 -3788
rect 14130 -3724 14296 -3716
rect 14130 -3792 14164 -3724
rect 14248 -3792 14296 -3724
rect 4652 -3796 4818 -3792
rect 14130 -3796 14296 -3792
rect 17274 -3724 17440 -3716
rect 17274 -3792 17308 -3724
rect 17392 -3792 17440 -3724
rect 20406 -3720 20572 -3712
rect 20406 -3788 20440 -3720
rect 20524 -3788 20572 -3720
rect 20406 -3792 20572 -3788
rect 23550 -3720 23716 -3712
rect 23550 -3788 23584 -3720
rect 23668 -3788 23716 -3720
rect 23550 -3792 23716 -3788
rect 17274 -3796 17440 -3792
<< via3 >>
rect 1702 22172 1802 22262
rect 1702 22170 1802 22172
rect 4846 22172 4946 22262
rect 4846 22170 4946 22172
rect 7978 22176 8078 22266
rect 7978 22174 8078 22176
rect 11122 22176 11222 22266
rect 11122 22174 11222 22176
rect 14324 22172 14424 22262
rect 14324 22170 14424 22172
rect 17468 22172 17568 22262
rect 17468 22170 17568 22172
rect 20600 22176 20700 22266
rect 20600 22174 20700 22176
rect 23744 22176 23844 22266
rect 23744 22174 23844 22176
rect 312 21169 389 21183
rect 312 21113 322 21169
rect 322 21113 378 21169
rect 378 21113 389 21169
rect 312 21100 389 21113
rect 22343 21024 22443 21034
rect 22343 20935 22354 21024
rect 22354 20935 22433 21024
rect 22433 20935 22443 21024
rect 22343 20925 22443 20935
rect 1716 19962 1722 20020
rect 1722 19962 1798 20020
rect 1798 19962 1800 20020
rect 1716 19952 1800 19962
rect 4860 19962 4866 20020
rect 4866 19962 4942 20020
rect 4942 19962 4944 20020
rect 4860 19952 4944 19962
rect 7992 19966 7998 20024
rect 7998 19966 8074 20024
rect 8074 19966 8076 20024
rect 7992 19956 8076 19966
rect 11136 19966 11142 20024
rect 11142 19966 11218 20024
rect 11218 19966 11220 20024
rect 11136 19956 11220 19966
rect 14338 19962 14344 20020
rect 14344 19962 14420 20020
rect 14420 19962 14422 20020
rect 14338 19952 14422 19962
rect 17482 19962 17488 20020
rect 17488 19962 17564 20020
rect 17564 19962 17566 20020
rect 17482 19952 17566 19962
rect 20614 19966 20620 20024
rect 20620 19966 20696 20024
rect 20696 19966 20698 20024
rect 20614 19956 20698 19966
rect 23758 19966 23764 20024
rect 23764 19966 23840 20024
rect 23840 19966 23842 20024
rect 23758 19956 23842 19966
rect 15204 17046 15326 17060
rect 15204 16955 15222 17046
rect 15222 16955 15312 17046
rect 15312 16955 15326 17046
rect 15204 16940 15326 16955
rect 16406 16968 16470 17032
rect 17574 16968 17638 17032
rect 18744 16970 18808 17034
rect 19916 16970 19980 17034
rect 21084 16968 21148 17032
rect 22252 16970 22316 17034
rect 23420 16970 23484 17034
rect 3244 16837 3314 16841
rect 3244 16775 3250 16837
rect 3250 16775 3310 16837
rect 3310 16775 3314 16837
rect 3244 16769 3314 16775
rect 4692 16837 4762 16841
rect 4692 16775 4698 16837
rect 4698 16775 4758 16837
rect 4758 16775 4762 16837
rect 4692 16769 4762 16775
rect 6190 16839 6260 16843
rect 6190 16777 6196 16839
rect 6196 16777 6256 16839
rect 6256 16777 6260 16839
rect 6190 16771 6260 16777
rect 7638 16839 7708 16843
rect 7638 16777 7644 16839
rect 7644 16777 7704 16839
rect 7704 16777 7708 16839
rect 7638 16771 7708 16777
rect 9158 16837 9228 16841
rect 9158 16775 9164 16837
rect 9164 16775 9224 16837
rect 9224 16775 9228 16837
rect 9158 16769 9228 16775
rect 10606 16837 10676 16841
rect 10606 16775 10612 16837
rect 10612 16775 10672 16837
rect 10672 16775 10676 16837
rect 10606 16769 10676 16775
rect 12104 16839 12174 16843
rect 12104 16777 12110 16839
rect 12110 16777 12170 16839
rect 12170 16777 12174 16839
rect 12104 16771 12174 16777
rect 13552 16839 13622 16843
rect 13552 16777 13558 16839
rect 13558 16777 13618 16839
rect 13618 16777 13622 16839
rect 13552 16771 13622 16777
rect 3466 15631 3540 15637
rect 3466 15569 3472 15631
rect 3472 15569 3536 15631
rect 3536 15569 3540 15631
rect 4204 15034 4304 15124
rect 4204 15032 4304 15034
rect 4218 12824 4224 12882
rect 4224 12824 4300 12882
rect 4300 12824 4302 12882
rect 4218 12814 4302 12824
rect 4204 12300 4304 12390
rect 4204 12298 4304 12300
rect 4218 10090 4224 10148
rect 4224 10090 4300 10148
rect 4300 10090 4302 10148
rect 4218 10080 4302 10090
rect 4194 9568 4294 9658
rect 4194 9566 4294 9568
rect 4208 7358 4214 7416
rect 4214 7358 4290 7416
rect 4290 7358 4292 7416
rect 4208 7348 4292 7358
rect 3510 6702 3586 6704
rect 3510 6638 3586 6702
rect 4914 15631 4988 15637
rect 4914 15569 4920 15631
rect 4920 15569 4984 15631
rect 4984 15569 4988 15631
rect 6412 15633 6486 15639
rect 6412 15571 6418 15633
rect 6418 15571 6482 15633
rect 6482 15571 6486 15633
rect 5578 6704 5654 6706
rect 5578 6640 5654 6704
rect 7860 15633 7934 15639
rect 7860 15571 7866 15633
rect 7866 15571 7930 15633
rect 7930 15571 7934 15633
rect 7348 15034 7448 15124
rect 7348 15032 7448 15034
rect 7362 12824 7368 12882
rect 7368 12824 7444 12882
rect 7444 12824 7446 12882
rect 7362 12814 7446 12824
rect 7348 12300 7448 12390
rect 7348 12298 7448 12300
rect 7362 10090 7368 10148
rect 7368 10090 7444 10148
rect 7444 10090 7446 10148
rect 7362 10080 7446 10090
rect 7338 9568 7438 9658
rect 7338 9566 7438 9568
rect 7352 7358 7358 7416
rect 7358 7358 7434 7416
rect 7434 7358 7436 7416
rect 7352 7348 7436 7358
rect 7647 6702 7723 6704
rect 7647 6638 7723 6702
rect 9380 15631 9454 15637
rect 9380 15569 9386 15631
rect 9386 15569 9450 15631
rect 9450 15569 9454 15631
rect 10828 15631 10902 15637
rect 10828 15569 10834 15631
rect 10834 15569 10898 15631
rect 10898 15569 10902 15631
rect 12326 15633 12400 15639
rect 12326 15571 12332 15633
rect 12332 15571 12396 15633
rect 12396 15571 12400 15633
rect 13774 15633 13848 15639
rect 13774 15571 13780 15633
rect 13780 15571 13844 15633
rect 13844 15571 13848 15633
rect 14747 15719 14857 15729
rect 14747 15628 14757 15719
rect 14757 15628 14847 15719
rect 14847 15628 14857 15719
rect 14747 15618 14857 15628
rect 15915 15719 16025 15729
rect 15915 15628 15925 15719
rect 15925 15628 16015 15719
rect 16015 15628 16025 15719
rect 15915 15618 16025 15628
rect 10480 15038 10580 15128
rect 10480 15036 10580 15038
rect 10494 12828 10500 12886
rect 10500 12828 10576 12886
rect 10576 12828 10578 12886
rect 10494 12818 10578 12828
rect 10480 12304 10580 12394
rect 10480 12302 10580 12304
rect 10494 10094 10500 10152
rect 10500 10094 10576 10152
rect 10576 10094 10578 10152
rect 10494 10084 10578 10094
rect 10470 9572 10570 9662
rect 10470 9570 10570 9572
rect 10484 7362 10490 7420
rect 10490 7362 10566 7420
rect 10566 7362 10568 7420
rect 10484 7352 10568 7362
rect 9715 6704 9791 6706
rect 9715 6640 9791 6704
rect 11784 6704 11860 6706
rect 11784 6640 11860 6704
rect 13624 15038 13724 15128
rect 13624 15036 13724 15038
rect 13638 12828 13644 12886
rect 13644 12828 13720 12886
rect 13720 12828 13722 12886
rect 13638 12818 13722 12828
rect 13624 12304 13724 12394
rect 13624 12302 13724 12304
rect 13638 10094 13644 10152
rect 13644 10094 13720 10152
rect 13720 10094 13722 10152
rect 13638 10084 13722 10094
rect 13614 9572 13714 9662
rect 13614 9570 13714 9572
rect 13628 7362 13634 7420
rect 13634 7362 13710 7420
rect 13710 7362 13712 7420
rect 13628 7352 13712 7362
rect 13852 6706 13928 6708
rect 13852 6642 13928 6706
rect 17083 15719 17193 15729
rect 17083 15628 17093 15719
rect 17093 15628 17183 15719
rect 17183 15628 17193 15719
rect 17083 15618 17193 15628
rect 18251 15719 18361 15729
rect 18251 15628 18261 15719
rect 18261 15628 18351 15719
rect 18351 15628 18361 15719
rect 18251 15618 18361 15628
rect 19425 15721 19535 15731
rect 19425 15630 19435 15721
rect 19435 15630 19525 15721
rect 19525 15630 19535 15721
rect 19425 15620 19535 15630
rect 20593 15721 20703 15731
rect 20593 15630 20603 15721
rect 20603 15630 20693 15721
rect 20693 15630 20703 15721
rect 20593 15620 20703 15630
rect 21761 15721 21871 15731
rect 21761 15630 21771 15721
rect 21771 15630 21861 15721
rect 21861 15630 21871 15721
rect 21761 15620 21871 15630
rect 22929 15721 23039 15731
rect 22929 15630 22939 15721
rect 22939 15630 23029 15721
rect 23029 15630 23039 15721
rect 22929 15620 23039 15630
rect 16826 15034 16926 15124
rect 16826 15032 16926 15034
rect 16840 12824 16846 12882
rect 16846 12824 16922 12882
rect 16922 12824 16924 12882
rect 16840 12814 16924 12824
rect 16826 12300 16926 12390
rect 16826 12298 16926 12300
rect 16840 10090 16846 10148
rect 16846 10090 16922 10148
rect 16922 10090 16924 10148
rect 16840 10080 16924 10090
rect 16816 9568 16916 9658
rect 16816 9566 16916 9568
rect 16830 7358 16836 7416
rect 16836 7358 16912 7416
rect 16912 7358 16914 7416
rect 16830 7348 16914 7358
rect 15921 6704 15997 6706
rect 15921 6640 15997 6704
rect 19970 15034 20070 15124
rect 19970 15032 20070 15034
rect 23102 15038 23202 15128
rect 23102 15036 23202 15038
rect 26246 15038 26346 15128
rect 26246 15036 26346 15038
rect 19984 12824 19990 12882
rect 19990 12824 20066 12882
rect 20066 12824 20068 12882
rect 19984 12814 20068 12824
rect 23116 12828 23122 12886
rect 23122 12828 23198 12886
rect 23198 12828 23200 12886
rect 23116 12818 23200 12828
rect 26260 12828 26266 12886
rect 26266 12828 26342 12886
rect 26342 12828 26344 12886
rect 26260 12818 26344 12828
rect 19970 12300 20070 12390
rect 19970 12298 20070 12300
rect 23102 12304 23202 12394
rect 23102 12302 23202 12304
rect 26246 12304 26346 12394
rect 26246 12302 26346 12304
rect 19984 10090 19990 10148
rect 19990 10090 20066 10148
rect 20066 10090 20068 10148
rect 19984 10080 20068 10090
rect 23116 10094 23122 10152
rect 23122 10094 23198 10152
rect 23198 10094 23200 10152
rect 23116 10084 23200 10094
rect 26260 10094 26266 10152
rect 26266 10094 26342 10152
rect 26342 10094 26344 10152
rect 26260 10084 26344 10094
rect 19960 9568 20060 9658
rect 19960 9566 20060 9568
rect 23092 9572 23192 9662
rect 23092 9570 23192 9572
rect 26236 9572 26336 9662
rect 26236 9570 26336 9572
rect 19974 7358 19980 7416
rect 19980 7358 20056 7416
rect 20056 7358 20058 7416
rect 19974 7348 20058 7358
rect 23106 7362 23112 7420
rect 23112 7362 23188 7420
rect 23188 7362 23190 7420
rect 23106 7352 23190 7362
rect 26250 7362 26256 7420
rect 26256 7362 26332 7420
rect 26332 7362 26334 7420
rect 26250 7352 26334 7362
rect 17989 6706 18065 6708
rect 17989 6642 18065 6706
rect 19569 6763 19679 6777
rect 19569 6679 19577 6763
rect 19577 6679 19671 6763
rect 19671 6679 19679 6763
rect 19569 6669 19679 6679
rect 20307 6761 20417 6775
rect 20307 6677 20315 6761
rect 20315 6677 20409 6761
rect 20409 6677 20417 6761
rect 20307 6667 20417 6677
rect 21045 6761 21155 6775
rect 21045 6677 21053 6761
rect 21053 6677 21147 6761
rect 21147 6677 21155 6761
rect 21045 6667 21155 6677
rect 21787 6761 21897 6775
rect 21787 6677 21795 6761
rect 21795 6677 21889 6761
rect 21889 6677 21897 6761
rect 21787 6667 21897 6677
rect 22527 6761 22637 6775
rect 22527 6677 22535 6761
rect 22535 6677 22629 6761
rect 22629 6677 22637 6761
rect 22527 6667 22637 6677
rect 23265 6761 23375 6775
rect 23265 6677 23273 6761
rect 23273 6677 23367 6761
rect 23367 6677 23375 6761
rect 23265 6667 23375 6677
rect 24003 6761 24113 6775
rect 24003 6677 24011 6761
rect 24011 6677 24105 6761
rect 24105 6677 24113 6761
rect 24003 6667 24113 6677
rect 24741 6761 24851 6775
rect 24741 6677 24749 6761
rect 24749 6677 24843 6761
rect 24843 6677 24851 6761
rect 24741 6667 24851 6677
rect 19509 5865 19611 5885
rect 19509 5807 19525 5865
rect 19525 5807 19591 5865
rect 19591 5807 19611 5865
rect 19509 5785 19611 5807
rect 20247 5863 20349 5883
rect 20247 5805 20263 5863
rect 20263 5805 20329 5863
rect 20329 5805 20349 5863
rect 20247 5783 20349 5805
rect 20985 5863 21087 5883
rect 20985 5805 21001 5863
rect 21001 5805 21067 5863
rect 21067 5805 21087 5863
rect 20985 5783 21087 5805
rect 21727 5863 21829 5883
rect 21727 5805 21743 5863
rect 21743 5805 21809 5863
rect 21809 5805 21829 5863
rect 21727 5783 21829 5805
rect 22467 5863 22569 5883
rect 22467 5805 22483 5863
rect 22483 5805 22549 5863
rect 22549 5805 22569 5863
rect 22467 5783 22569 5805
rect 23205 5863 23307 5883
rect 23205 5805 23221 5863
rect 23221 5805 23287 5863
rect 23287 5805 23307 5863
rect 23205 5783 23307 5805
rect 23943 5863 24045 5883
rect 23943 5805 23959 5863
rect 23959 5805 24025 5863
rect 24025 5805 24045 5863
rect 23943 5783 24045 5805
rect 24681 5863 24783 5883
rect 24681 5805 24697 5863
rect 24697 5805 24763 5863
rect 24763 5805 24783 5863
rect 24681 5783 24783 5805
rect 3448 4472 3542 4482
rect 3448 4402 3458 4472
rect 3458 4402 3530 4472
rect 3530 4402 3542 4472
rect 3448 4394 3542 4402
rect 5516 4474 5610 4484
rect 5516 4404 5526 4474
rect 5526 4404 5598 4474
rect 5598 4404 5610 4474
rect 5516 4396 5610 4404
rect 7585 4472 7679 4482
rect 7585 4402 7595 4472
rect 7595 4402 7667 4472
rect 7667 4402 7679 4472
rect 7585 4394 7679 4402
rect 9653 4474 9747 4484
rect 9653 4404 9663 4474
rect 9663 4404 9735 4474
rect 9735 4404 9747 4474
rect 9653 4396 9747 4404
rect 11722 4474 11816 4484
rect 11722 4404 11732 4474
rect 11732 4404 11804 4474
rect 11804 4404 11816 4474
rect 11722 4396 11816 4404
rect 13790 4476 13884 4486
rect 13790 4406 13800 4476
rect 13800 4406 13872 4476
rect 13872 4406 13884 4476
rect 13790 4398 13884 4406
rect 15859 4474 15953 4484
rect 15859 4404 15869 4474
rect 15869 4404 15941 4474
rect 15941 4404 15953 4474
rect 15859 4396 15953 4404
rect 17927 4476 18021 4486
rect 17927 4406 17937 4476
rect 17937 4406 18009 4476
rect 18009 4406 18021 4476
rect 17927 4398 18021 4406
rect 1496 2320 1596 2410
rect 1496 2318 1596 2320
rect 4640 2320 4740 2410
rect 4640 2318 4740 2320
rect 7772 2324 7872 2414
rect 7772 2322 7872 2324
rect 10916 2324 11016 2414
rect 10916 2322 11016 2324
rect 14118 2320 14218 2410
rect 14118 2318 14218 2320
rect 17262 2320 17362 2410
rect 17262 2318 17362 2320
rect 20394 2324 20494 2414
rect 20394 2322 20494 2324
rect 23538 2324 23638 2414
rect 23538 2322 23638 2324
rect 1510 110 1516 168
rect 1516 110 1592 168
rect 1592 110 1594 168
rect 1510 100 1594 110
rect 4654 110 4660 168
rect 4660 110 4736 168
rect 4736 110 4738 168
rect 4654 100 4738 110
rect 7786 114 7792 172
rect 7792 114 7868 172
rect 7868 114 7870 172
rect 7786 104 7870 114
rect 10930 114 10936 172
rect 10936 114 11012 172
rect 11012 114 11014 172
rect 10930 104 11014 114
rect 14132 110 14138 168
rect 14138 110 14214 168
rect 14214 110 14216 168
rect 14132 100 14216 110
rect 17276 110 17282 168
rect 17282 110 17358 168
rect 17358 110 17360 168
rect 17276 100 17360 110
rect 20408 114 20414 172
rect 20414 114 20490 172
rect 20490 114 20492 172
rect 20408 104 20492 114
rect 23552 114 23558 172
rect 23558 114 23634 172
rect 23634 114 23636 172
rect 23552 104 23636 114
rect 1528 -1572 1628 -1482
rect 1528 -1574 1628 -1572
rect 4672 -1572 4772 -1482
rect 4672 -1574 4772 -1572
rect 7804 -1568 7904 -1478
rect 7804 -1570 7904 -1568
rect 10948 -1568 11048 -1478
rect 10948 -1570 11048 -1568
rect 14150 -1572 14250 -1482
rect 14150 -1574 14250 -1572
rect 17294 -1572 17394 -1482
rect 17294 -1574 17394 -1572
rect 20426 -1568 20526 -1478
rect 20426 -1570 20526 -1568
rect 23570 -1568 23670 -1478
rect 23570 -1570 23670 -1568
rect 1542 -3782 1548 -3724
rect 1548 -3782 1624 -3724
rect 1624 -3782 1626 -3724
rect 1542 -3792 1626 -3782
rect 4686 -3782 4692 -3724
rect 4692 -3782 4768 -3724
rect 4768 -3782 4770 -3724
rect 4686 -3792 4770 -3782
rect 7818 -3778 7824 -3720
rect 7824 -3778 7900 -3720
rect 7900 -3778 7902 -3720
rect 7818 -3788 7902 -3778
rect 10962 -3778 10968 -3720
rect 10968 -3778 11044 -3720
rect 11044 -3778 11046 -3720
rect 10962 -3788 11046 -3778
rect 14164 -3782 14170 -3724
rect 14170 -3782 14246 -3724
rect 14246 -3782 14248 -3724
rect 14164 -3792 14248 -3782
rect 17308 -3782 17314 -3724
rect 17314 -3782 17390 -3724
rect 17390 -3782 17392 -3724
rect 17308 -3792 17392 -3782
rect 20440 -3778 20446 -3720
rect 20446 -3778 20522 -3720
rect 20522 -3778 20524 -3720
rect 20440 -3788 20524 -3778
rect 23584 -3778 23590 -3720
rect 23590 -3778 23666 -3720
rect 23666 -3778 23668 -3720
rect 23584 -3788 23668 -3778
<< metal4 >>
rect 846 22266 24776 22372
rect 846 22262 7978 22266
rect 846 22170 1702 22262
rect 1802 22170 4846 22262
rect 4946 22174 7978 22262
rect 8078 22174 11122 22266
rect 11222 22262 20600 22266
rect 11222 22174 14324 22262
rect 4946 22170 14324 22174
rect 14424 22170 17468 22262
rect 17568 22174 20600 22262
rect 20700 22174 23744 22266
rect 23844 22174 24776 22266
rect 17568 22170 24776 22174
rect 846 22138 24776 22170
rect 302 21183 390 21184
rect 302 21100 312 21183
rect 389 21100 390 21183
rect 302 20031 390 21100
rect 22333 21034 22454 21035
rect 22333 20925 22343 21034
rect 22443 20925 22454 21034
rect 22333 20032 22454 20925
rect 826 20031 24200 20032
rect 302 20024 24200 20031
rect 302 20020 7992 20024
rect 302 19952 1716 20020
rect 1800 19952 4860 20020
rect 4944 19956 7992 20020
rect 8076 19956 11136 20024
rect 11220 20020 20614 20024
rect 11220 19956 14338 20020
rect 4944 19952 14338 19956
rect 14422 19952 17482 20020
rect 17566 19956 20614 20020
rect 20698 19956 23758 20024
rect 23842 19956 24200 20024
rect 17566 19952 24200 19956
rect 302 19852 24200 19952
rect 13839 17060 23616 17126
rect 13839 16940 15204 17060
rect 15326 17034 23616 17060
rect 15326 17032 18744 17034
rect 15326 16968 16406 17032
rect 16470 16968 17574 17032
rect 17638 16970 18744 17032
rect 18808 16970 19916 17034
rect 19980 17032 22252 17034
rect 19980 16970 21084 17032
rect 17638 16968 21084 16970
rect 21148 16970 22252 17032
rect 22316 16970 23420 17034
rect 23484 16970 23616 17034
rect 21148 16968 23616 16970
rect 15326 16940 23616 16968
rect 13839 16930 23616 16940
rect 13839 16899 14695 16930
rect 2783 16843 14695 16899
rect 2783 16841 6190 16843
rect 2783 16769 3244 16841
rect 3314 16769 4692 16841
rect 4762 16771 6190 16841
rect 6260 16771 7638 16843
rect 7708 16841 12104 16843
rect 7708 16771 9158 16841
rect 4762 16769 9158 16771
rect 9228 16769 10606 16841
rect 10676 16771 12104 16841
rect 12174 16771 13552 16843
rect 13622 16771 14695 16843
rect 10676 16769 14695 16771
rect 2783 16742 14695 16769
rect 2783 16741 14022 16742
rect 2783 15231 3099 16741
rect 3348 15231 27278 15234
rect 2778 15128 27278 15231
rect 2778 15124 10480 15128
rect 2778 15088 4204 15124
rect 2770 15032 4204 15088
rect 4304 15032 7348 15124
rect 7448 15036 10480 15124
rect 10580 15036 13624 15128
rect 13724 15124 23102 15128
rect 13724 15036 16826 15124
rect 7448 15032 16826 15036
rect 16926 15032 19970 15124
rect 20070 15036 23102 15124
rect 23202 15036 26246 15128
rect 26346 15036 27278 15128
rect 20070 15032 27278 15036
rect 2770 15000 27278 15032
rect 2770 14998 3459 15000
rect 2770 12498 3058 14998
rect 3348 12498 27278 12500
rect 2770 12394 27278 12498
rect 2770 12390 10480 12394
rect 2770 12298 4204 12390
rect 4304 12298 7348 12390
rect 7448 12302 10480 12390
rect 10580 12302 13624 12394
rect 13724 12390 23102 12394
rect 13724 12302 16826 12390
rect 7448 12298 16826 12302
rect 16926 12298 19970 12390
rect 20070 12302 23102 12390
rect 23202 12302 26246 12394
rect 26346 12302 27278 12394
rect 20070 12298 27278 12302
rect 2770 12266 27278 12298
rect 2770 12263 3569 12266
rect 2770 9775 3058 12263
rect 2770 9768 3533 9775
rect 2770 9662 27268 9768
rect 2770 9658 10470 9662
rect 2770 9566 4194 9658
rect 4294 9566 7338 9658
rect 7438 9570 10470 9658
rect 10570 9570 13614 9662
rect 13714 9658 23092 9662
rect 13714 9570 16816 9658
rect 7438 9566 16816 9570
rect 16916 9566 19960 9658
rect 20060 9570 23092 9658
rect 23192 9570 26236 9662
rect 26336 9570 27268 9662
rect 20060 9566 27268 9570
rect 2770 9540 27268 9566
rect 2770 6840 3058 9540
rect 3338 9534 27268 9540
rect 18684 6851 19442 6852
rect 18684 6840 25039 6851
rect 2666 6777 25039 6840
rect 2666 6708 19569 6777
rect 2666 6706 13852 6708
rect 2666 6704 5578 6706
rect 2666 6638 3510 6704
rect 3586 6640 5578 6704
rect 5654 6704 9715 6706
rect 5654 6640 7647 6704
rect 3586 6638 7647 6640
rect 7723 6640 9715 6704
rect 9791 6640 11784 6706
rect 11860 6642 13852 6706
rect 13928 6706 17989 6708
rect 13928 6642 15921 6706
rect 11860 6640 15921 6642
rect 15997 6642 17989 6706
rect 18065 6669 19569 6708
rect 19679 6775 25039 6777
rect 19679 6669 20307 6775
rect 18065 6667 20307 6669
rect 20417 6667 21045 6775
rect 21155 6667 21787 6775
rect 21897 6667 22527 6775
rect 22637 6667 23265 6775
rect 23375 6667 24003 6775
rect 24113 6667 24741 6775
rect 24851 6667 25039 6775
rect 18065 6661 25039 6667
rect 18065 6642 19442 6661
rect 15997 6640 19442 6642
rect 7723 6638 19442 6640
rect 2666 6596 19442 6638
rect 2770 6587 3058 6596
rect 18684 6594 19442 6596
rect 19422 5751 19440 5941
rect 19676 5751 19683 5941
rect 20161 5751 20174 5941
rect 20410 5751 20423 5941
rect 20899 5751 20922 5941
rect 21158 5751 21159 5941
rect 21641 5751 21663 5941
rect 21899 5751 21902 5941
rect 22381 5751 22394 5941
rect 22630 5751 22643 5941
rect 23119 5751 23133 5941
rect 23369 5751 23380 5941
rect 23856 5751 23879 5941
rect 24115 5751 24117 5941
rect 24593 5751 24606 5941
rect 24842 5751 24855 5941
rect 3373 4298 3379 4488
rect 3615 4298 3625 4488
rect 5440 4298 5446 4490
rect 5682 4298 5692 4490
rect 7508 4298 7519 4488
rect 7755 4298 7763 4488
rect 9577 4298 9587 4490
rect 9823 4298 9831 4490
rect 11645 4298 11660 4490
rect 11896 4298 11898 4490
rect 13712 4298 13724 4492
rect 13960 4298 13968 4492
rect 15782 4298 15787 4490
rect 16023 4298 16036 4490
rect 17850 4298 17860 4492
rect 18096 4298 18105 4492
rect 640 2414 24570 2520
rect 640 2410 7772 2414
rect 640 2318 1496 2410
rect 1596 2318 4640 2410
rect 4740 2322 7772 2410
rect 7872 2322 10916 2414
rect 11016 2410 20394 2414
rect 11016 2322 14118 2410
rect 4740 2318 14118 2322
rect 14218 2318 17262 2410
rect 17362 2322 20394 2410
rect 20494 2322 23538 2414
rect 23638 2322 24570 2414
rect 17362 2318 24570 2322
rect 640 2286 24570 2318
rect 620 172 23994 180
rect 620 168 7786 172
rect 620 100 1510 168
rect 1594 100 4654 168
rect 4738 104 7786 168
rect 7870 104 10930 172
rect 11014 168 20408 172
rect 11014 104 14132 168
rect 4738 100 14132 104
rect 14216 100 17276 168
rect 17360 104 20408 168
rect 20492 104 23552 172
rect 23636 104 23994 172
rect 17360 100 23994 104
rect 620 0 23994 100
rect 672 -1478 24602 -1372
rect 672 -1482 7804 -1478
rect 672 -1574 1528 -1482
rect 1628 -1574 4672 -1482
rect 4772 -1570 7804 -1482
rect 7904 -1570 10948 -1478
rect 11048 -1482 20426 -1478
rect 11048 -1570 14150 -1482
rect 4772 -1574 14150 -1570
rect 14250 -1574 17294 -1482
rect 17394 -1570 20426 -1482
rect 20526 -1570 23570 -1478
rect 23670 -1570 24602 -1478
rect 17394 -1574 24602 -1570
rect 672 -1606 24602 -1574
rect 652 -3720 24026 -3712
rect 652 -3724 7818 -3720
rect 652 -3792 1542 -3724
rect 1626 -3792 4686 -3724
rect 4770 -3788 7818 -3724
rect 7902 -3788 10962 -3720
rect 11046 -3724 20440 -3720
rect 11046 -3788 14164 -3724
rect 4770 -3792 14164 -3788
rect 14248 -3792 17308 -3724
rect 17392 -3788 20440 -3724
rect 20524 -3788 23584 -3720
rect 23668 -3788 24026 -3720
rect 17392 -3792 24026 -3788
rect 652 -3892 24026 -3792
<< via4 >>
rect 3387 15637 3623 15730
rect 3387 15569 3466 15637
rect 3466 15569 3540 15637
rect 3540 15569 3623 15637
rect 3387 15494 3623 15569
rect 4836 15637 5072 15715
rect 4836 15569 4914 15637
rect 4914 15569 4988 15637
rect 4988 15569 5072 15637
rect 4836 15479 5072 15569
rect 6331 15639 6567 15724
rect 6331 15571 6412 15639
rect 6412 15571 6486 15639
rect 6486 15571 6567 15639
rect 6331 15488 6567 15571
rect 7780 15639 8016 15719
rect 7780 15571 7860 15639
rect 7860 15571 7934 15639
rect 7934 15571 8016 15639
rect 7780 15483 8016 15571
rect 9299 15637 9535 15719
rect 9299 15569 9380 15637
rect 9380 15569 9454 15637
rect 9454 15569 9535 15637
rect 9299 15483 9535 15569
rect 10747 15637 10983 15715
rect 10747 15569 10828 15637
rect 10828 15569 10902 15637
rect 10902 15569 10983 15637
rect 10747 15479 10983 15569
rect 12242 15639 12478 15730
rect 14678 15729 14914 15746
rect 12242 15571 12326 15639
rect 12326 15571 12400 15639
rect 12400 15571 12478 15639
rect 12242 15494 12478 15571
rect 13691 15639 13927 15724
rect 13691 15571 13774 15639
rect 13774 15571 13848 15639
rect 13848 15571 13927 15639
rect 13691 15488 13927 15571
rect 14678 15618 14747 15729
rect 14747 15618 14857 15729
rect 14857 15618 14914 15729
rect 14678 15510 14914 15618
rect 15850 15729 16086 15759
rect 15850 15618 15915 15729
rect 15915 15618 16025 15729
rect 16025 15618 16086 15729
rect 15850 15523 16086 15618
rect 17024 15729 17260 15746
rect 17024 15618 17083 15729
rect 17083 15618 17193 15729
rect 17193 15618 17260 15729
rect 17024 15510 17260 15618
rect 18188 15729 18424 15788
rect 18188 15618 18251 15729
rect 18251 15618 18361 15729
rect 18361 15618 18424 15729
rect 18188 15552 18424 15618
rect 19358 15731 19594 15786
rect 19358 15620 19425 15731
rect 19425 15620 19535 15731
rect 19535 15620 19594 15731
rect 19358 15550 19594 15620
rect 20527 15731 20763 15752
rect 20527 15620 20593 15731
rect 20593 15620 20703 15731
rect 20703 15620 20763 15731
rect 20527 15516 20763 15620
rect 21705 15731 21941 15764
rect 21705 15620 21761 15731
rect 21761 15620 21871 15731
rect 21871 15620 21941 15731
rect 21705 15528 21941 15620
rect 22870 15731 23106 15748
rect 22870 15620 22929 15731
rect 22929 15620 23039 15731
rect 23039 15620 23106 15731
rect 22870 15512 23106 15620
rect 4146 12882 4382 12922
rect 4146 12814 4218 12882
rect 4218 12814 4302 12882
rect 4302 12814 4382 12882
rect 4146 12686 4382 12814
rect 7283 12882 7519 12908
rect 7283 12814 7362 12882
rect 7362 12814 7446 12882
rect 7446 12814 7519 12882
rect 7283 12672 7519 12814
rect 10419 12886 10655 12926
rect 10419 12818 10494 12886
rect 10494 12818 10578 12886
rect 10578 12818 10655 12886
rect 10419 12690 10655 12818
rect 13570 12886 13806 12917
rect 13570 12818 13638 12886
rect 13638 12818 13722 12886
rect 13722 12818 13806 12886
rect 13570 12681 13806 12818
rect 16760 12882 16996 12930
rect 16760 12814 16840 12882
rect 16840 12814 16924 12882
rect 16924 12814 16996 12882
rect 16760 12694 16996 12814
rect 19906 12882 20142 12926
rect 19906 12814 19984 12882
rect 19984 12814 20068 12882
rect 20068 12814 20142 12882
rect 19906 12690 20142 12814
rect 23024 12886 23260 12935
rect 23024 12818 23116 12886
rect 23116 12818 23200 12886
rect 23200 12818 23260 12886
rect 23024 12699 23260 12818
rect 26179 12886 26415 12908
rect 26179 12818 26260 12886
rect 26260 12818 26344 12886
rect 26344 12818 26415 12886
rect 26179 12672 26415 12818
rect 4157 10148 4393 10207
rect 4157 10080 4218 10148
rect 4218 10080 4302 10148
rect 4302 10080 4393 10148
rect 4157 9971 4393 10080
rect 7297 10148 7533 10193
rect 7297 10080 7362 10148
rect 7362 10080 7446 10148
rect 7446 10080 7533 10148
rect 7297 9957 7533 10080
rect 10419 10152 10655 10185
rect 10419 10084 10494 10152
rect 10494 10084 10578 10152
rect 10578 10084 10655 10152
rect 10419 9949 10655 10084
rect 13575 10152 13811 10189
rect 13575 10084 13638 10152
rect 13638 10084 13722 10152
rect 13722 10084 13811 10152
rect 13575 9953 13811 10084
rect 16772 10148 17008 10185
rect 16772 10080 16840 10148
rect 16840 10080 16924 10148
rect 16924 10080 17008 10148
rect 16772 9949 17008 10080
rect 19905 10148 20141 10185
rect 19905 10080 19984 10148
rect 19984 10080 20068 10148
rect 20068 10080 20141 10148
rect 19905 9949 20141 10080
rect 23038 10152 23274 10194
rect 23038 10084 23116 10152
rect 23116 10084 23200 10152
rect 23200 10084 23274 10152
rect 23038 9958 23274 10084
rect 26170 10152 26406 10185
rect 26170 10084 26260 10152
rect 26260 10084 26344 10152
rect 26344 10084 26406 10152
rect 26170 9949 26406 10084
rect 4133 7416 4369 7456
rect 4133 7348 4208 7416
rect 4208 7348 4292 7416
rect 4292 7348 4369 7416
rect 4133 7220 4369 7348
rect 7287 7416 7523 7447
rect 7287 7348 7352 7416
rect 7352 7348 7436 7416
rect 7436 7348 7523 7416
rect 7287 7211 7523 7348
rect 10418 7420 10654 7447
rect 10418 7352 10484 7420
rect 10484 7352 10568 7420
rect 10568 7352 10654 7420
rect 10418 7211 10654 7352
rect 13549 7420 13785 7447
rect 13549 7352 13628 7420
rect 13628 7352 13712 7420
rect 13712 7352 13785 7420
rect 13549 7211 13785 7352
rect 16758 7416 16994 7442
rect 16758 7348 16830 7416
rect 16830 7348 16914 7416
rect 16914 7348 16994 7416
rect 16758 7206 16994 7348
rect 19899 7416 20135 7461
rect 19899 7348 19974 7416
rect 19974 7348 20058 7416
rect 20058 7348 20135 7416
rect 19899 7225 20135 7348
rect 23034 7420 23270 7447
rect 23034 7352 23106 7420
rect 23106 7352 23190 7420
rect 23190 7352 23270 7420
rect 23034 7211 23270 7352
rect 26174 7420 26410 7465
rect 26174 7352 26250 7420
rect 26250 7352 26334 7420
rect 26334 7352 26410 7420
rect 26174 7229 26410 7352
rect 19440 5885 19676 5960
rect 19440 5785 19509 5885
rect 19509 5785 19611 5885
rect 19611 5785 19676 5885
rect 19440 5724 19676 5785
rect 20174 5883 20410 5958
rect 20174 5783 20247 5883
rect 20247 5783 20349 5883
rect 20349 5783 20410 5883
rect 20174 5722 20410 5783
rect 20922 5883 21158 5956
rect 20922 5783 20985 5883
rect 20985 5783 21087 5883
rect 21087 5783 21158 5883
rect 20922 5720 21158 5783
rect 21663 5883 21899 5951
rect 21663 5783 21727 5883
rect 21727 5783 21829 5883
rect 21829 5783 21899 5883
rect 21663 5715 21899 5783
rect 22394 5883 22630 5962
rect 22394 5783 22467 5883
rect 22467 5783 22569 5883
rect 22569 5783 22630 5883
rect 22394 5726 22630 5783
rect 23133 5883 23369 5962
rect 23133 5783 23205 5883
rect 23205 5783 23307 5883
rect 23307 5783 23369 5883
rect 23133 5726 23369 5783
rect 23879 5883 24115 5960
rect 23879 5783 23943 5883
rect 23943 5783 24045 5883
rect 24045 5783 24115 5883
rect 23879 5724 24115 5783
rect 24606 5883 24842 5958
rect 24606 5783 24681 5883
rect 24681 5783 24783 5883
rect 24783 5783 24842 5883
rect 24606 5722 24842 5783
rect 3379 4482 3615 4515
rect 3379 4394 3448 4482
rect 3448 4394 3542 4482
rect 3542 4394 3615 4482
rect 3379 4279 3615 4394
rect 5446 4484 5682 4524
rect 5446 4396 5516 4484
rect 5516 4396 5610 4484
rect 5610 4396 5682 4484
rect 5446 4288 5682 4396
rect 7519 4482 7755 4529
rect 7519 4394 7585 4482
rect 7585 4394 7679 4482
rect 7679 4394 7755 4482
rect 7519 4293 7755 4394
rect 9587 4484 9823 4522
rect 9587 4396 9653 4484
rect 9653 4396 9747 4484
rect 9747 4396 9823 4484
rect 9587 4286 9823 4396
rect 11660 4484 11896 4515
rect 11660 4396 11722 4484
rect 11722 4396 11816 4484
rect 11816 4396 11896 4484
rect 11660 4279 11896 4396
rect 13724 4486 13960 4519
rect 13724 4398 13790 4486
rect 13790 4398 13884 4486
rect 13884 4398 13960 4486
rect 13724 4283 13960 4398
rect 15787 4484 16023 4519
rect 15787 4396 15859 4484
rect 15859 4396 15953 4484
rect 15953 4396 16023 4484
rect 15787 4283 16023 4396
rect 17860 4486 18096 4531
rect 17860 4398 17927 4486
rect 17927 4398 18021 4486
rect 18021 4398 18096 4486
rect 17860 4295 18096 4398
<< metal5 >>
rect 3203 15788 26656 15955
rect 3203 15759 18188 15788
rect 3203 15746 15850 15759
rect 3203 15730 14678 15746
rect 3203 15494 3387 15730
rect 3623 15724 12242 15730
rect 3623 15715 6331 15724
rect 3623 15494 4836 15715
rect 3203 15479 4836 15494
rect 5072 15488 6331 15715
rect 6567 15719 12242 15724
rect 6567 15488 7780 15719
rect 5072 15483 7780 15488
rect 8016 15483 9299 15719
rect 9535 15715 12242 15719
rect 9535 15483 10747 15715
rect 5072 15479 10747 15483
rect 10983 15494 12242 15715
rect 12478 15724 14678 15730
rect 12478 15494 13691 15724
rect 10983 15488 13691 15494
rect 13927 15510 14678 15724
rect 14914 15523 15850 15746
rect 16086 15746 18188 15759
rect 16086 15523 17024 15746
rect 14914 15510 17024 15523
rect 17260 15552 18188 15746
rect 18424 15786 26656 15788
rect 18424 15552 19358 15786
rect 17260 15550 19358 15552
rect 19594 15764 26656 15786
rect 19594 15752 21705 15764
rect 19594 15550 20527 15752
rect 17260 15516 20527 15550
rect 20763 15528 21705 15752
rect 21941 15748 26656 15764
rect 21941 15528 22870 15748
rect 20763 15516 22870 15528
rect 17260 15512 22870 15516
rect 23106 15512 26656 15748
rect 17260 15510 26656 15512
rect 13927 15488 26656 15510
rect 10983 15479 26656 15488
rect 3203 12935 26656 15479
rect 3203 12930 23024 12935
rect 3203 12926 16760 12930
rect 3203 12922 10419 12926
rect 3203 12686 4146 12922
rect 4382 12908 10419 12922
rect 4382 12686 7283 12908
rect 3203 12672 7283 12686
rect 7519 12690 10419 12908
rect 10655 12917 16760 12926
rect 10655 12690 13570 12917
rect 7519 12681 13570 12690
rect 13806 12694 16760 12917
rect 16996 12926 23024 12930
rect 16996 12694 19906 12926
rect 13806 12690 19906 12694
rect 20142 12699 23024 12926
rect 23260 12908 26656 12935
rect 23260 12699 26179 12908
rect 20142 12690 26179 12699
rect 13806 12681 26179 12690
rect 7519 12672 26179 12681
rect 26415 12672 26656 12908
rect 3203 10207 26656 12672
rect 3203 9971 4157 10207
rect 4393 10194 26656 10207
rect 4393 10193 23038 10194
rect 4393 9971 7297 10193
rect 3203 9957 7297 9971
rect 7533 10189 23038 10193
rect 7533 10185 13575 10189
rect 7533 9957 10419 10185
rect 3203 9949 10419 9957
rect 10655 9953 13575 10185
rect 13811 10185 23038 10189
rect 13811 9953 16772 10185
rect 10655 9949 16772 9953
rect 17008 9949 19905 10185
rect 20141 9958 23038 10185
rect 23274 10185 26656 10194
rect 23274 9958 26170 10185
rect 20141 9949 26170 9958
rect 26406 9949 26656 10185
rect 3203 7465 26656 9949
rect 3203 7461 26174 7465
rect 3203 7456 19899 7461
rect 3203 7220 4133 7456
rect 4369 7447 19899 7456
rect 4369 7220 7287 7447
rect 3203 7211 7287 7220
rect 7523 7211 10418 7447
rect 10654 7211 13549 7447
rect 13785 7442 19899 7447
rect 13785 7211 16758 7442
rect 3203 7206 16758 7211
rect 16994 7225 19899 7442
rect 20135 7447 26174 7461
rect 20135 7225 23034 7447
rect 16994 7211 23034 7225
rect 23270 7229 26174 7447
rect 26410 7229 26656 7465
rect 23270 7211 26656 7229
rect 16994 7206 26656 7211
rect 3203 5962 26656 7206
rect 3203 5960 22394 5962
rect 3203 5724 19440 5960
rect 19676 5958 22394 5960
rect 19676 5724 20174 5958
rect 3203 5722 20174 5724
rect 20410 5956 22394 5958
rect 20410 5722 20922 5956
rect 3203 5720 20922 5722
rect 21158 5951 22394 5956
rect 21158 5720 21663 5951
rect 3203 5715 21663 5720
rect 21899 5726 22394 5951
rect 22630 5726 23133 5962
rect 23369 5960 26656 5962
rect 23369 5726 23879 5960
rect 21899 5724 23879 5726
rect 24115 5958 26656 5960
rect 24115 5724 24606 5958
rect 21899 5722 24606 5724
rect 24842 5722 26656 5958
rect 21899 5715 26656 5722
rect 3203 4531 26656 5715
rect 3203 4529 17860 4531
rect 3203 4524 7519 4529
rect 3203 4515 5446 4524
rect 3203 4279 3379 4515
rect 3615 4288 5446 4515
rect 5682 4293 7519 4524
rect 7755 4522 17860 4529
rect 7755 4293 9587 4522
rect 5682 4288 9587 4293
rect 3615 4286 9587 4288
rect 9823 4519 17860 4522
rect 9823 4515 13724 4519
rect 9823 4286 11660 4515
rect 3615 4279 11660 4286
rect 11896 4283 13724 4515
rect 13960 4283 15787 4519
rect 16023 4295 17860 4519
rect 18096 4295 26656 4531
rect 16023 4283 26656 4295
rect 11896 4279 26656 4283
rect 3203 3832 26656 4279
use aritmetic_unit_pex  aritmetic_unit_pex_0
timestamp 1736796407
transform 1 0 33758 0 1 -3087
box -4203 -805 39597 29436
<< labels >>
flabel metal4 12520 22154 12882 22318 1 FreeSerif 960 0 0 0 shifter_unit_0.VDD
flabel metal4 12492 19860 12878 19988 1 FreeSerif 960 0 0 0 shifter_unit_0.VSS
flabel metal1 25605 21157 25681 21237 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[7]
flabel metal1 25633 20796 25675 20864 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[6]
flabel metal1 25631 20667 25676 20727 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[5]
flabel metal1 25624 20502 25677 20571 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[4]
flabel metal1 25617 20349 25678 20425 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[3]
flabel metal1 25609 20207 25684 20290 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[2]
flabel metal1 25606 20075 25679 20152 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[1]
flabel metal1 25617 19806 25673 19873 1 FreeSerif 720 0 0 0 shifter_unit_0.Y[0]
flabel metal1 64 21221 130 21297 1 FreeSerif 720 0 0 0 shifter_unit_0.dir
flabel metal1 67 20939 136 21009 1 FreeSerif 720 0 0 0 shifter_unit_0.A[1]
flabel metal1 69 20711 133 20761 1 FreeSerif 720 0 0 0 shifter_unit_0.A[2]
flabel metal1 68 20575 130 20627 1 FreeSerif 720 0 0 0 shifter_unit_0.A[3]
flabel metal1 68 20465 118 20515 1 FreeSerif 720 0 0 0 shifter_unit_0.A[4]
flabel metal1 75 20099 121 20147 1 FreeSerif 720 0 0 0 shifter_unit_0.A[6]
flabel metal1 65 20336 121 20392 1 FreeSerif 720 0 0 0 shifter_unit_0.A[5]
flabel metal1 77 19883 150 19918 1 FreeSerif 720 0 0 0 shifter_unit_0.A[7]
flabel metal1 64 21382 146 21436 1 FreeSerif 720 0 0 0 shifter_unit_0.A[0]
flabel metal5 20062 4001 22229 4739 1 FreeSerif 3200 0 0 0 logic_unit_0.VSS
flabel metal4 13900 16767 14605 17092 1 FreeSerif 1600 0 0 0 logic_unit_0.VDD
flabel metal1 408 5639 450 5688 1 FreeSerif 640 0 0 0 logic_unit_0.A[0]
flabel metal1 406 5845 455 5898 1 FreeSerif 640 0 0 0 logic_unit_0.A[1]
flabel metal1 410 6033 468 6087 1 FreeSerif 640 0 0 0 logic_unit_0.A[2]
flabel metal1 408 6340 467 6396 1 FreeSerif 640 0 0 0 logic_unit_0.A[4]
flabel metal1 406 6189 470 6243 1 FreeSerif 640 0 0 0 logic_unit_0.A[3]
flabel metal1 406 6500 468 6558 1 FreeSerif 640 0 0 0 logic_unit_0.A[5]
flabel metal1 408 6809 465 6861 1 FreeSerif 720 0 0 0 logic_unit_0.A[6]
flabel metal1 408 7100 468 7153 1 FreeSerif 720 0 0 0 logic_unit_0.A[7]
flabel metal1 128 15454 166 15502 1 FreeSerif 720 0 0 0 logic_unit_0.B[0]
flabel metal1 129 15829 190 15875 1 FreeSerif 720 0 0 0 logic_unit_0.B[1]
flabel metal1 128 17619 188 17678 1 FreeSerif 720 0 0 0 logic_unit_0.B[2]
flabel metal1 127 17816 187 17875 1 FreeSerif 720 0 0 0 logic_unit_0.B[3]
flabel metal1 129 18000 189 18059 1 FreeSerif 720 0 0 0 logic_unit_0.B[4]
flabel metal1 129 18187 189 18246 1 FreeSerif 720 0 0 0 logic_unit_0.B[5]
flabel metal1 130 18377 190 18436 1 FreeSerif 720 0 0 0 logic_unit_0.B[6]
flabel metal1 131 18579 190 18634 1 FreeSerif 720 0 0 0 logic_unit_0.B[7]
flabel metal1 103 11353 173 11425 1 FreeSerif 720 0 0 0 logic_unit_0.opcode[1]
flabel metal1 101 11027 179 11095 1 FreeSerif 720 0 0 0 logic_unit_0.opcode[0]
flabel metal1 27954 11231 28043 11361 1 FreeSerif 720 0 0 0 logic_unit_0.Y[7]
flabel metal1 27996 10872 28044 10934 1 FreeSerif 720 0 0 0 logic_unit_0.Y[6]
flabel metal1 27991 10681 28044 10743 1 FreeSerif 720 0 0 0 logic_unit_0.Y[5]
flabel metal1 27991 10459 28042 10521 1 FreeSerif 720 0 0 0 logic_unit_0.Y[4]
flabel metal1 27986 10268 28041 10332 1 FreeSerif 720 0 0 0 logic_unit_0.Y[3]
flabel metal1 27986 9927 28042 9991 1 FreeSerif 720 0 0 0 logic_unit_0.Y[2]
flabel metal1 27990 9755 28043 9816 1 FreeSerif 720 0 0 0 logic_unit_0.Y[1]
flabel metal1 27990 9395 28048 9460 1 FreeSerif 720 0 0 0 logic_unit_0.Y[0]
<< end >>
