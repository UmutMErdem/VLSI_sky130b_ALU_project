magic
tech sky130B
magscale 1 2
timestamp 1736110742
<< nwell >>
rect 458 1226 1372 1504
rect 888 418 1372 1226
<< psubdiff >>
rect 538 82 734 112
rect 538 16 578 82
rect 696 16 734 82
rect 538 -32 734 16
<< nsubdiff >>
rect 978 1426 1244 1464
rect 978 1354 1034 1426
rect 1178 1354 1244 1426
rect 978 1324 1244 1354
<< psubdiffcont >>
rect 578 16 696 82
<< nsubdiffcont >>
rect 1034 1354 1178 1426
<< poly >>
rect 400 1348 466 1364
rect 400 1314 416 1348
rect 450 1344 466 1348
rect 450 1314 950 1344
rect 400 1301 950 1314
rect 400 1298 466 1301
rect 400 1249 466 1256
rect 906 1249 950 1301
rect 400 1240 848 1249
rect 400 1206 416 1240
rect 450 1208 848 1240
rect 906 1208 1202 1249
rect 450 1207 584 1208
rect 450 1206 466 1207
rect 400 1190 466 1206
rect 552 681 613 770
rect 462 628 613 681
rect 462 410 522 628
rect 906 586 966 771
rect 580 535 966 586
rect 580 408 640 535
rect 695 477 761 493
rect 695 443 711 477
rect 745 443 761 477
rect 695 427 761 443
rect 698 172 758 194
rect 981 172 1041 194
rect 1099 172 1159 194
rect 1217 172 1277 194
rect 698 131 1277 172
<< polycont >>
rect 416 1314 450 1348
rect 416 1206 450 1240
rect 711 443 745 477
<< locali >>
rect 1002 1426 1206 1438
rect 1002 1354 1034 1426
rect 1178 1354 1206 1426
rect 1002 1352 1064 1354
rect 1144 1352 1206 1354
rect 400 1314 416 1348
rect 450 1314 466 1348
rect 1002 1336 1206 1352
rect 400 1206 416 1240
rect 450 1206 466 1240
rect 695 443 711 477
rect 745 443 761 477
rect 560 86 702 98
rect 560 82 600 86
rect 666 82 702 86
rect 560 16 578 82
rect 696 16 702 82
rect 560 -10 702 16
<< viali >>
rect 1064 1354 1144 1424
rect 1064 1352 1144 1354
rect 416 1314 450 1348
rect 416 1206 450 1240
rect 711 443 745 477
rect 600 82 666 86
rect 600 16 666 82
<< metal1 >>
rect 366 1348 466 1450
rect 366 1314 416 1348
rect 450 1314 466 1348
rect 1052 1424 1156 1430
rect 1052 1352 1064 1424
rect 1144 1352 1156 1424
rect 1052 1346 1156 1352
rect 366 1288 466 1314
rect 1087 1290 1122 1346
rect 366 1240 466 1260
rect 366 1206 416 1240
rect 450 1206 466 1240
rect 366 1108 466 1206
rect 624 1249 894 1277
rect 624 1184 658 1249
rect 860 1184 894 1249
rect 978 1249 1248 1290
rect 978 1180 1012 1249
rect 1214 1180 1248 1249
rect 506 745 540 816
rect 742 745 776 816
rect 506 717 776 745
rect 860 746 894 816
rect 1096 746 1130 816
rect 860 717 1130 746
rect 506 669 540 717
rect 506 639 569 669
rect 534 547 569 639
rect 1214 604 1248 788
rect 534 511 761 547
rect 534 364 569 511
rect 695 477 761 511
rect 695 443 711 477
rect 745 443 761 477
rect 1042 535 1139 586
rect 1214 550 1323 604
rect 1042 468 1099 535
rect 695 437 761 443
rect 936 432 1205 468
rect 936 394 969 432
rect 1172 397 1205 432
rect 1289 383 1323 550
rect 787 249 952 337
rect 416 165 450 218
rect 652 165 686 214
rect 416 126 686 165
rect 1053 166 1086 213
rect 1289 166 1322 213
rect 1053 130 1322 166
rect 616 98 650 126
rect 594 86 672 98
rect 594 16 600 86
rect 666 16 672 86
rect 594 4 672 16
<< via1 >>
rect 1078 1353 1130 1405
rect 607 29 659 81
<< metal2 >>
rect 1056 1426 1146 1436
rect 1056 1325 1146 1335
rect 591 99 681 109
rect 591 -2 681 8
<< via2 >>
rect 1056 1405 1146 1426
rect 1056 1353 1078 1405
rect 1078 1353 1130 1405
rect 1130 1353 1146 1405
rect 1056 1335 1146 1353
rect 591 81 681 99
rect 591 29 607 81
rect 607 29 659 81
rect 659 29 681 81
rect 591 8 681 29
<< metal3 >>
rect 1028 1320 1038 1440
rect 1160 1320 1170 1440
rect 571 -2 581 109
rect 691 -2 701 109
<< via3 >>
rect 1038 1426 1160 1440
rect 1038 1335 1056 1426
rect 1056 1335 1146 1426
rect 1146 1335 1160 1426
rect 1038 1320 1160 1335
rect 581 99 691 109
rect 581 8 591 99
rect 591 8 681 99
rect 681 8 691 99
rect 581 -2 691 8
<< metal4 >>
rect 954 1440 1258 1504
rect 954 1320 1038 1440
rect 1160 1320 1258 1440
rect 954 1310 1258 1320
rect 580 109 692 110
rect 580 98 581 109
rect 522 -2 581 98
rect 691 98 692 109
rect 691 -2 752 98
rect 522 -64 752 -2
use sky130_fd_pr__nfet_01v8_CLVMSK  sky130_fd_pr__nfet_01v8_CLVMSK_0
timestamp 1734818450
transform 1 0 610 0 1 304
box -206 -126 206 126
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_0
timestamp 1734818450
transform 1 0 877 0 1 987
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_0
timestamp 1734818450
transform 1 0 1129 0 1 304
box -242 -162 242 162
<< labels >>
flabel metal1 1049 541 1132 580 1 FreeSans 240 0 0 0 OUT
port 6 n
flabel metal4 1024 1320 1188 1432 1 FreeSerif 560 0 0 0 VDD
port 9 n
flabel metal4 548 -22 720 88 1 FreeSerif 560 0 0 0 VSS
port 10 n
flabel metal1 366 1110 464 1208 1 FreeSerif 480 0 0 0 A
port 14 n
flabel metal1 368 1378 466 1446 1 FreeSerif 480 0 0 0 B
port 15 n
<< end >>
