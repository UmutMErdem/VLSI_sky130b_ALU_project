* NGSPICE file created from carry_ripple_adder_pex.ext - technology: sky130B

.subckt carry_ripple_adder A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7] B[0],B[1],B[2],B[3],B[4],B[5],B[6],B[7] carry_in VDD VSS Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7] carry_out

X0 VDD.t151 a_7564_3012# a_8154_2575# w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X1 a_22002_2394# B[3].t0 VDD.t425 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X2 a_19659_n3206# a_19657_n3503.t4 VDD.t200 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X3 a_17433_4533# a_14688_2570# a_17551_4533# w_17397_4471# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X4 VDD.t81 a_1046_1411# a_1636_974# w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X5 VDD.t308 a_15222_n1096# a_15282_n1070# w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X6 VDD.t137 a_4101_n969# a_2130_n1097# w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X7 VDD.t9 a_20593_n1089# a_20653_n1063# w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X8 VSS.t156 B[0].t0 a_1274_4028# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X9 a_9749_1676# A[1].t0 VSS.t62 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X10 a_4741_n4834# a_52_n3507.t4 VSS.t84 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X11 a_4087_n2619# a_52_n3507.t5 a_4736_n3230# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X12 a_21660_n1723# a_21735_n1093# VSS.t68 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X13 a_3244_4537# a_1636_974# a_3362_4537# w_3208_4475# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X14 a_17551_4533# a_16555_3946# VDD.t478 w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X15 a_5134_1679# carry_in.t0 VDD.t354 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X16 VSS.t154 a_4087_n2619# a_1342_n1093# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X17 a_23706_n965# B[4].t0 VDD.t342 w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X18 Y[7].t3 a_54_n3210# a_594_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X19 VSS.t157 B[0].t1 a_2397_2398# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X20 a_7559_1408# A[1].t1 VDD.t232 w_7405_1346# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X21 a_5134_1679# carry_in.t1 VSS.t110 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X22 VDD.t414 a_19657_n3503.t5 a_19659_n3206# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X23 VDD.t477 a_16555_3946# a_17551_4533# w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X24 VDD.t64 a_9455_1702.t8 a_11235_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X25 a_18181_1671# a_11163_3955.t4 VDD.t16 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X26 a_24681_969# a_22547_1701# Y[3].t3 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X27 Y[7].t0 a_949_n3236.t8 a_948_n4635# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X28 a_17842_n1579# B[5].t0 VSS.t139 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X29 a_21232_4224# a_20642_4661# VDD.t325 w_20488_4599# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X30 a_17342_2390# a_15989_1697# VDD.t484 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X31 VDD.t117 a_14084_4657# a_14674_4220# w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X32 VSS.t2 a_9042_n1101# a_8613_n1731# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X33 a_9050_n3907# a_9462_n3933# a_7507_n3240.t2 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X34 a_7801_2375# a_4650_3958.t4 a_7564_3012# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X35 VDD.t34 A[2].t0 a_16283_1671# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X36 VSS.t101 a_4650_3958.t5 a_11589_970# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X37 a_4722_1705# a_2942_1705.t8 VDD.t432 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X38 a_21246_2574# a_20656_3011# VDD.t379 w_20502_2949# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X39 VDD.t124 B[2].t0 a_15444_2390# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X40 a_2492_n3903# A[7].t0 VDD.t18 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X41 a_9455_1702.t2 a_8910_2395# a_9337_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X42 a_7471_n1727# a_7900_n1097# a_7606_n1071# w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X43 a_988_n1093# a_2055_n1727# VDD.t198 w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X44 VDD.t86 A[4].t0 a_21557_n3206# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X45 a_712_n4635# a_1006_n3929# Y[7].t7 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X46 a_10659_n973# B[6].t0 VDD.t314 w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X47 a_7152_n3907# a_6612_n3214# Y[6].t2 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X48 VDD.t253 B[0].t2 a_1037_4665# w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X49 VDD.t297 B[7].t0 a_4087_n2619# w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X50 a_2942_1705.t6 a_3236_1679# a_2824_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X51 VDD.t262 A[3].t0 a_20651_1407# w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X52 a_9875_4534# a_8140_4225# VDD.t239 w_9721_4472# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X53 VDD.t17 a_11163_3955.t5 a_17769_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X54 VDD.t197 a_2055_n1727# a_988_n1093# w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X55 a_21557_n3206# A[4].t1 VDD.t10 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X56 VDD.t224 B[0].t3 a_1051_3015# w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X57 Y[6].t1 a_6612_n3214# a_7152_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X58 VDD.t204 B[6].t1 a_9462_n3933# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X59 VDD.t65 a_9455_1702.t9 a_10808_2395# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X60 a_4087_n2619# B[7].t1 VDD.t159 w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X61 a_16283_1671# A[2].t1 VSS.t44 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X62 VDD.t136 a_4101_n969# a_2130_n1097# w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 a_13686_n3902# a_14041_n3235# VDD.t6 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X64 a_15871_1697.t5 B[2].t1 VDD.t125 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X65 a_6612_n3214# a_6610_n3511.t4 VDD.t92 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X66 VDD.t443 a_17697_3950.t4 a_20651_1407# w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X67 VDD.t407 a_17193_n968# a_15222_n1096# w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X68 Y[0].t0 a_4295_2398# a_4840_973# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X69 a_988_n1093# a_2055_n1727# VDD.t196 w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X70 VDD.t11 A[4].t2 a_21557_n3206# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X71 VDD.t12 A[4].t3 a_22097_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X72 VDD.t50 A[6].t0 a_8510_n3214# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X73 VDD.t181 a_1627_4228# a_3362_4537# w_3208_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X74 a_17769_1697# a_18181_1671# Y[2].t6 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X75 a_7152_n3907# a_7564_n3933# Y[6].t6 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X76 a_9462_n3933# B[6].t2 VDD.t319 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X77 a_4101_n969# B[7].t2 VDD.t160 w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X78 a_19657_n3503.t3 a_23991_4537# VDD.t261 w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X79 a_1046_1411# A[0].t0 VDD.t450 w_892_1349# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X80 a_17193_n968# A[5].t0 VDD.t268 w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X81 VDD.t403 a_913_n1723# carry_out.t3 w_819_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X82 a_5134_1679# carry_in.t2 VDD.t362 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X83 VDD.t61 a_52_n3507.t6 a_4087_n2619# w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X84 a_23706_n965# A[4].t4 VDD.t386 w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X85 VSS.t90 a_15576_n1096# a_15147_n1726# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X86 VDD.t5 a_14041_n3235# a_13686_n3902# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X87 VDD.t338 a_4650_3958.t6 a_7559_1408# w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X88 a_17828_n3229# B[5].t1 VSS.t73 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X89 VDD.t442 A[0].t1 a_3236_1679# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X90 VDD.t111 a_4650_3958.t7 a_11235_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X91 VDD.t84 a_22849_4533# a_23113_3950# w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X92 VDD.t225 B[0].t4 a_2397_2398# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X93 a_22097_n3899# A[4].t5 VDD.t387 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X94 Y[6].t5 a_7564_n3933# a_7152_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X95 a_4504_4541# a_3508_3954# VDD.t207 w_4350_4479# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X96 VDD.t212 B[2].t2 a_15444_2390# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X97 VDD.t248 A[3].t1 a_22429_1701.t8 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X98 VDD.t347 B[1].t0 a_7550_4662# w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X99 VDD.t383 a_14098_3007# a_14688_2570# w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X100 Y[0].t3 a_4295_2398# a_4722_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X101 a_17833_n4833# a_13144_n3506.t4 VSS.t80 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X102 a_17179_n2618# a_13144_n3506.t5 a_17828_n3229# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X103 a_7152_n3907# a_6610_n3511.t5 VDD.t340 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X104 VSS.t98 a_17179_n2618# a_14434_n1092# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X105 a_11017_4538# a_10021_3951# VDD.t26 w_10863_4476# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X106 VDD.t131 a_949_n3236.t9 a_594_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X107 VDD.t343 B[4].t1 a_22097_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X108 VDD.t190 B[6].t3 a_9050_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X109 VDD.t206 a_3508_3954# a_4504_4541# w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X110 a_9455_1702.t1 a_8910_2395# a_9337_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X111 a_2942_973# a_3236_1679# VSS.t118 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X112 a_10645_n2623# B[6].t4 VDD.t191 w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X113 VDD.t490 a_1037_4665# a_1627_4228# w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X114 a_10021_3951# a_9757_4534# VSS.t79 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X115 VDD.t112 a_4650_3958.t8 a_7564_3012# w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X116 VDD.t451 a_17433_4533# a_17697_3950.t3 w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X117 a_22509_n3925# B[4].t2 VSS.t105 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X118 a_17184_n4222# A[5].t1 a_17833_n4833# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X119 a_2824_1705# B[0].t5 VDD.t358 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X120 a_22097_n3899# B[4].t3 VDD.t280 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X121 a_9050_n3907# B[6].t5 VDD.t171 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X122 VSS.t30 A[7].t1 a_1952_n3210# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X123 VDD.t334 a_4092_n4223# a_2484_n1097# w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X124 a_1046_1411# A[0].t2 VDD.t201 w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X125 a_2190_n1071# a_2130_n1097# VDD.t357 w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X126 VDD.t233 A[1].t2 a_9749_1676# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X127 VSS.t6 B[1].t1 a_7787_4025# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X128 a_15584_n3902.t5 A[5].t2 VDD.t236 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X129 a_9757_4534# a_8149_971# a_9875_4534# w_9721_4472# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X130 a_15871_1697.t11 A[2].t2 VDD.t146 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X131 a_13804_n4634# a_14098_n3928# Y[5].t1 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X132 a_14080_n1092# a_15147_n1726# VDD.t211 w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X133 a_15989_1697# a_15444_2390# a_15871_1697.t2 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X134 a_2904_n3929# B[7].t3 VDD.t287 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X135 a_20199_n3899# a_19657_n3503.t6 VDD.t415 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X136 a_23692_n2615# B[4].t4 VDD.t281 w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X137 a_20642_4661# A[3].t2 VDD.t249 w_20488_4599# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X138 VDD.t172 B[6].t6 a_9050_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X139 a_15871_1697.t1 a_15444_2390# a_15989_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X140 a_24327_1701.t2 a_24739_1675# Y[3].t2 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X141 VSS.t40 a_4101_n969# a_2130_n1097# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X142 a_594_n3903# a_1006_n3929# Y[7].t6 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X143 a_14084_4657# A[2].t3 VDD.t147 w_13930_4595# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X144 VDD.t220 a_22547_1701# a_24327_1701.t5 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X145 a_22429_1701.t5 a_22002_2394# a_22547_1701# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X146 VDD.t210 a_15147_n1726# a_14080_n1092# w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X147 VSS.t135 a_21232_4224# a_22849_4533# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X148 VSS.t117 a_19659_n3206# a_20317_n4631# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X149 a_16555_3946# a_16291_4529# VDD.t21 w_16255_4467# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X150 Y[3].t5 a_23900_2394# a_24445_969# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X151 a_24739_1675# a_17697_3950.t5 VSS.t43 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X152 VDD.t282 B[4].t5 a_23692_n2615# w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X153 a_6610_n3511.t3 a_14005_n1722# VDD.t390 w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X154 VDD.t175 a_7559_1408# a_8149_971# w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X155 a_21232_4224# a_20642_4661# VDD.t324 w_20488_4599# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X156 a_17179_n2618# B[5].t2 VDD.t255 w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X157 VDD.t275 a_9757_4534# a_10021_3951# w_9721_4472# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X158 a_10650_n4227# a_6610_n3511.t6 VDD.t341 w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X159 a_21232_4224# a_20642_4661# VSS.t96 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X160 a_23113_3950# a_22849_4533# VSS.t22 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X161 VDD.t176 B[3].t1 a_20656_3011# w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X162 Y[7].t5 a_1006_n3929# a_594_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X163 a_7606_n1071# a_7900_n1097# a_7471_n1727# w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X164 a_20653_n1063# a_20947_n1089# a_20518_n1719# w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X165 VDD.t373 a_10659_n973# a_8688_n1101# w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X166 a_1636_974# a_1046_1411# VSS.t21 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X167 a_11589_970# a_9455_1702.t10 Y[1].t0 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X168 a_20611_n3925# a_20554_n3232.t8 VDD.t318 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X169 a_14080_n1092# a_15147_n1726# VDD.t209 w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X170 VDD.t247 a_4386_4541# a_4650_3958.t3 w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X171 a_24109_4537# a_21246_2574# a_23991_4537# w_23955_4475# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X172 a_20879_4024# A[3].t3 a_20642_4661# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X173 a_20553_n4631# a_19657_n3503.t7 VSS.t103 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X174 VDD.t128 A[7].t2 a_4092_n4223# w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X175 a_22967_4533# a_21241_970# a_22849_4533# w_22813_4471# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X176 VDD.t234 A[1].t3 a_9337_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X177 a_14683_966# a_14093_1403# VDD.t158 w_13939_1341# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X178 a_23692_n2615# B[4].t6 VDD.t309 w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X179 VDD.t392 a_14005_n1722# a_6610_n3511.t2 w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X180 a_8140_4225# a_7550_4662# VDD.t230 w_7396_4600# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X181 a_9455_1702.t7 a_9749_1676# a_9337_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X182 VDD.t182 a_13144_n3506.t6 a_17179_n2618# w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X183 VDD.t202 a_6610_n3511.t7 a_10650_n4227# w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X184 a_21795_n1067# a_22089_n1093# a_21660_n1723# w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X185 a_22849_4533# a_21241_970# a_22967_4533# w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X186 VDD.t164 B[1].t2 a_7564_3012# w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X187 VDD.t363 carry_in.t3 a_4722_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X188 a_9337_1702# B[1].t3 VDD.t303 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X189 a_24739_1675# a_17697_3950.t6 VDD.t145 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X190 a_594_n3903# a_1006_n3929# Y[7].t4 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X191 a_17769_1697# a_15989_1697# VDD.t487 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X192 a_7471_n1727# a_7900_n1097# a_7606_n1071# w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X193 a_20518_n1719# a_20947_n1089# a_20653_n1063# w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X194 VDD.t463 a_20554_n3232.t9 a_20611_n3925# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X195 VDD.t165 a_7507_n3240.t8 a_7564_n3933# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X196 a_6610_n3511.t1 a_14005_n1722# VDD.t391 w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X197 VDD.t219 a_22547_1701# a_23900_2394# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X198 VDD.t74 a_14080_n1092# a_14140_n1066# w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X199 a_1037_4665# A[0].t3 VDD.t454 w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X200 a_2824_1705# A[0].t4 VDD.t40 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X201 a_1046_1411# carry_in.t4 VDD.t364 w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X202 a_17184_n4222# A[5].t3 VDD.t87 w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X203 VDD.t502 a_1051_3015# a_1641_2578# w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X204 a_10650_n4227# a_6610_n3511.t8 VDD.t203 w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X205 a_21660_n1723# a_22089_n1093# a_21795_n1067# w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X206 a_23697_n4219# a_19657_n3503.t8 VDD.t416 w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X207 a_21735_n1093# a_23706_n965# VDD.t278 w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X208 VDD.t129 A[7].t3 a_1952_n3210# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X209 a_20611_n3925# a_20554_n3232.t10 VDD.t185 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X210 a_7564_n3933# a_7507_n3240.t9 VDD.t166 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X211 VDD.t186 A[7].t4 a_4101_n969# w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X212 VDD.t256 B[5].t3 a_17193_n968# w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X213 Y[1].t3 a_10808_2395# a_11235_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X214 carry_out.t2 a_913_n1723# VDD.t402 w_819_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X215 VDD.t459 a_23692_n2615# a_20947_n1089# w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X216 VDD.t195 B[1].t4 a_8910_2395# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X217 a_8149_971# a_7559_1408# VSS.t50 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X218 a_14084_4657# B[2].t3 VDD.t213 w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X219 VDD.t444 a_17697_3950.t7 a_24327_1701.t11 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X220 Y[4].t3 a_19659_n3206# a_20199_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X221 VSS.t25 a_15044_n3209# a_15702_n4634# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X222 a_11235_1702# a_11647_1676# Y[1].t7 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X223 a_15282_n1070# a_15222_n1096# VDD.t307 w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X224 a_16291_4529# a_14683_966# VSS.t7 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X225 a_22547_969# a_22841_1675# VSS.t138 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X226 VDD.t401 a_17184_n4222# a_15576_n1096# w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X227 a_1641_2578# a_1051_3015# VSS.t159 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X228 a_8910_2395# B[1].t5 VDD.t134 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X229 VSS.t4 A[5].t4 a_15044_n3209# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X230 a_20653_n1063# a_20593_n1089# VDD.t8 w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X231 a_4092_n4223# A[7].t5 a_4741_n4834# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X232 VSS.t99 a_4092_n4223# a_2484_n1097# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X233 a_52_n3507.t3 a_7471_n1727# VDD.t398 w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X234 a_22429_1701.t2 B[3].t2 VDD.t177 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X235 a_14098_3007# a_11163_3955.t6 VDD.t430 w_13944_2945# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X236 a_1048_n1067# a_988_n1093# VDD.t367 w_819_n1712# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X237 a_15996_n3928# B[5].t4 VDD.t188 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X238 a_949_n3236.t7 a_1952_n3210# a_2492_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X239 VSS.t8 A[2].t4 a_16225_965# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X240 a_20199_n3899# a_19659_n3206# Y[4].t2 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X241 a_15147_n1726# a_15576_n1096# a_15282_n1070# w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X242 a_4504_4541# a_1641_2578# a_4386_4541# w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X243 a_7546_n1097# a_8613_n1731# VDD.t370 w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X244 VSS.t155 B[0].t6 a_1288_2378# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X245 Y[0].t2 a_4295_2398# a_4722_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X246 a_14683_966# a_14093_1403# VDD.t157 w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X247 a_20593_n1089# a_21660_n1723# VDD.t328 w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X248 a_20518_n1719# a_20947_n1089# a_20653_n1063# w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X249 a_11017_4538# a_8154_2575# a_10899_4538# w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X250 a_24109_4537# a_23113_3950# VDD.t96 w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X251 VSS.t100 carry_in.t5 a_1283_774# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X252 VSS.t134 a_17193_n968# a_15222_n1096# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X253 a_1037_4665# A[0].t5 VDD.t305 w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X254 a_4650_3958.t0 a_4386_4541# VSS.t70 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X255 a_9337_1702# B[1].t6 VDD.t384 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X256 VSS.t114 A[0].t6 a_3178_973# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X257 a_8140_4225# a_7550_4662# VDD.t229 w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X258 a_3508_3954# a_3244_4537# VDD.t54 w_3208_4475# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X259 VSS.t150 a_16555_3946# a_17433_4533# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X260 a_4722_1705# a_5134_1679# Y[0].t6 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X261 a_16409_4529# a_14683_966# a_16291_4529# w_16255_4467# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X262 VDD.t189 B[5].t5 a_15996_n3928# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X263 a_2824_1705# a_2397_2398# a_2942_1705.t2 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X264 a_24739_1675# a_17697_3950.t8 VDD.t445 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X265 Y[4].t1 a_19659_n3206# a_20199_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X266 VSS.t88 a_20518_n1719# a_13144_n3506.t0 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X267 a_11647_1676# a_4650_3958.t9 VDD.t113 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X268 a_22089_n1093# a_23697_n4219# VDD.t163 w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X269 a_15282_n1070# a_15576_n1096# a_15147_n1726# w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X270 VDD.t369 a_8613_n1731# a_7546_n1097# w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X271 VSS.t51 a_1627_4228# a_3244_4537# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X272 a_8748_n1075# a_8688_n1101# VDD.t294 w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X273 a_10808_2395# a_9455_1702.t11 VDD.t473 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X274 VDD.t138 A[3].t4 a_22841_1675# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X275 a_11647_1676# a_4650_3958.t10 VSS.t63 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X276 a_8154_2575# a_7564_3012# VDD.t150 w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X277 Y[5].t4 a_14098_n3928# a_13686_n3902# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X278 VSS.t9 a_2942_1705.t9 a_4295_2398# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X279 VSS.t140 a_11163_3955.t7 a_14330_766# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X280 Y[2].t3 a_17342_2390# a_17887_965# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X281 a_20518_n1719# a_20593_n1089# VSS.t1 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X282 a_7471_n1727# a_7546_n1097# VSS.t42 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X283 Y[1].t4 a_10808_2395# a_11353_970# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X284 VDD.t162 a_23697_n4219# a_22089_n1093# w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X285 a_1274_4028# A[0].t7 a_1037_4665# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X286 a_3362_4537# a_1636_974# a_3244_4537# w_3208_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X287 VDD.t476 a_16555_3946# a_17551_4533# w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X288 Y[3].t4 a_23900_2394# a_24327_1701.t8 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X289 VDD.t310 B[4].t7 a_23706_n965# w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X290 VDD.t235 A[1].t4 a_7559_1408# w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X291 a_20642_4661# A[3].t5 VDD.t470 w_20488_4599# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X292 a_13686_n3902# a_14098_n3928# Y[5].t3 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X293 VDD.t469 A[5].t5 a_17193_n968# w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X294 a_15871_1697.t8 a_16283_1671# a_15989_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X295 a_21241_970# a_20651_1407# VSS.t28 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X296 VDD.t431 a_11163_3955.t8 a_18181_1671# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X297 a_4295_2398# a_2942_1705.t10 VDD.t38 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X298 a_7559_1408# a_4650_3958.t11 VDD.t222 w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X299 VSS.t55 a_20947_n1089# a_20518_n1719# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X300 VSS.t18 a_7900_n1097# a_7471_n1727# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X301 VDD.t323 a_20642_4661# a_21232_4224# w_20488_4599# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X302 a_11163_3955.t0 a_10899_4538# VSS.t158 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X303 a_14674_4220# a_14084_4657# VDD.t116 w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X304 carry_out.t1 a_913_n1723# VDD.t404 w_819_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X305 VDD.t429 A[5].t6 a_15044_n3209# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X306 VDD.t62 a_52_n3507.t7 a_4087_n2619# w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X307 VSS.t74 a_22089_n1093# a_21660_n1723# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X308 a_16283_1671# A[2].t5 VDD.t32 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X309 VDD.t33 A[2].t6 a_14093_1403# w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X310 a_14098_3007# B[2].t4 VDD.t214 w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X311 VDD.t246 a_4386_4541# a_4650_3958.t2 w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X312 VDD.t496 a_4087_n2619# a_1342_n1093# w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X313 a_1037_4665# B[0].t7 VDD.t22 w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X314 a_15989_965# a_16283_1671# VSS.t95 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X315 a_21246_2574# a_20656_3011# VDD.t378 w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X316 a_17193_n968# A[5].t7 a_17842_n1579# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X317 VSS.t136 B[2].t5 a_15444_2390# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X318 VDD.t412 B[6].t7 a_10645_n2623# w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X319 a_10659_n973# A[6].t1 VDD.t433 w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X320 a_15044_n3209# A[5].t8 VDD.t351 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X321 a_2824_1705# a_3236_1679# a_2942_1705.t5 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X322 VDD.t336 carry_in.t6 a_4722_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X323 a_9337_1702# A[1].t5 VDD.t374 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X324 VDD.t187 A[7].t6 a_4092_n4223# w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X325 VDD.t238 a_8140_4225# a_9875_4534# w_9721_4472# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X326 a_16409_4529# a_14674_4220# VDD.t395 w_16255_4467# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X327 a_24346_n4830# a_19657_n3503.t9 VSS.t102 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X328 a_1051_3015# carry_in.t7 VDD.t337 w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X329 VSS.t148 A[3].t6 a_22783_969# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X330 VSS.t132 a_17184_n4222# a_15576_n1096# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X331 VSS.t126 a_1952_n3210# a_2610_n4635# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X332 a_8154_2575# a_7564_3012# VDD.t149 w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X333 a_11647_1676# a_4650_3958.t12 VDD.t223 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X334 a_14041_n3235# a_15044_n3209# a_15584_n3902.t2 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X335 VSS.t141 A[6].t2 a_8510_n3214# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X336 VDD.t467 A[7].t7 a_2492_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X337 VDD.t345 a_17697_3950.t9 a_20651_1407# w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X338 VDD.t142 a_11163_3955.t9 a_17769_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X339 a_10645_n2623# B[6].t8 VDD.t413 w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X340 VDD.t23 B[0].t8 a_1051_3015# w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X341 a_17769_1697# a_17342_2390# Y[2].t2 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X342 a_2130_n1097# a_4101_n969# VDD.t135 w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X343 VDD.t411 B[2].t6 a_15871_1697.t4 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X344 a_20651_1407# a_17697_3950.t10 VDD.t346 w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X345 a_24341_n3226# B[4].t8 VSS.t92 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X346 VSS.t48 a_23697_n4219# a_22089_n1093# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X347 a_3362_4537# a_1636_974# a_3244_4537# w_3208_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X348 Y[2].t1 a_17342_2390# a_17769_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X349 VDD.t288 B[7].t4 a_4101_n969# w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X350 a_2846_n4635# A[7].t8 VSS.t147 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X351 VDD.t260 a_23991_4537# a_19657_n3503.t2 w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X352 VDD.t311 B[4].t9 a_22097_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X353 a_15584_n3902.t1 a_15044_n3209# a_14041_n3235# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X354 Y[1].t2 a_10808_2395# a_11235_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X355 VSS.t36 B[3].t3 a_20893_2374# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X356 Y[3].t6 a_23900_2394# a_24327_1701.t7 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X357 VDD.t356 a_2130_n1097# a_2190_n1071# w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X358 VDD.t388 A[4].t6 a_23706_n965# w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X359 VDD.t180 a_1627_4228# a_3362_4537# w_3208_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X360 VDD.t300 a_6610_n3511.t9 a_10645_n2623# w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X361 a_3236_1679# A[0].t8 VDD.t339 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X362 a_14674_4220# a_14084_4657# VDD.t115 w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X363 VDD.t69 B[7].t5 a_2904_n3929# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X364 a_9455_970# a_9749_1676# VSS.t121 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X365 a_20656_3011# a_17697_3950.t11 VDD.t471 w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X366 a_3236_1679# A[0].t9 VSS.t72 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X367 VDD.t417 a_19657_n3503.t10 a_20199_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X368 VDD.t301 a_6610_n3511.t10 a_6612_n3214# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X369 VDD.t83 a_22849_4533# a_23113_3950# w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X370 VDD.t43 a_4650_3958.t13 a_11235_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X371 VSS.t76 B[1].t7 a_7801_2375# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X372 a_2190_n1071# a_2130_n1097# VDD.t355 w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X373 VDD.t46 B[0].t9 a_2397_2398# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X374 a_14330_766# A[2].t7 a_14093_1403# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X375 a_10645_n2623# a_6610_n3511.t11 VDD.t130 w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X376 a_7550_4662# A[1].t6 VDD.t375 w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X377 VDD.t143 a_11163_3955.t10 a_14093_1403# w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X378 a_22429_1701.t7 A[3].t7 VDD.t455 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X379 a_14683_966# a_14093_1403# VSS.t47 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X380 a_14688_2570# a_14098_3007# VDD.t382 w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X381 VDD.t366 a_988_n1093# a_1048_n1067# w_819_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X382 a_16225_965# B[2].t7 a_15989_1697# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X383 a_2904_n3929# B[7].t6 VSS.t14 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X384 a_4087_n2619# a_52_n3507.t8 VDD.t63 w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X385 a_2904_n3929# B[7].t7 VDD.t352 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X386 a_9337_1702# a_8910_2395# a_9455_1702.t0 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X387 a_20199_n3899# a_19657_n3503.t11 VDD.t418 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X388 a_17179_n2618# a_13144_n3506.t7 VDD.t199 w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X389 a_1283_774# A[0].t10 a_1046_1411# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X390 a_20554_n3232.t7 B[4].t10 a_22451_n4631# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X391 VSS.t66 a_8140_4225# a_9757_4534# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X392 a_2824_1705# B[0].t10 VDD.t47 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X393 a_7564_3012# a_4650_3958.t14 VDD.t44 w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X394 a_3178_973# B[0].t11 a_2942_1705.t7 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X395 a_2055_n1727# a_2484_n1097# a_2190_n1071# w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X396 a_7152_n3907# a_7564_n3933# Y[6].t4 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X397 a_594_n3903# a_52_n3507.t9 VDD.t100 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X398 a_1048_n1067# a_988_n1093# VDD.t365 w_819_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X399 a_9050_n3907# A[6].t3 VDD.t312 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X400 a_8140_4225# a_7550_4662# VSS.t64 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X401 VDD.t88 B[0].t12 a_2824_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X402 VSS.t29 B[2].t8 a_14335_2370# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X403 VDD.t237 a_8140_4225# a_9875_4534# w_9721_4472# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X404 a_4092_n4223# A[7].t9 VDD.t468 w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X405 VDD.t267 A[0].t11 a_1046_1411# w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X406 VDD.t461 a_20554_n3232.t11 a_20199_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X407 VDD.t167 a_7507_n3240.t10 a_7152_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X408 VDD.t85 a_13144_n3506.t8 a_17179_n2618# w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X409 a_21246_2574# a_20656_3011# VSS.t122 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X410 a_22215_n4631# a_22509_n3925# a_20554_n3232.t3 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X411 a_7787_4025# A[1].t7 a_7550_4662# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X412 a_9875_4534# a_8149_971# a_9757_4534# w_9721_4472# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X413 a_21241_970# a_20651_1407# VDD.t123 w_20497_1345# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X414 a_913_n1723# a_1342_n1093# a_1048_n1067# w_819_n1712# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X415 a_20611_n3925# a_20554_n3232.t12 VSS.t52 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X416 VDD.t331 a_17179_n2618# a_14434_n1092# w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X417 VSS.t61 a_22547_1701# a_23900_2394# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X418 Y[2].t5 a_18181_1671# a_17769_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X419 VSS.t94 B[1].t8 a_8910_2395# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X420 a_15222_n1096# a_17193_n968# VDD.t406 w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X421 a_20199_n3899# a_20554_n3232.t13 VDD.t75 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X422 a_7152_n3907# a_7507_n3240.t11 VDD.t118 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X423 Y[3].t1 a_24739_1675# a_24327_1701.t1 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X424 VDD.t259 a_23991_4537# a_19657_n3503.t1 w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X425 VDD.t231 A[5].t9 a_17184_n4222# w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X426 VDD.t313 A[6].t4 a_10650_n4227# w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X427 VDD.t497 a_10899_4538# a_11163_3955.t3 w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X428 VDD.t419 a_19657_n3503.t12 a_23697_n4219# w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X429 a_2484_n1097# a_4092_n4223# VDD.t333 w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X430 VDD.t295 A[2].t8 a_14084_4657# w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X431 a_19657_n3503.t0 a_23991_4537# VSS.t75 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X432 a_24327_1701.t4 a_22547_1701# VDD.t216 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X433 a_4101_n969# A[7].t10 a_4750_n1580# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X434 a_13686_n3902# a_13144_n3506.t9 VDD.t320 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X435 a_15871_1697.t7 a_16283_1671# a_15989_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X436 a_14321_4020# A[2].t9 a_14084_4657# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X437 VDD.t20 a_16291_4529# a_16555_3946# w_16255_4467# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X438 a_22849_4533# a_21241_970# VSS.t65 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X439 a_1048_n1067# a_1342_n1093# a_913_n1723# w_819_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X440 a_1952_n3210# A[7].t11 VDD.t106 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X441 a_14434_n1092# a_17179_n2618# VDD.t330 w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X442 VDD.t51 A[5].t10 a_15584_n3902.t4 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X443 a_8149_971# a_7559_1408# VDD.t174 w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X444 a_1006_n3929# a_949_n3236.t10 VDD.t285 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X445 VDD.t178 B[3].t4 a_20642_4661# w_20488_4599# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X446 a_22429_1701.t11 a_22841_1675# a_22547_1701# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X447 VDD.t263 a_20554_n3232.t14 a_20199_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X448 VDD.t119 a_7507_n3240.t12 a_7152_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X449 a_20656_3011# a_17697_3950.t12 VDD.t472 w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X450 a_10650_n4227# A[6].t5 VDD.t55 w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X451 a_4722_1705# a_4295_2398# Y[0].t1 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X452 a_23697_n4219# a_19657_n3503.t13 VDD.t420 w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X453 VSS.t112 a_8510_n3214# a_9168_n4639# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X454 a_8688_n1101# a_10659_n973# VDD.t372 w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X455 a_23991_4537# a_21246_2574# a_24109_4537# w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X456 VDD.t274 a_9757_4534# a_10021_3951# w_9721_4472# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X457 a_15938_n4634# A[5].t11 VSS.t49 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X458 VDD.t107 A[7].t12 a_1952_n3210# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X459 VDD.t144 a_11163_3955.t11 a_14093_1403# w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X460 a_15584_n3902.t3 A[5].t12 VDD.t304 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X461 a_9337_1702# a_9749_1676# a_9455_1702.t6 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X462 VDD.t286 a_949_n3236.t11 a_1006_n3929# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X463 VSS.t149 a_9455_1702.t12 a_10808_2395# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X464 a_4722_1705# carry_in.t8 VDD.t321 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X465 a_2942_1705.t1 a_2397_2398# a_2824_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X466 VDD.t397 a_7471_n1727# a_52_n3507.t2 w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X467 VDD.t56 A[6].t6 a_10650_n4227# w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X468 VDD.t218 a_22547_1701# a_23900_2394# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X469 a_9404_n4639# A[6].t7 VSS.t108 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X470 a_2492_n3903# a_1952_n3210# a_949_n3236.t6 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X471 a_14041_n3235# B[5].t6 a_15938_n4634# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X472 VDD.t410 a_21232_4224# a_22967_4533# w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X473 VDD.t453 a_17433_4533# a_17697_3950.t2 w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X474 a_23900_2394# a_22547_1701# VDD.t217 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X475 a_22783_969# B[3].t5 a_22547_1701# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X476 a_22097_n3899# a_22509_n3925# a_20554_n3232.t6 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X477 VDD.t327 a_21660_n1723# a_20593_n1089# w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X478 Y[4].t0 a_20554_n3232.t15 a_20553_n4631# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X479 VDD.t421 a_19657_n3503.t14 a_23692_n2615# w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X480 a_15996_n3928# B[5].t7 VSS.t69 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X481 VDD.t277 a_23706_n965# a_21735_n1093# w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X482 a_1636_974# a_1046_1411# VDD.t80 w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X483 a_7507_n3240.t4 B[6].t9 a_9404_n4639# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X484 a_949_n3236.t5 a_1952_n3210# a_2492_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X485 a_15996_n3928# B[5].t8 VDD.t243 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X486 VSS.t83 a_54_n3210# a_712_n4635# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X487 VDD.t192 B[3].t6 a_22002_2394# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X488 a_21241_970# a_20651_1407# VDD.t122 w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X489 a_17193_n968# B[5].t9 VDD.t244 w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X490 VSS.t24 a_52_n3507.t10 a_54_n3210# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X491 a_20554_n3232.t5 a_22509_n3925# a_22097_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X492 a_20593_n1089# a_21660_n1723# VDD.t326 w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X493 a_7546_n1097# a_8613_n1731# VDD.t368 w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X494 a_11299_n4838# a_6610_n3511.t12 VSS.t31 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X495 a_24355_n1576# B[4].t11 VSS.t93 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X496 a_4840_973# a_5134_1679# VSS.t81 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X497 VSS.t5 a_10021_3951# a_10899_4538# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X498 a_1051_3015# carry_in.t9 VDD.t322 w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X499 a_24327_1701.t3 a_22547_1701# VDD.t221 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X500 a_14140_n1066# a_14080_n1092# VDD.t73 w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X501 VDD.t126 B[2].t9 a_14084_4657# w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X502 a_2942_1705.t3 a_2397_2398# a_2942_973# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X503 VSS.t53 a_2055_n1727# a_988_n1093# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X504 Y[1].t6 a_11647_1676# a_11235_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X505 a_9168_n4639# a_9462_n3933# a_7507_n3240.t3 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X506 VDD.t499 a_10899_4538# a_11163_3955.t2 w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X507 a_11235_1702# a_9455_1702.t13 VDD.t97 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X508 VSS.t11 a_4650_3958.t15 a_7796_771# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X509 a_8613_n1731# a_9042_n1101# a_8748_n1075# w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X510 VSS.t119 A[1].t8 a_9691_970# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X511 a_10650_n4227# A[6].t8 a_11299_n4838# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X512 a_22097_n3899# a_22509_n3925# a_20554_n3232.t4 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X513 a_16555_3946# a_16291_4529# VSS.t3 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X514 VDD.t193 B[3].t7 a_22429_1701.t1 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X515 VSS.t137 a_10650_n4227# a_9042_n1101# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X516 a_11294_n3234# B[6].t10 VSS.t34 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X517 VSS.t82 a_23706_n965# a_21735_n1093# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X518 VDD.t349 a_11163_3955.t12 a_14098_3007# w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X519 VDD.t483 a_15989_1697# a_17342_2390# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X520 a_17887_965# a_18181_1671# VSS.t123 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X521 a_14005_n1722# a_14434_n1092# a_14140_n1066# w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X522 a_11017_4538# a_8154_2575# a_10899_4538# w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X523 a_22841_1675# A[3].t8 VSS.t143 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X524 a_2055_n1727# a_2130_n1097# VSS.t111 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X525 a_4386_4541# a_1641_2578# a_4504_4541# w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X526 a_7550_4662# A[1].t9 VDD.t250 w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X527 VDD.t194 B[3].t8 a_20656_3011# w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X528 a_15989_1697# a_15444_2390# a_15989_965# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X529 VSS.t85 a_13146_n3209# a_13804_n4634# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X530 a_1288_2378# carry_in.t10 a_1051_3015# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X531 VDD.t156 a_14093_1403# a_14683_966# w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X532 VSS.t133 a_913_n1723# carry_out.t0 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X533 a_9462_n3933# B[6].t11 VDD.t226 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X534 VDD.t95 a_23113_3950# a_24109_4537# w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X535 a_8748_n1075# a_9042_n1101# a_8613_n1731# w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X536 VDD.t353 B[7].t8 a_2492_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X537 a_10899_4538# a_8154_2575# a_11017_4538# w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X538 VSS.t17 a_13144_n3506.t10 a_13146_n3209# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X539 VSS.t104 a_19657_n3503.t15 a_19659_n3206# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X540 VDD.t458 a_23692_n2615# a_20947_n1089# w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X541 VSS.t57 a_3508_3954# a_4386_4541# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X542 a_15576_n1096# a_17184_n4222# VDD.t400 w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X543 VDD.t228 a_7550_4662# a_8140_4225# w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X544 a_16291_4529# a_14683_966# a_16409_4529# w_16255_4467# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X545 Y[0].t5 a_5134_1679# a_4722_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X546 a_10645_n2623# a_6610_n3511.t13 a_11294_n3234# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X547 VDD.t227 B[6].t12 a_10659_n973# w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X548 a_14140_n1066# a_14434_n1092# a_14005_n1722# w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X549 a_7606_n1071# a_7546_n1097# VDD.t141 w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X550 a_14098_n3928# a_14041_n3235# VDD.t3 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X551 a_20653_n1063# a_20593_n1089# VDD.t7 w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X552 a_3244_4537# a_1636_974# VSS.t46 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X553 VDD.t409 a_21232_4224# a_22967_4533# w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X554 a_14040_n4634# a_13144_n3506.t11 VSS.t129 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X555 VDD.t98 a_9455_1702.t14 a_10808_2395# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X556 a_913_n1723# a_988_n1093# VSS.t113 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X557 VDD.t0 A[0].t12 a_2824_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X558 a_18181_1671# a_11163_3955.t13 VSS.t107 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X559 a_15871_1697.t3 B[2].t10 VDD.t127 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X560 a_17769_1697# a_15989_1697# VDD.t486 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X561 VDD.t399 a_17184_n4222# a_15576_n1096# w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X562 VDD.t428 a_10650_n4227# a_9042_n1101# w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X563 a_21795_n1067# a_21735_n1093# VDD.t242 w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X564 a_14674_4220# a_14084_4657# VSS.t27 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X565 VDD.t272 A[5].t13 a_15044_n3209# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X566 a_14005_n1722# a_14434_n1092# a_14140_n1066# w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X567 VDD.t140 a_7546_n1097# a_7606_n1071# w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X568 VDD.t2 a_14041_n3235# a_14098_n3928# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X569 VSS.t13 a_10645_n2623# a_7900_n1097# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X570 VDD.t479 B[3].t9 a_22002_2394# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X571 a_17551_4533# a_14688_2570# a_17433_4533# w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X572 a_1636_974# a_1046_1411# VDD.t79 w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X573 a_20199_n3899# a_20611_n3925# Y[4].t6 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X574 a_7507_n3240.t7 a_8510_n3214# a_9050_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X575 a_15147_n1726# a_15576_n1096# a_15282_n1070# w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X576 VDD.t293 a_8688_n1101# a_8748_n1075# w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X577 a_2492_n3903# A[7].t13 VDD.t464 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X578 VDD.t283 carry_in.t11 a_5134_1679# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X579 VDD.t241 a_21735_n1093# a_21795_n1067# w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X580 VDD.t101 a_52_n3507.t11 a_54_n3210# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X581 VDD.t39 a_2942_1705.t11 a_4295_2398# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X582 VDD.t269 a_4650_3958.t16 a_7559_1408# w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X583 a_7606_n1071# a_7546_n1097# VDD.t139 w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X584 a_14098_n3928# a_14041_n3235# VDD.t1 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X585 a_24327_1701.t10 a_17697_3950.t13 VDD.t446 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X586 VDD.t66 B[2].t11 a_14084_4657# w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X587 a_11235_1702# a_9455_1702.t15 VDD.t99 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X588 a_2610_n4635# a_2904_n3929# a_949_n3236.t3 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X589 VDD.t254 B[1].t9 a_8910_2395# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X590 a_23692_n2615# a_19657_n3503.t16 a_24341_n3226# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X591 a_9050_n3907# a_8510_n3214# a_7507_n3240.t6 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X592 VDD.t265 A[3].t9 a_22429_1701.t6 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X593 VSS.t144 a_23692_n2615# a_20947_n1089# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X594 VDD.t447 a_17697_3950.t14 a_24327_1701.t9 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X595 VDD.t482 a_15989_1697# a_17342_2390# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X596 a_8748_n1075# a_8688_n1101# VDD.t292 w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X597 a_14041_n3235# a_15044_n3209# a_15584_n3902.t0 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X598 VDD.t70 B[7].t9 a_2492_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X599 a_21795_n1067# a_21735_n1093# VDD.t240 w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X600 a_14093_1403# A[2].t10 VDD.t108 w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X601 a_54_n3210# a_52_n3507.t12 VDD.t13 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X602 VDD.t205 a_3508_3954# a_4504_4541# w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X603 VDD.t102 A[6].t9 a_8510_n3214# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X604 VDD.t94 a_23113_3950# a_24109_4537# w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X605 VDD.t29 a_2942_1705.t12 a_4722_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X606 VDD.t377 a_20656_3011# a_21246_2574# w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X607 a_15444_2390# B[2].t12 VDD.t67 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X608 a_7507_n3240.t5 a_8510_n3214# a_9050_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X609 Y[7].t2 a_54_n3210# a_594_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X610 VSS.t58 a_15147_n1726# a_14080_n1092# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X611 VDD.t103 A[6].t10 a_10659_n973# w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X612 VDD.t25 a_10021_3951# a_11017_4538# w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X613 a_15584_n3902.t11 a_15996_n3928# a_14041_n3235# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X614 a_2492_n3903# B[7].t10 VDD.t71 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X615 a_2942_1705.t0 a_2397_2398# a_2824_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X616 a_1627_4228# a_1037_4665# VDD.t489 w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X617 a_4722_1705# a_2942_1705.t13 VDD.t30 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X618 VDD.t251 A[1].t10 a_9337_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X619 VDD.t376 a_13144_n3506.t12 a_13146_n3209# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X620 VDD.t77 a_6610_n3511.t14 a_10645_n2623# w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X621 VDD.t394 a_14674_4220# a_16409_4529# w_16255_4467# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X622 a_15584_n3902.t8 B[5].t10 VDD.t152 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X623 a_1627_4228# a_1037_4665# VSS.t152 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X624 a_3508_3954# a_3244_4537# VSS.t12 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X625 a_24445_969# a_24739_1675# VSS.t41 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X626 a_22097_n3899# A[4].t7 VDD.t183 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X627 a_8510_n3214# A[6].t11 VDD.t298 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X628 VDD.t284 carry_in.t12 a_1051_3015# w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X629 VDD.t270 a_4650_3958.t17 a_11647_1676# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X630 a_7564_n3933# a_7507_n3240.t13 VDD.t120 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X631 a_2824_1705# a_3236_1679# a_2942_1705.t4 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X632 VSS.t146 a_17697_3950.t15 a_20888_770# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X633 a_20651_1407# A[3].t10 VDD.t266 w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X634 a_22547_1701# a_22002_2394# a_22547_969# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X635 a_9050_n3907# a_9462_n3933# a_7507_n3240.t1 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X636 VSS.t115 a_8613_n1731# a_7546_n1097# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X637 a_17769_1697# a_11163_3955.t14 VDD.t350 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X638 a_9691_970# B[1].t10 a_9455_1702.t4 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X639 a_22841_1675# A[3].t11 VDD.t491 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X640 a_594_n3903# a_54_n3210# Y[7].t1 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X641 a_15147_n1726# a_15222_n1096# VSS.t91 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X642 a_1051_3015# B[0].t13 VDD.t89 w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X643 a_9749_1676# A[1].t11 VDD.t252 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X644 Y[2].t0 a_17342_2390# a_17769_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X645 a_1342_n1093# a_4087_n2619# VDD.t495 w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X646 VSS.t145 a_11163_3955.t15 a_18123_965# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X647 a_13146_n3209# a_13144_n3506.t13 VDD.t208 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X648 VSS.t128 a_14005_n1722# a_6610_n3511.t0 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X649 VDD.t153 B[5].t11 a_15584_n3902.t7 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X650 VDD.t299 A[6].t12 a_9050_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X651 VDD.t109 A[2].t11 a_15871_1697.t10 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X652 a_4101_n969# B[7].t11 VDD.t302 w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X653 a_23697_n4219# A[4].t8 a_24346_n4830# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X654 a_8613_n1731# a_8688_n1101# VSS.t89 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X655 a_7507_n3240.t0 a_9462_n3933# a_9050_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X656 a_20893_2374# a_17697_3950.t16 a_20656_3011# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X657 a_24327_1701.t6 a_23900_2394# Y[3].t7 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X658 VSS.t60 a_6610_n3511.t15 a_6612_n3214# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X659 Y[5].t7 a_13146_n3209# a_13686_n3902# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X660 a_3362_4537# a_1627_4228# VDD.t179 w_3208_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X661 VSS.t86 carry_in.t13 a_5076_973# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X662 VDD.t494 a_4087_n2619# a_1342_n1093# w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X663 VDD.t492 A[3].t12 a_20642_4661# w_20488_4599# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X664 VDD.t31 a_2942_1705.t14 a_4295_2398# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X665 a_22547_1701# a_22002_2394# a_22429_1701.t4 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X666 VDD.t503 a_13144_n3506.t14 a_13146_n3209# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X667 a_14005_n1722# a_14080_n1092# VSS.t15 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X668 VDD.t462 A[5].t14 a_17193_n968# w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X669 a_8154_2575# a_7564_3012# VSS.t45 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X670 VDD.t184 A[4].t9 a_23706_n965# w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X671 a_9050_n3907# A[6].t13 VDD.t316 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X672 a_7796_771# A[1].t12 a_7559_1408# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X673 Y[6].t0 a_6612_n3214# a_7152_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X674 a_23113_3950# a_22849_4533# VDD.t82 w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X675 a_11235_1702# a_4650_3958.t18 VDD.t271 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X676 a_2397_2398# B[0].t14 VDD.t90 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X677 a_13686_n3902# a_13146_n3209# Y[5].t6 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X678 a_949_n3236.t4 B[7].t12 a_2846_n4635# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X679 VDD.t434 A[1].t13 a_7550_4662# w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X680 a_14093_1403# A[2].t12 VDD.t110 w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X681 a_4087_n2619# B[7].t13 VDD.t264 w_3993_n2655# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X682 VDD.t68 B[2].t13 a_14098_3007# w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X683 a_11308_n1584# B[6].t13 VSS.t32 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X684 VDD.t332 a_4092_n4223# a_2484_n1097# w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X685 VSS.t78 a_14434_n1092# a_14005_n1722# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X686 a_16283_1671# A[2].t13 VDD.t35 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X687 a_9462_n3933# B[6].t14 VSS.t33 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X688 a_913_n1723# a_1342_n1093# a_1048_n1067# w_819_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X689 a_7550_4662# B[1].t11 VDD.t93 w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X690 a_14688_2570# a_14098_3007# VDD.t381 w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X691 VDD.t24 a_10021_3951# a_11017_4538# w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X692 a_9757_4534# a_8149_971# VSS.t16 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X693 Y[5].t5 a_13146_n3209# a_13686_n3902# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X694 VDD.t389 B[1].t12 a_7550_4662# w_7396_4600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X695 Y[5].t0 a_14041_n3235# a_14040_n4634# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X696 VDD.t317 A[6].t14 a_10659_n973# w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X697 VDD.t393 a_14674_4220# a_16409_4529# w_16255_4467# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X698 VDD.t4 a_14041_n3235# a_13686_n3902# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X699 a_10659_n973# A[6].t15 a_11308_n1584# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X700 a_14335_2370# a_11163_3955.t16 a_14098_3007# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X701 a_15702_n4634# a_15996_n3928# a_14041_n3235# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X702 a_4092_n4223# a_52_n3507.t13 VDD.t14 w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X703 VSS.t116 a_10659_n973# a_8688_n1101# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X704 VDD.t215 a_6610_n3511.t16 a_6612_n3214# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X705 a_1627_4228# a_1037_4665# VDD.t488 w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X706 a_7564_3012# a_4650_3958.t19 VDD.t296 w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X707 a_1006_n3929# a_949_n3236.t12 VSS.t87 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X708 VDD.t154 B[5].t12 a_15584_n3902.t6 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X709 a_1006_n3929# a_949_n3236.t13 VDD.t168 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X710 a_1641_2578# a_1051_3015# VDD.t501 w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X711 VDD.t91 A[0].t13 a_2824_1705# w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X712 VDD.t59 a_10645_n2623# a_7900_n1097# w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X713 VDD.t257 carry_in.t14 a_1046_1411# w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X714 a_9749_1676# A[1].t14 VDD.t435 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X715 VDD.t15 a_52_n3507.t14 a_4092_n4223# w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X716 a_2190_n1071# a_2484_n1097# a_2055_n1727# w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X717 a_7152_n3907# a_6610_n3511.t17 VDD.t474 w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X718 VSS.t131 a_7471_n1727# a_52_n3507.t0 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X719 VDD.t36 A[2].t14 a_15871_1697.t9 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X720 VSS.t39 a_21557_n3206# a_22215_n4631# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X721 VDD.t132 a_52_n3507.t15 a_594_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X722 a_23991_4537# a_21246_2574# VSS.t120 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X723 a_17551_4533# a_14688_2570# a_17433_4533# w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X724 a_24327_1701.t0 a_24739_1675# Y[3].t0 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X725 a_20317_n4631# a_20611_n3925# Y[4].t7 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X726 a_14084_4657# A[2].t15 VDD.t37 w_13930_4595# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X727 VDD.t480 B[3].t10 a_20642_4661# w_20488_4599# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X728 VSS.t23 a_23113_3950# a_23991_4537# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X729 a_23692_n2615# a_19657_n3503.t17 VDD.t422 w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X730 a_7900_n1097# a_10645_n2623# VDD.t58 w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X731 a_11235_1702# a_10808_2395# Y[1].t1 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X732 a_15989_1697# a_15444_2390# a_15871_1697.t0 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X733 a_949_n3236.t2 a_2904_n3929# a_2492_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X734 a_4092_n4223# a_52_n3507.t16 VDD.t133 w_3998_n4259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X735 a_20642_4661# B[3].t11 VDD.t481 w_20488_4599# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X736 a_2055_n1727# a_2484_n1097# a_2190_n1071# w_1961_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X737 a_948_n4635# a_52_n3507.t17 VSS.t35 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X738 VDD.t475 a_6610_n3511.t18 a_7152_n3907# w_6576_n3276# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X739 a_22547_1701# a_22002_2394# a_22429_1701.t3 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X740 a_22451_n4631# A[4].t10 VSS.t10 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X741 a_594_n3903# a_52_n3507.t18 VDD.t437 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X742 a_21660_n1723# a_22089_n1093# a_21795_n1067# w_21566_n1712# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X743 VDD.t448 a_17697_3950.t17 a_20656_3011# w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X744 a_3236_1679# A[0].t14 VDD.t45 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X745 a_8149_971# a_7559_1408# VDD.t173 w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X746 VDD.t371 a_10659_n973# a_8688_n1101# w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X747 a_10021_3951# a_9757_4534# VDD.t273 w_9721_4472# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X748 a_24109_4537# a_21246_2574# a_23991_4537# w_23955_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X749 VDD.t423 a_19657_n3503.t18 a_23692_n2615# w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X750 VDD.t57 a_10645_n2623# a_7900_n1097# w_10551_n2659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X751 a_2492_n3903# a_2904_n3929# a_949_n3236.t1 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X752 a_11353_970# a_11647_1676# VSS.t106 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X753 a_13144_n3506.t3 a_20518_n1719# VDD.t290 w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X754 a_14093_1403# a_11163_3955.t17 VDD.t460 w_13939_1341# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X755 VDD.t439 B[4].t12 a_22509_n3925# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X756 VDD.t380 a_13144_n3506.t15 a_13686_n3902# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X757 a_4650_3958.t1 a_4386_4541# VDD.t245 w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X758 VDD.t329 a_17179_n2618# a_14434_n1092# w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X759 VDD.t348 A[0].t15 a_1037_4665# w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X760 VSS.t38 B[3].t12 a_20879_4024# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X761 a_9337_1702# a_9749_1676# a_9455_1702.t5 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X762 VSS.t20 a_6612_n3214# a_7270_n4639# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X763 a_22967_4533# a_21241_970# a_22849_4533# w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X764 a_17697_3950.t1 a_17433_4533# VDD.t452 w_17397_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X765 a_7564_3012# B[1].t13 VDD.t344 w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X766 VDD.t114 B[1].t14 a_9337_1702# w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X767 VDD.t449 a_17697_3950.t18 a_24739_1675# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X768 VDD.t291 a_20518_n1719# a_13144_n3506.t2 w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X769 VDD.t53 a_3244_4537# a_3508_3954# w_3208_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X770 a_17433_4533# a_14688_2570# VSS.t56 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X771 VSS.t109 a_17697_3950.t19 a_24681_969# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X772 a_22509_n3925# B[4].t13 VDD.t440 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X773 VDD.t41 A[4].t11 a_23697_n4219# w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X774 a_13686_n3902# a_13144_n3506.t16 VDD.t279 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X775 a_20888_770# A[3].t13 a_20651_1407# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X776 a_8613_n1731# a_9042_n1101# a_8748_n1075# w_8519_n1720# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X777 a_17179_n2618# B[5].t13 VDD.t359 w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X778 VDD.t104 B[1].t15 a_7564_3012# w_7410_2950# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X779 a_20651_1407# A[3].t14 VDD.t148 w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X780 a_4750_n1580# B[7].t14 VSS.t77 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X781 a_9455_1702.t3 a_8910_2395# a_9455_970# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X782 VDD.t258 carry_in.t15 a_1046_1411# w_892_1349# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X783 a_22841_1675# A[3].t15 VDD.t456 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X784 a_1641_2578# a_1051_3015# VDD.t500 w_897_2953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X785 a_18123_965# a_15989_1697# Y[2].t7 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X786 a_20554_n3232.t2 a_21557_n3206# a_22097_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X787 a_7506_n4639# a_6610_n3511.t19 VSS.t71 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X788 VDD.t121 a_20651_1407# a_21241_970# w_20497_1345# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X789 a_13144_n3506.t1 a_20518_n1719# VDD.t289 w_20424_n1708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X790 VDD.t405 a_17193_n968# a_15222_n1096# w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X791 a_52_n3507.t1 a_7471_n1727# VDD.t396 w_7377_n1716# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X792 a_23697_n4219# A[4].t12 VDD.t42 w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X793 VDD.t276 a_23706_n965# a_21735_n1093# w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X794 a_17769_1697# a_18181_1671# Y[2].t4 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X795 VSS.t125 a_1342_n1093# a_913_n1723# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X796 a_4101_n969# A[7].t14 VDD.t465 w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X797 VDD.t360 B[5].t14 a_17179_n2618# w_17085_n2654# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X798 a_7559_1408# A[1].t15 VDD.t436 w_7405_1346# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X799 a_10899_4538# a_8154_2575# VSS.t67 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X800 a_17184_n4222# a_13144_n3506.t17 VDD.t76 w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X801 a_23706_n965# B[4].t14 VDD.t441 w_23612_n1001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X802 a_17193_n968# B[5].t15 VDD.t361 w_17099_n1004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X803 a_5076_973# a_2942_1705.t15 Y[0].t7 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X804 VSS.t37 B[3].t13 a_22002_2394# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X805 a_9042_n1101# a_10650_n4227# VDD.t427 w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X806 VSS.t127 B[2].t14 a_14321_4020# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X807 a_11235_1702# a_11647_1676# Y[1].t5 w_8873_2333# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X808 VDD.t466 A[7].t15 a_4101_n969# w_4007_n1005# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X809 a_14098_n3928# a_14041_n3235# VSS.t0 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X810 a_11163_3955.t1 a_10899_4538# VDD.t498 w_10863_4476# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X811 a_22097_n3899# a_21557_n3206# a_20554_n3232.t1 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X812 Y[6].t3 a_7507_n3240.t14 a_7506_n4639# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X813 a_22547_1701# a_22841_1675# a_22429_1701.t10 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X814 a_15989_1697# a_16283_1671# a_15871_1697.t6 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X815 VDD.t493 A[4].t13 a_23697_n4219# w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X816 a_2492_n3903# a_2904_n3929# a_949_n3236.t0 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X817 VSS.t130 a_14674_4220# a_16291_4529# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X818 a_18181_1671# a_11163_3955.t18 VDD.t48 w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X819 a_14098_3007# a_11163_3955.t19 VDD.t49 w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X820 a_22429_1701.t0 B[3].t14 VDD.t27 w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X821 Y[4].t5 a_20611_n3925# a_20199_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X822 a_22429_1701.t9 a_22841_1675# a_22547_1701# w_21965_2332# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X823 a_14688_2570# a_14098_3007# VSS.t124 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X824 VDD.t78 a_13144_n3506.t18 a_17184_n4222# w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X825 VDD.t19 a_16291_4529# a_16555_3946# w_16255_4467# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X826 a_7564_n3933# a_7507_n3240.t15 VSS.t54 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X827 VDD.t426 a_10650_n4227# a_9042_n1101# w_10556_n4263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X828 a_4504_4541# a_1641_2578# a_4386_4541# w_4350_4479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X829 VDD.t161 a_23697_n4219# a_22089_n1093# w_23603_n4255# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X830 VSS.t153 A[4].t14 a_21557_n3206# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X831 a_23706_n965# A[4].t15 a_24355_n1576# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X832 a_20656_3011# B[3].t15 VDD.t28 w_20502_2949# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X833 VDD.t385 B[2].t15 a_14098_3007# w_13944_2945# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X834 a_20554_n3232.t0 a_21557_n3206# a_22097_n3899# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X835 a_7270_n4639# a_7564_n3933# Y[6].t7 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X836 VSS.t151 a_15989_1697# a_17342_2390# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X837 a_4386_4541# a_1641_2578# VSS.t19 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X838 a_13686_n3902# a_14098_n3928# Y[5].t2 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X839 a_594_n3903# a_949_n3236.t14 VDD.t169 w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X840 a_14140_n1066# a_14080_n1092# VDD.t72 w_13911_n1711# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X841 a_16409_4529# a_14683_966# a_16291_4529# w_16255_4467# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X842 a_4722_1705# a_5134_1679# Y[0].t4 w_2360_2336# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X843 a_22509_n3925# B[4].t15 VDD.t335 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X844 a_20199_n3899# a_20611_n3925# Y[4].t4 w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X845 a_10659_n973# B[6].t15 VDD.t155 w_10565_n1009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X846 a_14041_n3235# a_15996_n3928# a_15584_n3902.t10 w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X847 a_17184_n4222# a_13144_n3506.t19 VDD.t105 w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X848 VDD.t60 B[0].t15 a_1037_4665# w_883_4603# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X849 VDD.t424 a_19657_n3503.t19 a_19659_n3206# w_19623_n3268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X850 VDD.t438 a_52_n3507.t19 a_54_n3210# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X851 VDD.t52 a_3244_4537# a_3508_3954# w_3208_4475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X852 a_22967_4533# a_21232_4224# VDD.t408 w_22813_4471# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X853 a_17697_3950.t0 a_17433_4533# VSS.t142 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X854 a_15282_n1070# a_15222_n1096# VDD.t306 w_15053_n1715# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X855 VSS.t26 a_2484_n1097# a_2055_n1727# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X856 a_9875_4534# a_8149_971# a_9757_4534# w_9721_4472# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X857 VDD.t170 a_949_n3236.t15 a_594_n3903# w_18_n3272# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X858 VDD.t485 a_15989_1697# a_17769_1697# w_15407_2328# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X859 a_4736_n3230# B[7].t15 VSS.t59 a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X860 VSS.t97 a_21660_n1723# a_20593_n1089# a_1596_n2079# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X861 a_15584_n3902.t9 a_15996_n3928# a_14041_n3235# w_13110_n3271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X862 a_20947_n1089# a_23692_n2615# VDD.t457 w_23598_n2651# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X863 VDD.t315 A[5].t15 a_17184_n4222# w_17090_n4258# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 VDD.n477 VDD.t250 30.163
R1 VDD.n183 VDD.t454 30.163
R2 VDD.n2 VDD.t37 30.163
R3 VDD.n61 VDD.t470 30.163
R4 VDD.n87 VDD.t471 30.163
R5 VDD.n79 VDD.t148 30.163
R6 VDD.n28 VDD.t49 30.163
R7 VDD.n20 VDD.t108 30.163
R8 VDD.n442 VDD.t322 30.163
R9 VDD.n187 VDD.t450 30.163
R10 VDD.n206 VDD.t466 30.163
R11 VDD.n263 VDD.t317 30.163
R12 VDD.n320 VDD.t462 30.163
R13 VDD.n377 VDD.t184 30.163
R14 VDD.n224 VDD.t77 30.163
R15 VDD.n234 VDD.t56 30.163
R16 VDD.n281 VDD.t85 30.163
R17 VDD.n291 VDD.t231 30.163
R18 VDD.n338 VDD.t423 30.163
R19 VDD.n348 VDD.t493 30.163
R20 VDD.n420 VDD.t62 30.163
R21 VDD.n430 VDD.t187 30.163
R22 VDD.n135 VDD.t44 30.163
R23 VDD.n127 VDD.t436 30.163
R24 VDD.n107 VDD.t219 28.664
R25 VDD.n112 VDD.t145 28.664
R26 VDD.n95 VDD.t479 28.664
R27 VDD.n100 VDD.t456 28.664
R28 VDD.n48 VDD.t482 28.664
R29 VDD.n53 VDD.t48 28.664
R30 VDD.n36 VDD.t212 28.664
R31 VDD.n41 VDD.t32 28.664
R32 VDD.n167 VDD.t31 28.664
R33 VDD.n172 VDD.t354 28.664
R34 VDD.n449 VDD.t46 28.664
R35 VDD.n454 VDD.t339 28.664
R36 VDD.n217 VDD.t50 28.664
R37 VDD.n212 VDD.t226 28.664
R38 VDD.n245 VDD.t301 28.664
R39 VDD.n240 VDD.t120 28.664
R40 VDD.n274 VDD.t272 28.664
R41 VDD.n269 VDD.t188 28.664
R42 VDD.n302 VDD.t503 28.664
R43 VDD.n297 VDD.t3 28.664
R44 VDD.n331 VDD.t11 28.664
R45 VDD.n326 VDD.t335 28.664
R46 VDD.n359 VDD.t414 28.664
R47 VDD.n354 VDD.t318 28.664
R48 VDD.n413 VDD.t107 28.664
R49 VDD.n408 VDD.t287 28.664
R50 VDD.n402 VDD.t438 28.664
R51 VDD.n397 VDD.t285 28.664
R52 VDD.n155 VDD.t65 28.664
R53 VDD.n160 VDD.t113 28.664
R54 VDD.n143 VDD.t254 28.664
R55 VDD.n148 VDD.t252 28.664
R56 VDD.n486 VDD.t274 28.57
R57 VDD.n492 VDD.t499 28.57
R58 VDD.n464 VDD.t52 28.57
R59 VDD.n470 VDD.t246 28.57
R60 VDD.n15 VDD.t453 28.57
R61 VDD.n10 VDD.t19 28.57
R62 VDD.n69 VDD.t83 28.57
R63 VDD.n74 VDD.t259 28.57
R64 VDD.n195 VDD.t402 28.57
R65 VDD.n201 VDD.t198 28.57
R66 VDD.n310 VDD.t390 28.57
R67 VDD.n315 VDD.t211 28.57
R68 VDD.n258 VDD.t370 28.57
R69 VDD.n253 VDD.t398 28.57
R70 VDD.n372 VDD.t328 28.57
R71 VDD.n367 VDD.t290 28.57
R72 VDD.n476 VDD.t375 28.565
R73 VDD.n476 VDD.t434 28.565
R74 VDD.n479 VDD.t229 28.565
R75 VDD.n479 VDD.t228 28.565
R76 VDD.n480 VDD.t230 28.565
R77 VDD.n480 VDD.t389 28.565
R78 VDD.n475 VDD.t93 28.565
R79 VDD.n475 VDD.t347 28.565
R80 VDD.n485 VDD.t273 28.565
R81 VDD.n485 VDD.t275 28.565
R82 VDD.n491 VDD.t498 28.565
R83 VDD.n491 VDD.t497 28.565
R84 VDD.n463 VDD.t54 28.565
R85 VDD.n463 VDD.t53 28.565
R86 VDD.n469 VDD.t245 28.565
R87 VDD.n469 VDD.t247 28.565
R88 VDD.n182 VDD.t305 28.565
R89 VDD.n182 VDD.t348 28.565
R90 VDD.n178 VDD.t488 28.565
R91 VDD.n178 VDD.t490 28.565
R92 VDD.n179 VDD.t489 28.565
R93 VDD.n179 VDD.t253 28.565
R94 VDD.n181 VDD.t22 28.565
R95 VDD.n181 VDD.t60 28.565
R96 VDD.n1 VDD.t147 28.565
R97 VDD.n1 VDD.t295 28.565
R98 VDD.n4 VDD.t115 28.565
R99 VDD.n4 VDD.t117 28.565
R100 VDD.n5 VDD.t116 28.565
R101 VDD.n5 VDD.t66 28.565
R102 VDD.n0 VDD.t213 28.565
R103 VDD.n0 VDD.t126 28.565
R104 VDD.n14 VDD.t452 28.565
R105 VDD.n14 VDD.t451 28.565
R106 VDD.n9 VDD.t21 28.565
R107 VDD.n9 VDD.t20 28.565
R108 VDD.n60 VDD.t249 28.565
R109 VDD.n60 VDD.t492 28.565
R110 VDD.n63 VDD.t325 28.565
R111 VDD.n63 VDD.t323 28.565
R112 VDD.n64 VDD.t324 28.565
R113 VDD.n64 VDD.t178 28.565
R114 VDD.n59 VDD.t481 28.565
R115 VDD.n59 VDD.t480 28.565
R116 VDD.n68 VDD.t82 28.565
R117 VDD.n68 VDD.t84 28.565
R118 VDD.n73 VDD.t261 28.565
R119 VDD.n73 VDD.t260 28.565
R120 VDD.n108 VDD.t217 28.565
R121 VDD.n108 VDD.t218 28.565
R122 VDD.n113 VDD.t445 28.565
R123 VDD.n113 VDD.t449 28.565
R124 VDD.n96 VDD.t425 28.565
R125 VDD.n96 VDD.t192 28.565
R126 VDD.n101 VDD.t491 28.565
R127 VDD.n101 VDD.t138 28.565
R128 VDD.n86 VDD.t472 28.565
R129 VDD.n86 VDD.t448 28.565
R130 VDD.n89 VDD.t378 28.565
R131 VDD.n89 VDD.t377 28.565
R132 VDD.n90 VDD.t379 28.565
R133 VDD.n90 VDD.t194 28.565
R134 VDD.n85 VDD.t28 28.565
R135 VDD.n85 VDD.t176 28.565
R136 VDD.n78 VDD.t266 28.565
R137 VDD.n78 VDD.t262 28.565
R138 VDD.n81 VDD.t122 28.565
R139 VDD.n81 VDD.t121 28.565
R140 VDD.n82 VDD.t123 28.565
R141 VDD.n82 VDD.t443 28.565
R142 VDD.n77 VDD.t346 28.565
R143 VDD.n77 VDD.t345 28.565
R144 VDD.n49 VDD.t484 28.565
R145 VDD.n49 VDD.t483 28.565
R146 VDD.n54 VDD.t16 28.565
R147 VDD.n54 VDD.t431 28.565
R148 VDD.n37 VDD.t67 28.565
R149 VDD.n37 VDD.t124 28.565
R150 VDD.n42 VDD.t35 28.565
R151 VDD.n42 VDD.t34 28.565
R152 VDD.n27 VDD.t430 28.565
R153 VDD.n27 VDD.t349 28.565
R154 VDD.n30 VDD.t381 28.565
R155 VDD.n30 VDD.t383 28.565
R156 VDD.n31 VDD.t382 28.565
R157 VDD.n31 VDD.t68 28.565
R158 VDD.n26 VDD.t214 28.565
R159 VDD.n26 VDD.t385 28.565
R160 VDD.n19 VDD.t110 28.565
R161 VDD.n19 VDD.t33 28.565
R162 VDD.n22 VDD.t157 28.565
R163 VDD.n22 VDD.t156 28.565
R164 VDD.n23 VDD.t158 28.565
R165 VDD.n23 VDD.t144 28.565
R166 VDD.n18 VDD.t460 28.565
R167 VDD.n18 VDD.t143 28.565
R168 VDD.n168 VDD.t38 28.565
R169 VDD.n168 VDD.t39 28.565
R170 VDD.n173 VDD.t362 28.565
R171 VDD.n173 VDD.t283 28.565
R172 VDD.n450 VDD.t90 28.565
R173 VDD.n450 VDD.t225 28.565
R174 VDD.n455 VDD.t45 28.565
R175 VDD.n455 VDD.t442 28.565
R176 VDD.n441 VDD.t337 28.565
R177 VDD.n441 VDD.t284 28.565
R178 VDD.n444 VDD.t500 28.565
R179 VDD.n444 VDD.t502 28.565
R180 VDD.n445 VDD.t501 28.565
R181 VDD.n445 VDD.t23 28.565
R182 VDD.n440 VDD.t89 28.565
R183 VDD.n440 VDD.t224 28.565
R184 VDD.n186 VDD.t201 28.565
R185 VDD.n186 VDD.t267 28.565
R186 VDD.n189 VDD.t79 28.565
R187 VDD.n189 VDD.t81 28.565
R188 VDD.n190 VDD.t80 28.565
R189 VDD.n190 VDD.t258 28.565
R190 VDD.n185 VDD.t364 28.565
R191 VDD.n185 VDD.t257 28.565
R192 VDD.n194 VDD.t404 28.565
R193 VDD.n194 VDD.t403 28.565
R194 VDD.n200 VDD.t196 28.565
R195 VDD.n200 VDD.t197 28.565
R196 VDD.n309 VDD.t391 28.565
R197 VDD.n309 VDD.t392 28.565
R198 VDD.n314 VDD.t209 28.565
R199 VDD.n314 VDD.t210 28.565
R200 VDD.n257 VDD.t368 28.565
R201 VDD.n257 VDD.t369 28.565
R202 VDD.n252 VDD.t396 28.565
R203 VDD.n252 VDD.t397 28.565
R204 VDD.n208 VDD.t135 28.565
R205 VDD.n208 VDD.t137 28.565
R206 VDD.n209 VDD.t302 28.565
R207 VDD.n209 VDD.t136 28.565
R208 VDD.n205 VDD.t465 28.565
R209 VDD.n205 VDD.t186 28.565
R210 VDD.n204 VDD.t160 28.565
R211 VDD.n204 VDD.t288 28.565
R212 VDD.n265 VDD.t372 28.565
R213 VDD.n265 VDD.t371 28.565
R214 VDD.n266 VDD.t155 28.565
R215 VDD.n266 VDD.t373 28.565
R216 VDD.n262 VDD.t433 28.565
R217 VDD.n262 VDD.t103 28.565
R218 VDD.n261 VDD.t314 28.565
R219 VDD.n261 VDD.t227 28.565
R220 VDD.n322 VDD.t406 28.565
R221 VDD.n322 VDD.t407 28.565
R222 VDD.n323 VDD.t244 28.565
R223 VDD.n323 VDD.t405 28.565
R224 VDD.n319 VDD.t268 28.565
R225 VDD.n319 VDD.t469 28.565
R226 VDD.n318 VDD.t361 28.565
R227 VDD.n318 VDD.t256 28.565
R228 VDD.n379 VDD.t278 28.565
R229 VDD.n379 VDD.t277 28.565
R230 VDD.n380 VDD.t441 28.565
R231 VDD.n380 VDD.t276 28.565
R232 VDD.n376 VDD.t386 28.565
R233 VDD.n376 VDD.t388 28.565
R234 VDD.n375 VDD.t342 28.565
R235 VDD.n375 VDD.t310 28.565
R236 VDD.n371 VDD.t326 28.565
R237 VDD.n371 VDD.t327 28.565
R238 VDD.n366 VDD.t289 28.565
R239 VDD.n366 VDD.t291 28.565
R240 VDD.n218 VDD.t298 28.565
R241 VDD.n218 VDD.t102 28.565
R242 VDD.n213 VDD.t319 28.565
R243 VDD.n213 VDD.t204 28.565
R244 VDD.n246 VDD.t92 28.565
R245 VDD.n246 VDD.t215 28.565
R246 VDD.n241 VDD.t166 28.565
R247 VDD.n241 VDD.t165 28.565
R248 VDD.n226 VDD.t58 28.565
R249 VDD.n226 VDD.t59 28.565
R250 VDD.n227 VDD.t191 28.565
R251 VDD.n227 VDD.t57 28.565
R252 VDD.n223 VDD.t130 28.565
R253 VDD.n223 VDD.t300 28.565
R254 VDD.n222 VDD.t413 28.565
R255 VDD.n222 VDD.t412 28.565
R256 VDD.n229 VDD.t427 28.565
R257 VDD.n229 VDD.t428 28.565
R258 VDD.n230 VDD.t341 28.565
R259 VDD.n230 VDD.t426 28.565
R260 VDD.n233 VDD.t55 28.565
R261 VDD.n233 VDD.t313 28.565
R262 VDD.n232 VDD.t203 28.565
R263 VDD.n232 VDD.t202 28.565
R264 VDD.n275 VDD.t351 28.565
R265 VDD.n275 VDD.t429 28.565
R266 VDD.n270 VDD.t243 28.565
R267 VDD.n270 VDD.t189 28.565
R268 VDD.n303 VDD.t208 28.565
R269 VDD.n303 VDD.t376 28.565
R270 VDD.n298 VDD.t1 28.565
R271 VDD.n298 VDD.t2 28.565
R272 VDD.n283 VDD.t330 28.565
R273 VDD.n283 VDD.t331 28.565
R274 VDD.n284 VDD.t359 28.565
R275 VDD.n284 VDD.t329 28.565
R276 VDD.n280 VDD.t199 28.565
R277 VDD.n280 VDD.t182 28.565
R278 VDD.n279 VDD.t255 28.565
R279 VDD.n279 VDD.t360 28.565
R280 VDD.n286 VDD.t400 28.565
R281 VDD.n286 VDD.t401 28.565
R282 VDD.n287 VDD.t76 28.565
R283 VDD.n287 VDD.t399 28.565
R284 VDD.n290 VDD.t87 28.565
R285 VDD.n290 VDD.t315 28.565
R286 VDD.n289 VDD.t105 28.565
R287 VDD.n289 VDD.t78 28.565
R288 VDD.n332 VDD.t10 28.565
R289 VDD.n332 VDD.t86 28.565
R290 VDD.n327 VDD.t440 28.565
R291 VDD.n327 VDD.t439 28.565
R292 VDD.n360 VDD.t200 28.565
R293 VDD.n360 VDD.t424 28.565
R294 VDD.n355 VDD.t185 28.565
R295 VDD.n355 VDD.t463 28.565
R296 VDD.n340 VDD.t457 28.565
R297 VDD.n340 VDD.t458 28.565
R298 VDD.n341 VDD.t281 28.565
R299 VDD.n341 VDD.t459 28.565
R300 VDD.n337 VDD.t422 28.565
R301 VDD.n337 VDD.t421 28.565
R302 VDD.n336 VDD.t309 28.565
R303 VDD.n336 VDD.t282 28.565
R304 VDD.n343 VDD.t163 28.565
R305 VDD.n343 VDD.t161 28.565
R306 VDD.n344 VDD.t416 28.565
R307 VDD.n344 VDD.t162 28.565
R308 VDD.n347 VDD.t42 28.565
R309 VDD.n347 VDD.t41 28.565
R310 VDD.n346 VDD.t420 28.565
R311 VDD.n346 VDD.t419 28.565
R312 VDD.n414 VDD.t106 28.565
R313 VDD.n414 VDD.t129 28.565
R314 VDD.n409 VDD.t352 28.565
R315 VDD.n409 VDD.t69 28.565
R316 VDD.n403 VDD.t13 28.565
R317 VDD.n403 VDD.t101 28.565
R318 VDD.n398 VDD.t168 28.565
R319 VDD.n398 VDD.t286 28.565
R320 VDD.n422 VDD.t495 28.565
R321 VDD.n422 VDD.t496 28.565
R322 VDD.n423 VDD.t264 28.565
R323 VDD.n423 VDD.t494 28.565
R324 VDD.n419 VDD.t63 28.565
R325 VDD.n419 VDD.t61 28.565
R326 VDD.n418 VDD.t159 28.565
R327 VDD.n418 VDD.t297 28.565
R328 VDD.n425 VDD.t333 28.565
R329 VDD.n425 VDD.t334 28.565
R330 VDD.n426 VDD.t14 28.565
R331 VDD.n426 VDD.t332 28.565
R332 VDD.n429 VDD.t468 28.565
R333 VDD.n429 VDD.t128 28.565
R334 VDD.n428 VDD.t133 28.565
R335 VDD.n428 VDD.t15 28.565
R336 VDD.n156 VDD.t473 28.565
R337 VDD.n156 VDD.t98 28.565
R338 VDD.n161 VDD.t223 28.565
R339 VDD.n161 VDD.t270 28.565
R340 VDD.n144 VDD.t134 28.565
R341 VDD.n144 VDD.t195 28.565
R342 VDD.n149 VDD.t435 28.565
R343 VDD.n149 VDD.t233 28.565
R344 VDD.n134 VDD.t296 28.565
R345 VDD.n134 VDD.t112 28.565
R346 VDD.n137 VDD.t149 28.565
R347 VDD.n137 VDD.t151 28.565
R348 VDD.n138 VDD.t150 28.565
R349 VDD.n138 VDD.t104 28.565
R350 VDD.n133 VDD.t344 28.565
R351 VDD.n133 VDD.t164 28.565
R352 VDD.n126 VDD.t232 28.565
R353 VDD.n126 VDD.t235 28.565
R354 VDD.n129 VDD.t173 28.565
R355 VDD.n129 VDD.t175 28.565
R356 VDD.n130 VDD.t174 28.565
R357 VDD.n130 VDD.t338 28.565
R358 VDD.n125 VDD.t222 28.565
R359 VDD.n125 VDD.t269 28.565
R360 VDD.n487 VDD.t237 14.284
R361 VDD.n493 VDD.t24 14.284
R362 VDD.n465 VDD.t180 14.284
R363 VDD.n471 VDD.t206 14.284
R364 VDD.n16 VDD.t477 14.284
R365 VDD.n11 VDD.t393 14.284
R366 VDD.n70 VDD.t409 14.284
R367 VDD.n75 VDD.t94 14.284
R368 VDD.n107 VDD.t216 14.284
R369 VDD.n112 VDD.t447 14.284
R370 VDD.n95 VDD.t27 14.284
R371 VDD.n100 VDD.t248 14.284
R372 VDD.n48 VDD.t487 14.284
R373 VDD.n53 VDD.t142 14.284
R374 VDD.n36 VDD.t127 14.284
R375 VDD.n41 VDD.t36 14.284
R376 VDD.n167 VDD.t432 14.284
R377 VDD.n172 VDD.t363 14.284
R378 VDD.n449 VDD.t47 14.284
R379 VDD.n454 VDD.t0 14.284
R380 VDD.n196 VDD.t367 14.284
R381 VDD.n202 VDD.t357 14.284
R382 VDD.n311 VDD.t72 14.284
R383 VDD.n316 VDD.t306 14.284
R384 VDD.n259 VDD.t294 14.284
R385 VDD.n254 VDD.t141 14.284
R386 VDD.n373 VDD.t242 14.284
R387 VDD.n368 VDD.t7 14.284
R388 VDD.n217 VDD.t312 14.284
R389 VDD.n212 VDD.t172 14.284
R390 VDD.n245 VDD.t474 14.284
R391 VDD.n240 VDD.t119 14.284
R392 VDD.n274 VDD.t236 14.284
R393 VDD.n269 VDD.t153 14.284
R394 VDD.n302 VDD.t320 14.284
R395 VDD.n297 VDD.t5 14.284
R396 VDD.n331 VDD.t183 14.284
R397 VDD.n326 VDD.t311 14.284
R398 VDD.n359 VDD.t415 14.284
R399 VDD.n354 VDD.t263 14.284
R400 VDD.n413 VDD.t18 14.284
R401 VDD.n408 VDD.t353 14.284
R402 VDD.n402 VDD.t100 14.284
R403 VDD.n397 VDD.t170 14.284
R404 VDD.n155 VDD.t97 14.284
R405 VDD.n160 VDD.t43 14.284
R406 VDD.n143 VDD.t303 14.284
R407 VDD.n148 VDD.t234 14.284
R408 VDD.n484 VDD.t239 14.282
R409 VDD.n484 VDD.t238 14.282
R410 VDD.n490 VDD.t26 14.282
R411 VDD.n490 VDD.t25 14.282
R412 VDD.n462 VDD.t179 14.282
R413 VDD.n462 VDD.t181 14.282
R414 VDD.n468 VDD.t207 14.282
R415 VDD.n468 VDD.t205 14.282
R416 VDD.n13 VDD.t478 14.282
R417 VDD.n13 VDD.t476 14.282
R418 VDD.n8 VDD.t395 14.282
R419 VDD.n8 VDD.t394 14.282
R420 VDD.n67 VDD.t408 14.282
R421 VDD.n67 VDD.t410 14.282
R422 VDD.n72 VDD.t96 14.282
R423 VDD.n72 VDD.t95 14.282
R424 VDD.n106 VDD.t221 14.282
R425 VDD.n106 VDD.t220 14.282
R426 VDD.n111 VDD.t446 14.282
R427 VDD.n111 VDD.t444 14.282
R428 VDD.n94 VDD.t177 14.282
R429 VDD.n94 VDD.t193 14.282
R430 VDD.n99 VDD.t455 14.282
R431 VDD.n99 VDD.t265 14.282
R432 VDD.n47 VDD.t486 14.282
R433 VDD.n47 VDD.t485 14.282
R434 VDD.n52 VDD.t350 14.282
R435 VDD.n52 VDD.t17 14.282
R436 VDD.n35 VDD.t125 14.282
R437 VDD.n35 VDD.t411 14.282
R438 VDD.n40 VDD.t146 14.282
R439 VDD.n40 VDD.t109 14.282
R440 VDD.n166 VDD.t30 14.282
R441 VDD.n166 VDD.t29 14.282
R442 VDD.n171 VDD.t321 14.282
R443 VDD.n171 VDD.t336 14.282
R444 VDD.n448 VDD.t358 14.282
R445 VDD.n448 VDD.t88 14.282
R446 VDD.n453 VDD.t40 14.282
R447 VDD.n453 VDD.t91 14.282
R448 VDD.n193 VDD.t365 14.282
R449 VDD.n193 VDD.t366 14.282
R450 VDD.n199 VDD.t355 14.282
R451 VDD.n199 VDD.t356 14.282
R452 VDD.n308 VDD.t73 14.282
R453 VDD.n308 VDD.t74 14.282
R454 VDD.n313 VDD.t307 14.282
R455 VDD.n313 VDD.t308 14.282
R456 VDD.n256 VDD.t292 14.282
R457 VDD.n256 VDD.t293 14.282
R458 VDD.n251 VDD.t139 14.282
R459 VDD.n251 VDD.t140 14.282
R460 VDD.n370 VDD.t240 14.282
R461 VDD.n370 VDD.t241 14.282
R462 VDD.n365 VDD.t8 14.282
R463 VDD.n365 VDD.t9 14.282
R464 VDD.n216 VDD.t316 14.282
R465 VDD.n216 VDD.t299 14.282
R466 VDD.n211 VDD.t171 14.282
R467 VDD.n211 VDD.t190 14.282
R468 VDD.n244 VDD.t340 14.282
R469 VDD.n244 VDD.t475 14.282
R470 VDD.n239 VDD.t118 14.282
R471 VDD.n239 VDD.t167 14.282
R472 VDD.n273 VDD.t304 14.282
R473 VDD.n273 VDD.t51 14.282
R474 VDD.n268 VDD.t152 14.282
R475 VDD.n268 VDD.t154 14.282
R476 VDD.n301 VDD.t279 14.282
R477 VDD.n301 VDD.t380 14.282
R478 VDD.n296 VDD.t6 14.282
R479 VDD.n296 VDD.t4 14.282
R480 VDD.n330 VDD.t387 14.282
R481 VDD.n330 VDD.t12 14.282
R482 VDD.n325 VDD.t280 14.282
R483 VDD.n325 VDD.t343 14.282
R484 VDD.n358 VDD.t418 14.282
R485 VDD.n358 VDD.t417 14.282
R486 VDD.n353 VDD.t75 14.282
R487 VDD.n353 VDD.t461 14.282
R488 VDD.n412 VDD.t464 14.282
R489 VDD.n412 VDD.t467 14.282
R490 VDD.n407 VDD.t71 14.282
R491 VDD.n407 VDD.t70 14.282
R492 VDD.n401 VDD.t437 14.282
R493 VDD.n401 VDD.t132 14.282
R494 VDD.n396 VDD.t169 14.282
R495 VDD.n396 VDD.t131 14.282
R496 VDD.n154 VDD.t99 14.282
R497 VDD.n154 VDD.t64 14.282
R498 VDD.n159 VDD.t271 14.282
R499 VDD.n159 VDD.t111 14.282
R500 VDD.n142 VDD.t384 14.282
R501 VDD.n142 VDD.t114 14.282
R502 VDD.n147 VDD.t374 14.282
R503 VDD.n147 VDD.t251 14.282
R504 VDD.n116 VDD.n110 4.276
R505 VDD.n104 VDD.n98 4.276
R506 VDD.n57 VDD.n51 4.276
R507 VDD.n45 VDD.n39 4.276
R508 VDD.n176 VDD.n170 4.276
R509 VDD.n458 VDD.n452 4.276
R510 VDD.n221 VDD.n215 4.276
R511 VDD.n249 VDD.n243 4.276
R512 VDD.n278 VDD.n272 4.276
R513 VDD.n306 VDD.n300 4.276
R514 VDD.n335 VDD.n329 4.276
R515 VDD.n363 VDD.n357 4.276
R516 VDD.n417 VDD.n411 4.276
R517 VDD.n406 VDD.n400 4.276
R518 VDD.n164 VDD.n158 4.276
R519 VDD.n152 VDD.n146 4.276
R520 VDD.n109 VDD.n108 2.451
R521 VDD.n97 VDD.n96 2.451
R522 VDD.n50 VDD.n49 2.451
R523 VDD.n38 VDD.n37 2.451
R524 VDD.n169 VDD.n168 2.451
R525 VDD.n451 VDD.n450 2.451
R526 VDD.n214 VDD.n213 2.451
R527 VDD.n242 VDD.n241 2.451
R528 VDD.n271 VDD.n270 2.451
R529 VDD.n299 VDD.n298 2.451
R530 VDD.n328 VDD.n327 2.451
R531 VDD.n356 VDD.n355 2.451
R532 VDD.n410 VDD.n409 2.451
R533 VDD.n399 VDD.n398 2.451
R534 VDD.n157 VDD.n156 2.451
R535 VDD.n145 VDD.n144 2.451
R536 VDD.n114 VDD.n113 2.449
R537 VDD.n102 VDD.n101 2.449
R538 VDD.n55 VDD.n54 2.449
R539 VDD.n43 VDD.n42 2.449
R540 VDD.n174 VDD.n173 2.449
R541 VDD.n456 VDD.n455 2.449
R542 VDD.n219 VDD.n218 2.449
R543 VDD.n247 VDD.n246 2.449
R544 VDD.n276 VDD.n275 2.449
R545 VDD.n304 VDD.n303 2.449
R546 VDD.n333 VDD.n332 2.449
R547 VDD.n361 VDD.n360 2.449
R548 VDD.n415 VDD.n414 2.449
R549 VDD.n404 VDD.n403 2.449
R550 VDD.n162 VDD.n161 2.449
R551 VDD.n150 VDD.n149 2.449
R552 VDD.n487 VDD.n486 2.195
R553 VDD.n493 VDD.n492 2.195
R554 VDD.n465 VDD.n464 2.195
R555 VDD.n471 VDD.n470 2.195
R556 VDD.n16 VDD.n15 2.195
R557 VDD.n11 VDD.n10 2.195
R558 VDD.n70 VDD.n69 2.195
R559 VDD.n75 VDD.n74 2.195
R560 VDD.n196 VDD.n195 2.195
R561 VDD.n202 VDD.n201 2.195
R562 VDD.n311 VDD.n310 2.195
R563 VDD.n316 VDD.n315 2.195
R564 VDD.n259 VDD.n258 2.195
R565 VDD.n254 VDD.n253 2.195
R566 VDD.n373 VDD.n372 2.195
R567 VDD.n368 VDD.n367 2.195
R568 VDD.n494 VDD.n490 1.72
R569 VDD.n472 VDD.n468 1.72
R570 VDD.n17 VDD.n13 1.72
R571 VDD.n76 VDD.n72 1.72
R572 VDD.n197 VDD.n193 1.72
R573 VDD.n312 VDD.n308 1.72
R574 VDD.n255 VDD.n251 1.72
R575 VDD.n369 VDD.n365 1.72
R576 VDD.n488 VDD.n484 1.698
R577 VDD.n466 VDD.n462 1.698
R578 VDD.n12 VDD.n8 1.698
R579 VDD.n71 VDD.n67 1.698
R580 VDD.n203 VDD.n199 1.698
R581 VDD.n317 VDD.n313 1.698
R582 VDD.n260 VDD.n256 1.698
R583 VDD.n374 VDD.n370 1.698
R584 VDD.n486 VDD.n485 1.651
R585 VDD.n492 VDD.n491 1.651
R586 VDD.n464 VDD.n463 1.651
R587 VDD.n470 VDD.n469 1.651
R588 VDD.n15 VDD.n14 1.651
R589 VDD.n10 VDD.n9 1.651
R590 VDD.n69 VDD.n68 1.651
R591 VDD.n74 VDD.n73 1.651
R592 VDD.n195 VDD.n194 1.651
R593 VDD.n201 VDD.n200 1.651
R594 VDD.n310 VDD.n309 1.651
R595 VDD.n315 VDD.n314 1.651
R596 VDD.n258 VDD.n257 1.651
R597 VDD.n253 VDD.n252 1.651
R598 VDD.n372 VDD.n371 1.651
R599 VDD.n367 VDD.n366 1.651
R600 VDD.n481 VDD.n479 1.564
R601 VDD.n180 VDD.n178 1.564
R602 VDD.n6 VDD.n4 1.564
R603 VDD.n65 VDD.n63 1.564
R604 VDD.n91 VDD.n89 1.564
R605 VDD.n83 VDD.n81 1.564
R606 VDD.n32 VDD.n30 1.564
R607 VDD.n24 VDD.n22 1.564
R608 VDD.n446 VDD.n444 1.564
R609 VDD.n191 VDD.n189 1.564
R610 VDD.n210 VDD.n208 1.564
R611 VDD.n267 VDD.n265 1.564
R612 VDD.n324 VDD.n322 1.564
R613 VDD.n381 VDD.n379 1.564
R614 VDD.n228 VDD.n226 1.564
R615 VDD.n231 VDD.n229 1.564
R616 VDD.n285 VDD.n283 1.564
R617 VDD.n288 VDD.n286 1.564
R618 VDD.n342 VDD.n340 1.564
R619 VDD.n345 VDD.n343 1.564
R620 VDD.n424 VDD.n422 1.564
R621 VDD.n427 VDD.n425 1.564
R622 VDD.n139 VDD.n137 1.564
R623 VDD.n131 VDD.n129 1.564
R624 VDD.n110 VDD.n106 0.922
R625 VDD.n115 VDD.n111 0.922
R626 VDD.n98 VDD.n94 0.922
R627 VDD.n103 VDD.n99 0.922
R628 VDD.n51 VDD.n47 0.922
R629 VDD.n56 VDD.n52 0.922
R630 VDD.n39 VDD.n35 0.922
R631 VDD.n44 VDD.n40 0.922
R632 VDD.n170 VDD.n166 0.922
R633 VDD.n175 VDD.n171 0.922
R634 VDD.n452 VDD.n448 0.922
R635 VDD.n457 VDD.n453 0.922
R636 VDD.n220 VDD.n216 0.922
R637 VDD.n215 VDD.n211 0.922
R638 VDD.n248 VDD.n244 0.922
R639 VDD.n243 VDD.n239 0.922
R640 VDD.n277 VDD.n273 0.922
R641 VDD.n272 VDD.n268 0.922
R642 VDD.n305 VDD.n301 0.922
R643 VDD.n300 VDD.n296 0.922
R644 VDD.n334 VDD.n330 0.922
R645 VDD.n329 VDD.n325 0.922
R646 VDD.n362 VDD.n358 0.922
R647 VDD.n357 VDD.n353 0.922
R648 VDD.n416 VDD.n412 0.922
R649 VDD.n411 VDD.n407 0.922
R650 VDD.n405 VDD.n401 0.922
R651 VDD.n400 VDD.n396 0.922
R652 VDD.n158 VDD.n154 0.922
R653 VDD.n163 VDD.n159 0.922
R654 VDD.n146 VDD.n142 0.922
R655 VDD.n151 VDD.n147 0.922
R656 VDD.n109 VDD.n107 0.921
R657 VDD.n114 VDD.n112 0.921
R658 VDD.n97 VDD.n95 0.921
R659 VDD.n102 VDD.n100 0.921
R660 VDD.n50 VDD.n48 0.921
R661 VDD.n55 VDD.n53 0.921
R662 VDD.n38 VDD.n36 0.921
R663 VDD.n43 VDD.n41 0.921
R664 VDD.n169 VDD.n167 0.921
R665 VDD.n174 VDD.n172 0.921
R666 VDD.n451 VDD.n449 0.921
R667 VDD.n456 VDD.n454 0.921
R668 VDD.n219 VDD.n217 0.921
R669 VDD.n214 VDD.n212 0.921
R670 VDD.n247 VDD.n245 0.921
R671 VDD.n242 VDD.n240 0.921
R672 VDD.n276 VDD.n274 0.921
R673 VDD.n271 VDD.n269 0.921
R674 VDD.n304 VDD.n302 0.921
R675 VDD.n299 VDD.n297 0.921
R676 VDD.n333 VDD.n331 0.921
R677 VDD.n328 VDD.n326 0.921
R678 VDD.n361 VDD.n359 0.921
R679 VDD.n356 VDD.n354 0.921
R680 VDD.n415 VDD.n413 0.921
R681 VDD.n410 VDD.n408 0.921
R682 VDD.n404 VDD.n402 0.921
R683 VDD.n399 VDD.n397 0.921
R684 VDD.n157 VDD.n155 0.921
R685 VDD.n162 VDD.n160 0.921
R686 VDD.n145 VDD.n143 0.921
R687 VDD.n150 VDD.n148 0.921
R688 VDD.n488 VDD.n487 0.806
R689 VDD.n466 VDD.n465 0.806
R690 VDD.n12 VDD.n11 0.806
R691 VDD.n71 VDD.n70 0.806
R692 VDD.n203 VDD.n202 0.806
R693 VDD.n317 VDD.n316 0.806
R694 VDD.n260 VDD.n259 0.806
R695 VDD.n374 VDD.n373 0.806
R696 VDD.n494 VDD.n493 0.778
R697 VDD.n472 VDD.n471 0.778
R698 VDD.n17 VDD.n16 0.778
R699 VDD.n76 VDD.n75 0.778
R700 VDD.n197 VDD.n196 0.778
R701 VDD.n312 VDD.n311 0.778
R702 VDD.n255 VDD.n254 0.778
R703 VDD.n369 VDD.n368 0.778
R704 VDD.n477 VDD.n476 0.747
R705 VDD.n481 VDD.n480 0.747
R706 VDD.n183 VDD.n182 0.747
R707 VDD.n180 VDD.n179 0.747
R708 VDD.n2 VDD.n1 0.747
R709 VDD.n6 VDD.n5 0.747
R710 VDD.n61 VDD.n60 0.747
R711 VDD.n65 VDD.n64 0.747
R712 VDD.n87 VDD.n86 0.747
R713 VDD.n91 VDD.n90 0.747
R714 VDD.n79 VDD.n78 0.747
R715 VDD.n83 VDD.n82 0.747
R716 VDD.n28 VDD.n27 0.747
R717 VDD.n32 VDD.n31 0.747
R718 VDD.n20 VDD.n19 0.747
R719 VDD.n24 VDD.n23 0.747
R720 VDD.n442 VDD.n441 0.747
R721 VDD.n446 VDD.n445 0.747
R722 VDD.n187 VDD.n186 0.747
R723 VDD.n191 VDD.n190 0.747
R724 VDD.n210 VDD.n209 0.747
R725 VDD.n206 VDD.n205 0.747
R726 VDD.n267 VDD.n266 0.747
R727 VDD.n263 VDD.n262 0.747
R728 VDD.n324 VDD.n323 0.747
R729 VDD.n320 VDD.n319 0.747
R730 VDD.n381 VDD.n380 0.747
R731 VDD.n377 VDD.n376 0.747
R732 VDD.n228 VDD.n227 0.747
R733 VDD.n224 VDD.n223 0.747
R734 VDD.n231 VDD.n230 0.747
R735 VDD.n234 VDD.n233 0.747
R736 VDD.n285 VDD.n284 0.747
R737 VDD.n281 VDD.n280 0.747
R738 VDD.n288 VDD.n287 0.747
R739 VDD.n291 VDD.n290 0.747
R740 VDD.n342 VDD.n341 0.747
R741 VDD.n338 VDD.n337 0.747
R742 VDD.n345 VDD.n344 0.747
R743 VDD.n348 VDD.n347 0.747
R744 VDD.n424 VDD.n423 0.747
R745 VDD.n420 VDD.n419 0.747
R746 VDD.n427 VDD.n426 0.747
R747 VDD.n430 VDD.n429 0.747
R748 VDD.n135 VDD.n134 0.747
R749 VDD.n139 VDD.n138 0.747
R750 VDD.n127 VDD.n126 0.747
R751 VDD.n131 VDD.n130 0.747
R752 VDD.n478 VDD.n475 0.689
R753 VDD.n184 VDD.n181 0.689
R754 VDD.n3 VDD.n0 0.689
R755 VDD.n62 VDD.n59 0.689
R756 VDD.n88 VDD.n85 0.689
R757 VDD.n80 VDD.n77 0.689
R758 VDD.n29 VDD.n26 0.689
R759 VDD.n21 VDD.n18 0.689
R760 VDD.n443 VDD.n440 0.689
R761 VDD.n188 VDD.n185 0.689
R762 VDD.n207 VDD.n204 0.689
R763 VDD.n264 VDD.n261 0.689
R764 VDD.n321 VDD.n318 0.689
R765 VDD.n378 VDD.n375 0.689
R766 VDD.n225 VDD.n222 0.689
R767 VDD.n235 VDD.n232 0.689
R768 VDD.n282 VDD.n279 0.689
R769 VDD.n292 VDD.n289 0.689
R770 VDD.n339 VDD.n336 0.689
R771 VDD.n349 VDD.n346 0.689
R772 VDD.n421 VDD.n418 0.689
R773 VDD.n431 VDD.n428 0.689
R774 VDD.n136 VDD.n133 0.689
R775 VDD.n128 VDD.n125 0.689
R776 VDD.n110 VDD.n109 0.686
R777 VDD.n115 VDD.n114 0.686
R778 VDD.n98 VDD.n97 0.686
R779 VDD.n103 VDD.n102 0.686
R780 VDD.n51 VDD.n50 0.686
R781 VDD.n56 VDD.n55 0.686
R782 VDD.n39 VDD.n38 0.686
R783 VDD.n44 VDD.n43 0.686
R784 VDD.n170 VDD.n169 0.686
R785 VDD.n175 VDD.n174 0.686
R786 VDD.n452 VDD.n451 0.686
R787 VDD.n457 VDD.n456 0.686
R788 VDD.n220 VDD.n219 0.686
R789 VDD.n215 VDD.n214 0.686
R790 VDD.n248 VDD.n247 0.686
R791 VDD.n243 VDD.n242 0.686
R792 VDD.n277 VDD.n276 0.686
R793 VDD.n272 VDD.n271 0.686
R794 VDD.n305 VDD.n304 0.686
R795 VDD.n300 VDD.n299 0.686
R796 VDD.n334 VDD.n333 0.686
R797 VDD.n329 VDD.n328 0.686
R798 VDD.n362 VDD.n361 0.686
R799 VDD.n357 VDD.n356 0.686
R800 VDD.n416 VDD.n415 0.686
R801 VDD.n411 VDD.n410 0.686
R802 VDD.n405 VDD.n404 0.686
R803 VDD.n400 VDD.n399 0.686
R804 VDD.n158 VDD.n157 0.686
R805 VDD.n163 VDD.n162 0.686
R806 VDD.n146 VDD.n145 0.686
R807 VDD.n151 VDD.n150 0.686
R808 VDD.n478 VDD.n477 0.59
R809 VDD.n184 VDD.n183 0.59
R810 VDD.n3 VDD.n2 0.59
R811 VDD.n62 VDD.n61 0.59
R812 VDD.n88 VDD.n87 0.59
R813 VDD.n80 VDD.n79 0.59
R814 VDD.n29 VDD.n28 0.59
R815 VDD.n21 VDD.n20 0.59
R816 VDD.n443 VDD.n442 0.59
R817 VDD.n188 VDD.n187 0.59
R818 VDD.n207 VDD.n206 0.59
R819 VDD.n264 VDD.n263 0.59
R820 VDD.n321 VDD.n320 0.59
R821 VDD.n378 VDD.n377 0.59
R822 VDD.n225 VDD.n224 0.59
R823 VDD.n235 VDD.n234 0.59
R824 VDD.n282 VDD.n281 0.59
R825 VDD.n292 VDD.n291 0.59
R826 VDD.n339 VDD.n338 0.59
R827 VDD.n349 VDD.n348 0.59
R828 VDD.n421 VDD.n420 0.59
R829 VDD.n431 VDD.n430 0.59
R830 VDD.n136 VDD.n135 0.59
R831 VDD.n128 VDD.n127 0.59
R832 VDD.n482 VDD.n481 0.451
R833 VDD.n461 VDD.n180 0.451
R834 VDD.n7 VDD.n6 0.451
R835 VDD.n66 VDD.n65 0.451
R836 VDD.n92 VDD.n91 0.451
R837 VDD.n84 VDD.n83 0.451
R838 VDD.n33 VDD.n32 0.451
R839 VDD.n25 VDD.n24 0.451
R840 VDD.n447 VDD.n446 0.451
R841 VDD.n192 VDD.n191 0.451
R842 VDD.n394 VDD.n210 0.451
R843 VDD.n390 VDD.n267 0.451
R844 VDD.n386 VDD.n324 0.451
R845 VDD.n382 VDD.n381 0.451
R846 VDD.n237 VDD.n228 0.451
R847 VDD.n236 VDD.n231 0.451
R848 VDD.n294 VDD.n285 0.451
R849 VDD.n293 VDD.n288 0.451
R850 VDD.n351 VDD.n342 0.451
R851 VDD.n350 VDD.n345 0.451
R852 VDD.n433 VDD.n424 0.451
R853 VDD.n432 VDD.n427 0.451
R854 VDD.n140 VDD.n139 0.451
R855 VDD.n132 VDD.n131 0.451
R856 VDD.n93 VDD.n84 0.276
R857 VDD.n34 VDD.n25 0.276
R858 VDD.n141 VDD.n132 0.276
R859 VDD.n237 VDD.n236 0.272
R860 VDD.n294 VDD.n293 0.272
R861 VDD.n351 VDD.n350 0.272
R862 VDD.n433 VDD.n432 0.272
R863 VDD.n395 VDD.n203 0.254
R864 VDD.n387 VDD.n317 0.254
R865 VDD.n391 VDD.n260 0.254
R866 VDD.n383 VDD.n374 0.254
R867 VDD.n489 VDD.n488 0.253
R868 VDD.n467 VDD.n466 0.253
R869 VDD.n123 VDD.n12 0.253
R870 VDD.n119 VDD.n71 0.253
R871 VDD.n198 VDD.n197 0.242
R872 VDD.n388 VDD.n312 0.242
R873 VDD.n392 VDD.n255 0.242
R874 VDD.n384 VDD.n369 0.242
R875 VDD.n495 VDD.n494 0.241
R876 VDD.n473 VDD.n472 0.241
R877 VDD.n122 VDD.n17 0.241
R878 VDD.n118 VDD.n76 0.241
R879 VDD.n116 VDD.n115 0.179
R880 VDD.n104 VDD.n103 0.179
R881 VDD.n57 VDD.n56 0.179
R882 VDD.n45 VDD.n44 0.179
R883 VDD.n176 VDD.n175 0.179
R884 VDD.n458 VDD.n457 0.179
R885 VDD.n221 VDD.n220 0.179
R886 VDD.n249 VDD.n248 0.179
R887 VDD.n278 VDD.n277 0.179
R888 VDD.n306 VDD.n305 0.179
R889 VDD.n335 VDD.n334 0.179
R890 VDD.n363 VDD.n362 0.179
R891 VDD.n417 VDD.n416 0.179
R892 VDD.n406 VDD.n405 0.179
R893 VDD.n164 VDD.n163 0.179
R894 VDD.n152 VDD.n151 0.179
R895 VDD.n435 VDD.n434 0.177
R896 VDD.n436 VDD.n435 0.176
R897 VDD.n250 VDD.n238 0.174
R898 VDD.n307 VDD.n295 0.174
R899 VDD.n364 VDD.n352 0.174
R900 VDD.n117 VDD.n105 0.174
R901 VDD.n58 VDD.n46 0.174
R902 VDD.n459 VDD.n177 0.174
R903 VDD.n165 VDD.n153 0.174
R904 VDD.n460 VDD.n459 0.172
R905 VDD.n121 VDD.n120 0.164
R906 VDD.n120 VDD.n119 0.163
R907 VDD.n483 VDD.n474 0.162
R908 VDD.n394 VDD.n393 0.162
R909 VDD.n105 VDD.n93 0.161
R910 VDD.n46 VDD.n34 0.161
R911 VDD.n153 VDD.n141 0.161
R912 VDD.n390 VDD.n389 0.161
R913 VDD.n467 VDD.n461 0.161
R914 VDD.n395 VDD.n394 0.161
R915 VDD.n489 VDD.n483 0.16
R916 VDD.n386 VDD.n385 0.16
R917 VDD.n383 VDD.n382 0.16
R918 VDD.n124 VDD.n123 0.159
R919 VDD.n238 VDD.n237 0.159
R920 VDD.n295 VDD.n294 0.159
R921 VDD.n352 VDD.n351 0.159
R922 VDD.n434 VDD.n433 0.159
R923 VDD.n387 VDD.n386 0.158
R924 VDD.n391 VDD.n390 0.158
R925 VDD.n118 VDD.n117 0.153
R926 VDD.n105 VDD.n104 0.142
R927 VDD.n46 VDD.n45 0.142
R928 VDD.n459 VDD.n458 0.142
R929 VDD.n153 VDD.n152 0.142
R930 VDD.n117 VDD.n116 0.141
R931 VDD.n58 VDD.n57 0.141
R932 VDD.n177 VDD.n176 0.141
R933 VDD.n238 VDD.n221 0.141
R934 VDD.n250 VDD.n249 0.141
R935 VDD.n295 VDD.n278 0.141
R936 VDD.n307 VDD.n306 0.141
R937 VDD.n352 VDD.n335 0.141
R938 VDD.n364 VDD.n363 0.141
R939 VDD.n434 VDD.n417 0.141
R940 VDD.n435 VDD.n406 0.141
R941 VDD.n165 VDD.n164 0.141
R942 VDD.n121 VDD.n58 0.129
R943 VDD.n393 VDD.n250 0.129
R944 VDD.n474 VDD.n177 0.129
R945 VDD.n496 VDD.n165 0.129
R946 VDD.n389 VDD.n307 0.128
R947 VDD.n385 VDD.n364 0.128
R948 VDD VDD.n124 0.114
R949 VDD.n461 VDD.n460 0.109
R950 VDD.n439 VDD.n438 0.108
R951 VDD.n460 VDD.n439 0.082
R952 VDD.n119 VDD.n118 0.078
R953 VDD.n495 VDD.n489 0.075
R954 VDD.n473 VDD.n467 0.075
R955 VDD.n123 VDD.n122 0.075
R956 VDD.n384 VDD.n383 0.073
R957 VDD.n388 VDD.n387 0.073
R958 VDD.n392 VDD.n391 0.073
R959 VDD.n437 VDD.n395 0.055
R960 VDD VDD.n496 0.048
R961 VDD.n385 VDD.n384 0.023
R962 VDD.n389 VDD.n388 0.023
R963 VDD.n393 VDD.n392 0.023
R964 VDD.n122 VDD.n121 0.023
R965 VDD.n474 VDD.n473 0.023
R966 VDD.n460 VDD.n447 0.019
R967 VDD VDD.n495 0.019
R968 VDD.n482 VDD.n478 0.011
R969 VDD.n461 VDD.n184 0.011
R970 VDD.n7 VDD.n3 0.011
R971 VDD.n66 VDD.n62 0.011
R972 VDD.n92 VDD.n88 0.011
R973 VDD.n84 VDD.n80 0.011
R974 VDD.n33 VDD.n29 0.011
R975 VDD.n25 VDD.n21 0.011
R976 VDD.n447 VDD.n443 0.011
R977 VDD.n192 VDD.n188 0.011
R978 VDD.n394 VDD.n207 0.011
R979 VDD.n390 VDD.n264 0.011
R980 VDD.n386 VDD.n321 0.011
R981 VDD.n382 VDD.n378 0.011
R982 VDD.n237 VDD.n225 0.011
R983 VDD.n236 VDD.n235 0.011
R984 VDD.n294 VDD.n282 0.011
R985 VDD.n293 VDD.n292 0.011
R986 VDD.n351 VDD.n339 0.011
R987 VDD.n350 VDD.n349 0.011
R988 VDD.n433 VDD.n421 0.011
R989 VDD.n432 VDD.n431 0.011
R990 VDD.n140 VDD.n136 0.011
R991 VDD.n132 VDD.n128 0.011
R992 VDD.n439 VDD.n192 0.011
R993 VDD.n496 VDD 0.004
R994 VDD.n438 VDD.n198 0.002
R995 VDD.n438 VDD.n437 0.001
R996 VDD.n93 VDD.n92 0.001
R997 VDD.n34 VDD.n33 0.001
R998 VDD.n141 VDD.n140 0.001
R999 VDD.n483 VDD.n482 0.001
R1000 VDD.n124 VDD.n7 0.001
R1001 VDD.n120 VDD.n66 0.001
R1002 VDD.n436 VDD.n198 0.001
R1003 VDD.n437 VDD.n436 0.001
R1004 B[3].n7 B[3].n6 861.987
R1005 B[3].n6 B[3].n5 560.726
R1006 B[3].t12 B[3].t10 415.315
R1007 B[3].t3 B[3].t1 415.315
R1008 B[3].n2 B[3].t14 394.151
R1009 B[3].n5 B[3].t5 294.653
R1010 B[3].n1 B[3].t2 269.523
R1011 B[3].t14 B[3].n1 269.523
R1012 B[3].n9 B[3].t12 217.716
R1013 B[3].n8 B[3].t4 214.335
R1014 B[3].t10 B[3].n8 214.335
R1015 B[3].n0 B[3].t8 214.335
R1016 B[3].t1 B[3].n0 214.335
R1017 B[3].n7 B[3].t3 198.921
R1018 B[3].n3 B[3].t6 198.043
R1019 B[3].n1 B[3].t7 160.666
R1020 B[3].n5 B[3].t13 111.663
R1021 B[3].n4 B[3].n2 97.816
R1022 B[3].n3 B[3].t0 93.989
R1023 B[3].n8 B[3].t11 80.333
R1024 B[3].n2 B[3].t9 80.333
R1025 B[3].n0 B[3].t15 80.333
R1026 B[3].n6 B[3].n4 65.07
R1027 B[3].n9 B[3].n7 16.411
R1028 B[3].n4 B[3].n3 6.615
R1029 B[3] B[3].n9 0.453
R1030 a_19657_n3503.n6 a_19657_n3503.n5 501.28
R1031 a_19657_n3503.t16 a_19657_n3503.t14 437.233
R1032 a_19657_n3503.t9 a_19657_n3503.t13 415.315
R1033 a_19657_n3503.t5 a_19657_n3503.n3 313.873
R1034 a_19657_n3503.n5 a_19657_n3503.t7 294.986
R1035 a_19657_n3503.n2 a_19657_n3503.t11 272.288
R1036 a_19657_n3503.n6 a_19657_n3503.t4 236.009
R1037 a_19657_n3503.n9 a_19657_n3503.t16 216.627
R1038 a_19657_n3503.n7 a_19657_n3503.t9 216.111
R1039 a_19657_n3503.n8 a_19657_n3503.t18 214.686
R1040 a_19657_n3503.t14 a_19657_n3503.n8 214.686
R1041 a_19657_n3503.n1 a_19657_n3503.t8 214.335
R1042 a_19657_n3503.t13 a_19657_n3503.n1 214.335
R1043 a_19657_n3503.n4 a_19657_n3503.t19 190.152
R1044 a_19657_n3503.n4 a_19657_n3503.t5 190.152
R1045 a_19657_n3503.n2 a_19657_n3503.t10 160.666
R1046 a_19657_n3503.n3 a_19657_n3503.t6 160.666
R1047 a_19657_n3503.n7 a_19657_n3503.n6 148.428
R1048 a_19657_n3503.n5 a_19657_n3503.t15 110.859
R1049 a_19657_n3503.n3 a_19657_n3503.n2 96.129
R1050 a_19657_n3503.n8 a_19657_n3503.t17 80.333
R1051 a_19657_n3503.n1 a_19657_n3503.t12 80.333
R1052 a_19657_n3503.t4 a_19657_n3503.n4 80.333
R1053 a_19657_n3503.n0 a_19657_n3503.t2 28.57
R1054 a_19657_n3503.n11 a_19657_n3503.t1 28.565
R1055 a_19657_n3503.t3 a_19657_n3503.n11 28.565
R1056 a_19657_n3503.n0 a_19657_n3503.t0 17.638
R1057 a_19657_n3503.n10 a_19657_n3503.n9 10.943
R1058 a_19657_n3503.n9 a_19657_n3503.n7 2.923
R1059 a_19657_n3503.n11 a_19657_n3503.n10 0.69
R1060 a_19657_n3503.n10 a_19657_n3503.n0 0.6
R1061 B[0].n7 B[0].n6 861.987
R1062 B[0].n6 B[0].n5 560.726
R1063 B[0].t0 B[0].t15 415.315
R1064 B[0].t6 B[0].t3 415.315
R1065 B[0].n2 B[0].t10 394.151
R1066 B[0].n5 B[0].t11 294.653
R1067 B[0].n1 B[0].t5 269.523
R1068 B[0].t10 B[0].n1 269.523
R1069 B[0].n9 B[0].t0 217.716
R1070 B[0].n8 B[0].t2 214.335
R1071 B[0].t15 B[0].n8 214.335
R1072 B[0].n0 B[0].t8 214.335
R1073 B[0].t3 B[0].n0 214.335
R1074 B[0].n7 B[0].t6 198.921
R1075 B[0].n3 B[0].t4 198.043
R1076 B[0].n1 B[0].t12 160.666
R1077 B[0].n5 B[0].t1 111.663
R1078 B[0].n4 B[0].n2 97.816
R1079 B[0].n3 B[0].t14 93.989
R1080 B[0].n8 B[0].t7 80.333
R1081 B[0].n2 B[0].t9 80.333
R1082 B[0].n0 B[0].t13 80.333
R1083 B[0].n6 B[0].n4 65.07
R1084 B[0].n9 B[0].n7 16.411
R1085 B[0].n4 B[0].n3 6.615
R1086 B[0] B[0].n9 0.458
R1087 VSS.n156 VSS.t60 20.763
R1088 VSS.n136 VSS.t141 20.763
R1089 VSS.n145 VSS.t24 20.763
R1090 VSS.n140 VSS.t30 20.763
R1091 VSS.n127 VSS.t17 20.763
R1092 VSS.n1 VSS.t4 20.763
R1093 VSS.n108 VSS.t104 20.763
R1094 VSS.n111 VSS.t153 20.763
R1095 VSS.n7 VSS.t43 20.763
R1096 VSS.n88 VSS.t143 20.763
R1097 VSS.n70 VSS.t44 20.763
R1098 VSS.n19 VSS.t107 20.763
R1099 VSS.n63 VSS.t63 20.763
R1100 VSS.n54 VSS.t62 20.763
R1101 VSS.n34 VSS.t72 20.763
R1102 VSS.n29 VSS.t110 20.763
R1103 VSS.n157 VSS.t54 20.606
R1104 VSS.n137 VSS.t33 20.606
R1105 VSS.n146 VSS.t87 20.606
R1106 VSS.n141 VSS.t14 20.606
R1107 VSS.n128 VSS.t0 20.606
R1108 VSS.n2 VSS.t69 20.606
R1109 VSS.n109 VSS.t52 20.606
R1110 VSS.n112 VSS.t105 20.606
R1111 VSS.n8 VSS.t61 20.606
R1112 VSS.n89 VSS.t37 20.606
R1113 VSS.n71 VSS.t136 20.606
R1114 VSS.n20 VSS.t151 20.606
R1115 VSS.n64 VSS.t149 20.606
R1116 VSS.n55 VSS.t94 20.606
R1117 VSS.n35 VSS.t157 20.606
R1118 VSS.n30 VSS.t9 20.606
R1119 VSS.n134 VSS.t137 18.185
R1120 VSS.n169 VSS.t13 18.185
R1121 VSS.n168 VSS.t116 18.185
R1122 VSS.n138 VSS.t99 18.185
R1123 VSS.n151 VSS.t40 18.185
R1124 VSS.n3 VSS.t132 18.185
R1125 VSS.n5 VSS.t98 18.185
R1126 VSS.n4 VSS.t134 18.185
R1127 VSS.n106 VSS.t48 18.185
R1128 VSS.n105 VSS.t144 18.185
R1129 VSS.n101 VSS.t82 18.185
R1130 VSS.n13 VSS.t122 18.185
R1131 VSS.n84 VSS.t28 18.185
R1132 VSS.n85 VSS.t96 18.185
R1133 VSS.n23 VSS.t124 18.185
R1134 VSS.n66 VSS.t47 18.185
R1135 VSS.n67 VSS.t27 18.185
R1136 VSS.n26 VSS.t45 18.185
R1137 VSS.n50 VSS.t50 18.185
R1138 VSS.n51 VSS.t64 18.185
R1139 VSS.n38 VSS.t159 18.185
R1140 VSS.n37 VSS.t21 18.185
R1141 VSS.n39 VSS.t152 18.185
R1142 VSS.n152 VSS.t154 18.089
R1143 VSS.n93 VSS.t120 17.929
R1144 VSS.n80 VSS.t56 17.929
R1145 VSS.n59 VSS.t67 17.929
R1146 VSS.n46 VSS.t19 17.929
R1147 VSS.n12 VSS.t65 17.925
R1148 VSS.n77 VSS.t7 17.925
R1149 VSS.n25 VSS.t16 17.925
R1150 VSS.n43 VSS.t46 17.925
R1151 VSS.n163 VSS.t18 17.888
R1152 VSS.n143 VSS.t125 17.888
R1153 VSS.n123 VSS.t78 17.888
R1154 VSS.n103 VSS.t55 17.888
R1155 VSS.n166 VSS.t2 17.884
R1156 VSS.n149 VSS.t26 17.884
R1157 VSS.n120 VSS.t90 17.884
R1158 VSS.n100 VSS.t74 17.884
R1159 VSS.n162 VSS.t42 17.4
R1160 VSS.n162 VSS.t131 17.4
R1161 VSS.n165 VSS.t89 17.4
R1162 VSS.n165 VSS.t115 17.4
R1163 VSS.n142 VSS.t113 17.4
R1164 VSS.n142 VSS.t133 17.4
R1165 VSS.n148 VSS.t111 17.4
R1166 VSS.n148 VSS.t53 17.4
R1167 VSS.n122 VSS.t15 17.4
R1168 VSS.n122 VSS.t128 17.4
R1169 VSS.n119 VSS.t91 17.4
R1170 VSS.n119 VSS.t58 17.4
R1171 VSS.n102 VSS.t1 17.4
R1172 VSS.n102 VSS.t88 17.4
R1173 VSS.n99 VSS.t68 17.4
R1174 VSS.n99 VSS.t97 17.4
R1175 VSS.n92 VSS.t75 17.4
R1176 VSS.n92 VSS.t23 17.4
R1177 VSS.n11 VSS.t22 17.4
R1178 VSS.n11 VSS.t135 17.4
R1179 VSS.n79 VSS.t142 17.4
R1180 VSS.n79 VSS.t150 17.4
R1181 VSS.n76 VSS.t3 17.4
R1182 VSS.n76 VSS.t130 17.4
R1183 VSS.n58 VSS.t158 17.4
R1184 VSS.n58 VSS.t5 17.4
R1185 VSS.n24 VSS.t79 17.4
R1186 VSS.n24 VSS.t66 17.4
R1187 VSS.n42 VSS.t12 17.4
R1188 VSS.n42 VSS.t51 17.4
R1189 VSS.n45 VSS.t70 17.4
R1190 VSS.n45 VSS.t57 17.4
R1191 VSS.n134 VSS.t31 9.487
R1192 VSS.n169 VSS.t34 9.487
R1193 VSS.n168 VSS.t32 9.487
R1194 VSS.n138 VSS.t84 9.487
R1195 VSS.n151 VSS.t77 9.487
R1196 VSS.n3 VSS.t80 9.487
R1197 VSS.n5 VSS.t73 9.487
R1198 VSS.n4 VSS.t139 9.487
R1199 VSS.n106 VSS.t102 9.487
R1200 VSS.n105 VSS.t92 9.487
R1201 VSS.n101 VSS.t93 9.487
R1202 VSS.n13 VSS.t36 9.487
R1203 VSS.n84 VSS.t146 9.487
R1204 VSS.n85 VSS.t38 9.487
R1205 VSS.n23 VSS.t29 9.487
R1206 VSS.n66 VSS.t140 9.487
R1207 VSS.n67 VSS.t127 9.487
R1208 VSS.n26 VSS.t76 9.487
R1209 VSS.n50 VSS.t11 9.487
R1210 VSS.n51 VSS.t6 9.487
R1211 VSS.n38 VSS.t155 9.487
R1212 VSS.n37 VSS.t100 9.487
R1213 VSS.n39 VSS.t156 9.487
R1214 VSS.n152 VSS.t59 9.46
R1215 VSS.n155 VSS.t71 8.7
R1216 VSS.n155 VSS.t20 8.7
R1217 VSS.n135 VSS.t108 8.7
R1218 VSS.n135 VSS.t112 8.7
R1219 VSS.n144 VSS.t35 8.7
R1220 VSS.n144 VSS.t83 8.7
R1221 VSS.n139 VSS.t147 8.7
R1222 VSS.n139 VSS.t126 8.7
R1223 VSS.n126 VSS.t129 8.7
R1224 VSS.n126 VSS.t85 8.7
R1225 VSS.n0 VSS.t49 8.7
R1226 VSS.n0 VSS.t25 8.7
R1227 VSS.n107 VSS.t103 8.7
R1228 VSS.n107 VSS.t117 8.7
R1229 VSS.n110 VSS.t10 8.7
R1230 VSS.n110 VSS.t39 8.7
R1231 VSS.n6 VSS.t41 8.7
R1232 VSS.n6 VSS.t109 8.7
R1233 VSS.n87 VSS.t138 8.7
R1234 VSS.n87 VSS.t148 8.7
R1235 VSS.n69 VSS.t95 8.7
R1236 VSS.n69 VSS.t8 8.7
R1237 VSS.n18 VSS.t123 8.7
R1238 VSS.n18 VSS.t145 8.7
R1239 VSS.n62 VSS.t106 8.7
R1240 VSS.n62 VSS.t101 8.7
R1241 VSS.n53 VSS.t121 8.7
R1242 VSS.n53 VSS.t119 8.7
R1243 VSS.n33 VSS.t118 8.7
R1244 VSS.n33 VSS.t114 8.7
R1245 VSS.n28 VSS.t81 8.7
R1246 VSS.n28 VSS.t86 8.7
R1247 VSS.n156 VSS.n155 0.948
R1248 VSS.n136 VSS.n135 0.948
R1249 VSS.n145 VSS.n144 0.948
R1250 VSS.n140 VSS.n139 0.948
R1251 VSS.n127 VSS.n126 0.948
R1252 VSS.n1 VSS.n0 0.948
R1253 VSS.n108 VSS.n107 0.948
R1254 VSS.n111 VSS.n110 0.948
R1255 VSS.n7 VSS.n6 0.948
R1256 VSS.n88 VSS.n87 0.948
R1257 VSS.n70 VSS.n69 0.948
R1258 VSS.n19 VSS.n18 0.948
R1259 VSS.n63 VSS.n62 0.948
R1260 VSS.n54 VSS.n53 0.948
R1261 VSS.n34 VSS.n33 0.948
R1262 VSS.n29 VSS.n28 0.948
R1263 VSS.n163 VSS.n162 0.72
R1264 VSS.n166 VSS.n165 0.72
R1265 VSS.n143 VSS.n142 0.72
R1266 VSS.n149 VSS.n148 0.72
R1267 VSS.n123 VSS.n122 0.72
R1268 VSS.n120 VSS.n119 0.72
R1269 VSS.n103 VSS.n102 0.72
R1270 VSS.n100 VSS.n99 0.72
R1271 VSS.n93 VSS.n92 0.72
R1272 VSS.n12 VSS.n11 0.72
R1273 VSS.n80 VSS.n79 0.72
R1274 VSS.n77 VSS.n76 0.72
R1275 VSS.n59 VSS.n58 0.72
R1276 VSS.n25 VSS.n24 0.72
R1277 VSS.n43 VSS.n42 0.72
R1278 VSS.n46 VSS.n45 0.72
R1279 VSS.n153 VSS.n152 0.239
R1280 VSS.n49 VSS.n48 0.205
R1281 VSS.n49 VSS.n31 0.189
R1282 VSS.n147 VSS.n146 0.151
R1283 VSS.n98 VSS.n97 0.149
R1284 VSS.n90 VSS.n89 0.148
R1285 VSS.n56 VSS.n55 0.148
R1286 VSS.n160 VSS.n157 0.146
R1287 VSS.n167 VSS.n137 0.146
R1288 VSS.n150 VSS.n141 0.146
R1289 VSS.n131 VSS.n128 0.146
R1290 VSS.n121 VSS.n2 0.146
R1291 VSS.n114 VSS.n109 0.146
R1292 VSS.n114 VSS.n112 0.146
R1293 VSS.n96 VSS.n8 0.146
R1294 VSS.n72 VSS.n71 0.146
R1295 VSS.n21 VSS.n20 0.146
R1296 VSS.n65 VSS.n64 0.146
R1297 VSS.n36 VSS.n35 0.146
R1298 VSS.n31 VSS.n30 0.146
R1299 VSS.n147 VSS.n143 0.143
R1300 VSS.n164 VSS.n163 0.142
R1301 VSS.n124 VSS.n123 0.142
R1302 VSS.n104 VSS.n103 0.142
R1303 VSS.n94 VSS.n93 0.142
R1304 VSS.n81 VSS.n80 0.142
R1305 VSS.n60 VSS.n59 0.142
R1306 VSS.n47 VSS.n46 0.142
R1307 VSS.n167 VSS.n166 0.138
R1308 VSS.n150 VSS.n149 0.138
R1309 VSS.n121 VSS.n120 0.138
R1310 VSS.n104 VSS.n100 0.138
R1311 VSS.n91 VSS.n12 0.138
R1312 VSS.n78 VSS.n77 0.138
R1313 VSS.n57 VSS.n25 0.138
R1314 VSS.n44 VSS.n43 0.138
R1315 VSS.n171 VSS.n133 0.135
R1316 VSS.n117 VSS.n116 0.131
R1317 VSS.n157 VSS.n156 0.125
R1318 VSS.n137 VSS.n136 0.125
R1319 VSS.n146 VSS.n145 0.125
R1320 VSS.n141 VSS.n140 0.125
R1321 VSS.n128 VSS.n127 0.125
R1322 VSS.n2 VSS.n1 0.125
R1323 VSS.n109 VSS.n108 0.125
R1324 VSS.n112 VSS.n111 0.125
R1325 VSS.n8 VSS.n7 0.125
R1326 VSS.n89 VSS.n88 0.125
R1327 VSS.n71 VSS.n70 0.125
R1328 VSS.n20 VSS.n19 0.125
R1329 VSS.n64 VSS.n63 0.125
R1330 VSS.n55 VSS.n54 0.125
R1331 VSS.n35 VSS.n34 0.125
R1332 VSS.n30 VSS.n29 0.125
R1333 VSS.n116 VSS.n98 0.083
R1334 VSS.n68 VSS.n65 0.076
R1335 VSS.n154 VSS.n153 0.076
R1336 VSS.n86 VSS.n83 0.075
R1337 VSS VSS.n133 0.063
R1338 VSS VSS.n171 0.037
R1339 VSS.n170 VSS.n134 0.022
R1340 VSS.n153 VSS.n138 0.022
R1341 VSS.n118 VSS.n3 0.022
R1342 VSS.n104 VSS.n101 0.019
R1343 VSS.n159 VSS.n158 0.018
R1344 VSS.n130 VSS.n129 0.018
R1345 VSS.n10 VSS.n9 0.018
R1346 VSS.n170 VSS.n168 0.018
R1347 VSS.n153 VSS.n151 0.018
R1348 VSS.n118 VSS.n4 0.018
R1349 VSS.n114 VSS.n106 0.018
R1350 VSS.n170 VSS.n169 0.018
R1351 VSS.n118 VSS.n5 0.018
R1352 VSS.n115 VSS.n105 0.018
R1353 VSS.n40 VSS.n39 0.017
R1354 VSS.n86 VSS.n13 0.015
R1355 VSS.n86 VSS.n84 0.015
R1356 VSS.n86 VSS.n85 0.015
R1357 VSS.n68 VSS.n23 0.015
R1358 VSS.n68 VSS.n66 0.015
R1359 VSS.n68 VSS.n67 0.015
R1360 VSS.n52 VSS.n26 0.015
R1361 VSS.n52 VSS.n50 0.015
R1362 VSS.n52 VSS.n51 0.015
R1363 VSS.n40 VSS.n38 0.015
R1364 VSS.n40 VSS.n37 0.015
R1365 VSS.n160 VSS.n159 0.01
R1366 VSS.n131 VSS.n130 0.01
R1367 VSS.n96 VSS.n10 0.01
R1368 VSS.n15 VSS.n14 0.009
R1369 VSS.n115 VSS.n114 0.009
R1370 VSS.n41 VSS.n40 0.009
R1371 VSS.n116 VSS.n104 0.009
R1372 VSS.n31 VSS.n27 0.007
R1373 VSS.n153 VSS.n150 0.007
R1374 VSS.n170 VSS.n167 0.007
R1375 VSS.n57 VSS.n52 0.007
R1376 VSS.n78 VSS.n68 0.007
R1377 VSS.n91 VSS.n86 0.007
R1378 VSS.n121 VSS.n118 0.007
R1379 VSS.n150 VSS.n147 0.005
R1380 VSS.n167 VSS.n164 0.005
R1381 VSS.n47 VSS.n44 0.005
R1382 VSS.n60 VSS.n57 0.005
R1383 VSS.n81 VSS.n78 0.005
R1384 VSS.n94 VSS.n91 0.005
R1385 VSS.n124 VSS.n121 0.005
R1386 VSS.n61 VSS.n60 0.004
R1387 VSS.n17 VSS.n16 0.003
R1388 VSS.n16 VSS.n15 0.003
R1389 VSS.n116 VSS.n115 0.003
R1390 VSS.n133 VSS.n132 0.002
R1391 VSS.n41 VSS.n36 0.002
R1392 VSS.n164 VSS.n161 0.002
R1393 VSS.n48 VSS.n47 0.002
R1394 VSS.n82 VSS.n81 0.002
R1395 VSS.n95 VSS.n94 0.002
R1396 VSS.n114 VSS.n113 0.002
R1397 VSS.n125 VSS.n124 0.002
R1398 VSS.n73 VSS.n72 0.001
R1399 VSS.n75 VSS.n74 0.001
R1400 VSS.n65 VSS.n61 0.001
R1401 VSS.n171 VSS.n170 0.001
R1402 VSS.n161 VSS.n160 0.001
R1403 VSS.n52 VSS.n49 0.001
R1404 VSS.n83 VSS.n82 0.001
R1405 VSS.n96 VSS.n95 0.001
R1406 VSS.n118 VSS.n117 0.001
R1407 VSS.n131 VSS.n125 0.001
R1408 VSS.n44 VSS.n41 0.001
R1409 VSS.n83 VSS.n17 0.001
R1410 VSS.n44 VSS.n32 0.001
R1411 VSS.n97 VSS.n96 0.001
R1412 VSS.n160 VSS.n154 0.001
R1413 VSS.n132 VSS.n131 0.001
R1414 VSS.n78 VSS.n75 0.001
R1415 VSS.n78 VSS.n73 0.001
R1416 VSS.n91 VSS.n90 0.001
R1417 VSS.n57 VSS.n56 0.001
R1418 VSS.n22 VSS.n21 0.001
R1419 VSS.n83 VSS.n22 0.001
R1420 A[1].n4 A[1].n3 535.449
R1421 A[1].t7 A[1].t6 437.233
R1422 A[1].t12 A[1].t1 437.233
R1423 A[1].t11 A[1].n1 313.873
R1424 A[1].n3 A[1].t8 294.986
R1425 A[1].n0 A[1].t10 272.288
R1426 A[1].n4 A[1].t2 245.184
R1427 A[1].n6 A[1].t12 218.628
R1428 A[1].n8 A[1].t7 217.024
R1429 A[1].n7 A[1].t9 214.686
R1430 A[1].t6 A[1].n7 214.686
R1431 A[1].n5 A[1].t15 214.686
R1432 A[1].t1 A[1].n5 214.686
R1433 A[1].n2 A[1].t11 190.152
R1434 A[1].n2 A[1].t14 190.152
R1435 A[1].n0 A[1].t5 160.666
R1436 A[1].n1 A[1].t3 160.666
R1437 A[1].n3 A[1].t0 110.859
R1438 A[1].n1 A[1].n0 96.129
R1439 A[1].n7 A[1].t13 80.333
R1440 A[1].t2 A[1].n2 80.333
R1441 A[1].n5 A[1].t4 80.333
R1442 A[1].n6 A[1].n4 14.9
R1443 A[1].n8 A[1].n6 2.599
R1444 A[1] A[1].n8 0.288
R1445 a_52_n3507.n6 a_52_n3507.n5 501.28
R1446 a_52_n3507.t5 a_52_n3507.t6 437.233
R1447 a_52_n3507.t4 a_52_n3507.t16 415.315
R1448 a_52_n3507.t19 a_52_n3507.n3 313.873
R1449 a_52_n3507.n5 a_52_n3507.t17 294.986
R1450 a_52_n3507.n2 a_52_n3507.t18 272.288
R1451 a_52_n3507.n6 a_52_n3507.t12 236.009
R1452 a_52_n3507.n9 a_52_n3507.t5 216.627
R1453 a_52_n3507.n7 a_52_n3507.t4 216.111
R1454 a_52_n3507.n8 a_52_n3507.t7 214.686
R1455 a_52_n3507.t6 a_52_n3507.n8 214.686
R1456 a_52_n3507.n1 a_52_n3507.t13 214.335
R1457 a_52_n3507.t16 a_52_n3507.n1 214.335
R1458 a_52_n3507.n4 a_52_n3507.t11 190.152
R1459 a_52_n3507.n4 a_52_n3507.t19 190.152
R1460 a_52_n3507.n2 a_52_n3507.t15 160.666
R1461 a_52_n3507.n3 a_52_n3507.t9 160.666
R1462 a_52_n3507.n7 a_52_n3507.n6 148.428
R1463 a_52_n3507.n5 a_52_n3507.t10 110.859
R1464 a_52_n3507.n3 a_52_n3507.n2 96.129
R1465 a_52_n3507.n8 a_52_n3507.t8 80.333
R1466 a_52_n3507.n1 a_52_n3507.t14 80.333
R1467 a_52_n3507.t12 a_52_n3507.n4 80.333
R1468 a_52_n3507.n0 a_52_n3507.t1 28.57
R1469 a_52_n3507.n11 a_52_n3507.t2 28.565
R1470 a_52_n3507.t3 a_52_n3507.n11 28.565
R1471 a_52_n3507.n0 a_52_n3507.t0 17.638
R1472 a_52_n3507.n10 a_52_n3507.n9 5.638
R1473 a_52_n3507.n9 a_52_n3507.n7 2.923
R1474 a_52_n3507.n11 a_52_n3507.n10 0.693
R1475 a_52_n3507.n10 a_52_n3507.n0 0.597
R1476 carry_in.n5 carry_in.n4 501.28
R1477 carry_in.t10 carry_in.t7 437.233
R1478 carry_in.t5 carry_in.t14 415.315
R1479 carry_in.t0 carry_in.n2 313.873
R1480 carry_in.n4 carry_in.t13 294.986
R1481 carry_in.n1 carry_in.t6 272.288
R1482 carry_in.n5 carry_in.t11 236.01
R1483 carry_in.n8 carry_in.t10 216.627
R1484 carry_in.n6 carry_in.t5 216.111
R1485 carry_in.n7 carry_in.t9 214.686
R1486 carry_in.t7 carry_in.n7 214.686
R1487 carry_in.n0 carry_in.t15 214.335
R1488 carry_in.t14 carry_in.n0 214.335
R1489 carry_in.n3 carry_in.t0 190.152
R1490 carry_in.n3 carry_in.t2 190.152
R1491 carry_in.n1 carry_in.t8 160.666
R1492 carry_in.n2 carry_in.t3 160.666
R1493 carry_in.n6 carry_in.n5 148.428
R1494 carry_in.n4 carry_in.t1 110.859
R1495 carry_in.n2 carry_in.n1 96.129
R1496 carry_in.n7 carry_in.t12 80.333
R1497 carry_in.n0 carry_in.t4 80.333
R1498 carry_in.t11 carry_in.n3 80.333
R1499 carry_in.n8 carry_in.n6 2.923
R1500 carry_in carry_in.n8 0.735
R1501 B[4].n7 B[4].n6 861.987
R1502 B[4].n6 B[4].n5 560.726
R1503 B[4].t11 B[4].t0 415.315
R1504 B[4].t8 B[4].t6 415.315
R1505 B[4].n3 B[4].t9 394.151
R1506 B[4].n5 B[4].t10 294.653
R1507 B[4].n2 B[4].t1 269.523
R1508 B[4].t9 B[4].n2 269.523
R1509 B[4].n9 B[4].t11 217.716
R1510 B[4].n8 B[4].t14 214.335
R1511 B[4].t0 B[4].n8 214.335
R1512 B[4].n0 B[4].t4 214.335
R1513 B[4].t6 B[4].n0 214.335
R1514 B[4].n7 B[4].t8 198.921
R1515 B[4].n1 B[4].t13 198.043
R1516 B[4].n2 B[4].t3 160.666
R1517 B[4].n5 B[4].t2 111.663
R1518 B[4].n4 B[4].n3 97.816
R1519 B[4].n1 B[4].t12 93.989
R1520 B[4].n8 B[4].t7 80.333
R1521 B[4].n3 B[4].t15 80.333
R1522 B[4].n0 B[4].t5 80.333
R1523 B[4].n6 B[4].n4 65.07
R1524 B[4].n9 B[4].n7 16.411
R1525 B[4].n4 B[4].n1 6.615
R1526 B[4].n10 B[4].n9 0.433
R1527 B[4] B[4].n10 0.075
R1528 B[4].n10 B[4] 0.014
R1529 Y[7].n7 Y[7].n6 217.612
R1530 Y[7].n4 Y[7].n2 157.665
R1531 Y[7].n4 Y[7].n3 122.746
R1532 Y[7].n6 Y[7].n0 90.436
R1533 Y[7].n5 Y[7].n1 90.416
R1534 Y[7].n6 Y[7].n5 74.302
R1535 Y[7].n5 Y[7].n4 50.575
R1536 Y[7].n3 Y[7].t4 14.282
R1537 Y[7].n3 Y[7].t5 14.282
R1538 Y[7].n1 Y[7].t6 14.282
R1539 Y[7].n1 Y[7].t3 14.282
R1540 Y[7].n0 Y[7].t1 14.282
R1541 Y[7].n0 Y[7].t2 14.282
R1542 Y[7].n2 Y[7].t7 8.7
R1543 Y[7].n2 Y[7].t0 8.7
R1544 Y[7] Y[7].n7 0.04
R1545 Y[7].n7 Y[7] 0.04
R1546 a_9455_1702.n8 a_9455_1702.n6 552.333
R1547 a_9455_1702.n4 a_9455_1702.t13 394.151
R1548 a_9455_1702.n9 a_9455_1702.n8 342.688
R1549 a_9455_1702.n7 a_9455_1702.t10 294.653
R1550 a_9455_1702.n3 a_9455_1702.t15 269.523
R1551 a_9455_1702.t13 a_9455_1702.n3 269.523
R1552 a_9455_1702.n5 a_9455_1702.t14 198.043
R1553 a_9455_1702.n3 a_9455_1702.t8 160.666
R1554 a_9455_1702.n11 a_9455_1702.n0 157.665
R1555 a_9455_1702.n8 a_9455_1702.n7 126.566
R1556 a_9455_1702.n12 a_9455_1702.n11 122.999
R1557 a_9455_1702.n7 a_9455_1702.t12 111.663
R1558 a_9455_1702.n6 a_9455_1702.n4 97.816
R1559 a_9455_1702.n5 a_9455_1702.t11 93.989
R1560 a_9455_1702.n9 a_9455_1702.n2 90.436
R1561 a_9455_1702.n10 a_9455_1702.n1 90.416
R1562 a_9455_1702.n4 a_9455_1702.t9 80.333
R1563 a_9455_1702.n10 a_9455_1702.n9 74.302
R1564 a_9455_1702.n11 a_9455_1702.n10 50.575
R1565 a_9455_1702.n2 a_9455_1702.t5 14.282
R1566 a_9455_1702.n2 a_9455_1702.t7 14.282
R1567 a_9455_1702.n1 a_9455_1702.t6 14.282
R1568 a_9455_1702.n1 a_9455_1702.t1 14.282
R1569 a_9455_1702.n12 a_9455_1702.t0 14.282
R1570 a_9455_1702.t2 a_9455_1702.n12 14.282
R1571 a_9455_1702.n0 a_9455_1702.t4 8.7
R1572 a_9455_1702.n0 a_9455_1702.t3 8.7
R1573 a_9455_1702.n6 a_9455_1702.n5 6.615
R1574 a_11163_3955.n6 a_11163_3955.n5 501.28
R1575 a_11163_3955.t16 a_11163_3955.t6 437.233
R1576 a_11163_3955.t7 a_11163_3955.t10 415.315
R1577 a_11163_3955.t18 a_11163_3955.n3 313.873
R1578 a_11163_3955.n5 a_11163_3955.t15 294.986
R1579 a_11163_3955.n2 a_11163_3955.t5 272.288
R1580 a_11163_3955.n6 a_11163_3955.t8 236.01
R1581 a_11163_3955.n9 a_11163_3955.t16 216.627
R1582 a_11163_3955.n7 a_11163_3955.t7 216.111
R1583 a_11163_3955.n8 a_11163_3955.t19 214.686
R1584 a_11163_3955.t6 a_11163_3955.n8 214.686
R1585 a_11163_3955.n1 a_11163_3955.t11 214.335
R1586 a_11163_3955.t10 a_11163_3955.n1 214.335
R1587 a_11163_3955.n4 a_11163_3955.t18 190.152
R1588 a_11163_3955.n4 a_11163_3955.t4 190.152
R1589 a_11163_3955.n2 a_11163_3955.t14 160.666
R1590 a_11163_3955.n3 a_11163_3955.t9 160.666
R1591 a_11163_3955.n7 a_11163_3955.n6 148.428
R1592 a_11163_3955.n5 a_11163_3955.t13 110.859
R1593 a_11163_3955.n3 a_11163_3955.n2 96.129
R1594 a_11163_3955.n8 a_11163_3955.t12 80.333
R1595 a_11163_3955.n1 a_11163_3955.t17 80.333
R1596 a_11163_3955.t8 a_11163_3955.n4 80.333
R1597 a_11163_3955.t3 a_11163_3955.n11 28.57
R1598 a_11163_3955.n0 a_11163_3955.t2 28.565
R1599 a_11163_3955.n0 a_11163_3955.t1 28.565
R1600 a_11163_3955.n11 a_11163_3955.t0 17.638
R1601 a_11163_3955.n10 a_11163_3955.n9 5.6
R1602 a_11163_3955.n9 a_11163_3955.n7 2.923
R1603 a_11163_3955.n10 a_11163_3955.n0 0.69
R1604 a_11163_3955.n11 a_11163_3955.n10 0.6
R1605 Y[3].n7 Y[3].n6 217.612
R1606 Y[3].n4 Y[3].n2 157.665
R1607 Y[3].n4 Y[3].n3 122.999
R1608 Y[3].n6 Y[3].n0 90.436
R1609 Y[3].n5 Y[3].n1 90.416
R1610 Y[3].n6 Y[3].n5 74.302
R1611 Y[3].n5 Y[3].n4 50.575
R1612 Y[3].n0 Y[3].t2 14.282
R1613 Y[3].n0 Y[3].t1 14.282
R1614 Y[3].n1 Y[3].t0 14.282
R1615 Y[3].n1 Y[3].t6 14.282
R1616 Y[3].n3 Y[3].t7 14.282
R1617 Y[3].n3 Y[3].t4 14.282
R1618 Y[3].n2 Y[3].t3 8.7
R1619 Y[3].n2 Y[3].t5 8.7
R1620 Y[3] Y[3].n7 0.04
R1621 Y[3].n7 Y[3] 0.039
R1622 a_949_n3236.n8 a_949_n3236.n6 552.333
R1623 a_949_n3236.n5 a_949_n3236.t15 394.151
R1624 a_949_n3236.n9 a_949_n3236.n8 342.688
R1625 a_949_n3236.n7 a_949_n3236.t8 294.653
R1626 a_949_n3236.n4 a_949_n3236.t9 269.523
R1627 a_949_n3236.t15 a_949_n3236.n4 269.523
R1628 a_949_n3236.n3 a_949_n3236.t13 198.043
R1629 a_949_n3236.n4 a_949_n3236.t14 160.666
R1630 a_949_n3236.n11 a_949_n3236.n0 157.665
R1631 a_949_n3236.n8 a_949_n3236.n7 126.566
R1632 a_949_n3236.n12 a_949_n3236.n11 122.747
R1633 a_949_n3236.n7 a_949_n3236.t12 111.663
R1634 a_949_n3236.n6 a_949_n3236.n5 97.816
R1635 a_949_n3236.n3 a_949_n3236.t11 93.989
R1636 a_949_n3236.n9 a_949_n3236.n2 90.436
R1637 a_949_n3236.n10 a_949_n3236.n1 90.416
R1638 a_949_n3236.n5 a_949_n3236.t10 80.333
R1639 a_949_n3236.n10 a_949_n3236.n9 74.302
R1640 a_949_n3236.n11 a_949_n3236.n10 50.575
R1641 a_949_n3236.n1 a_949_n3236.t0 14.282
R1642 a_949_n3236.n1 a_949_n3236.t5 14.282
R1643 a_949_n3236.n2 a_949_n3236.t6 14.282
R1644 a_949_n3236.n2 a_949_n3236.t7 14.282
R1645 a_949_n3236.n12 a_949_n3236.t1 14.282
R1646 a_949_n3236.t2 a_949_n3236.n12 14.282
R1647 a_949_n3236.n0 a_949_n3236.t3 8.7
R1648 a_949_n3236.n0 a_949_n3236.t4 8.7
R1649 a_949_n3236.n6 a_949_n3236.n3 6.615
R1650 B[5].n7 B[5].n6 861.987
R1651 B[5].n6 B[5].n5 560.726
R1652 B[5].t0 B[5].t15 415.315
R1653 B[5].t1 B[5].t2 415.315
R1654 B[5].n3 B[5].t11 394.151
R1655 B[5].n5 B[5].t6 294.653
R1656 B[5].n2 B[5].t12 269.523
R1657 B[5].t11 B[5].n2 269.523
R1658 B[5].n9 B[5].t0 217.716
R1659 B[5].n8 B[5].t9 214.335
R1660 B[5].t15 B[5].n8 214.335
R1661 B[5].n0 B[5].t13 214.335
R1662 B[5].t2 B[5].n0 214.335
R1663 B[5].n7 B[5].t1 198.921
R1664 B[5].n1 B[5].t8 198.043
R1665 B[5].n2 B[5].t10 160.666
R1666 B[5].n5 B[5].t7 111.663
R1667 B[5].n4 B[5].n3 97.816
R1668 B[5].n1 B[5].t5 93.989
R1669 B[5].n8 B[5].t3 80.333
R1670 B[5].n3 B[5].t4 80.333
R1671 B[5].n0 B[5].t14 80.333
R1672 B[5].n6 B[5].n4 65.07
R1673 B[5].n9 B[5].n7 16.411
R1674 B[5].n4 B[5].n1 6.615
R1675 B[5].n10 B[5].n9 0.433
R1676 B[5] B[5].n10 0.077
R1677 B[5].n10 B[5] 0.011
R1678 a_7507_n3240.n8 a_7507_n3240.n6 552.333
R1679 a_7507_n3240.n5 a_7507_n3240.t12 394.151
R1680 a_7507_n3240.n9 a_7507_n3240.n8 342.688
R1681 a_7507_n3240.n7 a_7507_n3240.t14 294.653
R1682 a_7507_n3240.n4 a_7507_n3240.t10 269.523
R1683 a_7507_n3240.t12 a_7507_n3240.n4 269.523
R1684 a_7507_n3240.n3 a_7507_n3240.t9 198.043
R1685 a_7507_n3240.n4 a_7507_n3240.t11 160.666
R1686 a_7507_n3240.n11 a_7507_n3240.n0 157.665
R1687 a_7507_n3240.n8 a_7507_n3240.n7 126.566
R1688 a_7507_n3240.n12 a_7507_n3240.n11 122.747
R1689 a_7507_n3240.n7 a_7507_n3240.t15 111.663
R1690 a_7507_n3240.n6 a_7507_n3240.n5 97.816
R1691 a_7507_n3240.n3 a_7507_n3240.t8 93.989
R1692 a_7507_n3240.n9 a_7507_n3240.n2 90.436
R1693 a_7507_n3240.n10 a_7507_n3240.n1 90.416
R1694 a_7507_n3240.n5 a_7507_n3240.t13 80.333
R1695 a_7507_n3240.n10 a_7507_n3240.n9 74.302
R1696 a_7507_n3240.n11 a_7507_n3240.n10 50.575
R1697 a_7507_n3240.n1 a_7507_n3240.t1 14.282
R1698 a_7507_n3240.n1 a_7507_n3240.t5 14.282
R1699 a_7507_n3240.n2 a_7507_n3240.t6 14.282
R1700 a_7507_n3240.n2 a_7507_n3240.t7 14.282
R1701 a_7507_n3240.t2 a_7507_n3240.n12 14.282
R1702 a_7507_n3240.n12 a_7507_n3240.t0 14.282
R1703 a_7507_n3240.n0 a_7507_n3240.t3 8.7
R1704 a_7507_n3240.n0 a_7507_n3240.t4 8.7
R1705 a_7507_n3240.n6 a_7507_n3240.n3 6.615
R1706 a_4650_3958.n6 a_4650_3958.n5 501.28
R1707 a_4650_3958.t4 a_4650_3958.t19 437.233
R1708 a_4650_3958.t15 a_4650_3958.t16 415.315
R1709 a_4650_3958.t9 a_4650_3958.n3 313.873
R1710 a_4650_3958.n5 a_4650_3958.t5 294.986
R1711 a_4650_3958.n2 a_4650_3958.t7 272.288
R1712 a_4650_3958.n6 a_4650_3958.t17 236.01
R1713 a_4650_3958.n9 a_4650_3958.t4 216.627
R1714 a_4650_3958.n7 a_4650_3958.t15 216.111
R1715 a_4650_3958.n8 a_4650_3958.t14 214.686
R1716 a_4650_3958.t19 a_4650_3958.n8 214.686
R1717 a_4650_3958.n1 a_4650_3958.t6 214.335
R1718 a_4650_3958.t16 a_4650_3958.n1 214.335
R1719 a_4650_3958.n4 a_4650_3958.t9 190.152
R1720 a_4650_3958.n4 a_4650_3958.t12 190.152
R1721 a_4650_3958.n2 a_4650_3958.t18 160.666
R1722 a_4650_3958.n3 a_4650_3958.t13 160.666
R1723 a_4650_3958.n7 a_4650_3958.n6 148.428
R1724 a_4650_3958.n5 a_4650_3958.t10 110.859
R1725 a_4650_3958.n3 a_4650_3958.n2 96.129
R1726 a_4650_3958.n8 a_4650_3958.t8 80.333
R1727 a_4650_3958.n1 a_4650_3958.t11 80.333
R1728 a_4650_3958.t17 a_4650_3958.n4 80.333
R1729 a_4650_3958.t3 a_4650_3958.n11 28.57
R1730 a_4650_3958.n0 a_4650_3958.t2 28.565
R1731 a_4650_3958.n0 a_4650_3958.t1 28.565
R1732 a_4650_3958.n11 a_4650_3958.t0 17.638
R1733 a_4650_3958.n10 a_4650_3958.n9 5.375
R1734 a_4650_3958.n9 a_4650_3958.n7 2.923
R1735 a_4650_3958.n10 a_4650_3958.n0 0.69
R1736 a_4650_3958.n11 a_4650_3958.n10 0.6
R1737 A[2].n4 A[2].n3 535.449
R1738 A[2].t9 A[2].t3 437.233
R1739 A[2].t7 A[2].t12 437.233
R1740 A[2].t5 A[2].n1 313.873
R1741 A[2].n3 A[2].t4 294.986
R1742 A[2].n0 A[2].t11 272.288
R1743 A[2].n4 A[2].t0 245.184
R1744 A[2].n6 A[2].t7 218.628
R1745 A[2].n8 A[2].t9 217.024
R1746 A[2].n7 A[2].t15 214.686
R1747 A[2].t3 A[2].n7 214.686
R1748 A[2].n5 A[2].t10 214.686
R1749 A[2].t12 A[2].n5 214.686
R1750 A[2].n2 A[2].t5 190.152
R1751 A[2].n2 A[2].t13 190.152
R1752 A[2].n0 A[2].t2 160.666
R1753 A[2].n1 A[2].t14 160.666
R1754 A[2].n3 A[2].t1 110.859
R1755 A[2].n1 A[2].n0 96.129
R1756 A[2].n7 A[2].t8 80.333
R1757 A[2].t0 A[2].n2 80.333
R1758 A[2].n5 A[2].t6 80.333
R1759 A[2].n6 A[2].n4 14.9
R1760 A[2].n8 A[2].n6 2.599
R1761 A[2] A[2].n8 0.287
R1762 a_2942_1705.n8 a_2942_1705.n6 552.333
R1763 a_2942_1705.n4 a_2942_1705.t8 394.151
R1764 a_2942_1705.n9 a_2942_1705.n8 342.688
R1765 a_2942_1705.n7 a_2942_1705.t15 294.653
R1766 a_2942_1705.n3 a_2942_1705.t13 269.523
R1767 a_2942_1705.t8 a_2942_1705.n3 269.523
R1768 a_2942_1705.n5 a_2942_1705.t11 198.043
R1769 a_2942_1705.n3 a_2942_1705.t12 160.666
R1770 a_2942_1705.n11 a_2942_1705.n0 157.665
R1771 a_2942_1705.n8 a_2942_1705.n7 126.566
R1772 a_2942_1705.n12 a_2942_1705.n11 122.999
R1773 a_2942_1705.n7 a_2942_1705.t9 111.663
R1774 a_2942_1705.n6 a_2942_1705.n4 97.816
R1775 a_2942_1705.n5 a_2942_1705.t10 93.989
R1776 a_2942_1705.n9 a_2942_1705.n2 90.436
R1777 a_2942_1705.n10 a_2942_1705.n1 90.416
R1778 a_2942_1705.n4 a_2942_1705.t14 80.333
R1779 a_2942_1705.n10 a_2942_1705.n9 74.302
R1780 a_2942_1705.n11 a_2942_1705.n10 50.575
R1781 a_2942_1705.n2 a_2942_1705.t4 14.282
R1782 a_2942_1705.n2 a_2942_1705.t6 14.282
R1783 a_2942_1705.n1 a_2942_1705.t5 14.282
R1784 a_2942_1705.n1 a_2942_1705.t0 14.282
R1785 a_2942_1705.t2 a_2942_1705.n12 14.282
R1786 a_2942_1705.n12 a_2942_1705.t1 14.282
R1787 a_2942_1705.n0 a_2942_1705.t7 8.7
R1788 a_2942_1705.n0 a_2942_1705.t3 8.7
R1789 a_2942_1705.n6 a_2942_1705.n5 6.615
R1790 B[2].n7 B[2].n6 861.987
R1791 B[2].n6 B[2].n5 560.726
R1792 B[2].t14 B[2].t9 415.315
R1793 B[2].t8 B[2].t15 415.315
R1794 B[2].n2 B[2].t10 394.151
R1795 B[2].n5 B[2].t7 294.653
R1796 B[2].n1 B[2].t1 269.523
R1797 B[2].t10 B[2].n1 269.523
R1798 B[2].n9 B[2].t14 217.716
R1799 B[2].n8 B[2].t11 214.335
R1800 B[2].t9 B[2].n8 214.335
R1801 B[2].n0 B[2].t13 214.335
R1802 B[2].t15 B[2].n0 214.335
R1803 B[2].n7 B[2].t8 198.921
R1804 B[2].n3 B[2].t0 198.043
R1805 B[2].n1 B[2].t6 160.666
R1806 B[2].n5 B[2].t5 111.663
R1807 B[2].n4 B[2].n2 97.816
R1808 B[2].n3 B[2].t12 93.989
R1809 B[2].n8 B[2].t3 80.333
R1810 B[2].n2 B[2].t2 80.333
R1811 B[2].n0 B[2].t4 80.333
R1812 B[2].n6 B[2].n4 65.07
R1813 B[2].n9 B[2].n7 16.411
R1814 B[2].n4 B[2].n3 6.615
R1815 B[2] B[2].n9 0.454
R1816 A[7].n4 A[7].n3 535.449
R1817 A[7].t10 A[7].t4 437.233
R1818 A[7].t5 A[7].t2 437.233
R1819 A[7].t12 A[7].n1 313.873
R1820 A[7].n3 A[7].t8 294.986
R1821 A[7].n0 A[7].t13 272.288
R1822 A[7].n4 A[7].t11 245.184
R1823 A[7].n6 A[7].t5 218.627
R1824 A[7].n8 A[7].t10 217.023
R1825 A[7].n7 A[7].t15 214.686
R1826 A[7].t4 A[7].n7 214.686
R1827 A[7].n5 A[7].t6 214.686
R1828 A[7].t2 A[7].n5 214.686
R1829 A[7].n2 A[7].t3 190.152
R1830 A[7].n2 A[7].t12 190.152
R1831 A[7].n0 A[7].t7 160.666
R1832 A[7].n1 A[7].t0 160.666
R1833 A[7].n3 A[7].t1 110.859
R1834 A[7].n1 A[7].n0 96.129
R1835 A[7].n7 A[7].t14 80.333
R1836 A[7].t11 A[7].n2 80.333
R1837 A[7].n5 A[7].t9 80.333
R1838 A[7].n6 A[7].n4 14.9
R1839 A[7].n8 A[7].n6 2.599
R1840 A[7].n9 A[7].n8 0.224
R1841 A[7] A[7].n9 0.08
R1842 A[7].n9 A[7] 0.009
R1843 A[4].n4 A[4].n3 535.449
R1844 A[4].t15 A[4].t6 437.233
R1845 A[4].t8 A[4].t11 437.233
R1846 A[4].t2 A[4].n1 313.873
R1847 A[4].n3 A[4].t10 294.986
R1848 A[4].n0 A[4].t5 272.288
R1849 A[4].n4 A[4].t1 245.184
R1850 A[4].n6 A[4].t8 218.627
R1851 A[4].n8 A[4].t15 217.023
R1852 A[4].n7 A[4].t9 214.686
R1853 A[4].t6 A[4].n7 214.686
R1854 A[4].n5 A[4].t13 214.686
R1855 A[4].t11 A[4].n5 214.686
R1856 A[4].n2 A[4].t0 190.152
R1857 A[4].n2 A[4].t2 190.152
R1858 A[4].n0 A[4].t3 160.666
R1859 A[4].n1 A[4].t7 160.666
R1860 A[4].n3 A[4].t14 110.859
R1861 A[4].n1 A[4].n0 96.129
R1862 A[4].n7 A[4].t4 80.333
R1863 A[4].t1 A[4].n2 80.333
R1864 A[4].n5 A[4].t12 80.333
R1865 A[4].n6 A[4].n4 14.9
R1866 A[4].n8 A[4].n6 2.599
R1867 A[4].n9 A[4].n8 0.224
R1868 A[4] A[4].n9 0.081
R1869 A[4].n9 A[4] 0.008
R1870 B[6].n7 B[6].n6 861.987
R1871 B[6].n6 B[6].n5 560.726
R1872 B[6].t13 B[6].t0 415.315
R1873 B[6].t10 B[6].t8 415.315
R1874 B[6].n3 B[6].t6 394.151
R1875 B[6].n5 B[6].t9 294.653
R1876 B[6].n2 B[6].t3 269.523
R1877 B[6].t6 B[6].n2 269.523
R1878 B[6].n9 B[6].t13 217.716
R1879 B[6].n8 B[6].t15 214.335
R1880 B[6].t0 B[6].n8 214.335
R1881 B[6].n0 B[6].t4 214.335
R1882 B[6].t8 B[6].n0 214.335
R1883 B[6].n7 B[6].t10 198.921
R1884 B[6].n1 B[6].t2 198.043
R1885 B[6].n2 B[6].t5 160.666
R1886 B[6].n5 B[6].t14 111.663
R1887 B[6].n4 B[6].n3 97.816
R1888 B[6].n1 B[6].t1 93.989
R1889 B[6].n8 B[6].t12 80.333
R1890 B[6].n3 B[6].t11 80.333
R1891 B[6].n0 B[6].t7 80.333
R1892 B[6].n6 B[6].n4 65.07
R1893 B[6].n9 B[6].n7 16.411
R1894 B[6].n4 B[6].n1 6.615
R1895 B[6].n10 B[6].n9 0.433
R1896 B[6] B[6].n10 0.08
R1897 B[6].n10 B[6] 0.009
R1898 Y[6].n7 Y[6].n6 217.612
R1899 Y[6].n4 Y[6].n2 157.665
R1900 Y[6].n4 Y[6].n3 122.746
R1901 Y[6].n6 Y[6].n0 90.436
R1902 Y[6].n5 Y[6].n1 90.416
R1903 Y[6].n6 Y[6].n5 74.302
R1904 Y[6].n5 Y[6].n4 50.575
R1905 Y[6].n3 Y[6].t4 14.282
R1906 Y[6].n3 Y[6].t5 14.282
R1907 Y[6].n1 Y[6].t6 14.282
R1908 Y[6].n1 Y[6].t1 14.282
R1909 Y[6].n0 Y[6].t2 14.282
R1910 Y[6].n0 Y[6].t0 14.282
R1911 Y[6].n2 Y[6].t7 8.7
R1912 Y[6].n2 Y[6].t3 8.7
R1913 Y[6] Y[6].n7 0.04
R1914 Y[6].n7 Y[6] 0.04
R1915 B[7].n7 B[7].n6 861.987
R1916 B[7].n6 B[7].n5 560.726
R1917 B[7].t14 B[7].t2 415.315
R1918 B[7].t15 B[7].t1 415.315
R1919 B[7].n3 B[7].t8 394.151
R1920 B[7].n5 B[7].t12 294.653
R1921 B[7].n2 B[7].t9 269.523
R1922 B[7].t8 B[7].n2 269.523
R1923 B[7].n9 B[7].t14 217.716
R1924 B[7].n8 B[7].t11 214.335
R1925 B[7].t2 B[7].n8 214.335
R1926 B[7].n0 B[7].t13 214.335
R1927 B[7].t1 B[7].n0 214.335
R1928 B[7].n7 B[7].t15 198.921
R1929 B[7].n1 B[7].t7 198.043
R1930 B[7].n2 B[7].t10 160.666
R1931 B[7].n5 B[7].t6 111.663
R1932 B[7].n4 B[7].n3 97.816
R1933 B[7].n1 B[7].t5 93.989
R1934 B[7].n8 B[7].t4 80.333
R1935 B[7].n3 B[7].t3 80.333
R1936 B[7].n0 B[7].t0 80.333
R1937 B[7].n6 B[7].n4 65.07
R1938 B[7].n9 B[7].n7 16.411
R1939 B[7].n4 B[7].n1 6.615
R1940 B[7].n10 B[7].n9 0.433
R1941 B[7] B[7].n10 0.077
R1942 B[7].n10 B[7] 0.012
R1943 A[3].n4 A[3].n3 535.449
R1944 A[3].t3 A[3].t2 437.233
R1945 A[3].t13 A[3].t10 437.233
R1946 A[3].t15 A[3].n1 313.873
R1947 A[3].n3 A[3].t6 294.986
R1948 A[3].n0 A[3].t9 272.288
R1949 A[3].n4 A[3].t4 245.184
R1950 A[3].n6 A[3].t13 218.628
R1951 A[3].n8 A[3].t3 217.024
R1952 A[3].n7 A[3].t5 214.686
R1953 A[3].t2 A[3].n7 214.686
R1954 A[3].n5 A[3].t14 214.686
R1955 A[3].t10 A[3].n5 214.686
R1956 A[3].n2 A[3].t15 190.152
R1957 A[3].n2 A[3].t11 190.152
R1958 A[3].n0 A[3].t7 160.666
R1959 A[3].n1 A[3].t1 160.666
R1960 A[3].n3 A[3].t8 110.859
R1961 A[3].n1 A[3].n0 96.129
R1962 A[3].n7 A[3].t12 80.333
R1963 A[3].t4 A[3].n2 80.333
R1964 A[3].n5 A[3].t0 80.333
R1965 A[3].n6 A[3].n4 14.9
R1966 A[3].n8 A[3].n6 2.599
R1967 A[3] A[3].n8 0.287
R1968 a_15871_1697.n3 a_15871_1697.n1 267.767
R1969 a_15871_1697.n7 a_15871_1697.t8 16.058
R1970 a_15871_1697.t2 a_15871_1697.n9 16.058
R1971 a_15871_1697.n2 a_15871_1697.t10 14.282
R1972 a_15871_1697.n2 a_15871_1697.t5 14.282
R1973 a_15871_1697.n1 a_15871_1697.t9 14.282
R1974 a_15871_1697.n1 a_15871_1697.t11 14.282
R1975 a_15871_1697.n4 a_15871_1697.t4 14.282
R1976 a_15871_1697.n4 a_15871_1697.t3 14.282
R1977 a_15871_1697.n0 a_15871_1697.t0 14.282
R1978 a_15871_1697.n0 a_15871_1697.t1 14.282
R1979 a_15871_1697.n6 a_15871_1697.t6 14.282
R1980 a_15871_1697.n6 a_15871_1697.t7 14.282
R1981 a_15871_1697.n5 a_15871_1697.n4 1.511
R1982 a_15871_1697.n9 a_15871_1697.n0 0.999
R1983 a_15871_1697.n7 a_15871_1697.n6 0.999
R1984 a_15871_1697.n5 a_15871_1697.n3 0.669
R1985 a_15871_1697.n9 a_15871_1697.n8 0.575
R1986 a_15871_1697.n8 a_15871_1697.n5 0.227
R1987 a_15871_1697.n8 a_15871_1697.n7 0.2
R1988 a_15871_1697.n3 a_15871_1697.n2 0.001
R1989 a_6610_n3511.n6 a_6610_n3511.n5 501.28
R1990 a_6610_n3511.t13 a_6610_n3511.t9 437.233
R1991 a_6610_n3511.t12 a_6610_n3511.t8 415.315
R1992 a_6610_n3511.t10 a_6610_n3511.n3 313.873
R1993 a_6610_n3511.n5 a_6610_n3511.t19 294.986
R1994 a_6610_n3511.n2 a_6610_n3511.t5 272.288
R1995 a_6610_n3511.n6 a_6610_n3511.t4 236.009
R1996 a_6610_n3511.n9 a_6610_n3511.t13 216.627
R1997 a_6610_n3511.n7 a_6610_n3511.t12 216.111
R1998 a_6610_n3511.n8 a_6610_n3511.t14 214.686
R1999 a_6610_n3511.t9 a_6610_n3511.n8 214.686
R2000 a_6610_n3511.n1 a_6610_n3511.t6 214.335
R2001 a_6610_n3511.t8 a_6610_n3511.n1 214.335
R2002 a_6610_n3511.n4 a_6610_n3511.t16 190.152
R2003 a_6610_n3511.n4 a_6610_n3511.t10 190.152
R2004 a_6610_n3511.n2 a_6610_n3511.t18 160.666
R2005 a_6610_n3511.n3 a_6610_n3511.t17 160.666
R2006 a_6610_n3511.n7 a_6610_n3511.n6 148.428
R2007 a_6610_n3511.n5 a_6610_n3511.t15 110.859
R2008 a_6610_n3511.n3 a_6610_n3511.n2 96.129
R2009 a_6610_n3511.n8 a_6610_n3511.t11 80.333
R2010 a_6610_n3511.n1 a_6610_n3511.t7 80.333
R2011 a_6610_n3511.t4 a_6610_n3511.n4 80.333
R2012 a_6610_n3511.n0 a_6610_n3511.t1 28.57
R2013 a_6610_n3511.n11 a_6610_n3511.t2 28.565
R2014 a_6610_n3511.t3 a_6610_n3511.n11 28.565
R2015 a_6610_n3511.n0 a_6610_n3511.t0 17.638
R2016 a_6610_n3511.n10 a_6610_n3511.n9 5.589
R2017 a_6610_n3511.n9 a_6610_n3511.n7 2.923
R2018 a_6610_n3511.n11 a_6610_n3511.n10 0.693
R2019 a_6610_n3511.n10 a_6610_n3511.n0 0.597
R2020 a_17697_3950.n6 a_17697_3950.n5 501.28
R2021 a_17697_3950.t16 a_17697_3950.t12 437.233
R2022 a_17697_3950.t15 a_17697_3950.t9 415.315
R2023 a_17697_3950.t6 a_17697_3950.n3 313.873
R2024 a_17697_3950.n5 a_17697_3950.t19 294.986
R2025 a_17697_3950.n2 a_17697_3950.t7 272.288
R2026 a_17697_3950.n6 a_17697_3950.t18 236.01
R2027 a_17697_3950.n9 a_17697_3950.t16 216.627
R2028 a_17697_3950.n7 a_17697_3950.t15 216.111
R2029 a_17697_3950.n8 a_17697_3950.t11 214.686
R2030 a_17697_3950.t12 a_17697_3950.n8 214.686
R2031 a_17697_3950.n1 a_17697_3950.t4 214.335
R2032 a_17697_3950.t9 a_17697_3950.n1 214.335
R2033 a_17697_3950.n4 a_17697_3950.t6 190.152
R2034 a_17697_3950.n4 a_17697_3950.t8 190.152
R2035 a_17697_3950.n2 a_17697_3950.t13 160.666
R2036 a_17697_3950.n3 a_17697_3950.t14 160.666
R2037 a_17697_3950.n7 a_17697_3950.n6 148.428
R2038 a_17697_3950.n5 a_17697_3950.t5 110.859
R2039 a_17697_3950.n3 a_17697_3950.n2 96.129
R2040 a_17697_3950.n8 a_17697_3950.t17 80.333
R2041 a_17697_3950.n1 a_17697_3950.t10 80.333
R2042 a_17697_3950.t18 a_17697_3950.n4 80.333
R2043 a_17697_3950.t3 a_17697_3950.n11 28.57
R2044 a_17697_3950.n0 a_17697_3950.t2 28.565
R2045 a_17697_3950.n0 a_17697_3950.t1 28.565
R2046 a_17697_3950.n11 a_17697_3950.t0 17.638
R2047 a_17697_3950.n10 a_17697_3950.n9 5.767
R2048 a_17697_3950.n9 a_17697_3950.n7 2.923
R2049 a_17697_3950.n10 a_17697_3950.n0 0.69
R2050 a_17697_3950.n11 a_17697_3950.n10 0.6
R2051 Y[0].n7 Y[0].n6 208.992
R2052 Y[0].n4 Y[0].n2 157.665
R2053 Y[0].n4 Y[0].n3 122.999
R2054 Y[0].n6 Y[0].n0 90.436
R2055 Y[0].n5 Y[0].n1 90.416
R2056 Y[0].n6 Y[0].n5 74.302
R2057 Y[0].n5 Y[0].n4 50.575
R2058 Y[0].n0 Y[0].t6 14.282
R2059 Y[0].n0 Y[0].t5 14.282
R2060 Y[0].n1 Y[0].t4 14.282
R2061 Y[0].n1 Y[0].t2 14.282
R2062 Y[0].n3 Y[0].t1 14.282
R2063 Y[0].n3 Y[0].t3 14.282
R2064 Y[0].n2 Y[0].t7 8.7
R2065 Y[0].n2 Y[0].t0 8.7
R2066 Y[0].n8 Y[0].n7 8.62
R2067 Y[0] Y[0].n8 0.039
R2068 Y[0].n8 Y[0] 0.038
R2069 A[6].n4 A[6].n3 535.449
R2070 A[6].t15 A[6].t10 437.233
R2071 A[6].t8 A[6].t4 437.233
R2072 A[6].t0 A[6].n1 313.873
R2073 A[6].n3 A[6].t7 294.986
R2074 A[6].n0 A[6].t13 272.288
R2075 A[6].n4 A[6].t11 245.184
R2076 A[6].n6 A[6].t8 218.627
R2077 A[6].n8 A[6].t15 217.023
R2078 A[6].n7 A[6].t14 214.686
R2079 A[6].t10 A[6].n7 214.686
R2080 A[6].n5 A[6].t6 214.686
R2081 A[6].t4 A[6].n5 214.686
R2082 A[6].n2 A[6].t9 190.152
R2083 A[6].n2 A[6].t0 190.152
R2084 A[6].n0 A[6].t12 160.666
R2085 A[6].n1 A[6].t3 160.666
R2086 A[6].n3 A[6].t2 110.859
R2087 A[6].n1 A[6].n0 96.129
R2088 A[6].n7 A[6].t1 80.333
R2089 A[6].t11 A[6].n2 80.333
R2090 A[6].n5 A[6].t5 80.333
R2091 A[6].n6 A[6].n4 14.9
R2092 A[6].n8 A[6].n6 2.599
R2093 A[6].n9 A[6].n8 0.224
R2094 A[6] A[6].n9 0.082
R2095 A[6].n9 A[6] 0.007
R2096 Y[2].n7 Y[2].n6 217.612
R2097 Y[2].n4 Y[2].n2 157.665
R2098 Y[2].n4 Y[2].n3 122.999
R2099 Y[2].n6 Y[2].n0 90.436
R2100 Y[2].n5 Y[2].n1 90.416
R2101 Y[2].n6 Y[2].n5 74.302
R2102 Y[2].n5 Y[2].n4 50.575
R2103 Y[2].n0 Y[2].t4 14.282
R2104 Y[2].n0 Y[2].t5 14.282
R2105 Y[2].n1 Y[2].t6 14.282
R2106 Y[2].n1 Y[2].t1 14.282
R2107 Y[2].n3 Y[2].t2 14.282
R2108 Y[2].n3 Y[2].t0 14.282
R2109 Y[2].n2 Y[2].t7 8.7
R2110 Y[2].n2 Y[2].t3 8.7
R2111 Y[2] Y[2].n7 0.04
R2112 Y[2].n7 Y[2] 0.039
R2113 A[0].n4 A[0].n3 535.449
R2114 A[0].t7 A[0].t5 437.233
R2115 A[0].t10 A[0].t2 437.233
R2116 A[0].t8 A[0].n1 313.873
R2117 A[0].n3 A[0].t6 294.986
R2118 A[0].n0 A[0].t13 272.288
R2119 A[0].n4 A[0].t1 245.184
R2120 A[0].n6 A[0].t10 218.628
R2121 A[0].n8 A[0].t7 217.024
R2122 A[0].n7 A[0].t3 214.686
R2123 A[0].t5 A[0].n7 214.686
R2124 A[0].n5 A[0].t0 214.686
R2125 A[0].t2 A[0].n5 214.686
R2126 A[0].n2 A[0].t8 190.152
R2127 A[0].n2 A[0].t14 190.152
R2128 A[0].n0 A[0].t4 160.666
R2129 A[0].n1 A[0].t12 160.666
R2130 A[0].n3 A[0].t9 110.859
R2131 A[0].n1 A[0].n0 96.129
R2132 A[0].n7 A[0].t15 80.333
R2133 A[0].t1 A[0].n2 80.333
R2134 A[0].n5 A[0].t11 80.333
R2135 A[0].n6 A[0].n4 14.9
R2136 A[0].n8 A[0].n6 2.599
R2137 A[0] A[0].n8 0.289
R2138 A[5].n4 A[5].n3 535.449
R2139 A[5].t7 A[5].t5 437.233
R2140 A[5].t1 A[5].t15 437.233
R2141 A[5].t13 A[5].n1 313.873
R2142 A[5].n3 A[5].t11 294.986
R2143 A[5].n0 A[5].t12 272.288
R2144 A[5].n4 A[5].t8 245.184
R2145 A[5].n6 A[5].t1 218.627
R2146 A[5].n8 A[5].t7 217.023
R2147 A[5].n7 A[5].t14 214.686
R2148 A[5].t5 A[5].n7 214.686
R2149 A[5].n5 A[5].t9 214.686
R2150 A[5].t15 A[5].n5 214.686
R2151 A[5].n2 A[5].t6 190.152
R2152 A[5].n2 A[5].t13 190.152
R2153 A[5].n0 A[5].t10 160.666
R2154 A[5].n1 A[5].t2 160.666
R2155 A[5].n3 A[5].t4 110.859
R2156 A[5].n1 A[5].n0 96.129
R2157 A[5].n7 A[5].t0 80.333
R2158 A[5].t8 A[5].n2 80.333
R2159 A[5].n5 A[5].t3 80.333
R2160 A[5].n6 A[5].n4 14.9
R2161 A[5].n8 A[5].n6 2.599
R2162 A[5].n9 A[5].n8 0.224
R2163 A[5] A[5].n9 0.082
R2164 A[5].n9 A[5] 0.007
R2165 carry_out.n1 carry_out.t1 28.57
R2166 carry_out.n0 carry_out.t3 28.565
R2167 carry_out.n0 carry_out.t2 28.565
R2168 carry_out.n1 carry_out.t0 17.638
R2169 carry_out.n3 carry_out.n2 2.059
R2170 carry_out.n2 carry_out.n0 0.693
R2171 carry_out.n2 carry_out.n1 0.597
R2172 carry_out.n3 carry_out 0.13
R2173 carry_out carry_out.n3 0.074
R2174 a_22429_1701.n8 a_22429_1701.n0 267.767
R2175 a_22429_1701.n4 a_22429_1701.t4 16.058
R2176 a_22429_1701.n2 a_22429_1701.t9 16.058
R2177 a_22429_1701.n3 a_22429_1701.t3 14.282
R2178 a_22429_1701.n3 a_22429_1701.t5 14.282
R2179 a_22429_1701.n1 a_22429_1701.t10 14.282
R2180 a_22429_1701.n1 a_22429_1701.t11 14.282
R2181 a_22429_1701.n6 a_22429_1701.t1 14.282
R2182 a_22429_1701.n6 a_22429_1701.t0 14.282
R2183 a_22429_1701.n0 a_22429_1701.t8 14.282
R2184 a_22429_1701.n0 a_22429_1701.t7 14.282
R2185 a_22429_1701.n9 a_22429_1701.t6 14.282
R2186 a_22429_1701.t2 a_22429_1701.n9 14.282
R2187 a_22429_1701.n7 a_22429_1701.n6 1.511
R2188 a_22429_1701.n4 a_22429_1701.n3 0.999
R2189 a_22429_1701.n2 a_22429_1701.n1 0.999
R2190 a_22429_1701.n8 a_22429_1701.n7 0.669
R2191 a_22429_1701.n5 a_22429_1701.n4 0.575
R2192 a_22429_1701.n7 a_22429_1701.n5 0.227
R2193 a_22429_1701.n5 a_22429_1701.n2 0.2
R2194 a_22429_1701.n9 a_22429_1701.n8 0.001
R2195 B[1].n7 B[1].n6 861.987
R2196 B[1].n6 B[1].n5 560.726
R2197 B[1].t1 B[1].t0 415.315
R2198 B[1].t7 B[1].t2 415.315
R2199 B[1].n2 B[1].t3 394.151
R2200 B[1].n5 B[1].t10 294.653
R2201 B[1].n1 B[1].t6 269.523
R2202 B[1].t3 B[1].n1 269.523
R2203 B[1].n9 B[1].t1 217.716
R2204 B[1].n8 B[1].t12 214.335
R2205 B[1].t0 B[1].n8 214.335
R2206 B[1].n0 B[1].t15 214.335
R2207 B[1].t2 B[1].n0 214.335
R2208 B[1].n7 B[1].t7 198.921
R2209 B[1].n3 B[1].t4 198.043
R2210 B[1].n1 B[1].t14 160.666
R2211 B[1].n5 B[1].t8 111.663
R2212 B[1].n4 B[1].n2 97.816
R2213 B[1].n3 B[1].t5 93.989
R2214 B[1].n8 B[1].t11 80.333
R2215 B[1].n2 B[1].t9 80.333
R2216 B[1].n0 B[1].t13 80.333
R2217 B[1].n6 B[1].n4 65.07
R2218 B[1].n9 B[1].n7 16.411
R2219 B[1].n4 B[1].n3 6.615
R2220 B[1] B[1].n9 0.456
R2221 a_13144_n3506.n6 a_13144_n3506.n5 501.28
R2222 a_13144_n3506.t5 a_13144_n3506.t6 437.233
R2223 a_13144_n3506.t4 a_13144_n3506.t19 415.315
R2224 a_13144_n3506.t14 a_13144_n3506.n3 313.873
R2225 a_13144_n3506.n5 a_13144_n3506.t11 294.986
R2226 a_13144_n3506.n2 a_13144_n3506.t16 272.288
R2227 a_13144_n3506.n6 a_13144_n3506.t13 236.009
R2228 a_13144_n3506.n9 a_13144_n3506.t5 216.627
R2229 a_13144_n3506.n7 a_13144_n3506.t4 216.111
R2230 a_13144_n3506.n8 a_13144_n3506.t8 214.686
R2231 a_13144_n3506.t6 a_13144_n3506.n8 214.686
R2232 a_13144_n3506.n1 a_13144_n3506.t17 214.335
R2233 a_13144_n3506.t19 a_13144_n3506.n1 214.335
R2234 a_13144_n3506.n4 a_13144_n3506.t12 190.152
R2235 a_13144_n3506.n4 a_13144_n3506.t14 190.152
R2236 a_13144_n3506.n2 a_13144_n3506.t15 160.666
R2237 a_13144_n3506.n3 a_13144_n3506.t9 160.666
R2238 a_13144_n3506.n7 a_13144_n3506.n6 148.428
R2239 a_13144_n3506.n5 a_13144_n3506.t10 110.859
R2240 a_13144_n3506.n3 a_13144_n3506.n2 96.129
R2241 a_13144_n3506.n8 a_13144_n3506.t7 80.333
R2242 a_13144_n3506.n1 a_13144_n3506.t18 80.333
R2243 a_13144_n3506.t13 a_13144_n3506.n4 80.333
R2244 a_13144_n3506.n0 a_13144_n3506.t1 28.57
R2245 a_13144_n3506.n11 a_13144_n3506.t2 28.565
R2246 a_13144_n3506.t3 a_13144_n3506.n11 28.565
R2247 a_13144_n3506.n0 a_13144_n3506.t0 17.638
R2248 a_13144_n3506.n10 a_13144_n3506.n9 5.55
R2249 a_13144_n3506.n9 a_13144_n3506.n7 2.923
R2250 a_13144_n3506.n11 a_13144_n3506.n10 0.693
R2251 a_13144_n3506.n10 a_13144_n3506.n0 0.597
R2252 a_15584_n3902.n3 a_15584_n3902.n1 267.767
R2253 a_15584_n3902.n7 a_15584_n3902.t9 16.058
R2254 a_15584_n3902.t2 a_15584_n3902.n9 16.058
R2255 a_15584_n3902.n2 a_15584_n3902.t6 14.282
R2256 a_15584_n3902.n2 a_15584_n3902.t3 14.282
R2257 a_15584_n3902.n1 a_15584_n3902.t4 14.282
R2258 a_15584_n3902.n1 a_15584_n3902.t5 14.282
R2259 a_15584_n3902.n4 a_15584_n3902.t7 14.282
R2260 a_15584_n3902.n4 a_15584_n3902.t8 14.282
R2261 a_15584_n3902.n0 a_15584_n3902.t0 14.282
R2262 a_15584_n3902.n0 a_15584_n3902.t1 14.282
R2263 a_15584_n3902.n6 a_15584_n3902.t10 14.282
R2264 a_15584_n3902.n6 a_15584_n3902.t11 14.282
R2265 a_15584_n3902.n5 a_15584_n3902.n4 1.511
R2266 a_15584_n3902.n9 a_15584_n3902.n0 0.999
R2267 a_15584_n3902.n7 a_15584_n3902.n6 0.999
R2268 a_15584_n3902.n5 a_15584_n3902.n3 0.669
R2269 a_15584_n3902.n8 a_15584_n3902.n7 0.575
R2270 a_15584_n3902.n8 a_15584_n3902.n5 0.227
R2271 a_15584_n3902.n9 a_15584_n3902.n8 0.2
R2272 a_15584_n3902.n3 a_15584_n3902.n2 0.001
R2273 Y[5].n7 Y[5].n6 217.612
R2274 Y[5].n4 Y[5].n2 157.665
R2275 Y[5].n4 Y[5].n3 122.746
R2276 Y[5].n6 Y[5].n0 90.436
R2277 Y[5].n5 Y[5].n1 90.416
R2278 Y[5].n6 Y[5].n5 74.302
R2279 Y[5].n5 Y[5].n4 50.575
R2280 Y[5].n3 Y[5].t3 14.282
R2281 Y[5].n3 Y[5].t4 14.282
R2282 Y[5].n1 Y[5].t2 14.282
R2283 Y[5].n1 Y[5].t5 14.282
R2284 Y[5].n0 Y[5].t6 14.282
R2285 Y[5].n0 Y[5].t7 14.282
R2286 Y[5].n2 Y[5].t1 8.7
R2287 Y[5].n2 Y[5].t0 8.7
R2288 Y[5] Y[5].n7 0.041
R2289 Y[5].n7 Y[5] 0.039
R2290 a_24327_1701.n3 a_24327_1701.n1 267.767
R2291 a_24327_1701.n7 a_24327_1701.t8 16.058
R2292 a_24327_1701.t2 a_24327_1701.n9 16.058
R2293 a_24327_1701.n2 a_24327_1701.t11 14.282
R2294 a_24327_1701.n2 a_24327_1701.t3 14.282
R2295 a_24327_1701.n1 a_24327_1701.t9 14.282
R2296 a_24327_1701.n1 a_24327_1701.t10 14.282
R2297 a_24327_1701.n4 a_24327_1701.t5 14.282
R2298 a_24327_1701.n4 a_24327_1701.t4 14.282
R2299 a_24327_1701.n6 a_24327_1701.t7 14.282
R2300 a_24327_1701.n6 a_24327_1701.t6 14.282
R2301 a_24327_1701.n0 a_24327_1701.t1 14.282
R2302 a_24327_1701.n0 a_24327_1701.t0 14.282
R2303 a_24327_1701.n5 a_24327_1701.n4 1.511
R2304 a_24327_1701.n7 a_24327_1701.n6 0.999
R2305 a_24327_1701.n9 a_24327_1701.n0 0.999
R2306 a_24327_1701.n5 a_24327_1701.n3 0.669
R2307 a_24327_1701.n8 a_24327_1701.n7 0.575
R2308 a_24327_1701.n8 a_24327_1701.n5 0.227
R2309 a_24327_1701.n9 a_24327_1701.n8 0.2
R2310 a_24327_1701.n3 a_24327_1701.n2 0.001
R2311 Y[1].n7 Y[1].n6 217.612
R2312 Y[1].n4 Y[1].n2 157.665
R2313 Y[1].n4 Y[1].n3 122.999
R2314 Y[1].n6 Y[1].n0 90.436
R2315 Y[1].n5 Y[1].n1 90.416
R2316 Y[1].n6 Y[1].n5 74.302
R2317 Y[1].n5 Y[1].n4 50.575
R2318 Y[1].n0 Y[1].t7 14.282
R2319 Y[1].n0 Y[1].t6 14.282
R2320 Y[1].n1 Y[1].t5 14.282
R2321 Y[1].n1 Y[1].t3 14.282
R2322 Y[1].n3 Y[1].t1 14.282
R2323 Y[1].n3 Y[1].t2 14.282
R2324 Y[1].n2 Y[1].t0 8.7
R2325 Y[1].n2 Y[1].t4 8.7
R2326 Y[1] Y[1].n7 0.04
R2327 Y[1].n7 Y[1] 0.039
R2328 a_20554_n3232.n10 a_20554_n3232.n8 552.333
R2329 a_20554_n3232.n7 a_20554_n3232.t14 394.151
R2330 a_20554_n3232.n11 a_20554_n3232.n10 342.688
R2331 a_20554_n3232.n9 a_20554_n3232.t15 294.653
R2332 a_20554_n3232.n6 a_20554_n3232.t11 269.523
R2333 a_20554_n3232.t14 a_20554_n3232.n6 269.523
R2334 a_20554_n3232.n5 a_20554_n3232.t10 198.043
R2335 a_20554_n3232.n6 a_20554_n3232.t13 160.666
R2336 a_20554_n3232.n3 a_20554_n3232.n1 157.665
R2337 a_20554_n3232.n10 a_20554_n3232.n9 126.566
R2338 a_20554_n3232.n3 a_20554_n3232.n2 122.746
R2339 a_20554_n3232.n9 a_20554_n3232.t12 111.663
R2340 a_20554_n3232.n8 a_20554_n3232.n7 97.816
R2341 a_20554_n3232.n5 a_20554_n3232.t9 93.989
R2342 a_20554_n3232.n12 a_20554_n3232.n11 90.436
R2343 a_20554_n3232.n4 a_20554_n3232.n0 90.416
R2344 a_20554_n3232.n7 a_20554_n3232.t8 80.333
R2345 a_20554_n3232.n11 a_20554_n3232.n4 74.302
R2346 a_20554_n3232.n4 a_20554_n3232.n3 50.575
R2347 a_20554_n3232.n2 a_20554_n3232.t4 14.282
R2348 a_20554_n3232.n2 a_20554_n3232.t5 14.282
R2349 a_20554_n3232.n0 a_20554_n3232.t6 14.282
R2350 a_20554_n3232.n0 a_20554_n3232.t0 14.282
R2351 a_20554_n3232.n12 a_20554_n3232.t1 14.282
R2352 a_20554_n3232.t2 a_20554_n3232.n12 14.282
R2353 a_20554_n3232.n1 a_20554_n3232.t3 8.7
R2354 a_20554_n3232.n1 a_20554_n3232.t7 8.7
R2355 a_20554_n3232.n8 a_20554_n3232.n5 6.615
R2356 Y[4].n7 Y[4].n6 217.612
R2357 Y[4].n4 Y[4].n2 157.665
R2358 Y[4].n4 Y[4].n3 122.746
R2359 Y[4].n6 Y[4].n0 90.436
R2360 Y[4].n5 Y[4].n1 90.416
R2361 Y[4].n6 Y[4].n5 74.302
R2362 Y[4].n5 Y[4].n4 50.575
R2363 Y[4].n3 Y[4].t4 14.282
R2364 Y[4].n3 Y[4].t5 14.282
R2365 Y[4].n1 Y[4].t6 14.282
R2366 Y[4].n1 Y[4].t1 14.282
R2367 Y[4].n0 Y[4].t2 14.282
R2368 Y[4].n0 Y[4].t3 14.282
R2369 Y[4].n2 Y[4].t7 8.7
R2370 Y[4].n2 Y[4].t0 8.7
R2371 Y[4] Y[4].n7 0.041
R2372 Y[4].n7 Y[4] 0.039
C0 a_1636_974# w_2360_2336# 0.06fF
C1 a_15222_n1096# A[2] 0.00fF
C2 w_10556_n4263# a_9462_n3933# 0.04fF
C3 w_16255_4467# w_17397_4471# 0.03fF
C4 a_24341_n3226# a_23697_n4219# 0.01fF
C5 a_1636_974# a_3178_973# 0.01fF
C6 a_14688_2570# a_16409_4529# 0.02fF
C7 a_21241_970# a_24109_4537# 0.00fF
C8 a_4750_n1580# A[7] 0.00fF
C9 a_8149_971# a_7559_1408# 0.14fF
C10 w_23603_n4255# a_22509_n3925# 0.04fF
C11 w_17090_n4258# a_17184_n4222# 0.13fF
C12 w_13939_1341# a_14093_1403# 0.12fF
C13 a_21660_n1723# a_20653_n1063# 0.00fF
C14 w_7405_1346# a_7796_771# 0.00fF
C15 a_1641_2578# a_4295_2398# 0.00fF
C16 w_20497_1345# a_18181_1671# 0.00fF
C17 a_4722_1705# a_2397_2398# 0.00fF
C18 a_16225_965# a_15444_2390# 0.00fF
C19 a_14098_n3928# B[5] 0.00fF
C20 a_16555_3946# VDD 1.34fF
C21 a_24341_n3226# A[4] 0.01fF
C22 a_14335_2370# VSS 0.37fF
C23 a_9462_n3933# a_11299_n4838# 0.00fF
C24 a_21735_n1093# a_22547_1701# 0.00fF
C25 a_1627_4228# a_4504_4541# 0.01fF
C26 a_54_n3210# VDD 0.68fF
C27 a_15576_n1096# B[5] 0.13fF
C28 a_1048_n1067# a_2130_n1097# 0.01fF
C29 a_2824_1705# a_3236_1679# 0.14fF
C30 a_2397_2398# a_4295_2398# 0.00fF
C31 a_1342_n1093# a_2484_n1097# 0.12fF
C32 a_3236_1679# VDD 0.71fF
C33 a_1048_n1067# carry_out 0.09fF
C34 w_21965_2332# VSS 0.36fF
C35 VDD a_10645_n2623# 1.48fF
C36 a_22841_1675# a_22089_n1093# 0.00fF
C37 w_1961_n1716# w_819_n1712# 0.03fF
C38 a_16555_3946# a_17551_4533# 0.06fF
C39 a_9168_n4639# Y[6] 0.00fF
C40 a_20651_1407# a_20656_3011# 0.01fF
C41 a_20656_3011# a_21241_970# 0.03fF
C42 a_20947_n1089# VSS 0.87fF
C43 a_22783_969# VSS 0.42fF
C44 a_8910_2395# B[1] 0.60fF
C45 a_22841_1675# B[3] 0.01fF
C46 a_13686_n3902# a_15044_n3209# 0.02fF
C47 a_16283_1671# VDD 0.71fF
C48 a_20651_1407# B[3] 0.03fF
C49 a_20611_n3925# a_20553_n4631# 0.00fF
C50 a_21241_970# B[3] 0.13fF
C51 a_8154_2575# a_7550_4662# 0.00fF
C52 a_1342_n1093# a_1006_n3929# 0.00fF
C53 a_14321_4020# VSS 0.37fF
C54 B[7] a_4092_n4223# 0.03fF
C55 w_17085_n2654# VDD 0.37fF
C56 a_9875_4534# VSS 0.05fF
C57 w_10556_n4263# w_6576_n3276# 0.00fF
C58 w_18_n3272# a_712_n4635# 0.02fF
C59 a_21660_n1723# a_20518_n1719# 0.01fF
C60 a_21795_n1067# a_22089_n1093# 0.05fF
C61 a_3362_4537# a_3508_3954# 0.13fF
C62 w_9721_4472# a_8154_2575# 0.08fF
C63 a_2492_n3903# a_54_n3210# 0.00fF
C64 w_21965_2332# w_23955_4475# 0.02fF
C65 w_892_1349# w_897_2953# 0.02fF
C66 B[7] a_2846_n4635# 0.00fF
C67 a_22089_n1093# B[4] 0.13fF
C68 Y[5] A[5] 0.01fF
C69 w_19623_n3268# a_22089_n1093# 0.06fF
C70 w_6576_n3276# a_8688_n1101# 0.00fF
C71 a_9749_1676# a_11647_1676# 0.00fF
C72 a_17342_2390# a_17433_4533# 0.00fF
C73 w_13110_n3271# a_13804_n4634# 0.02fF
C74 a_17828_n3229# VDD 0.03fF
C75 w_18_n3272# a_2484_n1097# 0.06fF
C76 w_8873_2333# a_9455_970# 0.02fF
C77 a_18181_1671# a_18123_965# 0.00fF
C78 a_17842_n1579# a_15222_n1096# 0.00fF
C79 B[6] a_10650_n4227# 0.03fF
C80 a_14674_4220# VSS 0.39fF
C81 w_17099_n1004# a_15282_n1070# 0.00fF
C82 w_22813_4471# a_22967_4533# 0.08fF
C83 a_8140_4225# a_8154_2575# 0.04fF
C84 w_18_n3272# a_1006_n3929# 0.26fF
C85 a_5134_1679# a_5076_973# 0.00fF
C86 a_14688_2570# w_13930_4595# 0.00fF
C87 a_24445_969# A[3] 0.00fF
C88 a_1627_4228# a_1274_4028# 0.00fF
C89 a_2397_2398# a_2942_973# 0.02fF
C90 a_712_n4635# a_594_n3903# 0.01fF
C91 a_7564_3012# a_8154_2575# 0.11fF
C92 w_8873_2333# A[2] 0.01fF
C93 a_1283_774# VSS 0.37fF
C94 a_15938_n4634# a_15996_n3928# 0.00fF
C95 a_4386_4541# w_2360_2336# 0.04fF
C96 a_7559_1408# A[1] 0.22fF
C97 a_17887_965# VDD 0.01fF
C98 a_2824_1705# VSS 0.26fF
C99 w_7410_2950# a_7559_1408# 0.00fF
C100 a_7546_n1097# a_8748_n1075# 0.13fF
C101 VDD VSS 118.91fF
C102 w_3998_n4259# w_3993_n2655# 0.02fF
C103 VDD A[6] 1.30fF
C104 a_4087_n2619# VSS 0.26fF
C105 a_16225_965# a_16283_1671# 0.00fF
C106 a_15989_965# a_17342_2390# 0.01fF
C107 w_8873_2333# a_7801_2375# 0.00fF
C108 w_1961_n1716# a_2190_n1071# 0.09fF
C109 w_19623_n3268# a_20199_n3899# 0.32fF
C110 a_4101_n969# B[7] 0.09fF
C111 a_21557_n3206# w_21566_n1712# 0.00fF
C112 a_2055_n1727# VSS 0.66fF
C113 a_1046_1411# w_819_n1712# 0.00fF
C114 a_8149_971# w_7396_4600# 0.02fF
C115 w_13939_1341# B[2] 0.17fF
C116 a_17179_n2618# a_14434_n1092# 0.12fF
C117 a_14084_4657# VSS 0.19fF
C118 a_11235_1702# Y[1] 2.33fF
C119 a_9042_n1101# a_7900_n1097# 0.12fF
C120 a_17551_4533# VSS 0.05fF
C121 a_1006_n3929# a_594_n3903# 0.16fF
C122 a_2130_n1097# A[7] 0.01fF
C123 w_20502_2949# a_20651_1407# 0.00fF
C124 a_14688_2570# a_14335_2370# 0.00fF
C125 w_20502_2949# a_21241_970# 0.04fF
C126 w_883_4603# B[0] 0.14fF
C127 a_20317_n4631# VDD 0.00fF
C128 a_2492_n3903# VSS 0.25fF
C129 w_1961_n1716# a_1952_n3210# 0.00fF
C130 w_23955_4475# VDD 0.66fF
C131 a_23706_n965# VSS 0.24fF
C132 a_22841_1675# a_22547_1701# 0.17fF
C133 w_16255_4467# a_17433_4533# 0.03fF
C134 w_16255_4467# a_16291_4529# 0.20fF
C135 a_3244_4537# a_3362_4537# 1.20fF
C136 a_20651_1407# a_22547_1701# 0.01fF
C137 a_21241_970# a_22547_1701# 0.04fF
C138 a_1641_2578# a_1046_1411# 0.01fF
C139 a_22967_4533# a_23991_4537# 0.02fF
C140 w_10863_4476# a_10021_3951# 0.29fF
C141 a_4840_973# Y[0] 0.43fF
C142 a_5076_973# carry_in 0.01fF
C143 a_17769_1697# Y[2] 2.33fF
C144 a_16225_965# VSS 0.42fF
C145 a_11647_1676# A[2] 0.01fF
C146 a_10899_4538# a_11017_4538# 1.20fF
C147 w_21965_2332# a_20656_3011# 0.02fF
C148 a_2397_2398# a_1046_1411# 0.02fF
C149 a_22089_n1093# a_20947_n1089# 0.12fF
C150 w_21965_2332# B[3] 0.43fF
C151 w_2360_2336# a_5076_973# 0.00fF
C152 a_1641_2578# w_4350_4479# 0.12fF
C153 a_3362_4537# a_4504_4541# 0.01fF
C154 a_22089_n1093# a_22783_969# 0.00fF
C155 w_23598_n2651# a_21735_n1093# 0.01fF
C156 w_8519_n1720# B[6] 0.00fF
C157 a_15444_2390# a_17342_2390# 0.00fF
C158 a_20593_n1089# VSS 0.44fF
C159 w_8519_n1720# a_8748_n1075# 0.09fF
C160 w_7377_n1716# a_8613_n1731# 0.01fF
C161 B[3] a_22783_969# 0.00fF
C162 w_883_4603# a_1051_3015# 0.00fF
C163 a_14093_1403# Y[1] 0.00fF
C164 a_10899_4538# a_8149_971# 0.01fF
C165 a_14688_2570# a_14674_4220# 0.04fF
C166 a_17179_n2618# a_17193_n968# 0.01fF
C167 w_15053_n1715# a_14683_966# 0.00fF
C168 w_22813_4471# VSS 0.15fF
C169 w_897_2953# VSS 0.17fF
C170 a_23697_n4219# VSS 0.31fF
C171 w_7396_4600# A[1] 0.06fF
C172 w_7396_4600# w_7410_2950# 0.01fF
C173 a_23900_2394# a_24681_969# 0.00fF
C174 a_9042_n1101# a_8510_n3214# 0.01fF
C175 w_8519_n1720# a_10659_n973# 0.00fF
C176 a_24109_4537# VDD 1.34fF
C177 A[4] VSS 1.90fF
C178 a_14688_2570# VDD 1.65fF
C179 a_15702_n4634# A[5] 0.10fF
C180 a_3362_4537# a_1627_4228# 0.04fF
C181 w_8873_2333# a_11235_1702# 0.35fF
C182 a_7796_771# B[1] 0.00fF
C183 VDD a_15996_n3928# 0.83fF
C184 a_14041_n3235# Y[5] 0.18fF
C185 a_15989_1697# a_18123_965# 0.00fF
C186 a_9337_1702# Y[1] 0.00fF
C187 w_22813_4471# w_23955_4475# 0.03fF
C188 a_14330_766# A[2] 0.01fF
C189 a_14688_2570# a_14084_4657# 0.00fF
C190 a_14688_2570# a_17551_4533# 0.04fF
C191 a_7546_n1097# a_7559_1408# 0.00fF
C192 a_4741_n4834# a_2484_n1097# 0.00fF
C193 a_4722_1705# a_3236_1679# 0.02fF
C194 a_9404_n4639# a_10650_n4227# 0.00fF
C195 a_1342_n1093# VDD 1.77fF
C196 a_20656_3011# VDD 1.47fF
C197 a_1342_n1093# a_4087_n2619# 0.12fF
C198 VDD Y[6] 0.08fF
C199 A[7] a_4736_n3230# 0.01fF
C200 a_20317_n4631# A[4] 0.00fF
C201 w_10556_n4263# a_11294_n3234# 0.00fF
C202 a_22089_n1093# VDD 1.32fF
C203 VDD B[3] 0.92fF
C204 B[0] carry_in 0.63fF
C205 w_892_1349# a_2942_973# 0.00fF
C206 A[0] Y[0] 0.01fF
C207 a_16555_3946# a_17342_2390# 0.00fF
C208 w_10556_n4263# a_9168_n4639# 0.00fF
C209 a_3236_1679# a_4295_2398# 0.20fF
C210 a_1342_n1093# a_2055_n1727# 0.04fF
C211 a_13146_n3209# a_13804_n4634# 0.02fF
C212 w_892_1349# w_1961_n1716# 0.00fF
C213 a_1048_n1067# a_913_n1723# 1.19fF
C214 a_1037_4665# A[0] 0.14fF
C215 a_11294_n3234# a_11299_n4838# 0.00fF
C216 w_2360_2336# B[0] 0.43fF
C217 a_20653_n1063# VSS 0.07fF
C218 w_13930_4595# A[2] 0.06fF
C219 a_4840_973# A[0] 0.00fF
C220 a_17769_1697# VDD 2.54fF
C221 a_3178_973# B[0] 0.00fF
C222 a_13686_n3902# w_13911_n1711# 0.00fF
C223 a_988_n1093# A[0] 0.00fF
C224 a_20611_n3925# a_22451_n4631# 0.00fF
C225 a_1342_n1093# a_2492_n3903# 0.03fF
C226 a_16283_1671# a_17342_2390# 0.20fF
C227 a_14140_n1066# A[2] 0.00fF
C228 a_23991_4537# VSS 0.62fF
C229 Y[3] VSS 0.23fF
C230 B[5] A[5] 1.71fF
C231 w_17090_n4258# w_13110_n3271# 0.00fF
C232 w_18_n3272# VDD 1.02fF
C233 w_17085_n2654# a_17179_n2618# 0.13fF
C234 a_16409_4529# a_14683_966# 0.05fF
C235 w_18_n3272# a_4087_n2619# 0.02fF
C236 a_11017_4538# VSS 0.05fF
C237 a_1037_4665# a_1636_974# 0.03fF
C238 a_23706_n965# a_22089_n1093# 0.03fF
C239 w_15407_2328# a_18181_1671# 0.20fF
C240 w_21965_2332# a_22547_1701# 0.58fF
C241 a_17833_n4833# B[5] 0.00fF
C242 a_21246_2574# A[3] 0.07fF
C243 a_17828_n3229# a_17179_n2618# 0.38fF
C244 a_11235_1702# a_11647_1676# 0.15fF
C245 w_13110_n3271# a_14040_n4634# 0.00fF
C246 a_9042_n1101# a_9462_n3933# 0.10fF
C247 w_23612_n1001# a_23692_n2615# 0.00fF
C248 a_20199_n3899# VDD 2.54fF
C249 Y[2] A[2] 0.01fF
C250 w_18_n3272# a_2055_n1727# 0.02fF
C251 a_9749_1676# VDD 0.71fF
C252 a_22547_1701# a_22783_969# 0.36fF
C253 a_15222_n1096# B[2] 0.00fF
C254 a_4750_n1580# a_2130_n1097# 0.00fF
C255 w_23612_n1001# a_24355_n1576# 0.00fF
C256 w_10565_n1009# a_10645_n2623# 0.00fF
C257 w_17099_n1004# VDD 0.38fF
C258 a_1636_974# a_988_n1093# 0.00fF
C259 a_4722_1705# VSS 0.22fF
C260 a_14098_n3928# A[5] 0.04fF
C261 a_8149_971# VSS 1.12fF
C262 B[7] a_1952_n3210# 0.01fF
C263 w_23955_4475# a_23991_4537# 0.21fF
C264 a_20518_n1719# VSS 0.64fF
C265 w_22813_4471# a_24109_4537# 0.01fF
C266 carry_in a_1051_3015# 0.14fF
C267 a_14335_2370# A[2] 0.01fF
C268 w_18_n3272# a_2492_n3903# 0.27fF
C269 a_15576_n1096# A[5] 0.14fF
C270 a_594_n3903# VDD 2.55fF
C271 a_3236_1679# a_2942_973# 0.02fF
C272 w_2360_2336# a_1051_3015# 0.02fF
C273 w_7377_n1716# VDD 0.67fF
C274 a_4295_2398# VSS 0.46fF
C275 a_14330_766# a_14683_966# 0.00fF
C276 a_15576_n1096# a_17833_n4833# 0.00fF
C277 a_22089_n1093# a_20593_n1089# 0.03fF
C278 a_8688_n1101# a_8613_n1731# 0.14fF
C279 a_17179_n2618# VSS 0.26fF
C280 carry_in a_2484_n1097# 0.02fF
C281 w_3998_n4259# B[7] 0.17fF
C282 a_17887_965# a_17342_2390# 0.02fF
C283 w_20502_2949# VDD 0.37fF
C284 w_892_1349# a_1046_1411# 0.12fF
C285 w_8873_2333# a_9337_1702# 0.29fF
C286 a_17342_2390# VSS 0.46fF
C287 w_4007_n1005# a_2484_n1097# 0.02fF
C288 a_17184_n4222# a_15044_n3209# 0.00fF
C289 a_16555_3946# w_16255_4467# 0.23fF
C290 w_23612_n1001# a_21660_n1723# 0.01fF
C291 a_22089_n1093# a_23697_n4219# 0.14fF
C292 w_6576_n3276# a_9042_n1101# 0.06fF
C293 w_23598_n2651# B[4] 0.29fF
C294 A[7] a_4092_n4223# 0.18fF
C295 a_14321_4020# A[2] 0.00fF
C296 a_3178_973# a_2484_n1097# 0.00fF
C297 w_22813_4471# B[3] 0.00fF
C298 w_3993_n2655# VSS 0.17fF
C299 a_2492_n3903# a_594_n3903# 0.02fF
C300 a_22089_n1093# A[4] 0.14fF
C301 a_19659_n3206# VSS 0.36fF
C302 Y[4] A[5] 0.01fF
C303 A[7] a_2846_n4635# 0.00fF
C304 w_10551_n2659# a_11294_n3234# 0.00fF
C305 w_13930_4595# a_14683_966# 0.02fF
C306 a_22547_1701# VDD 0.23fF
C307 a_15222_n1096# B[5] 0.01fF
C308 w_7405_1346# B[1] 0.17fF
C309 w_10565_n1009# VSS 0.19fF
C310 w_10565_n1009# A[6] 0.07fF
C311 w_16255_4467# a_16283_1671# 0.00fF
C312 w_8873_2333# a_9691_970# 0.00fF
C313 VDD a_9455_970# 0.01fF
C314 a_21246_2574# a_20642_4661# 0.00fF
C315 a_7900_n1097# a_8510_n3214# 0.02fF
C316 a_7606_n1071# a_8613_n1731# 0.00fF
C317 a_7471_n1727# a_8748_n1075# 0.02fF
C318 a_14674_4220# A[2] 0.01fF
C319 w_13110_n3271# a_13686_n3902# 0.32fF
C320 a_15702_n4634# a_14041_n3235# 0.44fF
C321 a_1636_974# A[0] 0.17fF
C322 a_22215_n4631# a_21557_n3206# 0.02fF
C323 a_23991_4537# a_24109_4537# 1.20fF
C324 a_19659_n3206# a_20317_n4631# 0.02fF
C325 a_2942_973# VSS 0.68fF
C326 w_8873_2333# B[2] 0.00fF
C327 a_14080_n1092# a_15044_n3209# 0.00fF
C328 a_1288_2378# a_1274_4028# 0.00fF
C329 VDD A[2] 1.46fF
C330 A[1] VSS 1.99fF
C331 w_17397_4471# a_15989_1697# 0.01fF
C332 w_1961_n1716# VSS 0.24fF
C333 a_11647_1676# a_9337_1702# 0.00fF
C334 w_7410_2950# VSS 0.16fF
C335 a_7559_1408# a_8910_2395# 0.02fF
C336 a_21246_2574# a_23113_3950# 0.49fF
C337 a_20199_n3899# A[4] 0.02fF
C338 a_14335_2370# a_14683_966# 0.01fF
C339 a_3236_1679# a_1046_1411# 0.00fF
C340 a_22849_4533# a_21232_4224# 0.16fF
C341 a_15576_n1096# a_15222_n1096# 0.48fF
C342 a_22002_2394# a_21246_2574# 0.03fF
C343 a_7801_2375# VDD 0.02fF
C344 a_4101_n969# A[7] 0.14fF
C345 a_22089_n1093# a_20653_n1063# 0.00fF
C346 a_1048_n1067# w_819_n1712# 0.08fF
C347 a_4750_n1580# a_4736_n3230# 0.00fF
C348 a_7471_n1727# a_7152_n3907# 0.00fF
C349 a_14084_4657# A[2] 0.14fF
C350 a_2130_n1097# carry_out 0.00fF
C351 a_22841_1675# a_24445_969# 0.01fF
C352 w_883_4603# VDD 0.38fF
C353 a_14330_766# a_14093_1403# 0.38fF
C354 w_16255_4467# VSS 0.15fF
C355 a_24739_1675# a_24681_969# 0.00fF
C356 a_14321_4020# a_14683_966# 0.01fF
C357 w_23603_n4255# a_22215_n4631# 0.00fF
C358 w_15407_2328# a_15989_1697# 0.58fF
C359 a_14041_n3235# B[5] 0.17fF
C360 a_14688_2570# a_17342_2390# 0.00fF
C361 w_8873_2333# a_8140_4225# 0.00fF
C362 a_21557_n3206# B[4] 0.01fF
C363 VDD a_4741_n4834# 0.01fF
C364 a_15996_n3928# a_17179_n2618# 0.00fF
C365 a_10650_n4227# a_10645_n2623# 0.01fF
C366 a_20518_n1719# a_22089_n1093# 0.01fF
C367 a_7564_n3933# a_9050_n3907# 0.02fF
C368 w_19623_n3268# a_21557_n3206# 0.19fF
C369 a_5076_973# Y[0] 0.36fF
C370 w_10556_n4263# VDD 0.33fF
C371 a_7900_n1097# a_9462_n3933# 0.03fF
C372 w_23598_n2651# a_20947_n1089# 0.05fF
C373 a_16225_965# A[2] 0.01fF
C374 w_8873_2333# a_7564_3012# 0.02fF
C375 a_11647_1676# B[2] 0.00fF
C376 a_5134_1679# a_2824_1705# 0.00fF
C377 a_14674_4220# a_14683_966# 0.49fF
C378 a_5134_1679# VDD 0.69fF
C379 a_8688_n1101# VDD 0.97fF
C380 a_11299_n4838# VDD 0.01fF
C381 a_17842_n1579# VDD 0.02fF
C382 w_15053_n1715# B[5] 0.00fF
C383 a_1046_1411# VSS 0.27fF
C384 a_14140_n1066# a_14093_1403# 0.00fF
C385 A[7] a_7152_n3907# 0.00fF
C386 a_10899_4538# a_10808_2395# 0.00fF
C387 a_14041_n3235# a_14098_n3928# 0.59fF
C388 a_4840_973# a_5076_973# 0.04fF
C389 a_13146_n3209# a_14040_n4634# 0.00fF
C390 a_1048_n1067# a_2190_n1071# 0.01fF
C391 a_15576_n1096# a_14041_n3235# 0.04fF
C392 VDD a_14683_966# 1.34fF
C393 w_3993_n2655# a_1342_n1093# 0.05fF
C394 w_4350_4479# VSS 0.14fF
C395 a_20199_n3899# a_20518_n1719# 0.00fF
C396 a_1641_2578# a_3508_3954# 0.49fF
C397 a_17342_2390# a_17769_1697# 0.19fF
C398 a_8149_971# a_9749_1676# 0.01fF
C399 a_14335_2370# a_14093_1403# 0.01fF
C400 w_23603_n4255# B[4] 0.17fF
C401 a_15576_n1096# w_15053_n1715# 0.12fF
C402 w_6576_n3276# a_7900_n1097# 0.12fF
C403 a_17551_4533# a_14683_966# 0.00fF
C404 w_23603_n4255# w_19623_n3268# 0.00fF
C405 a_14084_4657# a_14683_966# 0.03fF
C406 a_4386_4541# a_1636_974# 0.01fF
C407 a_10650_n4227# VSS 0.31fF
C408 a_10650_n4227# A[6] 0.18fF
C409 a_7606_n1071# VDD 1.34fF
C410 a_20642_4661# A[3] 0.14fF
C411 w_20497_1345# a_20893_2374# 0.00fF
C412 a_11235_1702# VDD 2.54fF
C413 a_20879_4024# A[3] 0.00fF
C414 w_883_4603# w_897_2953# 0.01fF
C415 w_17099_n1004# a_17179_n2618# 0.00fF
C416 w_23598_n2651# VDD 0.37fF
C417 a_9042_n1101# a_11294_n3234# 0.01fF
C418 a_14330_766# B[2] 0.00fF
C419 a_9042_n1101# a_9168_n4639# 0.02fF
C420 a_8149_971# w_7377_n1716# 0.00fF
C421 w_1961_n1716# a_1342_n1093# 0.10fF
C422 a_13804_n4634# A[6] 0.00fF
C423 a_7546_n1097# A[6] 0.00fF
C424 a_13804_n4634# VSS 0.69fF
C425 Y[3] a_22547_1701# 0.18fF
C426 a_14688_2570# w_16255_4467# 0.08fF
C427 a_7546_n1097# VSS 0.44fF
C428 a_2610_n4635# a_2904_n3929# 0.02fF
C429 VDD Y[5] 0.08fF
C430 a_9462_n3933# a_8510_n3214# 0.07fF
C431 a_1283_774# carry_in 0.03fF
C432 a_23991_4537# a_22547_1701# 0.01fF
C433 a_2824_1705# carry_in 0.00fF
C434 a_15989_1697# a_17433_4533# 0.01fF
C435 VDD carry_in 1.30fF
C436 a_19659_n3206# a_20199_n3899# 0.17fF
C437 w_17090_n4258# a_14434_n1092# 0.01fF
C438 a_1037_4665# B[0] 0.10fF
C439 a_22002_2394# A[3] 0.11fF
C440 a_23113_3950# A[3] 0.00fF
C441 w_4007_n1005# VDD 0.38fF
C442 a_16225_965# a_14683_966# 0.01fF
C443 w_4007_n1005# a_4087_n2619# 0.00fF
C444 carry_in a_2055_n1727# 0.01fF
C445 a_8510_n3214# a_7270_n4639# 0.01fF
C446 a_7564_n3933# a_7506_n4639# 0.00fF
C447 w_2360_2336# a_2824_1705# 0.29fF
C448 a_2824_1705# a_3178_973# 0.00fF
C449 w_13939_1341# Y[1] 0.00fF
C450 w_2360_2336# VDD 0.93fF
C451 Y[1] a_11353_970# 0.43fF
C452 a_3178_973# VDD 0.00fF
C453 w_21965_2332# a_24445_969# 0.02fF
C454 a_5076_973# A[0] 0.00fF
C455 w_4007_n1005# a_2055_n1727# 0.01fF
C456 w_13930_4595# B[2] 0.14fF
C457 a_21557_n3206# a_20947_n1089# 0.02fF
C458 w_8873_2333# a_8154_2575# 0.14fF
C459 a_15938_n4634# a_15702_n4634# 0.04fF
C460 w_23598_n2651# a_23706_n965# 0.03fF
C461 B[7] VSS 0.78fF
C462 A[7] a_948_n4635# 0.00fF
C463 a_13146_n3209# a_13686_n3902# 0.17fF
C464 a_4750_n1580# a_4101_n969# 0.38fF
C465 w_10551_n2659# VDD 0.37fF
C466 a_8149_971# a_9455_970# 0.02fF
C467 a_15576_n1096# a_15282_n1070# 0.05fF
C468 w_19623_n3268# B[5] 0.00fF
C469 a_17833_n4833# A[5] 0.01fF
C470 a_20611_n3925# VSS 0.48fF
C471 a_7559_1408# a_7796_771# 0.38fF
C472 a_15989_965# a_15989_1697# 0.43fF
C473 a_14093_1403# VDD 1.38fF
C474 w_7396_4600# a_9757_4534# 0.01fF
C475 a_9749_1676# A[1] 0.81fF
C476 a_10808_2395# VSS 0.46fF
C477 a_22215_n4631# Y[4] 0.00fF
C478 w_6576_n3276# a_8510_n3214# 0.19fF
C479 w_23612_n1001# VSS 0.20fF
C480 a_16283_1671# a_18181_1671# 0.00fF
C481 a_3244_4537# a_1641_2578# 0.04fF
C482 a_20642_4661# a_20879_4024# 0.38fF
C483 a_9042_n1101# a_8613_n1731# 0.08fF
C484 A[7] a_1952_n3210# 0.80fF
C485 a_14335_2370# B[2] 0.03fF
C486 a_1037_4665# a_1051_3015# 0.01fF
C487 w_13110_n3271# a_15044_n3209# 0.19fF
C488 a_22451_n4631# a_22097_n3899# 0.00fF
C489 a_8149_971# a_7801_2375# 0.01fF
C490 a_22215_n4631# a_22509_n3925# 0.02fF
C491 a_20611_n3925# a_20317_n4631# 0.02fF
C492 w_8519_n1720# VSS 0.23fF
C493 w_3998_n4259# A[7] 0.13fF
C494 w_23603_n4255# a_20947_n1089# 0.01fF
C495 w_8519_n1720# A[6] 0.01fF
C496 w_7377_n1716# A[1] 0.02fF
C497 a_14080_n1092# w_13911_n1711# 0.29fF
C498 a_23692_n2615# a_22097_n3899# 0.00fF
C499 B[6] a_7564_n3933# 0.00fF
C500 a_1641_2578# a_4504_4541# 0.04fF
C501 w_13944_2945# VSS 0.16fF
C502 w_23598_n2651# a_23697_n4219# 0.00fF
C503 a_22841_1675# a_21246_2574# 0.02fF
C504 a_9337_1702# VDD 2.55fF
C505 a_17342_2390# A[2] 0.04fF
C506 VDD a_21557_n3206# 0.71fF
C507 a_21241_970# a_21246_2574# 0.12fF
C508 a_24445_969# VDD 0.01fF
C509 a_15938_n4634# B[5] 0.00fF
C510 a_20651_1407# a_21246_2574# 0.01fF
C511 w_20424_n1708# A[3] 0.03fF
C512 w_23598_n2651# A[4] 0.07fF
C513 a_14321_4020# B[2] 0.02fF
C514 a_21735_n1093# A[3] 0.00fF
C515 w_897_2953# carry_in 0.07fF
C516 A[0] B[0] 2.23fF
C517 a_988_n1093# a_2484_n1097# 0.03fF
C518 a_2130_n1097# a_913_n1723# 0.01fF
C519 a_17887_965# a_18181_1671# 0.02fF
C520 a_16225_965# a_14093_1403# 0.00fF
C521 carry_out a_913_n1723# 0.07fF
C522 a_18181_1671# VSS 0.36fF
C523 w_19623_n3268# Y[4] 0.15fF
C524 a_15222_n1096# A[5] 0.01fF
C525 a_15938_n4634# a_14098_n3928# 0.00fF
C526 w_8873_2333# a_11353_970# 0.02fF
C527 a_15989_1697# a_15444_2390# 0.09fF
C528 a_15576_n1096# a_15938_n4634# 0.01fF
C529 a_1641_2578# a_1627_4228# 0.04fF
C530 a_7152_n3907# a_7564_n3933# 0.16fF
C531 VDD a_9691_970# 0.00fF
C532 w_3208_4475# a_1037_4665# 0.00fF
C533 a_9875_4534# a_7550_4662# 0.00fF
C534 w_20424_n1708# w_21566_n1712# 0.03fF
C535 A[1] a_9455_970# 0.11fF
C536 a_10899_4538# a_9757_4534# 0.01fF
C537 a_6612_n3214# a_8510_n3214# 0.00fF
C538 a_988_n1093# a_1006_n3929# 0.00fF
C539 a_14005_n1722# a_13686_n3902# 0.00fF
C540 a_23900_2394# a_24739_1675# 0.08fF
C541 a_9875_4534# w_9721_4472# 0.08fF
C542 a_4722_1705# a_5134_1679# 0.15fF
C543 a_21735_n1093# w_21566_n1712# 0.21fF
C544 a_14674_4220# B[2] 0.01fF
C545 a_21660_n1723# a_22097_n3899# 0.01fF
C546 w_6576_n3276# a_9462_n3933# 0.25fF
C547 a_22509_n3925# B[4] 0.56fF
C548 a_15576_n1096# a_14140_n1066# 0.00fF
C549 a_1636_974# B[0] 0.13fF
C550 w_19623_n3268# a_22509_n3925# 0.25fF
C551 w_13110_n3271# a_17184_n4222# 0.00fF
C552 w_23603_n4255# VDD 0.33fF
C553 w_15407_2328# a_14098_3007# 0.02fF
C554 w_6576_n3276# a_7270_n4639# 0.02fF
C555 a_5134_1679# a_4295_2398# 0.08fF
C556 VDD B[2] 0.92fF
C557 a_4101_n969# a_2130_n1097# 0.12fF
C558 a_7900_n1097# a_11294_n3234# 0.00fF
C559 a_7801_2375# A[1] 0.01fF
C560 a_15702_n4634# VDD 0.00fF
C561 a_17842_n1579# a_17179_n2618# 0.00fF
C562 a_20888_770# A[3] 0.01fF
C563 a_8910_2395# VSS 0.48fF
C564 a_9875_4534# a_8140_4225# 0.04fF
C565 w_7410_2950# a_7801_2375# 0.00fF
C566 w_17090_n4258# w_17085_n2654# 0.02fF
C567 w_20424_n1708# A[5] 0.00fF
C568 A[0] a_1051_3015# 0.06fF
C569 a_1342_n1093# B[7] 0.06fF
C570 a_14084_4657# B[2] 0.10fF
C571 VDD a_7550_4662# 1.42fF
C572 a_21557_n3206# a_20593_n1089# 0.00fF
C573 w_17090_n4258# a_17828_n3229# 0.00fF
C574 A[7] Y[7] 0.01fF
C575 a_15044_n3209# a_15147_n1726# 0.00fF
C576 w_9721_4472# VDD 0.53fF
C577 w_16255_4467# A[2] 0.01fF
C578 w_13939_1341# a_11647_1676# 0.00fF
C579 w_7405_1346# a_7559_1408# 0.12fF
C580 a_23697_n4219# a_21557_n3206# 0.00fF
C581 a_16555_3946# a_15989_1697# 0.00fF
C582 A[0] a_2484_n1097# 0.00fF
C583 a_11647_1676# a_11353_970# 0.02fF
C584 w_23612_n1001# a_22089_n1093# 0.02fF
C585 w_10565_n1009# a_8688_n1101# 0.06fF
C586 w_13110_n3271# a_14080_n1092# 0.01fF
C587 a_1636_974# a_1051_3015# 0.03fF
C588 a_14688_2570# w_13944_2945# 0.05fF
C589 a_7787_4025# B[1] 0.02fF
C590 a_14041_n3235# A[5] 0.19fF
C591 a_9042_n1101# VDD 1.31fF
C592 a_21557_n3206# A[4] 0.80fF
C593 a_3508_3954# a_3236_1679# 0.00fF
C594 a_8140_4225# VDD 0.97fF
C595 a_24445_969# A[4] 0.00fF
C596 a_22002_2394# a_21735_n1093# 0.00fF
C597 a_4736_n3230# a_4092_n4223# 0.01fF
C598 w_18_n3272# B[7] 0.40fF
C599 a_4722_1705# carry_in 0.13fF
C600 w_17090_n4258# VSS 0.20fF
C601 a_16225_965# B[2] 0.00fF
C602 a_15989_1697# a_16283_1671# 0.17fF
C603 a_5134_1679# A[1] 0.01fF
C604 a_1048_n1067# VSS 0.06fF
C605 w_7377_n1716# a_7546_n1097# 0.29fF
C606 VDD B[5] 0.91fF
C607 a_7564_3012# VDD 1.47fF
C608 a_8688_n1101# A[1] 0.00fF
C609 w_2360_2336# a_4722_1705# 0.35fF
C610 a_14040_n4634# VSS 0.42fF
C611 a_2904_n3929# a_2484_n1097# 0.10fF
C612 w_15053_n1715# A[5] 0.01fF
C613 w_3208_4475# A[0] 0.01fF
C614 a_6612_n3214# a_7270_n4639# 0.02fF
C615 w_21965_2332# a_21246_2574# 0.14fF
C616 a_4295_2398# carry_in 0.03fF
C617 a_7900_n1097# a_8613_n1731# 0.04fF
C618 a_20199_n3899# a_20611_n3925# 0.16fF
C619 a_22841_1675# A[3] 0.81fF
C620 a_21241_970# A[3] 0.17fF
C621 a_9749_1676# a_10808_2395# 0.20fF
C622 w_2360_2336# a_4295_2398# 0.26fF
C623 a_7564_n3933# a_9404_n4639# 0.00fF
C624 a_20651_1407# A[3] 0.22fF
C625 a_8510_n3214# a_9168_n4639# 0.02fF
C626 VSS a_9757_4534# 0.65fF
C627 a_4295_2398# a_3178_973# 0.00fF
C628 a_2904_n3929# a_1006_n3929# 0.00fF
C629 w_23603_n4255# a_23697_n4219# 0.13fF
C630 VDD a_14098_n3928# 0.78fF
C631 a_22509_n3925# a_20947_n1089# 0.03fF
C632 A[7] a_54_n3210# 0.00fF
C633 a_15576_n1096# VDD 1.32fF
C634 w_13939_1341# a_14330_766# 0.00fF
C635 a_13146_n3209# a_15044_n3209# 0.00fF
C636 a_2130_n1097# w_819_n1712# 0.02fF
C637 w_3208_4475# a_1636_974# 0.12fF
C638 w_23603_n4255# A[4] 0.13fF
C639 w_3993_n2655# w_4007_n1005# 0.01fF
C640 w_6576_n3276# a_6612_n3214# 0.20fF
C641 carry_out w_819_n1712# 0.17fF
C642 a_18181_1671# B[3] 0.00fF
C643 a_22002_2394# a_20888_770# 0.00fF
C644 a_7471_n1727# VSS 0.63fF
C645 a_24445_969# Y[3] 0.43fF
C646 a_23900_2394# a_22547_969# 0.01fF
C647 a_20651_1407# w_21566_n1712# 0.00fF
C648 w_16255_4467# a_14683_966# 0.12fF
C649 a_7606_n1071# A[1] 0.00fF
C650 a_17887_965# a_15989_1697# 0.09fF
C651 a_21241_970# w_21566_n1712# 0.01fF
C652 a_15989_1697# VSS 0.54fF
C653 a_24341_n3226# a_24346_n4830# 0.00fF
C654 a_11235_1702# A[1] 0.02fF
C655 a_3508_3954# VSS 0.37fF
C656 a_9875_4534# a_8154_2575# 0.02fF
C657 a_17769_1697# a_18181_1671# 0.15fF
C658 a_3362_4537# a_1641_2578# 0.02fF
C659 w_21566_n1712# B[4] 0.00fF
C660 a_21795_n1067# w_21566_n1712# 0.09fF
C661 VDD Y[4] 0.08fF
C662 a_2942_973# carry_in 0.01fF
C663 a_2824_1705# Y[0] 0.00fF
C664 w_8873_2333# Y[1] 0.15fF
C665 VDD Y[0] 0.08fF
C666 w_13110_n3271# w_13911_n1711# 0.01fF
C667 a_21246_2574# VDD 1.65fF
C668 A[1] carry_in 0.08fF
C669 w_1961_n1716# carry_in 0.06fF
C670 a_8149_971# a_9337_1702# 0.05fF
C671 w_20424_n1708# a_21735_n1093# 0.02fF
C672 a_3244_4537# a_3236_1679# 0.00fF
C673 w_10565_n1009# w_10551_n2659# 0.01fF
C674 a_14080_n1092# a_15147_n1726# 0.09fF
C675 a_1037_4665# VDD 1.48fF
C676 w_7377_n1716# w_8519_n1720# 0.03fF
C677 a_15222_n1096# w_15053_n1715# 0.21fF
C678 w_2360_2336# a_2942_973# 0.02fF
C679 B[6] a_9050_n3907# 0.10fF
C680 a_3178_973# a_2942_973# 0.04fF
C681 w_23612_n1001# a_22547_1701# 0.00fF
C682 w_2360_2336# A[1] 0.01fF
C683 a_13686_n3902# VSS 0.21fF
C684 a_8510_n3214# a_8613_n1731# 0.00fF
C685 a_13686_n3902# A[6] 0.00fF
C686 a_988_n1093# a_1283_774# 0.00fF
C687 a_4840_973# VDD 0.01fF
C688 a_2130_n1097# a_2397_2398# 0.00fF
C689 a_10808_2395# a_9455_970# 0.01fF
C690 VDD a_22509_n3925# 0.83fF
C691 a_16225_965# a_15576_n1096# 0.00fF
C692 a_21241_970# a_20642_4661# 0.03fF
C693 a_988_n1093# VDD 1.34fF
C694 a_2610_n4635# a_712_n4635# 0.01fF
C695 a_2846_n4635# a_4092_n4223# 0.00fF
C696 a_11294_n3234# a_9462_n3933# 0.00fF
C697 A[7] VSS 1.74fF
C698 a_21241_970# a_20879_4024# 0.01fF
C699 VDD a_8154_2575# 1.65fF
C700 w_13939_1341# a_14335_2370# 0.00fF
C701 a_9462_n3933# a_9168_n4639# 0.02fF
C702 a_8149_971# a_9691_970# 0.01fF
C703 a_15044_n3209# a_14434_n1092# 0.02fF
C704 a_2130_n1097# a_2190_n1071# 0.05fF
C705 a_988_n1093# a_2055_n1727# 0.09fF
C706 a_2610_n4635# a_2484_n1097# 0.02fF
C707 w_17090_n4258# a_15996_n3928# 0.04fF
C708 w_19623_n3268# A[5] 0.01fF
C709 w_10556_n4263# a_10650_n4227# 0.13fF
C710 a_22002_2394# a_22841_1675# 0.08fF
C711 a_22841_1675# a_23113_3950# 0.00fF
C712 a_7796_771# VSS 0.38fF
C713 Y[2] A[3] 0.01fF
C714 a_19659_n3206# a_21557_n3206# 0.00fF
C715 a_7270_n4639# a_9168_n4639# 0.01fF
C716 a_11299_n4838# a_10650_n4227# 0.38fF
C717 a_22002_2394# a_20651_1407# 0.02fF
C718 a_21241_970# a_23113_3950# 0.03fF
C719 a_9749_1676# a_8910_2395# 0.08fF
C720 w_20497_1345# a_22547_969# 0.00fF
C721 w_3208_4475# a_4386_4541# 0.03fF
C722 a_7152_n3907# a_9050_n3907# 0.02fF
C723 w_20424_n1708# a_20888_770# 0.00fF
C724 a_22002_2394# a_21241_970# 0.10fF
C725 a_2610_n4635# a_1006_n3929# 0.01fF
C726 a_988_n1093# a_2492_n3903# 0.00fF
C727 a_10899_4538# w_10863_4476# 0.21fF
C728 a_11017_4538# w_9721_4472# 0.01fF
C729 a_14098_3007# a_15444_2390# 0.00fF
C730 a_1342_n1093# a_1048_n1067# 0.04fF
C731 a_11647_1676# Y[1] 0.15fF
C732 a_7546_n1097# a_8688_n1101# 0.07fF
C733 a_7900_n1097# VDD 1.77fF
C734 a_3244_4537# VSS 0.65fF
C735 a_1046_1411# carry_in 0.15fF
C736 w_6576_n3276# a_11294_n3234# 0.00fF
C737 w_21965_2332# A[3] 0.60fF
C738 w_6576_n3276# a_9168_n4639# 0.02fF
C739 a_15282_n1070# a_15222_n1096# 0.05fF
C740 B[7] a_4741_n4834# 0.00fF
C741 a_8149_971# a_7550_4662# 0.03fF
C742 w_13944_2945# A[2] 0.07fF
C743 a_22783_969# A[3] 0.01fF
C744 a_22097_n3899# VSS 0.24fF
C745 a_9337_1702# A[1] 0.24fF
C746 a_14688_2570# a_15989_1697# 0.01fF
C747 a_11017_4538# a_8140_4225# 0.01fF
C748 a_17342_2390# B[2] 0.00fF
C749 a_15938_n4634# A[5] 0.00fF
C750 a_10899_4538# a_10021_3951# 0.15fF
C751 w_2360_2336# a_1046_1411# 0.00fF
C752 a_24681_969# VSS 0.42fF
C753 a_8149_971# w_9721_4472# 0.12fF
C754 a_3178_973# a_1046_1411# 0.00fF
C755 a_4504_4541# VSS 0.05fF
C756 w_22813_4471# a_21246_2574# 0.08fF
C757 w_4350_4479# carry_in 0.00fF
C758 a_1283_774# A[0] 0.01fF
C759 a_7559_1408# B[1] 0.03fF
C760 w_20488_4599# a_22849_4533# 0.01fF
C761 a_2824_1705# A[0] 0.24fF
C762 w_15407_2328# a_18123_965# 0.00fF
C763 a_17184_n4222# a_14434_n1092# 0.01fF
C764 A[0] VDD 2.01fF
C765 a_1037_4665# w_897_2953# 0.02fF
C766 Y[4] A[4] 0.01fF
C767 a_11308_n1584# B[6] 0.02fF
C768 w_4350_4479# w_2360_2336# 0.01fF
C769 a_18181_1671# A[2] 0.00fF
C770 w_13911_n1711# a_15147_n1726# 0.01fF
C771 a_7606_n1071# a_7546_n1097# 0.05fF
C772 w_21566_n1712# a_20947_n1089# 0.10fF
C773 w_13939_1341# VDD 0.33fF
C774 a_23697_n4219# a_22509_n3925# 0.02fF
C775 a_8149_971# a_8140_4225# 0.49fF
C776 Y[5] a_10650_n4227# 0.00fF
C777 VDD a_11353_970# 0.01fF
C778 A[1] a_9691_970# 0.01fF
C779 a_8149_971# a_7564_3012# 0.03fF
C780 w_20488_4599# a_21232_4224# 0.06fF
C781 a_1636_974# a_1283_774# 0.00fF
C782 a_22509_n3925# A[4] 0.07fF
C783 a_1641_2578# a_1288_2378# 0.00fF
C784 a_8910_2395# a_9455_970# 0.02fF
C785 a_1636_974# a_2824_1705# 0.05fF
C786 a_11308_n1584# a_10659_n973# 0.38fF
C787 a_9749_1676# a_9757_4534# 0.00fF
C788 a_1636_974# VDD 1.43fF
C789 a_13804_n4634# Y[5] 0.44fF
C790 a_2904_n3929# VDD 0.83fF
C791 a_15996_n3928# a_13686_n3902# 0.00fF
C792 a_2904_n3929# a_4087_n2619# 0.00fF
C793 w_20424_n1708# a_20651_1407# 0.00fF
C794 a_22841_1675# a_21735_n1093# 0.00fF
C795 w_20424_n1708# a_21241_970# 0.00fF
C796 a_1627_4228# VSS 0.39fF
C797 a_1288_2378# a_2397_2398# 0.00fF
C798 a_15989_1697# a_17769_1697# 0.12fF
C799 w_13110_n3271# B[6] 0.00fF
C800 w_8519_n1720# a_8688_n1101# 0.21fF
C801 VDD A[3] 1.46fF
C802 a_17179_n2618# B[5] 0.18fF
C803 w_6576_n3276# a_8613_n1731# 0.02fF
C804 w_10551_n2659# a_10650_n4227# 0.00fF
C805 a_7152_n3907# a_7506_n4639# 0.00fF
C806 VDD a_8510_n3214# 0.71fF
C807 w_20424_n1708# a_21795_n1067# 0.01fF
C808 a_14080_n1092# a_14434_n1092# 0.49fF
C809 a_7801_2375# a_8910_2395# 0.00fF
C810 B[0] a_1051_3015# 0.18fF
C811 w_8873_2333# a_11647_1676# 0.20fF
C812 a_21795_n1067# a_21735_n1093# 0.05fF
C813 a_1342_n1093# A[7] 0.07fF
C814 w_20424_n1708# w_19623_n3268# 0.01fF
C815 a_21735_n1093# B[4] 0.01fF
C816 a_10808_2395# a_11235_1702# 0.19fF
C817 w_10565_n1009# a_9042_n1101# 0.02fF
C818 A[1] a_7550_4662# 0.14fF
C819 VSS a_1274_4028# 0.36fF
C820 a_9050_n3907# a_9404_n4639# 0.00fF
C821 w_13944_2945# a_14683_966# 0.04fF
C822 w_19623_n3268# a_21735_n1093# 0.00fF
C823 a_24346_n4830# VSS 0.38fF
C824 w_7410_2950# a_7550_4662# 0.02fF
C825 a_2904_n3929# a_2492_n3903# 0.16fF
C826 A[7] Y[6] 0.01fF
C827 a_22849_4533# a_22967_4533# 1.20fF
C828 B[7] carry_in 0.01fF
C829 w_10863_4476# VSS 0.14fF
C830 a_19659_n3206# B[5] 0.00fF
C831 VDD w_21566_n1712# 0.52fF
C832 w_9721_4472# A[1] 0.01fF
C833 a_21246_2574# a_23991_4537# 0.20fF
C834 w_16255_4467# B[2] 0.00fF
C835 w_23612_n1001# w_23598_n2651# 0.01fF
C836 a_14140_n1066# a_15222_n1096# 0.01fF
C837 a_15576_n1096# a_17179_n2618# 0.03fF
C838 w_13939_1341# a_16225_965# 0.00fF
C839 w_21965_2332# a_22002_2394# 0.26fF
C840 w_21965_2332# a_23113_3950# 0.01fF
C841 a_14005_n1722# a_14080_n1092# 0.14fF
C842 B[0] a_2484_n1097# 0.00fF
C843 w_7405_1346# VSS 0.20fF
C844 a_15282_n1070# w_15053_n1715# 0.09fF
C845 w_4007_n1005# B[7] 0.13fF
C846 w_3998_n4259# a_4736_n3230# 0.00fF
C847 w_819_n1712# a_913_n1723# 0.22fF
C848 a_22002_2394# a_22783_969# 0.00fF
C849 a_20651_1407# a_20888_770# 0.38fF
C850 a_4750_n1580# VSS 0.38fF
C851 w_7377_n1716# a_7471_n1727# 0.22fF
C852 w_8519_n1720# a_7606_n1071# 0.01fF
C853 w_7396_4600# B[1] 0.14fF
C854 a_9042_n1101# A[1] 0.00fF
C855 a_21241_970# a_20888_770# 0.00fF
C856 w_897_2953# A[0] 0.07fF
C857 a_8140_4225# A[1] 0.01fF
C858 a_10021_3951# VSS 0.37fF
C859 a_4722_1705# Y[0] 2.33fF
C860 w_18_n3272# A[7] 0.59fF
C861 a_22967_4533# a_21232_4224# 0.04fF
C862 a_8140_4225# w_7410_2950# 0.01fF
C863 a_10659_n973# B[6] 0.09fF
C864 a_11017_4538# a_8154_2575# 0.04fF
C865 a_10659_n973# a_8748_n1075# 0.00fF
C866 a_14098_3007# VSS 0.25fF
C867 a_7564_3012# A[1] 0.06fF
C868 VDD A[5] 1.30fF
C869 w_7410_2950# a_7564_3012# 0.13fF
C870 a_23706_n965# w_21566_n1712# 0.00fF
C871 w_3208_4475# B[0] 0.00fF
C872 w_13110_n3271# a_15147_n1726# 0.02fF
C873 a_8688_n1101# a_8910_2395# 0.00fF
C874 a_4295_2398# Y[0] 0.10fF
C875 a_4722_1705# a_4840_973# 0.01fF
C876 a_17833_n4833# VDD 0.01fF
C877 a_7564_n3933# VSS 0.48fF
C878 a_7564_n3933# A[6] 0.04fF
C879 a_20642_4661# VDD 1.42fF
C880 a_22089_n1093# a_22097_n3899# 0.05fF
C881 a_20593_n1089# A[3] 0.00fF
C882 VDD a_20879_4024# 0.02fF
C883 a_4386_4541# VDD 0.28fF
C884 a_8149_971# a_8154_2575# 0.12fF
C885 a_1636_974# w_897_2953# 0.04fF
C886 a_9462_n3933# VDD 0.83fF
C887 a_4295_2398# a_4840_973# 0.02fF
C888 a_15044_n3209# VSS 0.43fF
C889 A[7] a_594_n3903# 0.02fF
C890 w_22813_4471# A[3] 0.01fF
C891 a_2130_n1097# a_3236_1679# 0.00fF
C892 a_19659_n3206# Y[4] 0.16fF
C893 a_2610_n4635# VDD 0.00fF
C894 a_22002_2394# VDD 0.81fF
C895 VDD a_23113_3950# 1.33fF
C896 w_7377_n1716# A[7] 0.00fF
C897 a_15938_n4634# a_14041_n3235# 0.36fF
C898 VDD a_7270_n4639# 0.00fF
C899 w_17085_n2654# a_17184_n4222# 0.00fF
C900 w_21566_n1712# a_20593_n1089# 0.24fF
C901 w_13911_n1711# a_14434_n1092# 0.12fF
C902 a_913_n1723# a_2190_n1071# 0.02fF
C903 a_22215_n4631# B[4] 0.09fF
C904 w_7377_n1716# a_7796_771# 0.00fF
C905 w_15407_2328# w_17397_4471# 0.01fF
C906 a_15989_1697# A[2] 0.20fF
C907 w_13944_2945# a_14093_1403# 0.00fF
C908 w_19623_n3268# a_22215_n4631# 0.02fF
C909 a_17828_n3229# a_17184_n4222# 0.01fF
C910 a_20611_n3925# a_21557_n3206# 0.23fF
C911 a_1006_n3929# a_712_n4635# 0.02fF
C912 a_1952_n3210# a_4092_n4223# 0.00fF
C913 a_20199_n3899# a_22097_n3899# 0.02fF
C914 a_22841_1675# a_21241_970# 0.01fF
C915 a_11235_1702# a_8910_2395# 0.00fF
C916 a_10808_2395# a_9337_1702# 0.02fF
C917 a_22841_1675# a_20651_1407# 0.00fF
C918 a_8149_971# a_7900_n1097# 0.00fF
C919 w_20424_n1708# a_20947_n1089# 0.12fF
C920 a_2846_n4635# a_1952_n3210# 0.00fF
C921 a_2610_n4635# a_2492_n3903# 0.01fF
C922 a_21735_n1093# a_20947_n1089# 0.04fF
C923 a_21735_n1093# a_22783_969# 0.00fF
C924 a_14005_n1722# w_13911_n1711# 0.22fF
C925 a_14140_n1066# w_15053_n1715# 0.01fF
C926 a_20651_1407# a_21241_970# 0.14fF
C927 a_2942_973# Y[0] 0.00fF
C928 w_3998_n4259# a_4092_n4223# 0.13fF
C929 w_21566_n1712# A[4] 0.01fF
C930 w_23612_n1001# a_24445_969# 0.00fF
C931 w_6576_n3276# VDD 1.02fF
C932 a_22849_4533# VSS 0.65fF
C933 a_13804_n4634# a_15702_n4634# 0.01fF
C934 VDD Y[1] 0.08fF
C935 A[1] Y[0] 0.01fF
C936 a_3362_4537# VSS 0.05fF
C937 w_3998_n4259# a_2846_n4635# 0.00fF
C938 w_13110_n3271# a_13146_n3209# 0.20fF
C939 a_15222_n1096# VDD 0.97fF
C940 w_892_1349# a_1288_2378# 0.00fF
C941 a_20653_n1063# A[3] 0.00fF
C942 a_4840_973# a_2942_973# 0.01fF
C943 a_4722_1705# A[0] 0.02fF
C944 a_4101_n969# a_2190_n1071# 0.00fF
C945 a_17184_n4222# VSS 0.31fF
C946 a_5076_973# VDD 0.00fF
C947 w_1961_n1716# a_988_n1093# 0.24fF
C948 a_10808_2395# a_9691_970# 0.00fF
C949 a_4840_973# A[1] 0.00fF
C950 a_22089_n1093# a_24346_n4830# 0.00fF
C951 a_2130_n1097# VSS 0.49fF
C952 a_9042_n1101# a_10650_n4227# 0.14fF
C953 w_23955_4475# a_22849_4533# 0.01fF
C954 a_20893_2374# VSS 0.37fF
C955 w_22813_4471# a_20642_4661# 0.00fF
C956 a_21232_4224# VSS 0.39fF
C957 carry_out VSS 0.28fF
C958 Y[3] A[3] 0.01fF
C959 A[1] a_8154_2575# 0.07fF
C960 w_7410_2950# a_8154_2575# 0.05fF
C961 a_4295_2398# A[0] 0.04fF
C962 a_14688_2570# a_14098_3007# 0.11fF
C963 a_23900_2394# VSS 0.47fF
C964 B[6] a_13146_n3209# 0.00fF
C965 w_19623_n3268# B[4] 0.40fF
C966 B[6] a_9404_n4639# 0.00fF
C967 w_10565_n1009# a_7900_n1097# 0.00fF
C968 a_7471_n1727# a_8688_n1101# 0.01fF
C969 a_9042_n1101# a_7546_n1097# 0.03fF
C970 w_21566_n1712# a_20653_n1063# 0.01fF
C971 a_7801_2375# a_7796_771# 0.00fF
C972 w_20424_n1708# VDD 0.67fF
C973 a_24681_969# a_22547_1701# 0.00fF
C974 a_21735_n1093# VDD 0.97fF
C975 w_22813_4471# a_23113_3950# 0.23fF
C976 w_23955_4475# a_21232_4224# 0.02fF
C977 a_15282_n1070# a_14140_n1066# 0.01fF
C978 w_7396_4600# a_7787_4025# 0.00fF
C979 w_17397_4471# a_17433_4533# 0.21fF
C980 w_17397_4471# a_16291_4529# 0.01fF
C981 a_14040_n4634# Y[5] 0.36fF
C982 a_15989_1697# a_14683_966# 0.04fF
C983 w_13930_4595# a_16409_4529# 0.00fF
C984 a_1048_n1067# carry_in 0.02fF
C985 a_6612_n3214# VDD 0.69fF
C986 a_7564_n3933# Y[6] 0.10fF
C987 a_15996_n3928# a_15044_n3209# 0.07fF
C988 a_14080_n1092# VSS 0.44fF
C989 a_16225_965# a_15222_n1096# 0.00fF
C990 w_13110_n3271# a_14434_n1092# 0.12fF
C991 A[7] a_4741_n4834# 0.01fF
C992 w_7405_1346# a_9749_1676# 0.00fF
C993 w_13944_2945# B[2] 0.29fF
C994 a_9050_n3907# a_10645_n2623# 0.00fF
C995 VDD a_14041_n3235# 0.25fF
C996 a_13804_n4634# a_14098_n3928# 0.02fF
C997 a_8910_2395# a_9337_1702# 0.19fF
C998 a_20518_n1719# w_21566_n1712# 0.03fF
C999 a_20651_1407# Y[2] 0.00fF
C1000 w_10565_n1009# a_11353_970# 0.00fF
C1001 a_988_n1093# a_1046_1411# 0.00fF
C1002 a_7606_n1071# a_7471_n1727# 1.19fF
C1003 a_23706_n965# a_21735_n1093# 0.12fF
C1004 a_2942_973# A[0] 0.11fF
C1005 w_8873_2333# VDD 0.92fF
C1006 a_1283_774# B[0] 0.00fF
C1007 a_10021_3951# a_9749_1676# 0.00fF
C1008 B[1] VSS 0.78fF
C1009 a_2824_1705# B[0] 0.12fF
C1010 a_3244_4537# w_883_4603# 0.01fF
C1011 w_13110_n3271# a_14005_n1722# 0.05fF
C1012 B[0] VDD 1.07fF
C1013 a_22849_4533# a_24109_4537# 0.00fF
C1014 VDD a_20888_770# 0.01fF
C1015 VDD w_15053_n1715# 0.52fF
C1016 w_21965_2332# a_22841_1675# 0.19fF
C1017 w_7405_1346# w_7377_n1716# 0.00fF
C1018 w_20497_1345# VSS 0.20fF
C1019 a_16283_1671# a_18123_965# 0.00fF
C1020 a_14330_766# a_14140_n1066# 0.00fF
C1021 A[1] a_11353_970# 0.00fF
C1022 w_15407_2328# a_17433_4533# 0.04fF
C1023 w_15407_2328# a_16291_4529# 0.02fF
C1024 a_11589_970# VSS 0.42fF
C1025 w_819_n1712# a_2190_n1071# 0.01fF
C1026 w_21965_2332# a_20651_1407# 0.00fF
C1027 w_21965_2332# a_21241_970# 0.06fF
C1028 a_22841_1675# a_22783_969# 0.00fF
C1029 a_8910_2395# a_9691_970# 0.00fF
C1030 a_20518_n1719# A[5] 0.00fF
C1031 a_21241_970# a_20947_n1089# 0.00fF
C1032 a_20651_1407# a_22783_969# 0.00fF
C1033 a_1636_974# a_2942_973# 0.02fF
C1034 w_8519_n1720# a_9042_n1101# 0.12fF
C1035 a_21241_970# a_22783_969# 0.01fF
C1036 a_1636_974# w_1961_n1716# 0.00fF
C1037 w_20424_n1708# a_20593_n1089# 0.29fF
C1038 a_4736_n3230# VSS 0.37fF
C1039 a_3508_3954# w_2360_2336# 0.01fF
C1040 a_24109_4537# a_21232_4224# 0.01fF
C1041 a_23991_4537# a_23113_3950# 0.15fF
C1042 a_17184_n4222# a_15996_n3928# 0.02fF
C1043 a_21735_n1093# a_20593_n1089# 0.07fF
C1044 a_4386_4541# a_4722_1705# 0.00fF
C1045 a_1288_2378# VSS 0.37fF
C1046 a_21795_n1067# a_20947_n1089# 0.02fF
C1047 a_17179_n2618# A[5] 0.06fF
C1048 B[4] a_20947_n1089# 0.06fF
C1049 a_14330_766# a_14335_2370# 0.00fF
C1050 a_1641_2578# a_2397_2398# 0.03fF
C1051 a_22215_n4631# VDD 0.00fF
C1052 w_19623_n3268# a_20947_n1089# 0.12fF
C1053 a_9050_n3907# VSS 0.24fF
C1054 a_9050_n3907# A[6] 0.22fF
C1055 Y[5] a_13686_n3902# 2.32fF
C1056 w_7405_1346# a_9455_970# 0.00fF
C1057 a_1342_n1093# a_2130_n1097# 0.04fF
C1058 a_2824_1705# a_1051_3015# 0.00fF
C1059 a_4386_4541# a_4295_2398# 0.00fF
C1060 a_23692_n2615# a_24355_n1576# 0.00fF
C1061 VDD a_1051_3015# 1.49fF
C1062 a_7606_n1071# a_7796_771# 0.00fF
C1063 w_15407_2328# a_15989_965# 0.02fF
C1064 a_11647_1676# VDD 0.69fF
C1065 a_20893_2374# a_20656_3011# 0.38fF
C1066 a_21735_n1093# A[4] 0.01fF
C1067 a_15989_1697# a_14093_1403# 0.01fF
C1068 a_20656_3011# a_21232_4224# 0.01fF
C1069 a_1342_n1093# carry_out 0.01fF
C1070 a_1627_4228# w_883_4603# 0.05fF
C1071 a_712_n4635# VDD 0.00fF
C1072 a_14674_4220# a_16409_4529# 0.04fF
C1073 a_17887_965# a_18123_965# 0.04fF
C1074 a_20893_2374# B[3] 0.03fF
C1075 a_18123_965# VSS 0.42fF
C1076 A[7] carry_in 0.01fF
C1077 a_19659_n3206# A[5] 0.01fF
C1078 B[3] a_21232_4224# 0.01fF
C1079 w_10863_4476# A[2] 0.00fF
C1080 w_13911_n1711# VSS 0.22fF
C1081 a_1046_1411# A[0] 0.22fF
C1082 a_9337_1702# a_9757_4534# 0.01fF
C1083 w_13911_n1711# A[6] 0.00fF
C1084 a_23900_2394# B[3] 0.00fF
C1085 VDD a_2484_n1097# 1.32fF
C1086 a_20611_n3925# Y[4] 0.10fF
C1087 a_15282_n1070# VDD 1.32fF
C1088 a_4087_n2619# a_2484_n1097# 0.03fF
C1089 a_11294_n3234# VDD 0.03fF
C1090 a_11308_n1584# a_10645_n2623# 0.00fF
C1091 a_22841_1675# VDD 0.71fF
C1092 w_4007_n1005# A[7] 0.07fF
C1093 VDD a_9168_n4639# 0.00fF
C1094 w_7405_1346# a_7801_2375# 0.00fF
C1095 a_20651_1407# VDD 1.38fF
C1096 a_15147_n1726# a_14434_n1092# 0.04fF
C1097 a_16409_4529# VDD 1.31fF
C1098 a_7900_n1097# a_10650_n4227# 0.01fF
C1099 a_2484_n1097# a_2055_n1727# 0.08fF
C1100 a_21241_970# VDD 1.34fF
C1101 a_20593_n1089# a_20888_770# 0.00fF
C1102 w_18_n3272# a_2130_n1097# 0.00fF
C1103 w_883_4603# a_1274_4028# 0.00fF
C1104 w_897_2953# B[0] 0.29fF
C1105 a_20611_n3925# a_22509_n3925# 0.00fF
C1106 a_1952_n3210# a_948_n4635# 0.00fF
C1107 a_1006_n3929# VDD 0.78fF
C1108 a_9042_n1101# a_8910_2395# 0.00fF
C1109 a_1636_974# a_1046_1411# 0.14fF
C1110 w_18_n3272# carry_out 0.03fF
C1111 w_20424_n1708# a_20653_n1063# 0.08fF
C1112 a_7546_n1097# a_7900_n1097# 0.49fF
C1113 VDD B[4] 0.88fF
C1114 w_17090_n4258# a_15702_n4634# 0.00fF
C1115 a_14084_4657# a_16409_4529# 0.00fF
C1116 a_21795_n1067# VDD 1.32fF
C1117 a_16409_4529# a_17551_4533# 0.01fF
C1118 a_21735_n1093# a_20653_n1063# 0.01fF
C1119 a_16291_4529# a_17433_4533# 0.01fF
C1120 a_14098_3007# A[2] 0.06fF
C1121 a_14005_n1722# a_15147_n1726# 0.01fF
C1122 a_2492_n3903# a_2484_n1097# 0.05fF
C1123 a_7564_3012# a_8910_2395# 0.00fF
C1124 w_3208_4475# VDD 0.53fF
C1125 a_10808_2395# a_8154_2575# 0.00fF
C1126 a_20553_n4631# VSS 0.42fF
C1127 w_13930_4595# a_14321_4020# 0.00fF
C1128 w_19623_n3268# VDD 1.02fF
C1129 a_4722_1705# a_5076_973# 0.00fF
C1130 a_4386_4541# A[1] 0.00fF
C1131 a_15222_n1096# a_17179_n2618# 0.01fF
C1132 a_3244_4537# w_2360_2336# 0.02fF
C1133 w_4350_4479# a_1636_974# 0.00fF
C1134 a_14330_766# VDD 0.01fF
C1135 a_1006_n3929# a_2492_n3903# 0.02fF
C1136 a_4295_2398# a_5076_973# 0.00fF
C1137 w_15407_2328# a_15444_2390# 0.26fF
C1138 a_4092_n4223# VSS 0.31fF
C1139 carry_out a_594_n3903# 0.00fF
C1140 a_11308_n1584# VSS 0.38fF
C1141 a_11308_n1584# A[6] 0.00fF
C1142 w_13110_n3271# a_17828_n3229# 0.00fF
C1143 a_2846_n4635# VSS 0.42fF
C1144 a_20553_n4631# a_20317_n4631# 0.04fF
C1145 a_16555_3946# w_17397_4471# 0.29fF
C1146 a_14674_4220# w_13930_4595# 0.05fF
C1147 a_22215_n4631# a_23697_n4219# 0.00fF
C1148 a_913_n1723# VSS 0.63fF
C1149 a_21795_n1067# a_23706_n965# 0.00fF
C1150 B[6] a_10645_n2623# 0.18fF
C1151 a_7506_n4639# A[6] 0.00fF
C1152 w_20497_1345# a_20656_3011# 0.03fF
C1153 w_3998_n4259# a_1952_n3210# 0.00fF
C1154 w_7405_1346# a_5134_1679# 0.00fF
C1155 a_7506_n4639# VSS 0.42fF
C1156 w_20502_2949# a_20893_2374# 0.00fF
C1157 a_9757_4534# a_7550_4662# 0.01fF
C1158 a_23706_n965# B[4] 0.09fF
C1159 w_20502_2949# a_21232_4224# 0.01fF
C1160 VDD a_8613_n1731# 0.19fF
C1161 w_20424_n1708# a_20518_n1719# 0.22fF
C1162 w_21965_2332# a_22783_969# 0.00fF
C1163 a_7787_4025# VSS 0.37fF
C1164 a_24341_n3226# a_23692_n2615# 0.38fF
C1165 a_14335_2370# a_14321_4020# 0.00fF
C1166 w_897_2953# a_1051_3015# 0.13fF
C1167 a_20518_n1719# a_21735_n1093# 0.01fF
C1168 a_24739_1675# VSS 0.41fF
C1169 w_892_1349# w_819_n1712# 0.00fF
C1170 w_9721_4472# a_9757_4534# 0.20fF
C1171 w_20497_1345# B[3] 0.17fF
C1172 a_22215_n4631# A[4] 0.10fF
C1173 a_15147_n1726# a_17193_n968# 0.01fF
C1174 a_15938_n4634# VDD 0.00fF
C1175 w_13930_4595# VDD 0.39fF
C1176 a_15989_1697# B[2] 0.17fF
C1177 a_20653_n1063# a_20888_770# 0.00fF
C1178 a_24341_n3226# a_24355_n1576# 0.00fF
C1179 w_17090_n4258# B[5] 0.17fF
C1180 a_8510_n3214# a_10650_n4227# 0.00fF
C1181 a_1342_n1093# a_4736_n3230# 0.00fF
C1182 a_21241_970# a_20593_n1089# 0.00fF
C1183 a_10659_n973# a_10645_n2623# 0.01fF
C1184 a_14140_n1066# VDD 1.34fF
C1185 a_20651_1407# a_20593_n1089# 0.00fF
C1186 w_22813_4471# a_22841_1675# 0.00fF
C1187 w_13110_n3271# A[6] 0.01fF
C1188 w_13110_n3271# VSS 0.34fF
C1189 w_22813_4471# a_21241_970# 0.12fF
C1190 w_13930_4595# a_14084_4657# 0.12fF
C1191 a_7546_n1097# a_8510_n3214# 0.00fF
C1192 a_23900_2394# a_22547_1701# 0.62fF
C1193 a_8140_4225# a_9757_4534# 0.16fF
C1194 w_8519_n1720# a_7900_n1097# 0.10fF
C1195 VDD Y[2] 0.08fF
C1196 a_9050_n3907# Y[6] 0.00fF
C1197 A[1] Y[1] 0.01fF
C1198 a_9749_1676# B[1] 0.01fF
C1199 a_4101_n969# VSS 0.24fF
C1200 w_10863_4476# a_11235_1702# 0.00fF
C1201 a_21795_n1067# a_20593_n1089# 0.13fF
C1202 a_1627_4228# w_2360_2336# 0.00fF
C1203 w_8873_2333# a_8149_971# 0.06fF
C1204 a_14098_3007# a_14683_966# 0.03fF
C1205 w_15407_2328# a_16555_3946# 0.01fF
C1206 w_892_1349# a_1641_2578# 0.01fF
C1207 w_19623_n3268# a_20593_n1089# 0.01fF
C1208 a_14335_2370# VDD 0.02fF
C1209 a_10808_2395# a_11353_970# 0.02fF
C1210 a_9749_1676# a_11589_970# 0.00fF
C1211 w_17090_n4258# a_15576_n1096# 0.08fF
C1212 a_23697_n4219# B[4] 0.03fF
C1213 a_14040_n4634# a_14098_n3928# 0.00fF
C1214 carry_in a_1274_4028# 0.00fF
C1215 a_948_n4635# Y[7] 0.36fF
C1216 w_18_n3272# a_4736_n3230# 0.00fF
C1217 B[7] a_2904_n3929# 0.56fF
C1218 w_19623_n3268# a_23697_n4219# 0.00fF
C1219 B[6] VSS 0.77fF
C1220 w_892_1349# a_2397_2398# 0.04fF
C1221 a_7471_n1727# a_9042_n1101# 0.01fF
C1222 a_21557_n3206# a_22097_n3899# 0.16fF
C1223 a_8748_n1075# VSS 0.08fF
C1224 w_21965_2332# VDD 0.93fF
C1225 B[6] A[6] 1.71fF
C1226 B[4] A[4] 1.71fF
C1227 a_3362_4537# w_883_4603# 0.00fF
C1228 a_4295_2398# B[0] 0.00fF
C1229 a_4386_4541# w_4350_4479# 0.21fF
C1230 a_24445_969# a_24681_969# 0.04fF
C1231 a_14674_4220# a_14321_4020# 0.00fF
C1232 a_8910_2395# a_8154_2575# 0.03fF
C1233 w_15407_2328# a_16283_1671# 0.19fF
C1234 w_7405_1346# carry_in 0.00fF
C1235 VDD a_20947_n1089# 1.77fF
C1236 VDD a_22783_969# 0.00fF
C1237 w_19623_n3268# A[4] 0.59fF
C1238 w_17397_4471# VSS 0.14fF
C1239 a_17769_1697# a_18123_965# 0.00fF
C1240 w_20497_1345# w_20502_2949# 0.02fF
C1241 w_13939_1341# w_13944_2945# 0.02fF
C1242 a_10659_n973# VSS 0.23fF
C1243 a_1952_n3210# Y[7] 0.01fF
C1244 a_4750_n1580# carry_in 0.00fF
C1245 a_14321_4020# VDD 0.02fF
C1246 a_10659_n973# A[6] 0.14fF
C1247 a_9875_4534# VDD 1.31fF
C1248 w_17090_n4258# Y[4] 0.00fF
C1249 a_13804_n4634# A[5] 0.00fF
C1250 w_4007_n1005# a_4750_n1580# 0.00fF
C1251 a_22841_1675# Y[3] 0.01fF
C1252 a_9462_n3933# a_10650_n4227# 0.02fF
C1253 a_7152_n3907# VSS 0.21fF
C1254 a_14005_n1722# a_14434_n1092# 0.15fF
C1255 a_14080_n1092# A[2] 0.00fF
C1256 a_7152_n3907# A[6] 0.02fF
C1257 a_14084_4657# a_14321_4020# 0.38fF
C1258 a_9455_970# B[1] 0.09fF
C1259 a_21241_970# a_23991_4537# 0.01fF
C1260 a_23706_n965# a_20947_n1089# 0.00fF
C1261 a_21795_n1067# a_20653_n1063# 0.01fF
C1262 w_20497_1345# a_22547_1701# 0.01fF
C1263 a_15576_n1096# a_15989_1697# 0.00fF
C1264 w_23603_n4255# a_22097_n3899# 0.02fF
C1265 a_14674_4220# VDD 0.97fF
C1266 a_15989_965# a_15444_2390# 0.02fF
C1267 w_8519_n1720# a_8510_n3214# 0.00fF
C1268 a_1641_2578# a_3236_1679# 0.02fF
C1269 a_1342_n1093# a_4092_n4223# 0.01fF
C1270 a_4092_n4223# Y[6] 0.00fF
C1271 Y[5] a_15044_n3209# 0.01fF
C1272 a_1048_n1067# a_988_n1093# 0.05fF
C1273 a_948_n4635# a_54_n3210# 0.00fF
C1274 a_1342_n1093# a_913_n1723# 0.15fF
C1275 a_2397_2398# a_3236_1679# 0.08fF
C1276 w_15407_2328# a_17887_965# 0.02fF
C1277 a_2824_1705# VDD 2.55fF
C1278 a_2942_973# B[0] 0.09fF
C1279 w_15407_2328# VSS 0.34fF
C1280 w_8873_2333# A[1] 0.60fF
C1281 a_1283_774# VDD 0.02fF
C1282 VDD a_4087_n2619# 1.48fF
C1283 a_15147_n1726# VSS 0.66fF
C1284 a_14674_4220# a_17551_4533# 0.01fF
C1285 a_7506_n4639# Y[6] 0.36fF
C1286 a_16555_3946# a_17433_4533# 0.15fF
C1287 w_819_n1712# VSS 0.16fF
C1288 a_7801_2375# B[1] 0.03fF
C1289 a_22547_969# VSS 0.68fF
C1290 a_14674_4220# a_14084_4657# 0.10fF
C1291 a_16555_3946# a_16291_4529# 0.08fF
C1292 a_14098_3007# a_14093_1403# 0.01fF
C1293 a_13686_n3902# a_14098_n3928# 0.16fF
C1294 a_18181_1671# A[3] 0.01fF
C1295 a_20199_n3899# a_20553_n4631# 0.00fF
C1296 VDD a_2055_n1727# 0.19fF
C1297 a_8154_2575# a_9757_4534# 0.04fF
C1298 w_6576_n3276# a_10650_n4227# 0.00fF
C1299 w_13110_n3271# a_15996_n3928# 0.25fF
C1300 a_17193_n968# a_14434_n1092# 0.00fF
C1301 w_7405_1346# a_9337_1702# 0.01fF
C1302 a_20947_n1089# a_20593_n1089# 0.49fF
C1303 a_17551_4533# VDD 1.35fF
C1304 w_18_n3272# a_4092_n4223# 0.00fF
C1305 a_1952_n3210# a_54_n3210# 0.00fF
C1306 a_14084_4657# VDD 1.41fF
C1307 a_21795_n1067# a_20518_n1719# 0.02fF
C1308 B[7] a_2610_n4635# 0.09fF
C1309 w_19623_n3268# a_20518_n1719# 0.05fF
C1310 w_18_n3272# a_2846_n4635# 0.00fF
C1311 w_6576_n3276# a_7546_n1097# 0.01fF
C1312 a_16291_4529# a_16283_1671# 0.00fF
C1313 a_2492_n3903# a_4087_n2619# 0.00fF
C1314 w_18_n3272# a_913_n1723# 0.05fF
C1315 a_23697_n4219# a_20947_n1089# 0.01fF
C1316 w_3993_n2655# a_2484_n1097# 0.04fF
C1317 a_2492_n3903# VDD 2.56fF
C1318 a_10021_3951# a_9337_1702# 0.00fF
C1319 a_1342_n1093# a_4101_n969# 0.00fF
C1320 a_23706_n965# VDD 1.42fF
C1321 a_2492_n3903# a_2055_n1727# 0.01fF
C1322 A[4] a_20947_n1089# 0.07fF
C1323 a_22451_n4631# VSS 0.42fF
C1324 w_20488_4599# a_22967_4533# 0.00fF
C1325 a_1641_2578# VSS 0.87fF
C1326 a_14688_2570# w_17397_4471# 0.12fF
C1327 w_7405_1346# a_9691_970# 0.00fF
C1328 a_23692_n2615# VSS 0.26fF
C1329 a_14080_n1092# a_14683_966# 0.00fF
C1330 a_11647_1676# A[1] 0.00fF
C1331 w_23603_n4255# a_24346_n4830# 0.00fF
C1332 a_7559_1408# VSS 0.30fF
C1333 a_2130_n1097# carry_in 0.07fF
C1334 a_16225_965# VDD 0.00fF
C1335 a_2397_2398# VSS 0.48fF
C1336 a_948_n4635# VSS 0.42fF
C1337 w_6576_n3276# B[7] 0.00fF
C1338 a_5134_1679# B[1] 0.00fF
C1339 a_8688_n1101# B[1] 0.00fF
C1340 a_24355_n1576# VSS 0.38fF
C1341 a_1048_n1067# A[0] 0.00fF
C1342 a_594_n3903# a_913_n1723# 0.00fF
C1343 w_13911_n1711# A[2] 0.02fF
C1344 a_15989_965# a_16283_1671# 0.02fF
C1345 a_2942_973# a_2484_n1097# 0.00fF
C1346 a_18123_965# A[2] 0.00fF
C1347 w_4007_n1005# a_2130_n1097# 0.06fF
C1348 a_1046_1411# B[0] 0.03fF
C1349 a_13146_n3209# VSS 0.36fF
C1350 w_19623_n3268# a_19659_n3206# 0.20fF
C1351 a_13146_n3209# A[6] 0.01fF
C1352 w_1961_n1716# a_2484_n1097# 0.12fF
C1353 a_2190_n1071# VSS 0.08fF
C1354 a_9404_n4639# A[6] 0.00fF
C1355 a_2130_n1097# a_3178_973# 0.00fF
C1356 a_9404_n4639# VSS 0.42fF
C1357 a_4736_n3230# a_4741_n4834# 0.00fF
C1358 VDD a_20593_n1089# 1.33fF
C1359 a_10808_2395# Y[1] 0.10fF
C1360 a_7471_n1727# a_7900_n1097# 0.15fF
C1361 a_17433_4533# VSS 0.62fF
C1362 a_16291_4529# VSS 0.65fF
C1363 A[7] a_4840_973# 0.00fF
C1364 a_988_n1093# A[7] 0.00fF
C1365 a_20947_n1089# a_20653_n1063# 0.04fF
C1366 w_897_2953# VDD 0.37fF
C1367 a_23697_n4219# VDD 1.36fF
C1368 w_22813_4471# VDD 0.53fF
C1369 a_1952_n3210# VSS 0.43fF
C1370 w_21965_2332# Y[3] 0.15fF
C1371 w_9721_4472# w_10863_4476# 0.03fF
C1372 w_15407_2328# a_14688_2570# 0.14fF
C1373 w_17085_n2654# a_14434_n1092# 0.05fF
C1374 w_21965_2332# a_23991_4537# 0.04fF
C1375 w_17397_4471# a_17769_1697# 0.00fF
C1376 a_21660_n1723# VSS 0.66fF
C1377 a_7152_n3907# Y[6] 2.32fF
C1378 w_10556_n4263# a_9050_n3907# 0.02fF
C1379 VDD A[4] 1.25fF
C1380 a_14098_3007# B[2] 0.18fF
C1381 w_3998_n4259# VSS 0.21fF
C1382 a_17828_n3229# a_14434_n1092# 0.00fF
C1383 a_8688_n1101# a_9050_n3907# 0.00fF
C1384 a_13804_n4634# a_14041_n3235# 0.09fF
C1385 w_16255_4467# a_16409_4529# 0.08fF
C1386 a_24739_1675# a_22547_1701# 0.01fF
C1387 a_3244_4537# a_1037_4665# 0.01fF
C1388 a_22097_n3899# Y[4] 0.00fF
C1389 w_10565_n1009# a_8613_n1731# 0.01fF
C1390 a_3508_3954# A[0] 0.00fF
C1391 w_9721_4472# a_10021_3951# 0.23fF
C1392 w_10863_4476# a_8140_4225# 0.02fF
C1393 a_17342_2390# Y[2] 0.10fF
C1394 a_9875_4534# a_11017_4538# 0.01fF
C1395 a_15989_965# a_17887_965# 0.01fF
C1396 a_15989_965# VSS 0.68fF
C1397 a_54_n3210# Y[7] 0.16fF
C1398 a_1046_1411# a_1051_3015# 0.01fF
C1399 w_13939_1341# a_15989_1697# 0.01fF
C1400 a_11235_1702# a_11589_970# 0.00fF
C1401 w_15407_2328# B[3] 0.00fF
C1402 a_15702_n4634# a_15044_n3209# 0.02fF
C1403 B[7] a_6612_n3214# 0.00fF
C1404 a_20518_n1719# a_20947_n1089# 0.15fF
C1405 a_1342_n1093# w_819_n1712# 0.12fF
C1406 a_22089_n1093# a_22547_969# 0.00fF
C1407 carry_in B[1] 0.00fF
C1408 a_22097_n3899# a_22509_n3925# 0.16fF
C1409 w_23612_n1001# a_21735_n1093# 0.06fF
C1410 w_892_1349# a_3236_1679# 0.00fF
C1411 w_7405_1346# a_7564_3012# 0.03fF
C1412 a_15444_2390# a_16283_1671# 0.08fF
C1413 a_14434_n1092# VSS 0.87fF
C1414 B[3] a_22547_969# 0.09fF
C1415 a_23706_n965# A[4] 0.14fF
C1416 w_7377_n1716# a_8748_n1075# 0.01fF
C1417 a_3508_3954# a_1636_974# 0.03fF
C1418 a_8140_4225# a_10021_3951# 0.08fF
C1419 a_9875_4534# a_8149_971# 0.05fF
C1420 a_14080_n1092# a_14093_1403# 0.00fF
C1421 w_2360_2336# B[1] 0.00fF
C1422 w_13911_n1711# a_14683_966# 0.00fF
C1423 VDD a_20653_n1063# 1.34fF
C1424 w_15407_2328# a_17769_1697# 0.35fF
C1425 w_20488_4599# VSS 0.10fF
C1426 w_7396_4600# VSS 0.10fF
C1427 a_24341_n3226# VSS 0.37fF
C1428 a_7801_2375# a_7787_4025# 0.00fF
C1429 a_23900_2394# a_24445_969# 0.02fF
C1430 Y[3] VDD 0.07fF
C1431 w_17090_n4258# A[5] 0.13fF
C1432 a_14005_n1722# VSS 0.63fF
C1433 a_14005_n1722# A[6] 0.00fF
C1434 a_23991_4537# VDD 0.28fF
C1435 a_11017_4538# VDD 1.35fF
C1436 w_17090_n4258# a_17833_n4833# 0.00fF
C1437 w_17085_n2654# a_17193_n968# 0.03fF
C1438 a_14040_n4634# A[5] 0.00fF
C1439 w_18_n3272# w_819_n1712# 0.02fF
C1440 w_8873_2333# a_10808_2395# 0.26fF
C1441 w_7377_n1716# a_7152_n3907# 0.00fF
C1442 a_1037_4665# a_1627_4228# 0.10fF
C1443 a_1288_2378# carry_in 0.00fF
C1444 a_22089_n1093# a_22451_n4631# 0.01fF
C1445 a_4092_n4223# a_4741_n4834# 0.38fF
C1446 A[4] a_20593_n1089# 0.00fF
C1447 a_11294_n3234# a_10650_n4227# 0.01fF
C1448 a_14688_2570# a_17433_4533# 0.20fF
C1449 a_22089_n1093# a_23692_n2615# 0.03fF
C1450 w_17099_n1004# a_15147_n1726# 0.01fF
C1451 a_14688_2570# a_16291_4529# 0.04fF
C1452 w_2360_2336# a_1288_2378# 0.00fF
C1453 a_4722_1705# a_2824_1705# 0.02fF
C1454 a_4722_1705# VDD 2.54fF
C1455 a_8149_971# VDD 1.34fF
C1456 a_9168_n4639# a_10650_n4227# 0.00fF
C1457 a_15044_n3209# B[5] 0.01fF
C1458 a_22089_n1093# a_24355_n1576# 0.01fF
C1459 a_15444_2390# VSS 0.48fF
C1460 a_23697_n4219# A[4] 0.18fF
C1461 a_20518_n1719# VDD 0.27fF
C1462 Y[7] VSS 0.21fF
C1463 A[7] a_2904_n3929# 0.07fF
C1464 w_3208_4475# w_4350_4479# 0.03fF
C1465 a_15702_n4634# a_17184_n4222# 0.00fF
C1466 a_11308_n1584# a_8688_n1101# 0.00fF
C1467 a_16555_3946# a_16283_1671# 0.00fF
C1468 a_2824_1705# a_4295_2398# 0.02fF
C1469 a_1342_n1093# a_2190_n1071# 0.02fF
C1470 a_1037_4665# a_1274_4028# 0.38fF
C1471 a_3244_4537# A[0] 0.01fF
C1472 a_4295_2398# VDD 0.77fF
C1473 w_892_1349# VSS 0.17fF
C1474 a_594_n3903# w_819_n1712# 0.00fF
C1475 VDD a_17179_n2618# 1.48fF
C1476 w_7405_1346# Y[0] 0.00fF
C1477 a_17193_n968# VSS 0.23fF
C1478 a_9337_1702# B[1] 0.12fF
C1479 a_24346_n4830# a_22509_n3925# 0.00fF
C1480 a_14098_n3928# a_15044_n3209# 0.23fF
C1481 a_17342_2390# VDD 0.77fF
C1482 a_20611_n3925# a_22215_n4631# 0.01fF
C1483 a_15576_n1096# a_15044_n3209# 0.01fF
C1484 a_1342_n1093# a_1952_n3210# 0.02fF
C1485 a_22967_4533# VSS 0.05fF
C1486 a_20653_n1063# a_20593_n1089# 0.05fF
C1487 w_3993_n2655# VDD 0.37fF
C1488 w_3993_n2655# a_4087_n2619# 0.13fF
C1489 a_10899_4538# VSS 0.62fF
C1490 w_18_n3272# a_948_n4635# 0.00fF
C1491 w_10863_4476# a_8154_2575# 0.12fF
C1492 a_21660_n1723# a_22089_n1093# 0.08fF
C1493 a_4386_4541# a_3508_3954# 0.15fF
C1494 a_3244_4537# a_1636_974# 0.07fF
C1495 B[7] a_2484_n1097# 0.13fF
C1496 a_9749_1676# a_7559_1408# 0.00fF
C1497 a_17769_1697# a_17433_4533# 0.00fF
C1498 w_7405_1346# a_8154_2575# 0.01fF
C1499 w_3998_n4259# a_1342_n1093# 0.01fF
C1500 a_19659_n3206# VDD 0.69fF
C1501 a_10808_2395# a_11647_1676# 0.08fF
C1502 w_3998_n4259# Y[6] 0.00fF
C1503 a_14093_1403# w_13911_n1711# 0.00fF
C1504 a_22547_1701# a_22547_969# 0.43fF
C1505 w_10565_n1009# VDD 0.38fF
C1506 a_9691_970# B[1] 0.00fF
C1507 a_10021_3951# a_8154_2575# 0.48fF
C1508 a_17828_n3229# w_17085_n2654# 0.00fF
C1509 a_1636_974# a_4504_4541# 0.00fF
C1510 a_15996_n3928# a_14434_n1092# 0.03fF
C1511 a_16555_3946# VSS 0.37fF
C1512 a_13686_n3902# A[5] 0.02fF
C1513 w_22813_4471# a_23991_4537# 0.03fF
C1514 a_17184_n4222# B[5] 0.03fF
C1515 w_23955_4475# a_22967_4533# 0.01fF
C1516 w_18_n3272# a_1952_n3210# 0.19fF
C1517 B[7] a_1006_n3929# 0.00fF
C1518 a_24681_969# A[3] 0.00fF
C1519 w_10556_n4263# B[6] 0.17fF
C1520 a_54_n3210# VSS 0.33fF
C1521 a_948_n4635# a_594_n3903# 0.00fF
C1522 a_2824_1705# a_2942_973# 0.01fF
C1523 a_1627_4228# A[0] 0.01fF
C1524 w_15407_2328# A[2] 0.60fF
C1525 w_7377_n1716# a_7559_1408# 0.00fF
C1526 a_2942_973# VDD 0.01fF
C1527 w_1961_n1716# VDD 0.54fF
C1528 a_3236_1679# VSS 0.45fF
C1529 a_8688_n1101# B[6] 0.01fF
C1530 B[6] a_11299_n4838# 0.00fF
C1531 a_7546_n1097# a_8613_n1731# 0.09fF
C1532 a_8688_n1101# a_8748_n1075# 0.05fF
C1533 carry_in a_913_n1723# 0.01fF
C1534 VDD A[1] 1.46fF
C1535 w_3998_n4259# w_18_n3272# 0.00fF
C1536 a_10645_n2623# VSS 0.26fF
C1537 a_10645_n2623# A[6] 0.06fF
C1538 a_20518_n1719# a_20593_n1089# 0.14fF
C1539 a_16225_965# a_17342_2390# 0.00fF
C1540 w_7410_2950# VDD 0.37fF
C1541 a_17887_965# a_16283_1671# 0.01fF
C1542 w_8873_2333# a_8910_2395# 0.26fF
C1543 a_16283_1671# VSS 0.46fF
C1544 a_20611_n3925# B[4] 0.00fF
C1545 w_20488_4599# a_20656_3011# 0.00fF
C1546 w_19623_n3268# a_20611_n3925# 0.26fF
C1547 w_1961_n1716# a_2055_n1727# 0.21fF
C1548 a_14674_4220# w_16255_4467# 0.21fF
C1549 w_23612_n1001# a_21795_n1067# 0.00fF
C1550 w_6576_n3276# a_7471_n1727# 0.05fF
C1551 a_22089_n1093# a_24341_n3226# 0.01fF
C1552 a_15576_n1096# a_17184_n4222# 0.14fF
C1553 w_23612_n1001# B[4] 0.13fF
C1554 w_17085_n2654# VSS 0.17fF
C1555 w_20488_4599# B[3] 0.14fF
C1556 B[1] a_7550_4662# 0.10fF
C1557 A[0] a_1274_4028# 0.00fF
C1558 a_1952_n3210# a_594_n3903# 0.02fF
C1559 a_8688_n1101# a_10659_n973# 0.12fF
C1560 a_15222_n1096# a_15989_1697# 0.00fF
C1561 a_1627_4228# a_1636_974# 0.49fF
C1562 a_14688_2570# a_15444_2390# 0.03fF
C1563 w_9721_4472# B[1] 0.00fF
C1564 a_17828_n3229# VSS 0.37fF
C1565 A[7] a_2610_n4635# 0.10fF
C1566 w_10551_n2659# a_11308_n1584# 0.00fF
C1567 w_16255_4467# VDD 0.53fF
C1568 w_17397_4471# a_14683_966# 0.00fF
C1569 w_13110_n3271# Y[5] 0.15fF
C1570 a_7559_1408# a_9455_970# 0.00fF
C1571 a_21246_2574# a_22849_4533# 0.04fF
C1572 a_7900_n1097# a_7564_n3933# 0.00fF
C1573 w_17090_n4258# a_14041_n3235# 0.01fF
C1574 a_4101_n969# carry_in 0.01fF
C1575 a_9042_n1101# B[1] 0.00fF
C1576 a_7606_n1071# a_8748_n1075# 0.01fF
C1577 a_14040_n4634# a_14041_n3235# 0.00fF
C1578 w_16255_4467# a_14084_4657# 0.00fF
C1579 a_1037_4665# a_3362_4537# 0.00fF
C1580 w_16255_4467# a_17551_4533# 0.01fF
C1581 a_3244_4537# a_4386_4541# 0.01fF
C1582 a_1636_974# a_1274_4028# 0.01fF
C1583 a_8140_4225# B[1] 0.01fF
C1584 a_17184_n4222# Y[4] 0.00fF
C1585 w_4007_n1005# a_4101_n969# 0.13fF
C1586 w_17099_n1004# a_14434_n1092# 0.00fF
C1587 a_22967_4533# a_24109_4537# 0.01fF
C1588 a_20553_n4631# a_21557_n3206# 0.00fF
C1589 a_17887_965# VSS 0.69fF
C1590 a_14080_n1092# a_14098_n3928# 0.00fF
C1591 A[6] VSS 1.73fF
C1592 w_6576_n3276# A[7] 0.01fF
C1593 a_7564_3012# B[1] 0.18fF
C1594 a_1283_774# a_1046_1411# 0.38fF
C1595 a_7559_1408# a_7801_2375# 0.01fF
C1596 a_21246_2574# a_21232_4224# 0.04fF
C1597 a_15576_n1096# a_14080_n1092# 0.03fF
C1598 a_20893_2374# a_21246_2574# 0.00fF
C1599 a_19659_n3206# A[4] 0.00fF
C1600 a_1046_1411# VDD 1.44fF
C1601 a_20518_n1719# a_20653_n1063# 1.19fF
C1602 a_1641_2578# w_883_4603# 0.00fF
C1603 a_4386_4541# a_4504_4541# 1.20fF
C1604 a_23900_2394# a_21246_2574# 0.00fF
C1605 a_15444_2390# a_17769_1697# 0.00fF
C1606 w_13939_1341# a_14098_3007# 0.03fF
C1607 w_8873_2333# a_9757_4534# 0.02fF
C1608 w_8519_n1720# a_8613_n1731# 0.21fF
C1609 w_15407_2328# a_14683_966# 0.06fF
C1610 a_988_n1093# a_2130_n1097# 0.07fF
C1611 a_11017_4538# a_8149_971# 0.00fF
C1612 a_14688_2570# a_16555_3946# 0.48fF
C1613 a_16291_4529# A[2] 0.01fF
C1614 a_988_n1093# carry_out 0.05fF
C1615 w_18_n3272# Y[7] 0.15fF
C1616 w_23955_4475# VSS 0.14fF
C1617 a_20317_n4631# VSS 0.69fF
C1618 w_4350_4479# VDD 0.66fF
C1619 a_24739_1675# a_24445_969# 0.02fF
C1620 w_20502_2949# w_20488_4599# 0.01fF
C1621 w_13944_2945# w_13930_4595# 0.01fF
C1622 w_10551_n2659# B[6] 0.29fF
C1623 a_9042_n1101# a_9050_n3907# 0.05fF
C1624 a_14688_2570# a_16283_1671# 0.02fF
C1625 a_4386_4541# a_1627_4228# 0.01fF
C1626 a_20611_n3925# a_20947_n1089# 0.00fF
C1627 VDD a_10650_n4227# 1.36fF
C1628 a_7564_n3933# a_8510_n3214# 0.23fF
C1629 w_10551_n2659# a_10659_n973# 0.03fF
C1630 a_15989_965# A[2] 0.11fF
C1631 w_17099_n1004# a_17193_n968# 0.13fF
C1632 w_23612_n1001# a_20947_n1089# 0.00fF
C1633 a_594_n3903# Y[7] 2.32fF
C1634 a_4722_1705# a_4295_2398# 0.19fF
C1635 a_7546_n1097# VDD 1.33fF
C1636 a_13804_n4634# VDD 0.00fF
C1637 w_10556_n4263# a_13146_n3209# 0.00fF
C1638 A[7] a_6612_n3214# 0.01fF
C1639 w_13944_2945# a_14335_2370# 0.00fF
C1640 w_10556_n4263# a_9404_n4639# 0.00fF
C1641 a_14041_n3235# a_13686_n3902# 0.10fF
C1642 carry_in w_819_n1712# 0.06fF
C1643 a_1048_n1067# a_2484_n1097# 0.00fF
C1644 a_17828_n3229# a_15996_n3928# 0.00fF
C1645 a_18181_1671# Y[2] 0.15fF
C1646 w_20497_1345# a_21246_2574# 0.01fF
C1647 a_2130_n1097# A[0] 0.00fF
C1648 w_18_n3272# a_54_n3210# 0.20fF
C1649 w_3998_n4259# a_4741_n4834# 0.00fF
C1650 a_16283_1671# a_17769_1697# 0.02fF
C1651 w_897_2953# a_1046_1411# 0.00fF
C1652 B[7] a_4087_n2619# 0.18fF
C1653 a_15576_n1096# w_13911_n1711# 0.00fF
C1654 a_24109_4537# VSS 0.05fF
C1655 a_8154_2575# B[1] 0.07fF
C1656 B[7] VDD 0.91fF
C1657 a_16291_4529# a_14683_966# 0.07fF
C1658 a_14688_2570# VSS 0.87fF
C1659 w_13944_2945# a_14321_4020# 0.00fF
C1660 a_7787_4025# a_7550_4662# 0.38fF
C1661 a_17433_4533# a_14683_966# 0.01fF
C1662 a_3362_4537# a_1636_974# 0.05fF
C1663 a_7606_n1071# a_7559_1408# 0.00fF
C1664 a_21735_n1093# a_22097_n3899# 0.00fF
C1665 w_15407_2328# a_14093_1403# 0.00fF
C1666 w_23598_n2651# a_23692_n2615# 0.13fF
C1667 a_20611_n3925# VDD 0.78fF
C1668 a_22849_4533# A[3] 0.01fF
C1669 w_13110_n3271# a_15702_n4634# 0.02fF
C1670 a_15996_n3928# VSS 0.49fF
C1671 a_10808_2395# VDD 0.77fF
C1672 w_23598_n2651# a_24355_n1576# 0.00fF
C1673 w_23612_n1001# VDD 0.38fF
C1674 a_11308_n1584# a_9042_n1101# 0.01fF
C1675 a_1641_2578# carry_in 0.01fF
C1676 a_4722_1705# A[1] 0.00fF
C1677 a_20656_3011# VSS 0.25fF
C1678 a_8149_971# A[1] 0.17fF
C1679 a_15044_n3209# A[5] 0.80fF
C1680 a_22089_n1093# VSS 1.20fF
C1681 w_23955_4475# a_24109_4537# 0.09fF
C1682 a_54_n3210# a_594_n3903# 0.17fF
C1683 B[7] a_2492_n3903# 0.10fF
C1684 a_15444_2390# A[2] 0.11fF
C1685 a_1342_n1093# VSS 0.87fF
C1686 a_8149_971# w_7410_2950# 0.04fF
C1687 a_1641_2578# w_2360_2336# 0.14fF
C1688 Y[6] VSS 0.22fF
C1689 a_9462_n3933# a_7564_n3933# 0.00fF
C1690 Y[6] A[6] 0.01fF
C1691 a_7559_1408# carry_in 0.00fF
C1692 a_14674_4220# w_13944_2945# 0.01fF
C1693 B[3] VSS 0.78fF
C1694 a_2397_2398# carry_in 0.03fF
C1695 a_8140_4225# a_7787_4025# 0.00fF
C1696 w_17099_n1004# w_17085_n2654# 0.01fF
C1697 a_4295_2398# a_2942_973# 0.01fF
C1698 a_13146_n3209# Y[5] 0.16fF
C1699 a_20893_2374# A[3] 0.01fF
C1700 a_21232_4224# A[3] 0.01fF
C1701 a_15989_965# a_14683_966# 0.02fF
C1702 w_8519_n1720# VDD 0.53fF
C1703 w_2360_2336# a_2397_2398# 0.26fF
C1704 carry_in a_2190_n1071# 0.03fF
C1705 a_7564_3012# a_7787_4025# 0.00fF
C1706 a_23900_2394# A[3] 0.04fF
C1707 a_7564_n3933# a_7270_n4639# 0.02fF
C1708 w_13944_2945# VDD 0.37fF
C1709 a_2397_2398# a_3178_973# 0.00fF
C1710 a_17887_965# a_17769_1697# 0.01fF
C1711 w_17090_n4258# a_15938_n4634# 0.00fF
C1712 a_17769_1697# VSS 0.22fF
C1713 w_4007_n1005# a_2190_n1071# 0.00fF
C1714 w_23612_n1001# a_23706_n965# 0.13fF
C1715 a_24445_969# a_22547_969# 0.01fF
C1716 w_3208_4475# a_3508_3954# 0.23fF
C1717 a_10899_4538# A[2] 0.00fF
C1718 A[7] a_712_n4635# 0.00fF
C1719 w_18_n3272# VSS 0.32fF
C1720 a_14434_n1092# a_14683_966# 0.00fF
C1721 w_13944_2945# a_14084_4657# 0.02fF
C1722 A[7] a_2484_n1097# 0.14fF
C1723 a_20199_n3899# VSS 0.21fF
C1724 w_13110_n3271# B[5] 0.40fF
C1725 a_18181_1671# VDD 0.69fF
C1726 a_20553_n4631# Y[4] 0.36fF
C1727 a_9749_1676# VSS 0.46fF
C1728 w_6576_n3276# a_7564_n3933# 0.26fF
C1729 w_17099_n1004# a_17887_965# 0.00fF
C1730 w_17099_n1004# VSS 0.19fF
C1731 a_22849_4533# a_20642_4661# 0.01fF
C1732 a_7900_n1097# a_9050_n3907# 0.03fF
C1733 a_9042_n1101# B[6] 0.13fF
C1734 a_20611_n3925# a_20593_n1089# 0.00fF
C1735 a_7471_n1727# a_8613_n1731# 0.01fF
C1736 a_9042_n1101# a_8748_n1075# 0.05fF
C1737 A[7] a_1006_n3929# 0.04fF
C1738 a_17184_n4222# A[5] 0.18fF
C1739 a_16555_3946# A[2] 0.00fF
C1740 a_3362_4537# a_4386_4541# 0.02fF
C1741 w_13110_n3271# a_14098_n3928# 0.26fF
C1742 a_17833_n4833# a_17184_n4222# 0.38fF
C1743 a_22451_n4631# a_21557_n3206# 0.00fF
C1744 a_22215_n4631# a_22097_n3899# 0.01fF
C1745 a_594_n3903# VSS 0.21fF
C1746 a_11353_970# a_11589_970# 0.04fF
C1747 a_20199_n3899# a_20317_n4631# 0.01fF
C1748 w_15407_2328# B[2] 0.43fF
C1749 w_13110_n3271# a_15576_n1096# 0.06fF
C1750 a_1627_4228# B[0] 0.01fF
C1751 w_7377_n1716# VSS 0.22fF
C1752 a_1288_2378# A[0] 0.01fF
C1753 w_20502_2949# VSS 0.16fF
C1754 w_23598_n2651# a_24341_n3226# 0.00fF
C1755 a_9042_n1101# a_10659_n973# 0.03fF
C1756 a_22849_4533# a_23113_3950# 0.08fF
C1757 a_20611_n3925# A[4] 0.04fF
C1758 a_20642_4661# a_21232_4224# 0.10fF
C1759 w_7410_2950# A[1] 0.07fF
C1760 a_15444_2390# a_14683_966# 0.10fF
C1761 a_16283_1671# A[2] 0.81fF
C1762 w_4350_4479# a_4722_1705# 0.00fF
C1763 a_8910_2395# VDD 0.81fF
C1764 a_17842_n1579# a_17193_n968# 0.38fF
C1765 a_21232_4224# a_20879_4024# 0.00fF
C1766 a_20893_2374# a_20879_4024# 0.00fF
C1767 w_20497_1345# A[3] 0.19fF
C1768 w_23612_n1001# A[4] 0.07fF
C1769 a_15989_1697# Y[2] 0.18fF
C1770 B[0] a_1274_4028# 0.02fF
C1771 w_8873_2333# w_10863_4476# 0.01fF
C1772 a_988_n1093# a_913_n1723# 0.14fF
C1773 a_22841_1675# a_24681_969# 0.00fF
C1774 a_2904_n3929# a_4736_n3230# 0.00fF
C1775 a_15989_965# a_14093_1403# 0.00fF
C1776 w_7405_1346# w_8873_2333# 0.00fF
C1777 a_20893_2374# a_22002_2394# 0.00fF
C1778 a_1636_974# a_1288_2378# 0.01fF
C1779 a_22547_1701# VSS 0.54fF
C1780 a_21232_4224# a_23113_3950# 0.08fF
C1781 a_14080_n1092# A[5] 0.00fF
C1782 a_7559_1408# a_9691_970# 0.00fF
C1783 a_22002_2394# a_23900_2394# 0.00fF
C1784 a_23900_2394# a_23113_3950# 0.00fF
C1785 w_20497_1345# w_21566_n1712# 0.00fF
C1786 w_13939_1341# w_13911_n1711# 0.00fF
C1787 a_6612_n3214# a_7564_n3933# 0.07fF
C1788 a_9875_4534# a_9757_4534# 1.20fF
C1789 w_3208_4475# a_3244_4537# 0.20fF
C1790 a_9455_970# VSS 0.68fF
C1791 w_23603_n4255# a_22451_n4631# 0.00fF
C1792 a_21660_n1723# a_21557_n3206# 0.00fF
C1793 w_8873_2333# a_10021_3951# 0.01fF
C1794 a_22097_n3899# B[4] 0.10fF
C1795 a_8149_971# a_7546_n1097# 0.00fF
C1796 w_23603_n4255# a_23692_n2615# 0.03fF
C1797 a_1627_4228# a_1051_3015# 0.01fF
C1798 a_8510_n3214# a_9050_n3907# 0.16fF
C1799 a_20656_3011# B[3] 0.18fF
C1800 w_19623_n3268# a_22097_n3899# 0.27fF
C1801 w_10556_n4263# a_10645_n2623# 0.03fF
C1802 a_22089_n1093# B[3] 0.00fF
C1803 w_17090_n4258# VDD 0.33fF
C1804 w_23955_4475# a_22547_1701# 0.01fF
C1805 a_1048_n1067# a_1283_774# 0.00fF
C1806 a_17887_965# A[2] 0.00fF
C1807 VSS A[2] 1.98fF
C1808 a_5134_1679# a_3236_1679# 0.00fF
C1809 w_3208_4475# a_4504_4541# 0.01fF
C1810 a_16555_3946# a_14683_966# 0.03fF
C1811 a_2942_973# a_1046_1411# 0.00fF
C1812 a_1048_n1067# VDD 1.34fF
C1813 a_8688_n1101# a_10645_n2623# 0.01fF
C1814 a_14040_n4634# VDD 0.00fF
C1815 a_7801_2375# VSS 0.37fF
C1816 w_1961_n1716# a_1046_1411# 0.00fF
C1817 w_892_1349# carry_in 0.20fF
C1818 a_14041_n3235# a_15044_n3209# 0.18fF
C1819 a_10899_4538# a_11235_1702# 0.00fF
C1820 a_1048_n1067# a_2055_n1727# 0.00fF
C1821 a_1051_3015# a_1274_4028# 0.00fF
C1822 w_892_1349# w_2360_2336# 0.00fF
C1823 VDD a_9757_4534# 0.19fF
C1824 w_892_1349# a_3178_973# 0.00fF
C1825 w_17085_n2654# a_17842_n1579# 0.00fF
C1826 w_18_n3272# a_1342_n1093# 0.12fF
C1827 w_883_4603# VSS 0.09fF
C1828 w_4350_4479# A[1] 0.00fF
C1829 a_16283_1671# a_14683_966# 0.01fF
C1830 a_17828_n3229# a_17842_n1579# 0.00fF
C1831 a_15044_n3209# w_15053_n1715# 0.00fF
C1832 a_20611_n3925# a_20518_n1719# 0.00fF
C1833 a_15576_n1096# a_15147_n1726# 0.08fF
C1834 a_15444_2390# a_14093_1403# 0.02fF
C1835 w_3208_4475# a_1627_4228# 0.21fF
C1836 a_14080_n1092# a_15222_n1096# 0.07fF
C1837 a_4741_n4834# VSS 0.38fF
C1838 w_20497_1345# a_22002_2394# 0.04fF
C1839 a_3508_3954# a_2824_1705# 0.00fF
C1840 a_7471_n1727# VDD 0.27fF
C1841 a_3508_3954# VDD 1.34fF
C1842 a_15989_1697# VDD 0.23fF
C1843 w_3993_n2655# B[7] 0.29fF
C1844 a_2904_n3929# a_4092_n4223# 0.02fF
C1845 a_7564_3012# a_7559_1408# 0.01fF
C1846 w_10556_n4263# VSS 0.20fF
C1847 w_10556_n4263# A[6] 0.13fF
C1848 a_15989_965# B[2] 0.09fF
C1849 a_4750_n1580# a_2484_n1097# 0.01fF
C1850 a_5134_1679# VSS 0.36fF
C1851 a_8688_n1101# VSS 0.49fF
C1852 a_8149_971# w_8519_n1720# 0.00fF
C1853 a_9042_n1101# a_9404_n4639# 0.01fF
C1854 a_24346_n4830# B[4] 0.00fF
C1855 a_2846_n4635# a_2904_n3929# 0.00fF
C1856 a_8688_n1101# A[6] 0.01fF
C1857 a_11299_n4838# VSS 0.38fF
C1858 w_20502_2949# a_20656_3011# 0.13fF
C1859 a_17842_n1579# VSS 0.38fF
C1860 a_11299_n4838# A[6] 0.01fF
C1861 a_7546_n1097# A[1] 0.00fF
C1862 a_9462_n3933# a_9050_n3907# 0.16fF
C1863 a_7900_n1097# B[6] 0.06fF
C1864 a_3236_1679# carry_in 0.02fF
C1865 a_7900_n1097# a_8748_n1075# 0.02fF
C1866 a_19659_n3206# a_20611_n3925# 0.07fF
C1867 a_17184_n4222# a_14041_n3235# 0.01fF
C1868 w_20502_2949# B[3] 0.29fF
C1869 a_8510_n3214# a_7506_n4639# 0.00fF
C1870 a_7564_n3933# a_9168_n4639# 0.01fF
C1871 VSS a_14683_966# 1.12fF
C1872 w_2360_2336# a_3236_1679# 0.19fF
C1873 a_24739_1675# A[3] 0.00fF
C1874 a_3236_1679# a_3178_973# 0.00fF
C1875 w_23603_n4255# a_24341_n3226# 0.00fF
C1876 w_21965_2332# a_24681_969# 0.00fF
C1877 Y[1] a_11589_970# 0.36fF
C1878 VDD a_13686_n3902# 2.54fF
C1879 a_2130_n1097# B[0] 0.00fF
C1880 w_18_n3272# a_594_n3903# 0.34fF
C1881 a_22097_n3899# a_20947_n1089# 0.03fF
C1882 a_10659_n973# a_7900_n1097# 0.00fF
C1883 a_22089_n1093# a_22547_1701# 0.00fF
C1884 w_1961_n1716# B[7] 0.00fF
C1885 a_13146_n3209# a_14098_n3928# 0.07fF
C1886 a_988_n1093# w_819_n1712# 0.29fF
C1887 A[7] a_4087_n2619# 0.06fF
C1888 a_14688_2570# A[2] 0.07fF
C1889 A[7] VDD 1.30fF
C1890 a_20893_2374# a_20888_770# 0.00fF
C1891 a_22547_1701# B[3] 0.17fF
C1892 w_10551_n2659# a_10645_n2623# 0.13fF
C1893 a_7606_n1071# VSS 0.07fF
C1894 A[7] a_2055_n1727# 0.01fF
C1895 w_7396_4600# a_7550_4662# 0.12fF
C1896 a_7796_771# VDD 0.01fF
C1897 a_16225_965# a_15989_1697# 0.36fF
C1898 w_6576_n3276# a_9050_n3907# 0.27fF
C1899 a_10808_2395# A[1] 0.04fF
C1900 a_11235_1702# VSS 0.22fF
C1901 w_23598_n2651# VSS 0.17fF
C1902 a_17342_2390# a_18181_1671# 0.08fF
C1903 a_16283_1671# a_14093_1403# 0.00fF
C1904 a_1037_4665# a_1641_2578# 0.00fF
C1905 a_14080_n1092# a_14041_n3235# 0.00fF
C1906 w_20497_1345# w_20424_n1708# 0.00fF
C1907 A[7] a_2492_n3903# 0.22fF
C1908 Y[5] VSS 0.22fF
C1909 a_15444_2390# B[2] 0.60fF
C1910 Y[5] A[6] 0.01fF
C1911 a_7559_1408# Y[0] 0.00fF
C1912 a_8149_971# a_8910_2395# 0.10fF
C1913 a_22451_n4631# a_22509_n3925# 0.00fF
C1914 carry_in VSS 1.55fF
C1915 a_3244_4537# a_2824_1705# 0.01fF
C1916 B[5] a_14434_n1092# 0.06fF
C1917 a_3244_4537# VDD 0.19fF
C1918 a_14080_n1092# w_15053_n1715# 0.24fF
C1919 w_7396_4600# a_8140_4225# 0.05fF
C1920 a_23692_n2615# a_22509_n3925# 0.00fF
C1921 w_4007_n1005# VSS 0.22fF
C1922 a_15222_n1096# w_13911_n1711# 0.02fF
C1923 w_2360_2336# VSS 0.34fF
C1924 B[6] a_8510_n3214# 0.01fF
C1925 a_22841_1675# a_22849_4533# 0.00fF
C1926 VDD a_22097_n3899# 2.56fF
C1927 a_17769_1697# A[2] 0.02fF
C1928 a_9749_1676# a_9455_970# 0.02fF
C1929 a_3178_973# VSS 0.42fF
C1930 w_13930_4595# a_14098_3007# 0.00fF
C1931 w_17397_4471# A[3] 0.00fF
C1932 w_7396_4600# a_7564_3012# 0.00fF
C1933 a_15989_965# a_15576_n1096# 0.00fF
C1934 a_21241_970# a_22849_4533# 0.07fF
C1935 a_24681_969# VDD 0.00fF
C1936 a_2610_n4635# a_4092_n4223# 0.00fF
C1937 a_7559_1408# a_8154_2575# 0.01fF
C1938 VDD a_4504_4541# 1.35fF
C1939 w_10551_n2659# A[6] 0.07fF
C1940 w_8873_2333# B[1] 0.43fF
C1941 w_10551_n2659# VSS 0.17fF
C1942 a_2130_n1097# a_2484_n1097# 0.48fF
C1943 a_14098_n3928# a_14434_n1092# 0.00fF
C1944 a_988_n1093# a_2190_n1071# 0.13fF
C1945 a_2610_n4635# a_2846_n4635# 0.04fF
C1946 w_13110_n3271# A[5] 0.59fF
C1947 A[0] w_819_n1712# 0.03fF
C1948 carry_out a_2484_n1097# 0.00fF
C1949 a_15576_n1096# a_14434_n1092# 0.12fF
C1950 a_14093_1403# VSS 0.30fF
C1951 w_13939_1341# w_15407_2328# 0.00fF
C1952 a_7270_n4639# a_7506_n4639# 0.04fF
C1953 a_15938_n4634# a_15044_n3209# 0.00fF
C1954 a_20893_2374# a_20651_1407# 0.01fF
C1955 w_8873_2333# a_11589_970# 0.00fF
C1956 a_22841_1675# a_23900_2394# 0.20fF
C1957 a_6612_n3214# a_9050_n3907# 0.00fF
C1958 a_20893_2374# a_21241_970# 0.01fF
C1959 a_14688_2570# a_14683_966# 0.12fF
C1960 a_7152_n3907# a_8510_n3214# 0.02fF
C1961 a_11017_4538# a_9757_4534# 0.00fF
C1962 w_3208_4475# a_3362_4537# 0.08fF
C1963 a_21241_970# a_21232_4224# 0.49fF
C1964 a_988_n1093# a_1952_n3210# 0.00fF
C1965 a_14005_n1722# a_14098_n3928# 0.00fF
C1966 w_20497_1345# a_20888_770# 0.00fF
C1967 a_10899_4538# w_9721_4472# 0.03fF
C1968 a_9875_4534# w_10863_4476# 0.01fF
C1969 a_15576_n1096# a_14005_n1722# 0.01fF
C1970 a_14098_3007# a_14335_2370# 0.38fF
C1971 a_1627_4228# a_2824_1705# 0.00fF
C1972 w_17090_n4258# a_17179_n2618# 0.03fF
C1973 a_1636_974# w_819_n1712# 0.00fF
C1974 a_1627_4228# VDD 0.99fF
C1975 w_15407_2328# A[3] 0.01fF
C1976 a_1288_2378# B[0] 0.03fF
C1977 w_6576_n3276# a_7506_n4639# 0.00fF
C1978 a_15282_n1070# a_14080_n1092# 0.13fF
C1979 a_8149_971# a_9757_4534# 0.07fF
C1980 B[5] a_17193_n968# 0.09fF
C1981 a_21557_n3206# VSS 0.43fF
C1982 a_9337_1702# VSS 0.26fF
C1983 a_8910_2395# A[1] 0.11fF
C1984 a_22547_969# A[3] 0.11fF
C1985 a_1641_2578# A[0] 0.07fF
C1986 a_9875_4534# a_10021_3951# 0.13fF
C1987 a_16283_1671# B[2] 0.01fF
C1988 a_10899_4538# a_8140_4225# 0.01fF
C1989 a_14041_n3235# w_13911_n1711# 0.01fF
C1990 a_24445_969# VSS 0.70fF
C1991 B[6] a_9462_n3933# 0.56fF
C1992 w_20488_4599# a_21246_2574# 0.00fF
C1993 a_14098_3007# a_14321_4020# 0.00fF
C1994 a_15576_n1096# a_15444_2390# 0.00fF
C1995 VDD a_1274_4028# 0.02fF
C1996 a_2397_2398# A[0] 0.11fF
C1997 w_17090_n4258# a_19659_n3206# 0.00fF
C1998 a_22097_n3899# a_20593_n1089# 0.00fF
C1999 a_24346_n4830# VDD 0.01fF
C2000 w_10863_4476# VDD 0.66fF
C2001 w_13911_n1711# w_15053_n1715# 0.03fF
C2002 w_7405_1346# VDD 0.33fF
C2003 a_1641_2578# a_1636_974# 0.12fF
C2004 a_20317_n4631# a_21557_n3206# 0.01fF
C2005 a_11647_1676# a_11589_970# 0.00fF
C2006 a_15576_n1096# a_17193_n968# 0.03fF
C2007 a_8688_n1101# a_9749_1676# 0.00fF
C2008 a_15938_n4634# a_17184_n4222# 0.00fF
C2009 a_24341_n3226# a_22509_n3925# 0.00fF
C2010 a_9691_970# VSS 0.42fF
C2011 w_23598_n2651# a_22089_n1093# 0.04fF
C2012 w_17099_n1004# a_17842_n1579# 0.00fF
C2013 w_13110_n3271# a_15222_n1096# 0.00fF
C2014 a_14674_4220# a_14098_3007# 0.01fF
C2015 w_7396_4600# a_8154_2575# 0.00fF
C2016 a_22097_n3899# A[4] 0.22fF
C2017 a_4750_n1580# VDD 0.02fF
C2018 a_9042_n1101# a_10645_n2623# 0.03fF
C2019 w_20497_1345# a_22841_1675# 0.00fF
C2020 a_3508_3954# a_4295_2398# 0.00fF
C2021 a_4750_n1580# a_4087_n2619# 0.00fF
C2022 a_1636_974# a_2397_2398# 0.10fF
C2023 a_10021_3951# VDD 1.34fF
C2024 w_20497_1345# a_20651_1407# 0.12fF
C2025 a_7152_n3907# a_9462_n3933# 0.00fF
C2026 a_1342_n1093# carry_in 0.01fF
C2027 a_1288_2378# a_1051_3015# 0.38fF
C2028 a_14330_766# a_14080_n1092# 0.00fF
C2029 w_23603_n4255# VSS 0.21fF
C2030 w_20497_1345# a_21241_970# 0.09fF
C2031 a_15989_1697# a_17342_2390# 0.62fF
C2032 w_8519_n1720# a_7546_n1097# 0.24fF
C2033 w_1961_n1716# a_1048_n1067# 0.01fF
C2034 VSS B[2] 0.78fF
C2035 a_14098_3007# VDD 1.47fF
C2036 w_4007_n1005# a_1342_n1093# 0.00fF
C2037 w_6576_n3276# B[6] 0.40fF
C2038 w_7377_n1716# a_8688_n1101# 0.02fF
C2039 A[5] a_15147_n1726# 0.01fF
C2040 a_15702_n4634# VSS 0.68fF
C2041 a_4736_n3230# a_2484_n1097# 0.01fF
C2042 VDD a_7564_n3933# 0.78fF
C2043 w_21965_2332# a_22849_4533# 0.02fF
C2044 a_6612_n3214# a_7506_n4639# 0.00fF
C2045 a_7152_n3907# a_7270_n4639# 0.01fF
C2046 a_14688_2570# a_14093_1403# 0.01fF
C2047 w_17085_n2654# B[5] 0.29fF
C2048 a_14098_3007# a_14084_4657# 0.01fF
C2049 VSS a_7550_4662# 0.19fF
C2050 a_8510_n3214# a_9404_n4639# 0.00fF
C2051 a_17433_4533# A[3] 0.00fF
C2052 a_9050_n3907# a_9168_n4639# 0.01fF
C2053 a_9749_1676# a_11235_1702# 0.02fF
C2054 A[1] a_9757_4534# 0.01fF
C2055 a_2904_n3929# a_1952_n3210# 0.07fF
C2056 a_1627_4228# w_897_2953# 0.01fF
C2057 a_17828_n3229# B[5] 0.03fF
C2058 VDD a_15044_n3209# 0.71fF
C2059 w_9721_4472# VSS 0.15fF
C2060 a_21246_2574# a_22967_4533# 0.02fF
C2061 a_8149_971# a_7796_771# 0.00fF
C2062 a_14140_n1066# a_14080_n1092# 0.05fF
C2063 w_21965_2332# a_20893_2374# 0.00fF
C2064 w_13939_1341# a_15989_965# 0.00fF
C2065 w_21965_2332# a_21232_4224# 0.00fF
C2066 a_15282_n1070# w_13911_n1711# 0.01fF
C2067 w_3998_n4259# a_2904_n3929# 0.04fF
C2068 w_21965_2332# a_23900_2394# 0.26fF
C2069 a_15576_n1096# a_16283_1671# 0.00fF
C2070 w_6576_n3276# a_7152_n3907# 0.32fF
C2071 a_8688_n1101# a_9455_970# 0.00fF
C2072 a_22002_2394# a_22547_969# 0.02fF
C2073 a_23900_2394# a_22783_969# 0.00fF
C2074 a_24681_969# Y[3] 0.36fF
C2075 w_7377_n1716# a_7606_n1071# 0.08fF
C2076 a_9042_n1101# VSS 1.20fF
C2077 w_17085_n2654# a_15576_n1096# 0.04fF
C2078 w_897_2953# a_1274_4028# 0.00fF
C2079 a_9042_n1101# A[6] 0.14fF
C2080 w_13110_n3271# a_14041_n3235# 0.54fF
C2081 a_8140_4225# VSS 0.39fF
C2082 a_23697_n4219# a_24346_n4830# 0.38fF
C2083 w_3993_n2655# A[7] 0.07fF
C2084 a_10899_4538# a_8154_2575# 0.20fF
C2085 a_17828_n3229# a_15576_n1096# 0.01fF
C2086 a_7564_3012# VSS 0.25fF
C2087 a_4386_4541# a_1641_2578# 0.20fF
C2088 B[5] VSS 0.78fF
C2089 a_24346_n4830# A[4] 0.01fF
C2090 a_21660_n1723# w_21566_n1712# 0.21fF
C2091 a_3236_1679# Y[0] 0.01fF
C2092 a_22849_4533# VDD 0.19fF
C2093 a_22089_n1093# a_21557_n3206# 0.01fF
C2094 a_13146_n3209# A[5] 0.00fF
C2095 a_15222_n1096# a_15147_n1726# 0.14fF
C2096 a_3362_4537# VDD 1.31fF
C2097 A[2] a_14683_966# 0.17fF
C2098 a_3236_1679# a_4840_973# 0.01fF
C2099 a_9050_n3907# a_8613_n1731# 0.01fF
C2100 w_20497_1345# Y[2] 0.00fF
C2101 a_14330_766# w_13911_n1711# 0.00fF
C2102 a_14098_n3928# VSS 0.48fF
C2103 w_20488_4599# A[3] 0.06fF
C2104 VDD a_17184_n4222# 1.36fF
C2105 a_2130_n1097# a_4087_n2619# 0.01fF
C2106 a_15576_n1096# VSS 1.20fF
C2107 a_2130_n1097# VDD 0.97fF
C2108 a_4092_n4223# a_2484_n1097# 0.14fF
C2109 a_20893_2374# VDD 0.02fF
C2110 w_1961_n1716# A[7] 0.01fF
C2111 VDD a_21232_4224# 0.97fF
C2112 carry_out VDD 1.14fF
C2113 w_13939_1341# a_15444_2390# 0.04fF
C2114 a_14688_2570# B[2] 0.07fF
C2115 w_892_1349# A[0] 0.19fF
C2116 a_9462_n3933# a_9404_n4639# 0.00fF
C2117 a_23900_2394# VDD 0.77fF
C2118 a_11308_n1584# a_11294_n3234# 0.00fF
C2119 a_2130_n1097# a_2055_n1727# 0.14fF
C2120 a_6612_n3214# a_7152_n3907# 0.17fF
C2121 a_2846_n4635# a_2484_n1097# 0.01fF
C2122 a_913_n1723# a_2484_n1097# 0.01fF
C2123 carry_out a_2055_n1727# 0.00fF
C2124 a_11235_1702# A[2] 0.00fF
C2125 w_20497_1345# w_21965_2332# 0.00fF
C2126 a_7796_771# A[1] 0.01fF
C2127 a_19659_n3206# a_22097_n3899# 0.00fF
C2128 w_19623_n3268# a_20553_n4631# 0.00fF
C2129 a_20199_n3899# a_21557_n3206# 0.02fF
C2130 a_15702_n4634# a_15996_n3928# 0.02fF
C2131 a_22841_1675# a_24739_1675# 0.00fF
C2132 a_10808_2395# a_8910_2395# 0.00fF
C2133 w_20497_1345# a_22783_969# 0.00fF
C2134 a_9749_1676# a_9337_1702# 0.14fF
C2135 a_2846_n4635# a_1006_n3929# 0.00fF
C2136 a_2610_n4635# a_1952_n3210# 0.02fF
C2137 w_23603_n4255# a_22089_n1093# 0.08fF
C2138 a_2130_n1097# a_2492_n3903# 0.00fF
C2139 w_10556_n4263# a_11299_n4838# 0.00fF
C2140 a_11017_4538# w_10863_4476# 0.09fF
C2141 a_1006_n3929# a_913_n1723# 0.00fF
C2142 a_21735_n1093# a_22547_969# 0.00fF
C2143 a_14140_n1066# w_13911_n1711# 0.08fF
C2144 Y[4] VSS 0.22fF
C2145 w_892_1349# a_1636_974# 0.09fF
C2146 a_13804_n4634# a_14040_n4634# 0.04fF
C2147 a_21246_2574# VSS 0.87fF
C2148 Y[0] VSS 0.21fF
C2149 a_14080_n1092# VDD 1.33fF
C2150 a_7900_n1097# a_10645_n2623# 0.12fF
C2151 a_1037_4665# VSS 0.18fF
C2152 w_3998_n4259# a_2610_n4635# 0.00fF
C2153 Y[2] a_18123_965# 0.36fF
C2154 w_4350_4479# a_3508_3954# 0.29fF
C2155 A[5] a_14434_n1092# 0.07fF
C2156 w_6576_n3276# a_9404_n4639# 0.00fF
C2157 a_4840_973# VSS 0.69fF
C2158 a_4101_n969# a_2484_n1097# 0.03fF
C2159 a_22509_n3925# VSS 0.49fF
C2160 a_9749_1676# a_9691_970# 0.00fF
C2161 a_11017_4538# a_10021_3951# 0.06fF
C2162 a_988_n1093# VSS 0.42fF
C2163 a_8149_971# w_10863_4476# 0.00fF
C2164 a_20317_n4631# Y[4] 0.44fF
C2165 w_20488_4599# a_20642_4661# 0.13fF
C2166 w_23955_4475# a_21246_2574# 0.12fF
C2167 w_22813_4471# a_22849_4533# 0.20fF
C2168 w_883_4603# carry_in 0.00fF
C2169 a_8154_2575# VSS 0.87fF
C2170 a_3236_1679# A[0] 0.81fF
C2171 w_7405_1346# a_8149_971# 0.09fF
C2172 VDD B[1] 0.92fF
C2173 w_20488_4599# a_20879_4024# 0.00fF
C2174 B[6] a_11294_n3234# 0.03fF
C2175 a_14093_1403# A[2] 0.22fF
C2176 a_15996_n3928# B[5] 0.56fF
C2177 a_7606_n1071# a_8688_n1101# 0.01fF
C2178 a_21735_n1093# a_23692_n2615# 0.01fF
C2179 a_7471_n1727# a_7546_n1097# 0.14fF
C2180 w_15053_n1715# a_15147_n1726# 0.21fF
C2181 B[6] a_9168_n4639# 0.09fF
C2182 a_8149_971# a_10021_3951# 0.03fF
C2183 w_20497_1345# VDD 0.33fF
C2184 VDD a_11589_970# 0.00fF
C2185 a_24445_969# a_22547_1701# 0.09fF
C2186 a_21735_n1093# a_24355_n1576# 0.00fF
C2187 w_10556_n4263# Y[5] 0.00fF
C2188 w_13939_1341# a_16283_1671# 0.00fF
C2189 w_22813_4471# a_21232_4224# 0.21fF
C2190 a_9337_1702# a_9455_970# 0.01fF
C2191 a_1636_974# a_3236_1679# 0.01fF
C2192 w_17397_4471# a_16409_4529# 0.01fF
C2193 a_5134_1679# carry_in 0.96fF
C2194 a_4736_n3230# VDD 0.03fF
C2195 a_15996_n3928# a_14098_n3928# 0.00fF
C2196 a_4736_n3230# a_4087_n2619# 0.38fF
C2197 a_15989_965# a_15222_n1096# 0.00fF
C2198 a_7900_n1097# A[6] 0.07fF
C2199 a_1288_2378# a_1283_774# 0.00fF
C2200 w_9721_4472# a_9749_1676# 0.00fF
C2201 a_7900_n1097# VSS 0.87fF
C2202 a_15576_n1096# a_15996_n3928# 0.10fF
C2203 a_1288_2378# VDD 0.02fF
C2204 w_2360_2336# a_5134_1679# 0.20fF
C2205 w_3993_n2655# a_4750_n1580# 0.00fF
C2206 A[5] a_17193_n968# 0.14fF
C2207 a_1641_2578# B[0] 0.07fF
C2208 VDD a_9050_n3907# 2.56fF
C2209 a_13804_n4634# a_13686_n3902# 0.01fF
C2210 w_20424_n1708# a_21660_n1723# 0.01fF
C2211 w_10556_n4263# w_10551_n2659# 0.02fF
C2212 a_15222_n1096# a_14434_n1092# 0.04fF
C2213 a_21660_n1723# a_21735_n1093# 0.14fF
C2214 w_13110_n3271# a_15938_n4634# 0.00fF
C2215 a_13146_n3209# a_14041_n3235# 0.01fF
C2216 a_9455_970# a_9691_970# 0.04fF
C2217 w_8873_2333# a_7559_1408# 0.00fF
C2218 a_9042_n1101# a_9749_1676# 0.00fF
C2219 a_2610_n4635# Y[7] 0.00fF
C2220 a_2397_2398# B[0] 0.60fF
C2221 w_10551_n2659# a_8688_n1101# 0.01fF
C2222 a_3244_4537# w_4350_4479# 0.01fF
C2223 A[0] VSS 1.71fF
C2224 VDD w_13911_n1711# 0.67fF
C2225 a_20642_4661# a_22967_4533# 0.00fF
C2226 a_22849_4533# a_23991_4537# 0.01fF
C2227 a_21246_2574# a_24109_4537# 0.04fF
C2228 VDD a_18123_965# 0.00fF
C2229 a_14005_n1722# a_15222_n1096# 0.01fF
C2230 a_7546_n1097# a_7796_771# 0.00fF
C2231 a_15282_n1070# a_15147_n1726# 1.19fF
C2232 a_8748_n1075# a_8613_n1731# 1.19fF
C2233 w_7405_1346# A[1] 0.19fF
C2234 w_13939_1341# VSS 0.20fF
C2235 w_819_n1712# a_2484_n1097# 0.00fF
C2236 a_11353_970# VSS 0.69fF
C2237 w_3998_n4259# a_6612_n3214# 0.00fF
C2238 w_17099_n1004# B[5] 0.13fF
C2239 a_11353_970# A[6] 0.00fF
C2240 w_7405_1346# w_7410_2950# 0.02fF
C2241 w_21965_2332# a_24739_1675# 0.20fF
C2242 a_22841_1675# a_22547_969# 0.02fF
C2243 w_4350_4479# a_4504_4541# 0.09fF
C2244 w_7377_n1716# a_9042_n1101# 0.00fF
C2245 w_8519_n1720# a_7471_n1727# 0.03fF
C2246 a_20651_1407# a_22547_969# 0.00fF
C2247 a_14093_1403# a_14683_966# 0.14fF
C2248 a_21241_970# a_22547_969# 0.02fF
C2249 B[7] A[7] 1.71fF
C2250 a_22215_n4631# a_22451_n4631# 0.04fF
C2251 a_2904_n3929# VSS 0.49fF
C2252 a_10021_3951# A[1] 0.00fF
C2253 a_1636_974# VSS 1.12fF
C2254 a_20656_3011# a_21246_2574# 0.11fF
C2255 a_22967_4533# a_23113_3950# 0.13fF
C2256 a_23991_4537# a_21232_4224# 0.01fF
C2257 a_10659_n973# a_8613_n1731# 0.01fF
C2258 a_23900_2394# Y[3] 0.10fF
C2259 a_1641_2578# a_1051_3015# 0.11fF
C2260 a_23900_2394# a_23991_4537# 0.00fF
C2261 a_15222_n1096# a_15444_2390# 0.00fF
C2262 A[2] B[2] 2.23fF
C2263 a_21246_2574# B[3] 0.07fF
C2264 VSS A[3] 1.99fF
C2265 w_17099_n1004# a_15576_n1096# 0.02fF
C2266 a_20553_n4631# VDD 0.00fF
C2267 a_8510_n3214# VSS 0.43fF
C2268 a_8510_n3214# A[6] 0.80fF
C2269 a_22089_n1093# a_22509_n3925# 0.10fF
C2270 w_4007_n1005# carry_in 0.05fF
C2271 w_2360_2336# carry_in 0.39fF
C2272 a_1342_n1093# a_988_n1093# 0.49fF
C2273 a_2397_2398# a_1051_3015# 0.00fF
C2274 a_3178_973# carry_in 0.00fF
C2275 a_15222_n1096# a_17193_n968# 0.12fF
C2276 a_15989_1697# a_18181_1671# 0.01fF
C2277 w_17085_n2654# A[5] 0.07fF
C2278 a_712_n4635# a_948_n4635# 0.04fF
C2279 a_4092_n4223# VDD 1.36fF
C2280 a_1627_4228# w_4350_4479# 0.02fF
C2281 a_9462_n3933# a_10645_n2623# 0.00fF
C2282 a_4092_n4223# a_4087_n2619# 0.01fF
C2283 a_9042_n1101# a_9455_970# 0.00fF
C2284 a_14041_n3235# a_14434_n1092# 0.00fF
C2285 w_897_2953# a_1288_2378# 0.00fF
C2286 a_17828_n3229# A[5] 0.01fF
C2287 a_17184_n4222# a_17179_n2618# 0.01fF
C2288 w_21566_n1712# VSS 0.23fF
C2289 a_2397_2398# a_2484_n1097# 0.00fF
C2290 w_2360_2336# a_3178_973# 0.00fF
C2291 VDD a_913_n1723# 0.27fF
C2292 a_17828_n3229# a_17833_n4833# 0.00fF
C2293 a_11308_n1584# VDD 0.02fF
C2294 a_20199_n3899# Y[4] 2.32fF
C2295 a_2846_n4635# VDD 0.00fF
C2296 VDD a_7506_n4639# 0.00fF
C2297 a_8688_n1101# a_9691_970# 0.00fF
C2298 a_24739_1675# VDD 0.69fF
C2299 a_7787_4025# VDD 0.02fF
C2300 a_14005_n1722# a_14041_n3235# 0.01fF
C2301 a_2484_n1097# a_2190_n1071# 0.05fF
C2302 w_15053_n1715# a_14434_n1092# 0.10fF
C2303 a_913_n1723# a_2055_n1727# 0.01fF
C2304 a_22451_n4631# B[4] 0.00fF
C2305 w_18_n3272# a_988_n1093# 0.01fF
C2306 w_3993_n2655# a_2130_n1097# 0.01fF
C2307 w_3208_4475# a_1641_2578# 0.08fF
C2308 a_20199_n3899# a_22509_n3925# 0.00fF
C2309 a_20611_n3925# a_22097_n3899# 0.02fF
C2310 a_9168_n4639# a_9404_n4639# 0.04fF
C2311 a_1006_n3929# a_948_n4635# 0.00fF
C2312 a_1952_n3210# a_712_n4635# 0.01fF
C2313 a_23692_n2615# B[4] 0.18fF
C2314 w_19623_n3268# a_22451_n4631# 0.00fF
C2315 a_11235_1702# a_9337_1702# 0.02fF
C2316 w_19623_n3268# a_23692_n2615# 0.02fF
C2317 a_17887_965# A[5] 0.00fF
C2318 A[5] VSS 1.74fF
C2319 a_14140_n1066# a_15147_n1726# 0.00fF
C2320 a_16409_4529# a_17433_4533# 0.02fF
C2321 a_16291_4529# a_16409_4529# 1.20fF
C2322 a_24355_n1576# B[4] 0.02fF
C2323 a_2846_n4635# a_2492_n3903# 0.00fF
C2324 a_14005_n1722# w_15053_n1715# 0.03fF
C2325 a_1952_n3210# a_2484_n1097# 0.01fF
C2326 a_17833_n4833# VSS 0.38fF
C2327 w_6576_n3276# a_10645_n2623# 0.02fF
C2328 a_9749_1676# a_8154_2575# 0.02fF
C2329 w_13110_n3271# VDD 1.02fF
C2330 a_7564_3012# a_7801_2375# 0.38fF
C2331 a_20642_4661# VSS 0.20fF
C2332 w_15407_2328# Y[2] 0.15fF
C2333 w_13939_1341# a_14688_2570# 0.01fF
C2334 w_20502_2949# a_21246_2574# 0.05fF
C2335 a_20879_4024# VSS 0.37fF
C2336 a_4101_n969# VDD 1.42fF
C2337 a_4386_4541# VSS 0.62fF
C2338 a_4101_n969# a_4087_n2619# 0.01fF
C2339 w_3998_n4259# a_2484_n1097# 0.08fF
C2340 a_15222_n1096# a_16283_1671# 0.00fF
C2341 a_1006_n3929# a_1952_n3210# 0.23fF
C2342 B[2] a_14683_966# 0.13fF
C2343 a_9462_n3933# A[6] 0.07fF
C2344 a_3236_1679# a_5076_973# 0.00fF
C2345 w_15407_2328# a_14335_2370# 0.00fF
C2346 a_9462_n3933# VSS 0.49fF
C2347 a_4101_n969# a_2055_n1727# 0.01fF
C2348 a_2130_n1097# a_2942_973# 0.00fF
C2349 a_8149_971# B[1] 0.13fF
C2350 w_1961_n1716# a_2130_n1097# 0.21fF
C2351 a_20317_n4631# A[5] 0.00fF
C2352 a_2610_n4635# VSS 0.68fF
C2353 a_15576_n1096# A[2] 0.00fF
C2354 w_17085_n2654# a_15222_n1096# 0.01fF
C2355 a_14674_4220# w_17397_4471# 0.02fF
C2356 w_1961_n1716# carry_out 0.01fF
C2357 a_7270_n4639# VSS 0.69fF
C2358 a_7270_n4639# A[6] 0.00fF
C2359 a_21795_n1067# a_21660_n1723# 1.19fF
C2360 a_22002_2394# VSS 0.48fF
C2361 B[6] VDD 0.91fF
C2362 a_23113_3950# VSS 0.37fF
C2363 a_21246_2574# a_22547_1701# 0.01fF
C2364 w_892_1349# B[0] 0.17fF
C2365 VDD a_8748_n1075# 1.32fF
C2366 w_19623_n3268# a_21660_n1723# 0.02fF
C2367 w_21965_2332# a_22547_969# 0.02fF
C2368 w_10556_n4263# a_9042_n1101# 0.08fF
C2369 a_20553_n4631# A[4] 0.00fF
C2370 a_15282_n1070# a_14434_n1092# 0.02fF
C2371 w_23603_n4255# w_23598_n2651# 0.02fF
C2372 w_15053_n1715# a_17193_n968# 0.00fF
C2373 a_22547_969# a_22783_969# 0.04fF
C2374 a_9042_n1101# a_11299_n4838# 0.00fF
C2375 w_17397_4471# VDD 0.66fF
C2376 a_9042_n1101# a_8688_n1101# 0.48fF
C2377 a_8910_2395# a_7796_771# 0.00fF
C2378 a_1636_974# a_1342_n1093# 0.00fF
C2379 a_1342_n1093# a_2904_n3929# 0.03fF
C2380 w_8873_2333# a_10899_4538# 0.04fF
C2381 a_10659_n973# VDD 1.42fF
C2382 a_20656_3011# A[3] 0.06fF
C2383 a_22089_n1093# A[3] 0.00fF
C2384 w_23955_4475# a_23113_3950# 0.29fF
C2385 a_17842_n1579# B[5] 0.02fF
C2386 w_6576_n3276# VSS 0.34fF
C2387 w_6576_n3276# A[6] 0.59fF
C2388 a_15282_n1070# a_14005_n1722# 0.02fF
C2389 w_13930_4595# a_16291_4529# 0.01fF
C2390 w_20488_4599# a_21241_970# 0.02fF
C2391 w_17397_4471# a_17551_4533# 0.09fF
C2392 B[3] A[3] 2.23fF
C2393 Y[1] VSS 0.21fF
C2394 a_15702_n4634# Y[5] 0.00fF
C2395 a_7546_n1097# a_7564_n3933# 0.00fF
C2396 a_7152_n3907# VDD 2.54fF
C2397 w_7377_n1716# a_7900_n1097# 0.12fF
C2398 a_15222_n1096# VSS 0.49fF
C2399 a_8510_n3214# Y[6] 0.01fF
C2400 w_15407_2328# a_14674_4220# 0.00fF
C2401 a_4750_n1580# B[7] 0.02fF
C2402 a_5076_973# VSS 0.42fF
C2403 a_17769_1697# A[3] 0.00fF
C2404 a_14040_n4634# a_13686_n3902# 0.00fF
C2405 a_24341_n3226# B[4] 0.03fF
C2406 a_9749_1676# a_11353_970# 0.01fF
C2407 w_18_n3272# a_2904_n3929# 0.25fF
C2408 a_712_n4635# Y[7] 0.44fF
C2409 a_13804_n4634# a_15044_n3209# 0.01fF
C2410 w_3993_n2655# a_4736_n3230# 0.00fF
C2411 w_892_1349# a_1051_3015# 0.03fF
C2412 a_22089_n1093# w_21566_n1712# 0.12fF
C2413 w_19623_n3268# a_24341_n3226# 0.00fF
C2414 a_15576_n1096# a_17842_n1579# 0.01fF
C2415 a_7606_n1071# a_9042_n1101# 0.00fF
C2416 w_15407_2328# VDD 0.92fF
C2417 a_23692_n2615# a_20947_n1089# 0.12fF
C2418 a_10021_3951# a_10808_2395# 0.00fF
C2419 A[1] B[1] 2.23fF
C2420 a_3362_4537# w_4350_4479# 0.01fF
C2421 a_3236_1679# B[0] 0.01fF
C2422 a_1037_4665# w_883_4603# 0.12fF
C2423 a_7801_2375# a_8154_2575# 0.00fF
C2424 w_7410_2950# B[1] 0.29fF
C2425 a_1283_774# w_819_n1712# 0.00fF
C2426 VDD a_22547_969# 0.01fF
C2427 VDD w_819_n1712# 0.68fF
C2428 VDD a_15147_n1726# 0.19fF
C2429 a_15996_n3928# A[5] 0.07fF
C2430 a_14093_1403# B[2] 0.03fF
C2431 a_17342_2390# a_18123_965# 0.00fF
C2432 a_15282_n1070# a_17193_n968# 0.00fF
C2433 w_20424_n1708# VSS 0.22fF
C2434 a_17833_n4833# a_15996_n3928# 0.00fF
C2435 a_1006_n3929# Y[7] 0.10fF
C2436 A[1] a_11589_970# 0.00fF
C2437 w_819_n1712# a_2055_n1727# 0.01fF
C2438 a_21735_n1093# VSS 0.49fF
C2439 a_9337_1702# a_9691_970# 0.00fF
C2440 a_2904_n3929# a_594_n3903# 0.00fF
C2441 a_15989_965# Y[2] 0.00fF
C2442 a_5134_1679# Y[0] 0.15fF
C2443 a_6612_n3214# VSS 0.36fF
C2444 a_20656_3011# a_20642_4661# 0.01fF
C2445 a_14140_n1066# a_14434_n1092# 0.04fF
C2446 a_24109_4537# a_23113_3950# 0.06fF
C2447 a_6612_n3214# A[6] 0.00fF
C2448 a_20656_3011# a_20879_4024# 0.00fF
C2449 a_24739_1675# Y[3] 0.15fF
C2450 a_20642_4661# B[3] 0.10fF
C2451 a_21241_970# a_22967_4533# 0.05fF
C2452 w_13944_2945# a_14098_3007# 0.13fF
C2453 a_21660_n1723# a_20947_n1089# 0.04fF
C2454 w_23603_n4255# a_21557_n3206# 0.00fF
C2455 a_7471_n1727# A[7] 0.00fF
C2456 w_20502_2949# A[3] 0.07fF
C2457 a_14041_n3235# VSS 0.55fF
C2458 a_14330_766# a_15444_2390# 0.00fF
C2459 a_1641_2578# a_2824_1705# 0.03fF
C2460 w_10551_n2659# a_9042_n1101# 0.04fF
C2461 B[3] a_20879_4024# 0.02fF
C2462 a_22451_n4631# VDD 0.00fF
C2463 a_1641_2578# VDD 1.65fF
C2464 a_5134_1679# a_4840_973# 0.02fF
C2465 Y[5] a_14098_n3928# 0.10fF
C2466 a_712_n4635# a_54_n3210# 0.02fF
C2467 a_14140_n1066# a_14005_n1722# 1.19fF
C2468 a_23692_n2615# VDD 1.48fF
C2469 a_9455_970# a_11353_970# 0.01fF
C2470 a_2397_2398# a_1283_774# 0.00fF
C2471 a_2397_2398# a_2824_1705# 0.19fF
C2472 w_15407_2328# a_16225_965# 0.00fF
C2473 a_2397_2398# VDD 0.82fF
C2474 a_7559_1408# VDD 1.38fF
C2475 a_22002_2394# a_20656_3011# 0.00fF
C2476 w_8873_2333# VSS 0.34fF
C2477 a_22002_2394# a_22089_n1093# 0.00fF
C2478 B[0] VSS 0.62fF
C2479 a_948_n4635# VDD 0.00fF
C2480 a_8149_971# a_7787_4025# 0.01fF
C2481 a_16555_3946# a_16409_4529# 0.13fF
C2482 VDD a_24355_n1576# 0.02fF
C2483 a_7270_n4639# Y[6] 0.44fF
C2484 a_14674_4220# a_17433_4533# 0.01fF
C2485 w_15053_n1715# VSS 0.23fF
C2486 a_22002_2394# B[3] 0.60fF
C2487 a_20199_n3899# A[5] 0.00fF
C2488 a_20888_770# VSS 0.38fF
C2489 a_14674_4220# a_16291_4529# 0.16fF
C2490 a_3236_1679# a_2484_n1097# 0.00fF
C2491 a_22547_1701# A[3] 0.20fF
C2492 a_13146_n3209# VDD 0.69fF
C2493 a_11294_n3234# a_10645_n2623# 0.38fF
C2494 a_19659_n3206# a_20553_n4631# 0.00fF
C2495 VDD a_2190_n1071# 1.32fF
C2496 w_17099_n1004# A[5] 0.07fF
C2497 w_13939_1341# A[2] 0.19fF
C2498 a_11353_970# A[2] 0.00fF
C2499 VDD a_9404_n4639# 0.00fF
C2500 w_7405_1346# a_8910_2395# 0.04fF
C2501 w_3993_n2655# a_4092_n4223# 0.00fF
C2502 a_17433_4533# VDD 0.28fF
C2503 a_1006_n3929# a_54_n3210# 0.07fF
C2504 a_2190_n1071# a_2055_n1727# 1.19fF
C2505 a_16291_4529# VDD 0.19fF
C2506 a_3244_4537# a_3508_3954# 0.08fF
C2507 a_2130_n1097# B[7] 0.01fF
C2508 w_18_n3272# a_2610_n4635# 0.02fF
C2509 w_10556_n4263# a_7900_n1097# 0.01fF
C2510 w_883_4603# A[0] 0.06fF
C2511 a_23706_n965# a_23692_n2615# 0.01fF
C2512 a_1952_n3210# VDD 0.71fF
C2513 a_24341_n3226# a_20947_n1089# 0.00fF
C2514 w_6576_n3276# Y[6] 0.15fF
C2515 a_8140_4225# a_9337_1702# 0.00fF
C2516 a_8688_n1101# a_7900_n1097# 0.04fF
C2517 a_23706_n965# a_24355_n1576# 0.38fF
C2518 a_17433_4533# a_17551_4533# 1.20fF
C2519 a_16291_4529# a_17551_4533# 0.00fF
C2520 carry_in Y[0] 0.23fF
C2521 a_21660_n1723# VDD 0.19fF
C2522 w_3208_4475# a_3236_1679# 0.00fF
C2523 a_1952_n3210# a_2055_n1727# 0.00fF
C2524 a_16291_4529# a_14084_4657# 0.01fF
C2525 w_3998_n4259# VDD 0.33fF
C2526 a_3508_3954# a_4504_4541# 0.06fF
C2527 a_1288_2378# a_1046_1411# 0.01fF
C2528 w_3998_n4259# a_4087_n2619# 0.03fF
C2529 w_10565_n1009# a_11308_n1584# 0.00fF
C2530 w_13110_n3271# a_17179_n2618# 0.02fF
C2531 a_22215_n4631# VSS 0.68fF
C2532 a_7564_3012# a_9337_1702# 0.00fF
C2533 a_1037_4665# carry_in 0.00fF
C2534 a_9875_4534# w_7396_4600# 0.00fF
C2535 a_14335_2370# a_15444_2390# 0.00fF
C2536 w_20502_2949# a_20642_4661# 0.02fF
C2537 w_2360_2336# Y[0] 0.15fF
C2538 a_1051_3015# VSS 0.24fF
C2539 w_20502_2949# a_20879_4024# 0.00fF
C2540 a_4840_973# carry_in 0.12fF
C2541 a_11647_1676# VSS 0.36fF
C2542 w_883_4603# a_1636_974# 0.02fF
C2543 a_988_n1093# carry_in 0.02fF
C2544 a_1952_n3210# a_2492_n3903# 0.16fF
C2545 a_15989_965# VDD 0.01fF
C2546 a_5134_1679# A[0] 0.00fF
C2547 a_712_n4635# VSS 0.69fF
C2548 w_4007_n1005# a_4840_973# 0.00fF
C2549 a_9042_n1101# a_9691_970# 0.00fF
C2550 w_2360_2336# a_4840_973# 0.02fF
C2551 a_11294_n3234# VSS 0.37fF
C2552 a_11294_n3234# A[6] 0.01fF
C2553 w_1961_n1716# a_913_n1723# 0.03fF
C2554 w_3993_n2655# a_4101_n969# 0.03fF
C2555 a_15282_n1070# VSS 0.08fF
C2556 a_22451_n4631# a_23697_n4219# 0.00fF
C2557 a_22215_n4631# a_20317_n4631# 0.01fF
C2558 a_1641_2578# w_897_2953# 0.05fF
C2559 a_2484_n1097# VSS 1.21fF
C2560 w_3998_n4259# a_2492_n3903# 0.02fF
C2561 a_22841_1675# VSS 0.46fF
C2562 a_21660_n1723# a_23706_n965# 0.01fF
C2563 a_9168_n4639# VSS 0.68fF
C2564 a_9168_n4639# A[6] 0.10fF
C2565 w_20424_n1708# a_22089_n1093# 0.00fF
C2566 a_2904_n3929# a_4741_n4834# 0.00fF
C2567 VDD a_14434_n1092# 1.77fF
C2568 a_16409_4529# VSS 0.05fF
C2569 a_23697_n4219# a_23692_n2615# 0.01fF
C2570 a_7787_4025# A[1] 0.00fF
C2571 a_7606_n1071# a_7900_n1097# 0.04fF
C2572 a_20651_1407# VSS 0.30fF
C2573 a_9749_1676# Y[1] 0.01fF
C2574 a_21241_970# VSS 1.12fF
C2575 a_22089_n1093# a_21735_n1093# 0.48fF
C2576 w_9721_4472# a_7550_4662# 0.00fF
C2577 w_10863_4476# a_9757_4534# 0.01fF
C2578 w_7410_2950# a_7787_4025# 0.00fF
C2579 a_1627_4228# a_3508_3954# 0.08fF
C2580 a_22451_n4631# A[4] 0.00fF
C2581 w_7396_4600# VDD 0.39fF
C2582 a_21735_n1093# B[3] 0.00fF
C2583 a_24341_n3226# VDD 0.03fF
C2584 w_17099_n1004# a_15222_n1096# 0.06fF
C2585 a_1006_n3929# VSS 0.48fF
C2586 w_20488_4599# VDD 0.39fF
C2587 a_23692_n2615# A[4] 0.06fF
C2588 w_13939_1341# a_14683_966# 0.09fF
C2589 a_14041_n3235# a_15996_n3928# 0.10fF
C2590 a_6612_n3214# Y[6] 0.16fF
C2591 a_14005_n1722# VDD 0.27fF
C2592 a_21795_n1067# VSS 0.08fF
C2593 B[4] VSS 0.83fF
C2594 w_10556_n4263# a_8510_n3214# 0.00fF
C2595 Y[3] a_22547_969# 0.00fF
C2596 a_24355_n1576# A[4] 0.00fF
C2597 w_3208_4475# VSS 0.15fF
C2598 w_6576_n3276# w_7377_n1716# 0.01fF
C2599 a_22002_2394# a_22547_1701# 0.09fF
C2600 a_22547_1701# a_23113_3950# 0.00fF
C2601 a_15702_n4634# B[5] 0.09fF
C2602 w_19623_n3268# VSS 0.34fF
C2603 a_8140_4225# a_7550_4662# 0.10fF
C2604 a_10021_3951# a_9757_4534# 0.08fF
C2605 w_23955_4475# a_21241_970# 0.00fF
C2606 a_7546_n1097# a_9050_n3907# 0.00fF
C2607 w_10565_n1009# B[6] 0.14fF
C2608 w_10565_n1009# a_8748_n1075# 0.00fF
C2609 w_1961_n1716# a_4101_n969# 0.00fF
C2610 a_10808_2395# B[1] 0.00fF
C2611 a_21557_n3206# Y[4] 0.01fF
C2612 w_9721_4472# a_8140_4225# 0.21fF
C2613 a_21660_n1723# a_20593_n1089# 0.09fF
C2614 a_16283_1671# Y[2] 0.01fF
C2615 a_9875_4534# a_10899_4538# 0.02fF
C2616 a_15989_965# a_16225_965# 0.04fF
C2617 w_17090_n4258# a_15044_n3209# 0.00fF
C2618 w_20424_n1708# a_20199_n3899# 0.00fF
C2619 a_7564_3012# a_7550_4662# 0.01fF
C2620 a_14330_766# VSS 0.38fF
C2621 a_11235_1702# a_11353_970# 0.01fF
C2622 a_15444_2390# VDD 0.81fF
C2623 a_10808_2395# a_11589_970# 0.00fF
C2624 VDD Y[7] 0.07fF
C2625 B[7] a_4736_n3230# 0.03fF
C2626 a_14040_n4634# a_15044_n3209# 0.00fF
C2627 a_15702_n4634# a_14098_n3928# 0.01fF
C2628 a_3244_4537# a_4504_4541# 0.00fF
C2629 a_21557_n3206# a_22509_n3925# 0.07fF
C2630 A[0] carry_in 0.88fF
C2631 a_15576_n1096# B[2] 0.00fF
C2632 w_19623_n3268# a_20317_n4631# 0.02fF
C2633 w_10551_n2659# a_7900_n1097# 0.05fF
C2634 w_10565_n1009# a_10659_n973# 0.13fF
C2635 w_892_1349# a_1283_774# 0.00fF
C2636 w_892_1349# a_2824_1705# 0.01fF
C2637 a_15576_n1096# a_15702_n4634# 0.02fF
C2638 a_8613_n1731# VSS 0.66fF
C2639 B[3] a_20888_770# 0.00fF
C2640 w_892_1349# VDD 0.34fF
C2641 A[6] a_8613_n1731# 0.01fF
C2642 a_21660_n1723# A[4] 0.01fF
C2643 a_9337_1702# a_8154_2575# 0.03fF
C2644 w_2360_2336# A[0] 0.60fF
C2645 w_15407_2328# a_17342_2390# 0.26fF
C2646 VDD a_17193_n968# 1.42fF
C2647 a_15938_n4634# VSS 0.42fF
C2648 a_3178_973# A[0] 0.01fF
C2649 Y[1] a_9455_970# 0.00fF
C2650 w_13930_4595# VSS 0.10fF
C2651 a_8140_4225# a_7564_3012# 0.01fF
C2652 a_7471_n1727# a_7564_n3933# 0.00fF
C2653 a_14140_n1066# VSS 0.07fF
C2654 a_2492_n3903# Y[7] 0.00fF
C2655 a_10899_4538# VDD 0.28fF
C2656 a_1636_974# carry_in 0.11fF
C2657 a_22967_4533# VDD 1.31fF
C2658 a_17842_n1579# A[5] 0.00fF
C2659 w_8873_2333# a_9749_1676# 0.19fF
C2660 a_17887_965# Y[2] 0.43fF
C2661 a_3244_4537# a_1627_4228# 0.16fF
C2662 Y[2] VSS 0.21fF
C2663 Y[1] A[2] 0.01fF
C2664 a_22089_n1093# a_22215_n4631# 0.02fF
C2665 a_14674_4220# a_16555_3946# 0.08fF
C2666 Y[4] a_1596_n2079# 0.51fF
C2667 Y[5] a_1596_n2079# 0.51fF
C2668 Y[6] a_1596_n2079# 0.51fF
C2669 Y[7] a_1596_n2079# 0.53fF
C2670 A[4] a_1596_n2079# 3.91fF
C2671 B[4] a_1596_n2079# 3.24fF
C2672 A[5] a_1596_n2079# 3.80fF
C2673 B[5] a_1596_n2079# 3.24fF
C2674 A[6] a_1596_n2079# 3.81fF
C2675 B[6] a_1596_n2079# 3.24fF
C2676 carry_out a_1596_n2079# 0.44fF
C2677 A[7] a_1596_n2079# 3.82fF
C2678 B[7] a_1596_n2079# 3.24fF
C2679 Y[3] a_1596_n2079# 0.44fF
C2680 Y[2] a_1596_n2079# 0.44fF
C2681 Y[1] a_1596_n2079# 0.44fF
C2682 Y[0] a_1596_n2079# 0.44fF
C2683 carry_in a_1596_n2079# 5.32fF
C2684 B[3] a_1596_n2079# 3.75fF
C2685 A[3] a_1596_n2079# 4.11fF
C2686 B[2] a_1596_n2079# 3.75fF
C2687 A[2] a_1596_n2079# 4.10fF
C2688 VSS a_1596_n2079# 57.30fF
C2689 B[1] a_1596_n2079# 3.75fF
C2690 A[1] a_1596_n2079# 4.09fF
C2691 VDD a_1596_n2079# 52.01fF
C2692 B[0] a_1596_n2079# 3.79fF
C2693 A[0] a_1596_n2079# 4.40fF
C2694 a_24346_n4830# a_1596_n2079# 0.03fF
C2695 a_22451_n4631# a_1596_n2079# 0.02fF
C2696 a_22215_n4631# a_1596_n2079# 0.27fF
C2697 a_20553_n4631# a_1596_n2079# 0.02fF
C2698 a_17833_n4833# a_1596_n2079# 0.03fF
C2699 a_20317_n4631# a_1596_n2079# 0.32fF
C2700 a_23697_n4219# a_1596_n2079# 0.76fF
C2701 a_24341_n3226# a_1596_n2079# 0.03fF
C2702 a_15938_n4634# a_1596_n2079# 0.02fF
C2703 a_15702_n4634# a_1596_n2079# 0.27fF
C2704 a_14040_n4634# a_1596_n2079# 0.02fF
C2705 a_11299_n4838# a_1596_n2079# 0.03fF
C2706 a_13804_n4634# a_1596_n2079# 0.32fF
C2707 a_17184_n4222# a_1596_n2079# 0.76fF
C2708 a_22509_n3925# a_1596_n2079# 0.73fF
C2709 a_22097_n3899# a_1596_n2079# 0.24fF
C2710 a_21557_n3206# a_1596_n2079# 0.54fF
C2711 a_20611_n3925# a_1596_n2079# 0.63fF
C2712 a_20199_n3899# a_1596_n2079# 0.19fF
C2713 a_19659_n3206# a_1596_n2079# 0.64fF
C2714 a_17828_n3229# a_1596_n2079# 0.03fF
C2715 a_9404_n4639# a_1596_n2079# 0.02fF
C2716 a_9168_n4639# a_1596_n2079# 0.27fF
C2717 a_7506_n4639# a_1596_n2079# 0.02fF
C2718 a_7270_n4639# a_1596_n2079# 0.32fF
C2719 a_4741_n4834# a_1596_n2079# 0.03fF
C2720 a_10650_n4227# a_1596_n2079# 0.76fF
C2721 a_15996_n3928# a_1596_n2079# 0.73fF
C2722 a_15044_n3209# a_1596_n2079# 0.54fF
C2723 a_14098_n3928# a_1596_n2079# 0.63fF
C2724 a_13686_n3902# a_1596_n2079# 0.19fF
C2725 a_13146_n3209# a_1596_n2079# 0.64fF
C2726 a_11294_n3234# a_1596_n2079# 0.03fF
C2727 a_2846_n4635# a_1596_n2079# 0.02fF
C2728 a_2610_n4635# a_1596_n2079# 0.27fF
C2729 a_948_n4635# a_1596_n2079# 0.02fF
C2730 a_712_n4635# a_1596_n2079# 0.32fF
C2731 a_4092_n4223# a_1596_n2079# 0.76fF
C2732 a_9462_n3933# a_1596_n2079# 0.73fF
C2733 a_14041_n3235# a_1596_n2079# 1.31fF
C2734 a_9050_n3907# a_1596_n2079# 0.24fF
C2735 a_8510_n3214# a_1596_n2079# 0.54fF
C2736 a_7564_n3933# a_1596_n2079# 0.63fF
C2737 a_7152_n3907# a_1596_n2079# 0.19fF
C2738 a_6612_n3214# a_1596_n2079# 0.64fF
C2739 a_4736_n3230# a_1596_n2079# 0.03fF
C2740 a_2904_n3929# a_1596_n2079# 0.73fF
C2741 a_2492_n3903# a_1596_n2079# 0.25fF
C2742 a_1952_n3210# a_1596_n2079# 0.54fF
C2743 a_1006_n3929# a_1596_n2079# 0.63fF
C2744 a_594_n3903# a_1596_n2079# 0.22fF
C2745 a_54_n3210# a_1596_n2079# 0.69fF
C2746 a_23692_n2615# a_1596_n2079# 0.69fF
C2747 a_17179_n2618# a_1596_n2079# 0.69fF
C2748 a_10645_n2623# a_1596_n2079# 0.69fF
C2749 a_4087_n2619# a_1596_n2079# 0.69fF
C2750 a_24355_n1576# a_1596_n2079# 0.03fF
C2751 a_23706_n965# a_1596_n2079# 0.77fF
C2752 a_21660_n1723# a_1596_n2079# 0.62fF
C2753 a_21795_n1067# a_1596_n2079# 0.09fF
C2754 a_17842_n1579# a_1596_n2079# 0.03fF
C2755 a_22089_n1093# a_1596_n2079# 1.70fF
C2756 a_20518_n1719# a_1596_n2079# 0.45fF
C2757 a_20653_n1063# a_1596_n2079# 0.08fF
C2758 a_17193_n968# a_1596_n2079# 0.78fF
C2759 a_20947_n1089# a_1596_n2079# 1.57fF
C2760 a_15147_n1726# a_1596_n2079# 0.62fF
C2761 a_15282_n1070# a_1596_n2079# 0.09fF
C2762 a_11308_n1584# a_1596_n2079# 0.03fF
C2763 a_15576_n1096# a_1596_n2079# 1.70fF
C2764 a_14005_n1722# a_1596_n2079# 0.45fF
C2765 a_14140_n1066# a_1596_n2079# 0.08fF
C2766 a_10659_n973# a_1596_n2079# 0.78fF
C2767 a_21735_n1093# a_1596_n2079# 1.31fF
C2768 a_20593_n1089# a_1596_n2079# 0.65fF
C2769 a_14434_n1092# a_1596_n2079# 1.57fF
C2770 a_8613_n1731# a_1596_n2079# 0.62fF
C2771 a_8748_n1075# a_1596_n2079# 0.09fF
C2772 a_4750_n1580# a_1596_n2079# 0.03fF
C2773 a_9042_n1101# a_1596_n2079# 1.70fF
C2774 a_7471_n1727# a_1596_n2079# 0.44fF
C2775 a_7606_n1071# a_1596_n2079# 0.08fF
C2776 a_4101_n969# a_1596_n2079# 0.78fF
C2777 a_15222_n1096# a_1596_n2079# 1.31fF
C2778 a_14080_n1092# a_1596_n2079# 0.65fF
C2779 a_7900_n1097# a_1596_n2079# 1.57fF
C2780 a_2055_n1727# a_1596_n2079# 0.62fF
C2781 a_2190_n1071# a_1596_n2079# 0.09fF
C2782 a_2484_n1097# a_1596_n2079# 1.70fF
C2783 a_913_n1723# a_1596_n2079# 0.44fF
C2784 a_1048_n1067# a_1596_n2079# 0.08fF
C2785 a_8688_n1101# a_1596_n2079# 1.31fF
C2786 a_7546_n1097# a_1596_n2079# 0.65fF
C2787 a_1342_n1093# a_1596_n2079# 1.57fF
C2788 a_2130_n1097# a_1596_n2079# 1.31fF
C2789 a_988_n1093# a_1596_n2079# 0.65fF
C2790 a_24681_969# a_1596_n2079# 0.02fF
C2791 a_24445_969# a_1596_n2079# 0.32fF
C2792 a_22783_969# a_1596_n2079# 0.02fF
C2793 a_22547_969# a_1596_n2079# 0.27fF
C2794 a_20888_770# a_1596_n2079# 0.03fF
C2795 a_18123_965# a_1596_n2079# 0.02fF
C2796 a_17887_965# a_1596_n2079# 0.32fF
C2797 a_16225_965# a_1596_n2079# 0.02fF
C2798 a_15989_965# a_1596_n2079# 0.27fF
C2799 a_14330_766# a_1596_n2079# 0.03fF
C2800 a_20651_1407# a_1596_n2079# 0.74fF
C2801 a_24739_1675# a_1596_n2079# 0.67fF
C2802 a_23900_2394# a_1596_n2079# 0.59fF
C2803 a_22841_1675# a_1596_n2079# 0.59fF
C2804 a_22002_2394# a_1596_n2079# 0.70fF
C2805 a_20893_2374# a_1596_n2079# 0.03fF
C2806 a_11589_970# a_1596_n2079# 0.02fF
C2807 a_11353_970# a_1596_n2079# 0.32fF
C2808 a_9691_970# a_1596_n2079# 0.02fF
C2809 a_9455_970# a_1596_n2079# 0.27fF
C2810 a_7796_771# a_1596_n2079# 0.03fF
C2811 a_14093_1403# a_1596_n2079# 0.74fF
C2812 a_18181_1671# a_1596_n2079# 0.68fF
C2813 a_22547_1701# a_1596_n2079# 1.23fF
C2814 a_17769_1697# a_1596_n2079# 0.19fF
C2815 a_17342_2390# a_1596_n2079# 0.59fF
C2816 a_16283_1671# a_1596_n2079# 0.59fF
C2817 a_15444_2390# a_1596_n2079# 0.70fF
C2818 a_14335_2370# a_1596_n2079# 0.03fF
C2819 a_5076_973# a_1596_n2079# 0.02fF
C2820 a_4840_973# a_1596_n2079# 0.32fF
C2821 a_3178_973# a_1596_n2079# 0.02fF
C2822 a_2942_973# a_1596_n2079# 0.27fF
C2823 a_1283_774# a_1596_n2079# 0.03fF
C2824 a_7559_1408# a_1596_n2079# 0.74fF
C2825 a_11647_1676# a_1596_n2079# 0.68fF
C2826 a_15989_1697# a_1596_n2079# 1.23fF
C2827 a_11235_1702# a_1596_n2079# 0.19fF
C2828 a_10808_2395# a_1596_n2079# 0.59fF
C2829 a_9749_1676# a_1596_n2079# 0.59fF
C2830 a_9337_1702# a_1596_n2079# 0.25fF
C2831 a_8910_2395# a_1596_n2079# 0.70fF
C2832 a_7801_2375# a_1596_n2079# 0.03fF
C2833 a_1046_1411# a_1596_n2079# 0.74fF
C2834 a_5134_1679# a_1596_n2079# 0.67fF
C2835 a_20656_3011# a_1596_n2079# 0.69fF
C2836 a_4722_1705# a_1596_n2079# 0.19fF
C2837 a_4295_2398# a_1596_n2079# 0.59fF
C2838 a_3236_1679# a_1596_n2079# 0.59fF
C2839 a_2824_1705# a_1596_n2079# 0.25fF
C2840 a_2397_2398# a_1596_n2079# 0.70fF
C2841 a_1288_2378# a_1596_n2079# 0.03fF
C2842 a_14098_3007# a_1596_n2079# 0.69fF
C2843 a_7564_3012# a_1596_n2079# 0.69fF
C2844 a_1051_3015# a_1596_n2079# 0.69fF
C2845 a_20879_4024# a_1596_n2079# 0.03fF
C2846 a_24109_4537# a_1596_n2079# 0.09fF
C2847 a_23991_4537# a_1596_n2079# 0.43fF
C2848 a_22967_4533# a_1596_n2079# 0.09fF
C2849 a_14321_4020# a_1596_n2079# 0.03fF
C2850 a_20642_4661# a_1596_n2079# 0.78fF
C2851 a_22849_4533# a_1596_n2079# 0.64fF
C2852 a_21246_2574# a_1596_n2079# 1.47fF
C2853 a_17551_4533# a_1596_n2079# 0.09fF
C2854 a_17433_4533# a_1596_n2079# 0.43fF
C2855 a_16409_4529# a_1596_n2079# 0.09fF
C2856 a_7787_4025# a_1596_n2079# 0.03fF
C2857 a_14084_4657# a_1596_n2079# 0.77fF
C2858 a_16291_4529# a_1596_n2079# 0.63fF
C2859 a_21241_970# a_1596_n2079# 1.72fF
C2860 a_14688_2570# a_1596_n2079# 1.47fF
C2861 a_11017_4538# a_1596_n2079# 0.09fF
C2862 a_10899_4538# a_1596_n2079# 0.44fF
C2863 a_9875_4534# a_1596_n2079# 0.09fF
C2864 a_1274_4028# a_1596_n2079# 0.03fF
C2865 a_7550_4662# a_1596_n2079# 0.77fF
C2866 a_9757_4534# a_1596_n2079# 0.64fF
C2867 a_14683_966# a_1596_n2079# 1.71fF
C2868 a_23113_3950# a_1596_n2079# 0.67fF
C2869 a_21232_4224# a_1596_n2079# 1.35fF
C2870 a_8154_2575# a_1596_n2079# 1.48fF
C2871 a_4504_4541# a_1596_n2079# 0.09fF
C2872 a_4386_4541# a_1596_n2079# 0.43fF
C2873 a_3362_4537# a_1596_n2079# 0.09fF
C2874 a_1037_4665# a_1596_n2079# 0.77fF
C2875 a_3244_4537# a_1596_n2079# 0.63fF
C2876 a_8149_971# a_1596_n2079# 1.72fF
C2877 a_16555_3946# a_1596_n2079# 0.67fF
C2878 a_14674_4220# a_1596_n2079# 1.35fF
C2879 a_1641_2578# a_1596_n2079# 1.47fF
C2880 a_1636_974# a_1596_n2079# 1.71fF
C2881 a_10021_3951# a_1596_n2079# 0.67fF
C2882 a_8140_4225# a_1596_n2079# 1.35fF
C2883 a_3508_3954# a_1596_n2079# 0.67fF
C2884 a_1627_4228# a_1596_n2079# 1.35fF
C2885 w_23603_n4255# a_1596_n2079# 1.62fF
C2886 w_17090_n4258# a_1596_n2079# 1.62fF
C2887 w_10556_n4263# a_1596_n2079# 1.62fF
C2888 w_3998_n4259# a_1596_n2079# 1.62fF
C2889 w_19623_n3268# a_1596_n2079# 8.86fF
C2890 w_13110_n3271# a_1596_n2079# 8.86fF
C2891 w_6576_n3276# a_1596_n2079# 8.86fF
C2892 w_10551_n2659# a_1596_n2079# 1.63fF
C2893 w_18_n3272# a_1596_n2079# 8.87fF
C2894 w_3993_n2655# a_1596_n2079# 1.63fF
C2895 w_17085_n2654# a_1596_n2079# 1.63fF
C2896 w_23598_n2651# a_1596_n2079# 1.63fF
C2897 w_23612_n1001# a_1596_n2079# 1.65fF
C2898 w_17099_n1004# a_1596_n2079# 1.65fF
C2899 w_10565_n1009# a_1596_n2079# 1.65fF
C2900 w_4007_n1005# a_1596_n2079# 1.65fF
C2901 w_8519_n1720# a_1596_n2079# 2.69fF
C2902 w_7377_n1716# a_1596_n2079# 2.98fF
C2903 w_1961_n1716# a_1596_n2079# 2.69fF
C2904 w_819_n1712# a_1596_n2079# 2.98fF
C2905 w_15053_n1715# a_1596_n2079# 2.69fF
C2906 w_13911_n1711# a_1596_n2079# 2.98fF
C2907 w_21566_n1712# a_1596_n2079# 2.69fF
C2908 w_20424_n1708# a_1596_n2079# 2.98fF
C2909 w_20497_1345# a_1596_n2079# 1.62fF
C2910 w_13939_1341# a_1596_n2079# 1.62fF
C2911 w_7405_1346# a_1596_n2079# 1.62fF
C2912 w_892_1349# a_1596_n2079# 1.62fF
C2913 w_21965_2332# a_1596_n2079# 8.87fF
C2914 w_15407_2328# a_1596_n2079# 8.86fF
C2915 w_8873_2333# a_1596_n2079# 8.86fF
C2916 w_2360_2336# a_1596_n2079# 8.86fF
C2917 w_13944_2945# a_1596_n2079# 1.62fF
C2918 w_20502_2949# a_1596_n2079# 1.62fF
C2919 w_7410_2950# a_1596_n2079# 1.62fF
C2920 w_897_2953# a_1596_n2079# 1.62fF
C2921 w_20488_4599# a_1596_n2079# 1.65fF
C2922 w_13930_4595# a_1596_n2079# 1.65fF
C2923 w_17397_4471# a_1596_n2079# 2.98fF
C2924 w_16255_4467# a_1596_n2079# 2.70fF
C2925 w_23955_4475# a_1596_n2079# 2.98fF
C2926 w_22813_4471# a_1596_n2079# 2.70fF
C2927 w_7396_4600# a_1596_n2079# 1.65fF
C2928 w_10863_4476# a_1596_n2079# 2.99fF
C2929 w_9721_4472# a_1596_n2079# 2.70fF
C2930 w_883_4603# a_1596_n2079# 1.65fF
C2931 w_4350_4479# a_1596_n2079# 2.98fF
C2932 w_3208_4475# a_1596_n2079# 2.70fF
C2933 Y[4].t2 a_1596_n2079# 0.04fF
C2934 Y[4].t3 a_1596_n2079# 0.04fF
C2935 Y[4].n0 a_1596_n2079# 0.29fF $ **FLOATING
C2936 Y[4].t6 a_1596_n2079# 0.04fF
C2937 Y[4].t1 a_1596_n2079# 0.04fF
C2938 Y[4].n1 a_1596_n2079# 0.29fF $ **FLOATING
C2939 Y[4].t7 a_1596_n2079# 0.04fF
C2940 Y[4].t0 a_1596_n2079# 0.04fF
C2941 Y[4].n2 a_1596_n2079# 0.32fF $ **FLOATING
C2942 Y[4].t4 a_1596_n2079# 0.04fF
C2943 Y[4].t5 a_1596_n2079# 0.04fF
C2944 Y[4].n3 a_1596_n2079# 0.29fF $ **FLOATING
C2945 Y[4].n4 a_1596_n2079# 0.14fF $ **FLOATING
C2946 Y[4].n5 a_1596_n2079# 0.09fF $ **FLOATING
C2947 Y[4].n6 a_1596_n2079# 0.18fF $ **FLOATING
C2948 Y[4].n7 a_1596_n2079# 0.32fF $ **FLOATING
C2949 a_20554_n3232.t1 a_1596_n2079# 0.02fF
C2950 a_20554_n3232.t6 a_1596_n2079# 0.02fF
C2951 a_20554_n3232.t0 a_1596_n2079# 0.02fF
C2952 a_20554_n3232.n0 a_1596_n2079# 0.16fF $ **FLOATING
C2953 a_20554_n3232.t3 a_1596_n2079# 0.02fF
C2954 a_20554_n3232.t7 a_1596_n2079# 0.02fF
C2955 a_20554_n3232.n1 a_1596_n2079# 0.18fF $ **FLOATING
C2956 a_20554_n3232.t4 a_1596_n2079# 0.02fF
C2957 a_20554_n3232.t5 a_1596_n2079# 0.02fF
C2958 a_20554_n3232.n2 a_1596_n2079# 0.16fF $ **FLOATING
C2959 a_20554_n3232.n3 a_1596_n2079# 0.07fF $ **FLOATING
C2960 a_20554_n3232.n4 a_1596_n2079# 0.05fF $ **FLOATING
C2961 a_20554_n3232.t9 a_1596_n2079# 0.03fF
C2962 a_20554_n3232.t10 a_1596_n2079# 0.05fF
C2963 a_20554_n3232.n5 a_1596_n2079# 0.04fF $ **FLOATING
C2964 a_20554_n3232.t8 a_1596_n2079# 0.03fF
C2965 a_20554_n3232.t13 a_1596_n2079# 0.06fF
C2966 a_20554_n3232.t11 a_1596_n2079# 0.08fF
C2967 a_20554_n3232.n6 a_1596_n2079# 0.11fF $ **FLOATING
C2968 a_20554_n3232.t14 a_1596_n2079# 0.10fF
C2969 a_20554_n3232.n7 a_1596_n2079# 0.08fF $ **FLOATING
C2970 a_20554_n3232.n8 a_1596_n2079# 0.09fF $ **FLOATING
C2971 a_20554_n3232.t12 a_1596_n2079# 0.03fF
C2972 a_20554_n3232.t15 a_1596_n2079# 0.12fF
C2973 a_20554_n3232.n9 a_1596_n2079# 0.18fF $ **FLOATING
C2974 a_20554_n3232.n10 a_1596_n2079# 0.23fF $ **FLOATING
C2975 a_20554_n3232.n11 a_1596_n2079# 0.15fF $ **FLOATING
C2976 a_20554_n3232.n12 a_1596_n2079# 0.16fF $ **FLOATING
C2977 a_20554_n3232.t2 a_1596_n2079# 0.02fF
C2978 Y[1].t7 a_1596_n2079# 0.04fF
C2979 Y[1].t6 a_1596_n2079# 0.04fF
C2980 Y[1].n0 a_1596_n2079# 0.29fF $ **FLOATING
C2981 Y[1].t5 a_1596_n2079# 0.04fF
C2982 Y[1].t3 a_1596_n2079# 0.04fF
C2983 Y[1].n1 a_1596_n2079# 0.29fF $ **FLOATING
C2984 Y[1].t0 a_1596_n2079# 0.04fF
C2985 Y[1].t4 a_1596_n2079# 0.04fF
C2986 Y[1].n2 a_1596_n2079# 0.33fF $ **FLOATING
C2987 Y[1].t1 a_1596_n2079# 0.04fF
C2988 Y[1].t2 a_1596_n2079# 0.04fF
C2989 Y[1].n3 a_1596_n2079# 0.30fF $ **FLOATING
C2990 Y[1].n4 a_1596_n2079# 0.14fF $ **FLOATING
C2991 Y[1].n5 a_1596_n2079# 0.09fF $ **FLOATING
C2992 Y[1].n6 a_1596_n2079# 0.18fF $ **FLOATING
C2993 Y[1].n7 a_1596_n2079# 0.32fF $ **FLOATING
C2994 a_24327_1701.t1 a_1596_n2079# 0.06fF
C2995 a_24327_1701.t0 a_1596_n2079# 0.06fF
C2996 a_24327_1701.n0 a_1596_n2079# 0.45fF $ **FLOATING
C2997 a_24327_1701.t9 a_1596_n2079# 0.06fF
C2998 a_24327_1701.t10 a_1596_n2079# 0.06fF
C2999 a_24327_1701.n1 a_1596_n2079# 0.53fF $ **FLOATING
C3000 a_24327_1701.t11 a_1596_n2079# 0.06fF
C3001 a_24327_1701.t3 a_1596_n2079# 0.06fF
C3002 a_24327_1701.n2 a_1596_n2079# 0.12fF $ **FLOATING
C3003 a_24327_1701.n3 a_1596_n2079# 0.37fF $ **FLOATING
C3004 a_24327_1701.t5 a_1596_n2079# 0.06fF
C3005 a_24327_1701.t4 a_1596_n2079# 0.06fF
C3006 a_24327_1701.n4 a_1596_n2079# 0.48fF $ **FLOATING
C3007 a_24327_1701.n5 a_1596_n2079# 0.16fF $ **FLOATING
C3008 a_24327_1701.t7 a_1596_n2079# 0.06fF
C3009 a_24327_1701.t6 a_1596_n2079# 0.06fF
C3010 a_24327_1701.n6 a_1596_n2079# 0.45fF $ **FLOATING
C3011 a_24327_1701.t8 a_1596_n2079# 0.12fF
C3012 a_24327_1701.n7 a_1596_n2079# 0.71fF $ **FLOATING
C3013 a_24327_1701.n8 a_1596_n2079# 0.06fF $ **FLOATING
C3014 a_24327_1701.n9 a_1596_n2079# 0.69fF $ **FLOATING
C3015 a_24327_1701.t2 a_1596_n2079# 0.12fF
C3016 Y[5].t6 a_1596_n2079# 0.04fF
C3017 Y[5].t7 a_1596_n2079# 0.04fF
C3018 Y[5].n0 a_1596_n2079# 0.29fF $ **FLOATING
C3019 Y[5].t2 a_1596_n2079# 0.04fF
C3020 Y[5].t5 a_1596_n2079# 0.04fF
C3021 Y[5].n1 a_1596_n2079# 0.29fF $ **FLOATING
C3022 Y[5].t1 a_1596_n2079# 0.04fF
C3023 Y[5].t0 a_1596_n2079# 0.04fF
C3024 Y[5].n2 a_1596_n2079# 0.32fF $ **FLOATING
C3025 Y[5].t3 a_1596_n2079# 0.04fF
C3026 Y[5].t4 a_1596_n2079# 0.04fF
C3027 Y[5].n3 a_1596_n2079# 0.29fF $ **FLOATING
C3028 Y[5].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3029 Y[5].n5 a_1596_n2079# 0.09fF $ **FLOATING
C3030 Y[5].n6 a_1596_n2079# 0.18fF $ **FLOATING
C3031 Y[5].n7 a_1596_n2079# 0.32fF $ **FLOATING
C3032 a_15584_n3902.t0 a_1596_n2079# 0.06fF
C3033 a_15584_n3902.t1 a_1596_n2079# 0.06fF
C3034 a_15584_n3902.n0 a_1596_n2079# 0.45fF $ **FLOATING
C3035 a_15584_n3902.t4 a_1596_n2079# 0.06fF
C3036 a_15584_n3902.t5 a_1596_n2079# 0.06fF
C3037 a_15584_n3902.n1 a_1596_n2079# 0.53fF $ **FLOATING
C3038 a_15584_n3902.t6 a_1596_n2079# 0.06fF
C3039 a_15584_n3902.t3 a_1596_n2079# 0.06fF
C3040 a_15584_n3902.n2 a_1596_n2079# 0.12fF $ **FLOATING
C3041 a_15584_n3902.n3 a_1596_n2079# 0.37fF $ **FLOATING
C3042 a_15584_n3902.t7 a_1596_n2079# 0.06fF
C3043 a_15584_n3902.t8 a_1596_n2079# 0.06fF
C3044 a_15584_n3902.n4 a_1596_n2079# 0.48fF $ **FLOATING
C3045 a_15584_n3902.n5 a_1596_n2079# 0.16fF $ **FLOATING
C3046 a_15584_n3902.t10 a_1596_n2079# 0.06fF
C3047 a_15584_n3902.t11 a_1596_n2079# 0.06fF
C3048 a_15584_n3902.n6 a_1596_n2079# 0.45fF $ **FLOATING
C3049 a_15584_n3902.t9 a_1596_n2079# 0.12fF
C3050 a_15584_n3902.n7 a_1596_n2079# 0.71fF $ **FLOATING
C3051 a_15584_n3902.n8 a_1596_n2079# 0.06fF $ **FLOATING
C3052 a_15584_n3902.n9 a_1596_n2079# 0.69fF $ **FLOATING
C3053 a_15584_n3902.t2 a_1596_n2079# 0.12fF
C3054 a_13144_n3506.t2 a_1596_n2079# 0.02fF
C3055 a_13144_n3506.t0 a_1596_n2079# 0.02fF
C3056 a_13144_n3506.t1 a_1596_n2079# 0.02fF
C3057 a_13144_n3506.n0 a_1596_n2079# 0.26fF $ **FLOATING
C3058 a_13144_n3506.t18 a_1596_n2079# 0.04fF
C3059 a_13144_n3506.t17 a_1596_n2079# 0.07fF
C3060 a_13144_n3506.n1 a_1596_n2079# 0.08fF $ **FLOATING
C3061 a_13144_n3506.t19 a_1596_n2079# 0.13fF
C3062 a_13144_n3506.t4 a_1596_n2079# 0.13fF
C3063 a_13144_n3506.t9 a_1596_n2079# 0.09fF
C3064 a_13144_n3506.t15 a_1596_n2079# 0.09fF
C3065 a_13144_n3506.t16 a_1596_n2079# 0.12fF
C3066 a_13144_n3506.n2 a_1596_n2079# 0.11fF $ **FLOATING
C3067 a_13144_n3506.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3068 a_13144_n3506.t14 a_1596_n2079# 0.11fF
C3069 a_13144_n3506.t12 a_1596_n2079# 0.07fF
C3070 a_13144_n3506.n4 a_1596_n2079# 0.10fF $ **FLOATING
C3071 a_13144_n3506.t13 a_1596_n2079# 0.07fF
C3072 a_13144_n3506.t10 a_1596_n2079# 0.05fF
C3073 a_13144_n3506.t11 a_1596_n2079# 0.18fF
C3074 a_13144_n3506.n5 a_1596_n2079# 0.36fF $ **FLOATING
C3075 a_13144_n3506.n6 a_1596_n2079# 0.32fF $ **FLOATING
C3076 a_13144_n3506.n7 a_1596_n2079# 3.38fF $ **FLOATING
C3077 a_13144_n3506.t7 a_1596_n2079# 0.04fF
C3078 a_13144_n3506.t8 a_1596_n2079# 0.07fF
C3079 a_13144_n3506.n8 a_1596_n2079# 0.08fF $ **FLOATING
C3080 a_13144_n3506.t6 a_1596_n2079# 0.13fF
C3081 a_13144_n3506.t5 a_1596_n2079# 0.14fF
C3082 a_13144_n3506.n9 a_1596_n2079# 2.96fF $ **FLOATING
C3083 a_13144_n3506.n10 a_1596_n2079# 1.09fF $ **FLOATING
C3084 a_13144_n3506.n11 a_1596_n2079# 0.13fF $ **FLOATING
C3085 a_13144_n3506.t3 a_1596_n2079# 0.02fF
C3086 B[1].t13 a_1596_n2079# 0.04fF
C3087 B[1].t15 a_1596_n2079# 0.06fF
C3088 B[1].n0 a_1596_n2079# 0.07fF $ **FLOATING
C3089 B[1].t2 a_1596_n2079# 0.12fF
C3090 B[1].t7 a_1596_n2079# 0.12fF
C3091 B[1].t9 a_1596_n2079# 0.04fF
C3092 B[1].t14 a_1596_n2079# 0.08fF
C3093 B[1].t6 a_1596_n2079# 0.11fF
C3094 B[1].n1 a_1596_n2079# 0.14fF $ **FLOATING
C3095 B[1].t3 a_1596_n2079# 0.13fF
C3096 B[1].n2 a_1596_n2079# 0.10fF $ **FLOATING
C3097 B[1].t5 a_1596_n2079# 0.04fF
C3098 B[1].t4 a_1596_n2079# 0.06fF
C3099 B[1].n3 a_1596_n2079# 0.05fF $ **FLOATING
C3100 B[1].n4 a_1596_n2079# 0.03fF $ **FLOATING
C3101 B[1].t8 a_1596_n2079# 0.04fF
C3102 B[1].t10 a_1596_n2079# 0.16fF
C3103 B[1].n5 a_1596_n2079# 0.33fF $ **FLOATING
C3104 B[1].n6 a_1596_n2079# 0.38fF $ **FLOATING
C3105 B[1].n7 a_1596_n2079# 0.38fF $ **FLOATING
C3106 B[1].t11 a_1596_n2079# 0.04fF
C3107 B[1].t12 a_1596_n2079# 0.06fF
C3108 B[1].n8 a_1596_n2079# 0.07fF $ **FLOATING
C3109 B[1].t0 a_1596_n2079# 0.12fF
C3110 B[1].t1 a_1596_n2079# 0.13fF
C3111 B[1].n9 a_1596_n2079# 1.83fF $ **FLOATING
C3112 a_22429_1701.t6 a_1596_n2079# 0.06fF
C3113 a_22429_1701.t8 a_1596_n2079# 0.06fF
C3114 a_22429_1701.t7 a_1596_n2079# 0.06fF
C3115 a_22429_1701.n0 a_1596_n2079# 0.53fF $ **FLOATING
C3116 a_22429_1701.t10 a_1596_n2079# 0.06fF
C3117 a_22429_1701.t11 a_1596_n2079# 0.06fF
C3118 a_22429_1701.n1 a_1596_n2079# 0.45fF $ **FLOATING
C3119 a_22429_1701.t9 a_1596_n2079# 0.12fF
C3120 a_22429_1701.n2 a_1596_n2079# 0.69fF $ **FLOATING
C3121 a_22429_1701.t3 a_1596_n2079# 0.06fF
C3122 a_22429_1701.t5 a_1596_n2079# 0.06fF
C3123 a_22429_1701.n3 a_1596_n2079# 0.45fF $ **FLOATING
C3124 a_22429_1701.t4 a_1596_n2079# 0.12fF
C3125 a_22429_1701.n4 a_1596_n2079# 0.71fF $ **FLOATING
C3126 a_22429_1701.n5 a_1596_n2079# 0.06fF $ **FLOATING
C3127 a_22429_1701.t1 a_1596_n2079# 0.06fF
C3128 a_22429_1701.t0 a_1596_n2079# 0.06fF
C3129 a_22429_1701.n6 a_1596_n2079# 0.48fF $ **FLOATING
C3130 a_22429_1701.n7 a_1596_n2079# 0.16fF $ **FLOATING
C3131 a_22429_1701.n8 a_1596_n2079# 0.37fF $ **FLOATING
C3132 a_22429_1701.n9 a_1596_n2079# 0.12fF $ **FLOATING
C3133 a_22429_1701.t2 a_1596_n2079# 0.06fF
C3134 A[5].t2 a_1596_n2079# 0.04fF
C3135 A[5].t10 a_1596_n2079# 0.04fF
C3136 A[5].t12 a_1596_n2079# 0.05fF
C3137 A[5].n0 a_1596_n2079# 0.05fF $ **FLOATING
C3138 A[5].n1 a_1596_n2079# 0.05fF $ **FLOATING
C3139 A[5].t13 a_1596_n2079# 0.05fF
C3140 A[5].t6 a_1596_n2079# 0.03fF
C3141 A[5].n2 a_1596_n2079# 0.05fF $ **FLOATING
C3142 A[5].t8 a_1596_n2079# 0.04fF
C3143 A[5].t4 a_1596_n2079# 0.02fF
C3144 A[5].t11 a_1596_n2079# 0.08fF
C3145 A[5].n3 a_1596_n2079# 0.17fF $ **FLOATING
C3146 A[5].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3147 A[5].t3 a_1596_n2079# 0.02fF
C3148 A[5].t9 a_1596_n2079# 0.03fF
C3149 A[5].n5 a_1596_n2079# 0.04fF $ **FLOATING
C3150 A[5].t15 a_1596_n2079# 0.06fF
C3151 A[5].t1 a_1596_n2079# 0.07fF
C3152 A[5].n6 a_1596_n2079# 1.74fF $ **FLOATING
C3153 A[5].t0 a_1596_n2079# 0.02fF
C3154 A[5].t14 a_1596_n2079# 0.03fF
C3155 A[5].n7 a_1596_n2079# 0.04fF $ **FLOATING
C3156 A[5].t5 a_1596_n2079# 0.06fF
C3157 A[5].t7 a_1596_n2079# 0.06fF
C3158 A[5].n8 a_1596_n2079# 0.47fF $ **FLOATING
C3159 A[5].n9 a_1596_n2079# 0.10fF $ **FLOATING
C3160 A[0].t14 a_1596_n2079# 0.07fF
C3161 A[0].t12 a_1596_n2079# 0.09fF
C3162 A[0].t4 a_1596_n2079# 0.09fF
C3163 A[0].t13 a_1596_n2079# 0.12fF
C3164 A[0].n0 a_1596_n2079# 0.12fF $ **FLOATING
C3165 A[0].n1 a_1596_n2079# 0.11fF $ **FLOATING
C3166 A[0].t8 a_1596_n2079# 0.11fF
C3167 A[0].n2 a_1596_n2079# 0.10fF $ **FLOATING
C3168 A[0].t1 a_1596_n2079# 0.08fF
C3169 A[0].t9 a_1596_n2079# 0.05fF
C3170 A[0].t6 a_1596_n2079# 0.18fF
C3171 A[0].n3 a_1596_n2079# 0.38fF $ **FLOATING
C3172 A[0].n4 a_1596_n2079# 0.31fF $ **FLOATING
C3173 A[0].t11 a_1596_n2079# 0.04fF
C3174 A[0].t0 a_1596_n2079# 0.07fF
C3175 A[0].n5 a_1596_n2079# 0.08fF $ **FLOATING
C3176 A[0].t2 a_1596_n2079# 0.13fF
C3177 A[0].t10 a_1596_n2079# 0.15fF
C3178 A[0].n6 a_1596_n2079# 3.86fF $ **FLOATING
C3179 A[0].t15 a_1596_n2079# 0.04fF
C3180 A[0].t3 a_1596_n2079# 0.07fF
C3181 A[0].n7 a_1596_n2079# 0.08fF $ **FLOATING
C3182 A[0].t5 a_1596_n2079# 0.13fF
C3183 A[0].t7 a_1596_n2079# 0.14fF
C3184 A[0].n8 a_1596_n2079# 1.07fF $ **FLOATING
C3185 Y[2].t4 a_1596_n2079# 0.04fF
C3186 Y[2].t5 a_1596_n2079# 0.04fF
C3187 Y[2].n0 a_1596_n2079# 0.29fF $ **FLOATING
C3188 Y[2].t6 a_1596_n2079# 0.04fF
C3189 Y[2].t1 a_1596_n2079# 0.04fF
C3190 Y[2].n1 a_1596_n2079# 0.29fF $ **FLOATING
C3191 Y[2].t7 a_1596_n2079# 0.04fF
C3192 Y[2].t3 a_1596_n2079# 0.04fF
C3193 Y[2].n2 a_1596_n2079# 0.33fF $ **FLOATING
C3194 Y[2].t2 a_1596_n2079# 0.04fF
C3195 Y[2].t0 a_1596_n2079# 0.04fF
C3196 Y[2].n3 a_1596_n2079# 0.30fF $ **FLOATING
C3197 Y[2].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3198 Y[2].n5 a_1596_n2079# 0.09fF $ **FLOATING
C3199 Y[2].n6 a_1596_n2079# 0.18fF $ **FLOATING
C3200 Y[2].n7 a_1596_n2079# 0.32fF $ **FLOATING
C3201 A[6].t3 a_1596_n2079# 0.04fF
C3202 A[6].t12 a_1596_n2079# 0.04fF
C3203 A[6].t13 a_1596_n2079# 0.05fF
C3204 A[6].n0 a_1596_n2079# 0.05fF $ **FLOATING
C3205 A[6].n1 a_1596_n2079# 0.05fF $ **FLOATING
C3206 A[6].t0 a_1596_n2079# 0.05fF
C3207 A[6].t9 a_1596_n2079# 0.03fF
C3208 A[6].n2 a_1596_n2079# 0.05fF $ **FLOATING
C3209 A[6].t11 a_1596_n2079# 0.04fF
C3210 A[6].t2 a_1596_n2079# 0.02fF
C3211 A[6].t7 a_1596_n2079# 0.08fF
C3212 A[6].n3 a_1596_n2079# 0.17fF $ **FLOATING
C3213 A[6].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3214 A[6].t5 a_1596_n2079# 0.02fF
C3215 A[6].t6 a_1596_n2079# 0.03fF
C3216 A[6].n5 a_1596_n2079# 0.04fF $ **FLOATING
C3217 A[6].t4 a_1596_n2079# 0.06fF
C3218 A[6].t8 a_1596_n2079# 0.07fF
C3219 A[6].n6 a_1596_n2079# 1.74fF $ **FLOATING
C3220 A[6].t1 a_1596_n2079# 0.02fF
C3221 A[6].t14 a_1596_n2079# 0.03fF
C3222 A[6].n7 a_1596_n2079# 0.04fF $ **FLOATING
C3223 A[6].t10 a_1596_n2079# 0.06fF
C3224 A[6].t15 a_1596_n2079# 0.06fF
C3225 A[6].n8 a_1596_n2079# 0.47fF $ **FLOATING
C3226 A[6].n9 a_1596_n2079# 0.10fF $ **FLOATING
C3227 Y[0].t6 a_1596_n2079# 0.04fF
C3228 Y[0].t5 a_1596_n2079# 0.04fF
C3229 Y[0].n0 a_1596_n2079# 0.29fF $ **FLOATING
C3230 Y[0].t4 a_1596_n2079# 0.04fF
C3231 Y[0].t2 a_1596_n2079# 0.04fF
C3232 Y[0].n1 a_1596_n2079# 0.29fF $ **FLOATING
C3233 Y[0].t7 a_1596_n2079# 0.04fF
C3234 Y[0].t0 a_1596_n2079# 0.04fF
C3235 Y[0].n2 a_1596_n2079# 0.33fF $ **FLOATING
C3236 Y[0].t1 a_1596_n2079# 0.04fF
C3237 Y[0].t3 a_1596_n2079# 0.04fF
C3238 Y[0].n3 a_1596_n2079# 0.30fF $ **FLOATING
C3239 Y[0].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3240 Y[0].n5 a_1596_n2079# 0.09fF $ **FLOATING
C3241 Y[0].n6 a_1596_n2079# 0.17fF $ **FLOATING
C3242 Y[0].n7 a_1596_n2079# 0.21fF $ **FLOATING
C3243 Y[0].n8 a_1596_n2079# 0.12fF $ **FLOATING
C3244 a_17697_3950.t2 a_1596_n2079# 0.02fF
C3245 a_17697_3950.t1 a_1596_n2079# 0.02fF
C3246 a_17697_3950.n0 a_1596_n2079# 0.12fF $ **FLOATING
C3247 a_17697_3950.t10 a_1596_n2079# 0.04fF
C3248 a_17697_3950.t4 a_1596_n2079# 0.06fF
C3249 a_17697_3950.n1 a_1596_n2079# 0.08fF $ **FLOATING
C3250 a_17697_3950.t9 a_1596_n2079# 0.13fF
C3251 a_17697_3950.t15 a_1596_n2079# 0.13fF
C3252 a_17697_3950.t8 a_1596_n2079# 0.06fF
C3253 a_17697_3950.t14 a_1596_n2079# 0.09fF
C3254 a_17697_3950.t13 a_1596_n2079# 0.09fF
C3255 a_17697_3950.t7 a_1596_n2079# 0.11fF
C3256 a_17697_3950.n2 a_1596_n2079# 0.11fF $ **FLOATING
C3257 a_17697_3950.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3258 a_17697_3950.t6 a_1596_n2079# 0.10fF
C3259 a_17697_3950.n4 a_1596_n2079# 0.10fF $ **FLOATING
C3260 a_17697_3950.t18 a_1596_n2079# 0.07fF
C3261 a_17697_3950.t5 a_1596_n2079# 0.05fF
C3262 a_17697_3950.t19 a_1596_n2079# 0.17fF
C3263 a_17697_3950.n5 a_1596_n2079# 0.35fF $ **FLOATING
C3264 a_17697_3950.n6 a_1596_n2079# 0.31fF $ **FLOATING
C3265 a_17697_3950.n7 a_1596_n2079# 3.29fF $ **FLOATING
C3266 a_17697_3950.t17 a_1596_n2079# 0.04fF
C3267 a_17697_3950.t11 a_1596_n2079# 0.06fF
C3268 a_17697_3950.n8 a_1596_n2079# 0.08fF $ **FLOATING
C3269 a_17697_3950.t12 a_1596_n2079# 0.13fF
C3270 a_17697_3950.t16 a_1596_n2079# 0.13fF
C3271 a_17697_3950.n9 a_1596_n2079# 2.88fF $ **FLOATING
C3272 a_17697_3950.n10 a_1596_n2079# 1.03fF $ **FLOATING
C3273 a_17697_3950.t0 a_1596_n2079# 0.02fF
C3274 a_17697_3950.n11 a_1596_n2079# 0.26fF $ **FLOATING
C3275 a_17697_3950.t3 a_1596_n2079# 0.02fF
C3276 a_6610_n3511.t2 a_1596_n2079# 0.02fF
C3277 a_6610_n3511.t0 a_1596_n2079# 0.02fF
C3278 a_6610_n3511.t1 a_1596_n2079# 0.02fF
C3279 a_6610_n3511.n0 a_1596_n2079# 0.26fF $ **FLOATING
C3280 a_6610_n3511.t7 a_1596_n2079# 0.04fF
C3281 a_6610_n3511.t6 a_1596_n2079# 0.07fF
C3282 a_6610_n3511.n1 a_1596_n2079# 0.08fF $ **FLOATING
C3283 a_6610_n3511.t8 a_1596_n2079# 0.13fF
C3284 a_6610_n3511.t12 a_1596_n2079# 0.13fF
C3285 a_6610_n3511.t17 a_1596_n2079# 0.09fF
C3286 a_6610_n3511.t18 a_1596_n2079# 0.09fF
C3287 a_6610_n3511.t5 a_1596_n2079# 0.12fF
C3288 a_6610_n3511.n2 a_1596_n2079# 0.11fF $ **FLOATING
C3289 a_6610_n3511.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3290 a_6610_n3511.t10 a_1596_n2079# 0.11fF
C3291 a_6610_n3511.t16 a_1596_n2079# 0.07fF
C3292 a_6610_n3511.n4 a_1596_n2079# 0.10fF $ **FLOATING
C3293 a_6610_n3511.t4 a_1596_n2079# 0.07fF
C3294 a_6610_n3511.t15 a_1596_n2079# 0.05fF
C3295 a_6610_n3511.t19 a_1596_n2079# 0.18fF
C3296 a_6610_n3511.n5 a_1596_n2079# 0.36fF $ **FLOATING
C3297 a_6610_n3511.n6 a_1596_n2079# 0.32fF $ **FLOATING
C3298 a_6610_n3511.n7 a_1596_n2079# 3.39fF $ **FLOATING
C3299 a_6610_n3511.t11 a_1596_n2079# 0.04fF
C3300 a_6610_n3511.t14 a_1596_n2079# 0.07fF
C3301 a_6610_n3511.n8 a_1596_n2079# 0.08fF $ **FLOATING
C3302 a_6610_n3511.t9 a_1596_n2079# 0.13fF
C3303 a_6610_n3511.t13 a_1596_n2079# 0.14fF
C3304 a_6610_n3511.n9 a_1596_n2079# 2.98fF $ **FLOATING
C3305 a_6610_n3511.n10 a_1596_n2079# 1.10fF $ **FLOATING
C3306 a_6610_n3511.n11 a_1596_n2079# 0.13fF $ **FLOATING
C3307 a_6610_n3511.t3 a_1596_n2079# 0.02fF
C3308 a_15871_1697.t0 a_1596_n2079# 0.06fF
C3309 a_15871_1697.t1 a_1596_n2079# 0.06fF
C3310 a_15871_1697.n0 a_1596_n2079# 0.45fF $ **FLOATING
C3311 a_15871_1697.t9 a_1596_n2079# 0.06fF
C3312 a_15871_1697.t11 a_1596_n2079# 0.06fF
C3313 a_15871_1697.n1 a_1596_n2079# 0.53fF $ **FLOATING
C3314 a_15871_1697.t10 a_1596_n2079# 0.06fF
C3315 a_15871_1697.t5 a_1596_n2079# 0.06fF
C3316 a_15871_1697.n2 a_1596_n2079# 0.12fF $ **FLOATING
C3317 a_15871_1697.n3 a_1596_n2079# 0.37fF $ **FLOATING
C3318 a_15871_1697.t4 a_1596_n2079# 0.06fF
C3319 a_15871_1697.t3 a_1596_n2079# 0.06fF
C3320 a_15871_1697.n4 a_1596_n2079# 0.48fF $ **FLOATING
C3321 a_15871_1697.n5 a_1596_n2079# 0.16fF $ **FLOATING
C3322 a_15871_1697.t6 a_1596_n2079# 0.06fF
C3323 a_15871_1697.t7 a_1596_n2079# 0.06fF
C3324 a_15871_1697.n6 a_1596_n2079# 0.45fF $ **FLOATING
C3325 a_15871_1697.t8 a_1596_n2079# 0.12fF
C3326 a_15871_1697.n7 a_1596_n2079# 0.69fF $ **FLOATING
C3327 a_15871_1697.n8 a_1596_n2079# 0.06fF $ **FLOATING
C3328 a_15871_1697.n9 a_1596_n2079# 0.71fF $ **FLOATING
C3329 a_15871_1697.t2 a_1596_n2079# 0.12fF
C3330 A[3].t11 a_1596_n2079# 0.05fF
C3331 A[3].t1 a_1596_n2079# 0.07fF
C3332 A[3].t7 a_1596_n2079# 0.07fF
C3333 A[3].t9 a_1596_n2079# 0.09fF
C3334 A[3].n0 a_1596_n2079# 0.09fF $ **FLOATING
C3335 A[3].n1 a_1596_n2079# 0.08fF $ **FLOATING
C3336 A[3].t15 a_1596_n2079# 0.08fF
C3337 A[3].n2 a_1596_n2079# 0.08fF $ **FLOATING
C3338 A[3].t4 a_1596_n2079# 0.06fF
C3339 A[3].t8 a_1596_n2079# 0.04fF
C3340 A[3].t6 a_1596_n2079# 0.13fF
C3341 A[3].n3 a_1596_n2079# 0.28fF $ **FLOATING
C3342 A[3].n4 a_1596_n2079# 0.23fF $ **FLOATING
C3343 A[3].t0 a_1596_n2079# 0.03fF
C3344 A[3].t14 a_1596_n2079# 0.05fF
C3345 A[3].n5 a_1596_n2079# 0.06fF $ **FLOATING
C3346 A[3].t10 a_1596_n2079# 0.10fF
C3347 A[3].t13 a_1596_n2079# 0.11fF
C3348 A[3].n6 a_1596_n2079# 2.84fF $ **FLOATING
C3349 A[3].t12 a_1596_n2079# 0.03fF
C3350 A[3].t5 a_1596_n2079# 0.05fF
C3351 A[3].n7 a_1596_n2079# 0.06fF $ **FLOATING
C3352 A[3].t2 a_1596_n2079# 0.10fF
C3353 A[3].t3 a_1596_n2079# 0.10fF
C3354 A[3].n8 a_1596_n2079# 0.79fF $ **FLOATING
C3355 B[7].t0 a_1596_n2079# 0.02fF
C3356 B[7].t13 a_1596_n2079# 0.04fF
C3357 B[7].n0 a_1596_n2079# 0.04fF $ **FLOATING
C3358 B[7].t1 a_1596_n2079# 0.07fF
C3359 B[7].t15 a_1596_n2079# 0.07fF
C3360 B[7].t5 a_1596_n2079# 0.02fF
C3361 B[7].t7 a_1596_n2079# 0.04fF
C3362 B[7].n1 a_1596_n2079# 0.03fF $ **FLOATING
C3363 B[7].t3 a_1596_n2079# 0.02fF
C3364 B[7].t10 a_1596_n2079# 0.05fF
C3365 B[7].t9 a_1596_n2079# 0.06fF
C3366 B[7].n2 a_1596_n2079# 0.08fF $ **FLOATING
C3367 B[7].t8 a_1596_n2079# 0.07fF
C3368 B[7].n3 a_1596_n2079# 0.06fF $ **FLOATING
C3369 B[7].n4 a_1596_n2079# 0.02fF $ **FLOATING
C3370 B[7].t6 a_1596_n2079# 0.03fF
C3371 B[7].t12 a_1596_n2079# 0.09fF
C3372 B[7].n5 a_1596_n2079# 0.19fF $ **FLOATING
C3373 B[7].n6 a_1596_n2079# 0.22fF $ **FLOATING
C3374 B[7].n7 a_1596_n2079# 0.22fF $ **FLOATING
C3375 B[7].t4 a_1596_n2079# 0.02fF
C3376 B[7].t11 a_1596_n2079# 0.04fF
C3377 B[7].n8 a_1596_n2079# 0.04fF $ **FLOATING
C3378 B[7].t2 a_1596_n2079# 0.07fF
C3379 B[7].t14 a_1596_n2079# 0.07fF
C3380 B[7].n9 a_1596_n2079# 1.04fF $ **FLOATING
C3381 B[7].n10 a_1596_n2079# 0.22fF $ **FLOATING
C3382 Y[6].t2 a_1596_n2079# 0.04fF
C3383 Y[6].t0 a_1596_n2079# 0.04fF
C3384 Y[6].n0 a_1596_n2079# 0.29fF $ **FLOATING
C3385 Y[6].t6 a_1596_n2079# 0.04fF
C3386 Y[6].t1 a_1596_n2079# 0.04fF
C3387 Y[6].n1 a_1596_n2079# 0.29fF $ **FLOATING
C3388 Y[6].t7 a_1596_n2079# 0.04fF
C3389 Y[6].t3 a_1596_n2079# 0.04fF
C3390 Y[6].n2 a_1596_n2079# 0.32fF $ **FLOATING
C3391 Y[6].t4 a_1596_n2079# 0.04fF
C3392 Y[6].t5 a_1596_n2079# 0.04fF
C3393 Y[6].n3 a_1596_n2079# 0.29fF $ **FLOATING
C3394 Y[6].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3395 Y[6].n5 a_1596_n2079# 0.09fF $ **FLOATING
C3396 Y[6].n6 a_1596_n2079# 0.18fF $ **FLOATING
C3397 Y[6].n7 a_1596_n2079# 0.32fF $ **FLOATING
C3398 B[6].t7 a_1596_n2079# 0.02fF
C3399 B[6].t4 a_1596_n2079# 0.04fF
C3400 B[6].n0 a_1596_n2079# 0.04fF $ **FLOATING
C3401 B[6].t8 a_1596_n2079# 0.07fF
C3402 B[6].t10 a_1596_n2079# 0.07fF
C3403 B[6].t1 a_1596_n2079# 0.02fF
C3404 B[6].t2 a_1596_n2079# 0.04fF
C3405 B[6].n1 a_1596_n2079# 0.03fF $ **FLOATING
C3406 B[6].t11 a_1596_n2079# 0.02fF
C3407 B[6].t5 a_1596_n2079# 0.05fF
C3408 B[6].t3 a_1596_n2079# 0.06fF
C3409 B[6].n2 a_1596_n2079# 0.08fF $ **FLOATING
C3410 B[6].t6 a_1596_n2079# 0.07fF
C3411 B[6].n3 a_1596_n2079# 0.06fF $ **FLOATING
C3412 B[6].n4 a_1596_n2079# 0.02fF $ **FLOATING
C3413 B[6].t14 a_1596_n2079# 0.03fF
C3414 B[6].t9 a_1596_n2079# 0.09fF
C3415 B[6].n5 a_1596_n2079# 0.19fF $ **FLOATING
C3416 B[6].n6 a_1596_n2079# 0.22fF $ **FLOATING
C3417 B[6].n7 a_1596_n2079# 0.22fF $ **FLOATING
C3418 B[6].t12 a_1596_n2079# 0.02fF
C3419 B[6].t15 a_1596_n2079# 0.04fF
C3420 B[6].n8 a_1596_n2079# 0.04fF $ **FLOATING
C3421 B[6].t0 a_1596_n2079# 0.07fF
C3422 B[6].t13 a_1596_n2079# 0.07fF
C3423 B[6].n9 a_1596_n2079# 1.04fF $ **FLOATING
C3424 B[6].n10 a_1596_n2079# 0.22fF $ **FLOATING
C3425 A[4].t7 a_1596_n2079# 0.04fF
C3426 A[4].t3 a_1596_n2079# 0.04fF
C3427 A[4].t5 a_1596_n2079# 0.05fF
C3428 A[4].n0 a_1596_n2079# 0.05fF $ **FLOATING
C3429 A[4].n1 a_1596_n2079# 0.05fF $ **FLOATING
C3430 A[4].t2 a_1596_n2079# 0.05fF
C3431 A[4].t0 a_1596_n2079# 0.03fF
C3432 A[4].n2 a_1596_n2079# 0.05fF $ **FLOATING
C3433 A[4].t1 a_1596_n2079# 0.04fF
C3434 A[4].t14 a_1596_n2079# 0.02fF
C3435 A[4].t10 a_1596_n2079# 0.08fF
C3436 A[4].n3 a_1596_n2079# 0.17fF $ **FLOATING
C3437 A[4].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3438 A[4].t12 a_1596_n2079# 0.02fF
C3439 A[4].t13 a_1596_n2079# 0.03fF
C3440 A[4].n5 a_1596_n2079# 0.04fF $ **FLOATING
C3441 A[4].t11 a_1596_n2079# 0.06fF
C3442 A[4].t8 a_1596_n2079# 0.07fF
C3443 A[4].n6 a_1596_n2079# 1.79fF $ **FLOATING
C3444 A[4].t4 a_1596_n2079# 0.02fF
C3445 A[4].t9 a_1596_n2079# 0.03fF
C3446 A[4].n7 a_1596_n2079# 0.04fF $ **FLOATING
C3447 A[4].t6 a_1596_n2079# 0.06fF
C3448 A[4].t15 a_1596_n2079# 0.06fF
C3449 A[4].n8 a_1596_n2079# 0.48fF $ **FLOATING
C3450 A[4].n9 a_1596_n2079# 0.10fF $ **FLOATING
C3451 A[7].t0 a_1596_n2079# 0.04fF
C3452 A[7].t7 a_1596_n2079# 0.04fF
C3453 A[7].t13 a_1596_n2079# 0.05fF
C3454 A[7].n0 a_1596_n2079# 0.05fF $ **FLOATING
C3455 A[7].n1 a_1596_n2079# 0.05fF $ **FLOATING
C3456 A[7].t12 a_1596_n2079# 0.05fF
C3457 A[7].t3 a_1596_n2079# 0.03fF
C3458 A[7].n2 a_1596_n2079# 0.05fF $ **FLOATING
C3459 A[7].t11 a_1596_n2079# 0.04fF
C3460 A[7].t1 a_1596_n2079# 0.02fF
C3461 A[7].t8 a_1596_n2079# 0.08fF
C3462 A[7].n3 a_1596_n2079# 0.17fF $ **FLOATING
C3463 A[7].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3464 A[7].t9 a_1596_n2079# 0.02fF
C3465 A[7].t6 a_1596_n2079# 0.03fF
C3466 A[7].n5 a_1596_n2079# 0.04fF $ **FLOATING
C3467 A[7].t2 a_1596_n2079# 0.06fF
C3468 A[7].t5 a_1596_n2079# 0.07fF
C3469 A[7].n6 a_1596_n2079# 1.75fF $ **FLOATING
C3470 A[7].t14 a_1596_n2079# 0.02fF
C3471 A[7].t15 a_1596_n2079# 0.03fF
C3472 A[7].n7 a_1596_n2079# 0.04fF $ **FLOATING
C3473 A[7].t4 a_1596_n2079# 0.06fF
C3474 A[7].t10 a_1596_n2079# 0.06fF
C3475 A[7].n8 a_1596_n2079# 0.47fF $ **FLOATING
C3476 A[7].n9 a_1596_n2079# 0.10fF $ **FLOATING
C3477 B[2].t4 a_1596_n2079# 0.04fF
C3478 B[2].t13 a_1596_n2079# 0.06fF
C3479 B[2].n0 a_1596_n2079# 0.07fF $ **FLOATING
C3480 B[2].t15 a_1596_n2079# 0.12fF
C3481 B[2].t8 a_1596_n2079# 0.12fF
C3482 B[2].t2 a_1596_n2079# 0.04fF
C3483 B[2].t6 a_1596_n2079# 0.08fF
C3484 B[2].t1 a_1596_n2079# 0.11fF
C3485 B[2].n1 a_1596_n2079# 0.14fF $ **FLOATING
C3486 B[2].t10 a_1596_n2079# 0.13fF
C3487 B[2].n2 a_1596_n2079# 0.10fF $ **FLOATING
C3488 B[2].t12 a_1596_n2079# 0.04fF
C3489 B[2].t0 a_1596_n2079# 0.06fF
C3490 B[2].n3 a_1596_n2079# 0.05fF $ **FLOATING
C3491 B[2].n4 a_1596_n2079# 0.03fF $ **FLOATING
C3492 B[2].t5 a_1596_n2079# 0.04fF
C3493 B[2].t7 a_1596_n2079# 0.16fF
C3494 B[2].n5 a_1596_n2079# 0.33fF $ **FLOATING
C3495 B[2].n6 a_1596_n2079# 0.38fF $ **FLOATING
C3496 B[2].n7 a_1596_n2079# 0.38fF $ **FLOATING
C3497 B[2].t3 a_1596_n2079# 0.04fF
C3498 B[2].t11 a_1596_n2079# 0.06fF
C3499 B[2].n8 a_1596_n2079# 0.07fF $ **FLOATING
C3500 B[2].t9 a_1596_n2079# 0.12fF
C3501 B[2].t14 a_1596_n2079# 0.13fF
C3502 B[2].n9 a_1596_n2079# 1.82fF $ **FLOATING
C3503 a_2942_1705.t7 a_1596_n2079# 0.02fF
C3504 a_2942_1705.t3 a_1596_n2079# 0.02fF
C3505 a_2942_1705.n0 a_1596_n2079# 0.18fF $ **FLOATING
C3506 a_2942_1705.t5 a_1596_n2079# 0.02fF
C3507 a_2942_1705.t0 a_1596_n2079# 0.02fF
C3508 a_2942_1705.n1 a_1596_n2079# 0.16fF $ **FLOATING
C3509 a_2942_1705.t4 a_1596_n2079# 0.02fF
C3510 a_2942_1705.t6 a_1596_n2079# 0.02fF
C3511 a_2942_1705.n2 a_1596_n2079# 0.16fF $ **FLOATING
C3512 a_2942_1705.t14 a_1596_n2079# 0.03fF
C3513 a_2942_1705.t12 a_1596_n2079# 0.06fF
C3514 a_2942_1705.t13 a_1596_n2079# 0.08fF
C3515 a_2942_1705.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3516 a_2942_1705.t8 a_1596_n2079# 0.10fF
C3517 a_2942_1705.n4 a_1596_n2079# 0.08fF $ **FLOATING
C3518 a_2942_1705.t10 a_1596_n2079# 0.03fF
C3519 a_2942_1705.t11 a_1596_n2079# 0.05fF
C3520 a_2942_1705.n5 a_1596_n2079# 0.04fF $ **FLOATING
C3521 a_2942_1705.n6 a_1596_n2079# 0.09fF $ **FLOATING
C3522 a_2942_1705.t9 a_1596_n2079# 0.03fF
C3523 a_2942_1705.t15 a_1596_n2079# 0.12fF
C3524 a_2942_1705.n7 a_1596_n2079# 0.18fF $ **FLOATING
C3525 a_2942_1705.n8 a_1596_n2079# 0.23fF $ **FLOATING
C3526 a_2942_1705.n9 a_1596_n2079# 0.15fF $ **FLOATING
C3527 a_2942_1705.n10 a_1596_n2079# 0.05fF $ **FLOATING
C3528 a_2942_1705.n11 a_1596_n2079# 0.07fF $ **FLOATING
C3529 a_2942_1705.t1 a_1596_n2079# 0.02fF
C3530 a_2942_1705.n12 a_1596_n2079# 0.16fF $ **FLOATING
C3531 a_2942_1705.t2 a_1596_n2079# 0.02fF
C3532 A[2].t13 a_1596_n2079# 0.05fF
C3533 A[2].t14 a_1596_n2079# 0.07fF
C3534 A[2].t2 a_1596_n2079# 0.07fF
C3535 A[2].t11 a_1596_n2079# 0.09fF
C3536 A[2].n0 a_1596_n2079# 0.09fF $ **FLOATING
C3537 A[2].n1 a_1596_n2079# 0.08fF $ **FLOATING
C3538 A[2].t5 a_1596_n2079# 0.08fF
C3539 A[2].n2 a_1596_n2079# 0.08fF $ **FLOATING
C3540 A[2].t0 a_1596_n2079# 0.06fF
C3541 A[2].t1 a_1596_n2079# 0.04fF
C3542 A[2].t4 a_1596_n2079# 0.13fF
C3543 A[2].n3 a_1596_n2079# 0.28fF $ **FLOATING
C3544 A[2].n4 a_1596_n2079# 0.23fF $ **FLOATING
C3545 A[2].t6 a_1596_n2079# 0.03fF
C3546 A[2].t10 a_1596_n2079# 0.05fF
C3547 A[2].n5 a_1596_n2079# 0.06fF $ **FLOATING
C3548 A[2].t12 a_1596_n2079# 0.10fF
C3549 A[2].t7 a_1596_n2079# 0.11fF
C3550 A[2].n6 a_1596_n2079# 2.83fF $ **FLOATING
C3551 A[2].t8 a_1596_n2079# 0.03fF
C3552 A[2].t15 a_1596_n2079# 0.05fF
C3553 A[2].n7 a_1596_n2079# 0.06fF $ **FLOATING
C3554 A[2].t3 a_1596_n2079# 0.10fF
C3555 A[2].t9 a_1596_n2079# 0.10fF
C3556 A[2].n8 a_1596_n2079# 0.79fF $ **FLOATING
C3557 a_4650_3958.t2 a_1596_n2079# 0.02fF
C3558 a_4650_3958.t1 a_1596_n2079# 0.02fF
C3559 a_4650_3958.n0 a_1596_n2079# 0.12fF $ **FLOATING
C3560 a_4650_3958.t11 a_1596_n2079# 0.04fF
C3561 a_4650_3958.t6 a_1596_n2079# 0.06fF
C3562 a_4650_3958.n1 a_1596_n2079# 0.08fF $ **FLOATING
C3563 a_4650_3958.t16 a_1596_n2079# 0.13fF
C3564 a_4650_3958.t15 a_1596_n2079# 0.13fF
C3565 a_4650_3958.t12 a_1596_n2079# 0.06fF
C3566 a_4650_3958.t13 a_1596_n2079# 0.09fF
C3567 a_4650_3958.t18 a_1596_n2079# 0.09fF
C3568 a_4650_3958.t7 a_1596_n2079# 0.11fF
C3569 a_4650_3958.n2 a_1596_n2079# 0.11fF $ **FLOATING
C3570 a_4650_3958.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3571 a_4650_3958.t9 a_1596_n2079# 0.10fF
C3572 a_4650_3958.n4 a_1596_n2079# 0.10fF $ **FLOATING
C3573 a_4650_3958.t17 a_1596_n2079# 0.07fF
C3574 a_4650_3958.t10 a_1596_n2079# 0.05fF
C3575 a_4650_3958.t5 a_1596_n2079# 0.17fF
C3576 a_4650_3958.n5 a_1596_n2079# 0.35fF $ **FLOATING
C3577 a_4650_3958.n6 a_1596_n2079# 0.31fF $ **FLOATING
C3578 a_4650_3958.n7 a_1596_n2079# 3.29fF $ **FLOATING
C3579 a_4650_3958.t8 a_1596_n2079# 0.04fF
C3580 a_4650_3958.t14 a_1596_n2079# 0.06fF
C3581 a_4650_3958.n8 a_1596_n2079# 0.08fF $ **FLOATING
C3582 a_4650_3958.t19 a_1596_n2079# 0.13fF
C3583 a_4650_3958.t4 a_1596_n2079# 0.13fF
C3584 a_4650_3958.n9 a_1596_n2079# 2.95fF $ **FLOATING
C3585 a_4650_3958.n10 a_1596_n2079# 1.08fF $ **FLOATING
C3586 a_4650_3958.t0 a_1596_n2079# 0.02fF
C3587 a_4650_3958.n11 a_1596_n2079# 0.25fF $ **FLOATING
C3588 a_4650_3958.t3 a_1596_n2079# 0.02fF
C3589 a_7507_n3240.t3 a_1596_n2079# 0.02fF
C3590 a_7507_n3240.t4 a_1596_n2079# 0.02fF
C3591 a_7507_n3240.n0 a_1596_n2079# 0.18fF $ **FLOATING
C3592 a_7507_n3240.t1 a_1596_n2079# 0.02fF
C3593 a_7507_n3240.t5 a_1596_n2079# 0.02fF
C3594 a_7507_n3240.n1 a_1596_n2079# 0.16fF $ **FLOATING
C3595 a_7507_n3240.t6 a_1596_n2079# 0.02fF
C3596 a_7507_n3240.t7 a_1596_n2079# 0.02fF
C3597 a_7507_n3240.n2 a_1596_n2079# 0.16fF $ **FLOATING
C3598 a_7507_n3240.t8 a_1596_n2079# 0.03fF
C3599 a_7507_n3240.t9 a_1596_n2079# 0.05fF
C3600 a_7507_n3240.n3 a_1596_n2079# 0.04fF $ **FLOATING
C3601 a_7507_n3240.t13 a_1596_n2079# 0.03fF
C3602 a_7507_n3240.t11 a_1596_n2079# 0.06fF
C3603 a_7507_n3240.t10 a_1596_n2079# 0.08fF
C3604 a_7507_n3240.n4 a_1596_n2079# 0.11fF $ **FLOATING
C3605 a_7507_n3240.t12 a_1596_n2079# 0.10fF
C3606 a_7507_n3240.n5 a_1596_n2079# 0.08fF $ **FLOATING
C3607 a_7507_n3240.n6 a_1596_n2079# 0.09fF $ **FLOATING
C3608 a_7507_n3240.t15 a_1596_n2079# 0.03fF
C3609 a_7507_n3240.t14 a_1596_n2079# 0.12fF
C3610 a_7507_n3240.n7 a_1596_n2079# 0.18fF $ **FLOATING
C3611 a_7507_n3240.n8 a_1596_n2079# 0.23fF $ **FLOATING
C3612 a_7507_n3240.n9 a_1596_n2079# 0.15fF $ **FLOATING
C3613 a_7507_n3240.n10 a_1596_n2079# 0.05fF $ **FLOATING
C3614 a_7507_n3240.n11 a_1596_n2079# 0.07fF $ **FLOATING
C3615 a_7507_n3240.t0 a_1596_n2079# 0.02fF
C3616 a_7507_n3240.n12 a_1596_n2079# 0.16fF $ **FLOATING
C3617 a_7507_n3240.t2 a_1596_n2079# 0.02fF
C3618 B[5].t14 a_1596_n2079# 0.02fF
C3619 B[5].t13 a_1596_n2079# 0.04fF
C3620 B[5].n0 a_1596_n2079# 0.04fF $ **FLOATING
C3621 B[5].t2 a_1596_n2079# 0.07fF
C3622 B[5].t1 a_1596_n2079# 0.07fF
C3623 B[5].t5 a_1596_n2079# 0.02fF
C3624 B[5].t8 a_1596_n2079# 0.04fF
C3625 B[5].n1 a_1596_n2079# 0.03fF $ **FLOATING
C3626 B[5].t4 a_1596_n2079# 0.02fF
C3627 B[5].t10 a_1596_n2079# 0.05fF
C3628 B[5].t12 a_1596_n2079# 0.06fF
C3629 B[5].n2 a_1596_n2079# 0.08fF $ **FLOATING
C3630 B[5].t11 a_1596_n2079# 0.07fF
C3631 B[5].n3 a_1596_n2079# 0.06fF $ **FLOATING
C3632 B[5].n4 a_1596_n2079# 0.02fF $ **FLOATING
C3633 B[5].t7 a_1596_n2079# 0.03fF
C3634 B[5].t6 a_1596_n2079# 0.09fF
C3635 B[5].n5 a_1596_n2079# 0.19fF $ **FLOATING
C3636 B[5].n6 a_1596_n2079# 0.22fF $ **FLOATING
C3637 B[5].n7 a_1596_n2079# 0.22fF $ **FLOATING
C3638 B[5].t3 a_1596_n2079# 0.02fF
C3639 B[5].t9 a_1596_n2079# 0.04fF
C3640 B[5].n8 a_1596_n2079# 0.04fF $ **FLOATING
C3641 B[5].t15 a_1596_n2079# 0.07fF
C3642 B[5].t0 a_1596_n2079# 0.07fF
C3643 B[5].n9 a_1596_n2079# 1.04fF $ **FLOATING
C3644 B[5].n10 a_1596_n2079# 0.22fF $ **FLOATING
C3645 a_949_n3236.t1 a_1596_n2079# 0.02fF
C3646 a_949_n3236.t3 a_1596_n2079# 0.02fF
C3647 a_949_n3236.t4 a_1596_n2079# 0.02fF
C3648 a_949_n3236.n0 a_1596_n2079# 0.18fF $ **FLOATING
C3649 a_949_n3236.t0 a_1596_n2079# 0.02fF
C3650 a_949_n3236.t5 a_1596_n2079# 0.02fF
C3651 a_949_n3236.n1 a_1596_n2079# 0.16fF $ **FLOATING
C3652 a_949_n3236.t6 a_1596_n2079# 0.02fF
C3653 a_949_n3236.t7 a_1596_n2079# 0.02fF
C3654 a_949_n3236.n2 a_1596_n2079# 0.16fF $ **FLOATING
C3655 a_949_n3236.t11 a_1596_n2079# 0.03fF
C3656 a_949_n3236.t13 a_1596_n2079# 0.05fF
C3657 a_949_n3236.n3 a_1596_n2079# 0.04fF $ **FLOATING
C3658 a_949_n3236.t10 a_1596_n2079# 0.03fF
C3659 a_949_n3236.t14 a_1596_n2079# 0.06fF
C3660 a_949_n3236.t9 a_1596_n2079# 0.08fF
C3661 a_949_n3236.n4 a_1596_n2079# 0.11fF $ **FLOATING
C3662 a_949_n3236.t15 a_1596_n2079# 0.10fF
C3663 a_949_n3236.n5 a_1596_n2079# 0.08fF $ **FLOATING
C3664 a_949_n3236.n6 a_1596_n2079# 0.09fF $ **FLOATING
C3665 a_949_n3236.t12 a_1596_n2079# 0.03fF
C3666 a_949_n3236.t8 a_1596_n2079# 0.12fF
C3667 a_949_n3236.n7 a_1596_n2079# 0.18fF $ **FLOATING
C3668 a_949_n3236.n8 a_1596_n2079# 0.23fF $ **FLOATING
C3669 a_949_n3236.n9 a_1596_n2079# 0.15fF $ **FLOATING
C3670 a_949_n3236.n10 a_1596_n2079# 0.05fF $ **FLOATING
C3671 a_949_n3236.n11 a_1596_n2079# 0.07fF $ **FLOATING
C3672 a_949_n3236.n12 a_1596_n2079# 0.16fF $ **FLOATING
C3673 a_949_n3236.t2 a_1596_n2079# 0.02fF
C3674 Y[3].t2 a_1596_n2079# 0.04fF
C3675 Y[3].t1 a_1596_n2079# 0.04fF
C3676 Y[3].n0 a_1596_n2079# 0.29fF $ **FLOATING
C3677 Y[3].t0 a_1596_n2079# 0.04fF
C3678 Y[3].t6 a_1596_n2079# 0.04fF
C3679 Y[3].n1 a_1596_n2079# 0.29fF $ **FLOATING
C3680 Y[3].t3 a_1596_n2079# 0.04fF
C3681 Y[3].t5 a_1596_n2079# 0.04fF
C3682 Y[3].n2 a_1596_n2079# 0.33fF $ **FLOATING
C3683 Y[3].t7 a_1596_n2079# 0.04fF
C3684 Y[3].t4 a_1596_n2079# 0.04fF
C3685 Y[3].n3 a_1596_n2079# 0.30fF $ **FLOATING
C3686 Y[3].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3687 Y[3].n5 a_1596_n2079# 0.09fF $ **FLOATING
C3688 Y[3].n6 a_1596_n2079# 0.18fF $ **FLOATING
C3689 Y[3].n7 a_1596_n2079# 0.32fF $ **FLOATING
C3690 a_11163_3955.t2 a_1596_n2079# 0.02fF
C3691 a_11163_3955.t1 a_1596_n2079# 0.02fF
C3692 a_11163_3955.n0 a_1596_n2079# 0.12fF $ **FLOATING
C3693 a_11163_3955.t17 a_1596_n2079# 0.04fF
C3694 a_11163_3955.t11 a_1596_n2079# 0.06fF
C3695 a_11163_3955.n1 a_1596_n2079# 0.08fF $ **FLOATING
C3696 a_11163_3955.t10 a_1596_n2079# 0.13fF
C3697 a_11163_3955.t7 a_1596_n2079# 0.13fF
C3698 a_11163_3955.t4 a_1596_n2079# 0.07fF
C3699 a_11163_3955.t9 a_1596_n2079# 0.09fF
C3700 a_11163_3955.t14 a_1596_n2079# 0.09fF
C3701 a_11163_3955.t5 a_1596_n2079# 0.11fF
C3702 a_11163_3955.n2 a_1596_n2079# 0.11fF $ **FLOATING
C3703 a_11163_3955.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3704 a_11163_3955.t18 a_1596_n2079# 0.10fF
C3705 a_11163_3955.n4 a_1596_n2079# 0.10fF $ **FLOATING
C3706 a_11163_3955.t8 a_1596_n2079# 0.07fF
C3707 a_11163_3955.t13 a_1596_n2079# 0.05fF
C3708 a_11163_3955.t15 a_1596_n2079# 0.17fF
C3709 a_11163_3955.n5 a_1596_n2079# 0.36fF $ **FLOATING
C3710 a_11163_3955.n6 a_1596_n2079# 0.31fF $ **FLOATING
C3711 a_11163_3955.n7 a_1596_n2079# 3.31fF $ **FLOATING
C3712 a_11163_3955.t12 a_1596_n2079# 0.04fF
C3713 a_11163_3955.t19 a_1596_n2079# 0.06fF
C3714 a_11163_3955.n8 a_1596_n2079# 0.08fF $ **FLOATING
C3715 a_11163_3955.t6 a_1596_n2079# 0.13fF
C3716 a_11163_3955.t16 a_1596_n2079# 0.13fF
C3717 a_11163_3955.n9 a_1596_n2079# 2.92fF $ **FLOATING
C3718 a_11163_3955.n10 a_1596_n2079# 1.07fF $ **FLOATING
C3719 a_11163_3955.t0 a_1596_n2079# 0.02fF
C3720 a_11163_3955.n11 a_1596_n2079# 0.26fF $ **FLOATING
C3721 a_11163_3955.t3 a_1596_n2079# 0.02fF
C3722 a_9455_1702.t0 a_1596_n2079# 0.02fF
C3723 a_9455_1702.t4 a_1596_n2079# 0.02fF
C3724 a_9455_1702.t3 a_1596_n2079# 0.02fF
C3725 a_9455_1702.n0 a_1596_n2079# 0.18fF $ **FLOATING
C3726 a_9455_1702.t6 a_1596_n2079# 0.02fF
C3727 a_9455_1702.t1 a_1596_n2079# 0.02fF
C3728 a_9455_1702.n1 a_1596_n2079# 0.16fF $ **FLOATING
C3729 a_9455_1702.t5 a_1596_n2079# 0.02fF
C3730 a_9455_1702.t7 a_1596_n2079# 0.02fF
C3731 a_9455_1702.n2 a_1596_n2079# 0.16fF $ **FLOATING
C3732 a_9455_1702.t9 a_1596_n2079# 0.03fF
C3733 a_9455_1702.t8 a_1596_n2079# 0.06fF
C3734 a_9455_1702.t15 a_1596_n2079# 0.08fF
C3735 a_9455_1702.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3736 a_9455_1702.t13 a_1596_n2079# 0.10fF
C3737 a_9455_1702.n4 a_1596_n2079# 0.08fF $ **FLOATING
C3738 a_9455_1702.t11 a_1596_n2079# 0.03fF
C3739 a_9455_1702.t14 a_1596_n2079# 0.05fF
C3740 a_9455_1702.n5 a_1596_n2079# 0.04fF $ **FLOATING
C3741 a_9455_1702.n6 a_1596_n2079# 0.09fF $ **FLOATING
C3742 a_9455_1702.t12 a_1596_n2079# 0.03fF
C3743 a_9455_1702.t10 a_1596_n2079# 0.12fF
C3744 a_9455_1702.n7 a_1596_n2079# 0.18fF $ **FLOATING
C3745 a_9455_1702.n8 a_1596_n2079# 0.23fF $ **FLOATING
C3746 a_9455_1702.n9 a_1596_n2079# 0.15fF $ **FLOATING
C3747 a_9455_1702.n10 a_1596_n2079# 0.05fF $ **FLOATING
C3748 a_9455_1702.n11 a_1596_n2079# 0.07fF $ **FLOATING
C3749 a_9455_1702.n12 a_1596_n2079# 0.16fF $ **FLOATING
C3750 a_9455_1702.t2 a_1596_n2079# 0.02fF
C3751 Y[7].t1 a_1596_n2079# 0.04fF
C3752 Y[7].t2 a_1596_n2079# 0.04fF
C3753 Y[7].n0 a_1596_n2079# 0.29fF $ **FLOATING
C3754 Y[7].t6 a_1596_n2079# 0.04fF
C3755 Y[7].t3 a_1596_n2079# 0.04fF
C3756 Y[7].n1 a_1596_n2079# 0.29fF $ **FLOATING
C3757 Y[7].t7 a_1596_n2079# 0.04fF
C3758 Y[7].t0 a_1596_n2079# 0.04fF
C3759 Y[7].n2 a_1596_n2079# 0.32fF $ **FLOATING
C3760 Y[7].t4 a_1596_n2079# 0.04fF
C3761 Y[7].t5 a_1596_n2079# 0.04fF
C3762 Y[7].n3 a_1596_n2079# 0.29fF $ **FLOATING
C3763 Y[7].n4 a_1596_n2079# 0.14fF $ **FLOATING
C3764 Y[7].n5 a_1596_n2079# 0.09fF $ **FLOATING
C3765 Y[7].n6 a_1596_n2079# 0.18fF $ **FLOATING
C3766 Y[7].n7 a_1596_n2079# 0.32fF $ **FLOATING
C3767 B[4].t5 a_1596_n2079# 0.02fF
C3768 B[4].t4 a_1596_n2079# 0.04fF
C3769 B[4].n0 a_1596_n2079# 0.04fF $ **FLOATING
C3770 B[4].t6 a_1596_n2079# 0.07fF
C3771 B[4].t8 a_1596_n2079# 0.07fF
C3772 B[4].t12 a_1596_n2079# 0.02fF
C3773 B[4].t13 a_1596_n2079# 0.04fF
C3774 B[4].n1 a_1596_n2079# 0.03fF $ **FLOATING
C3775 B[4].t15 a_1596_n2079# 0.02fF
C3776 B[4].t3 a_1596_n2079# 0.05fF
C3777 B[4].t1 a_1596_n2079# 0.06fF
C3778 B[4].n2 a_1596_n2079# 0.08fF $ **FLOATING
C3779 B[4].t9 a_1596_n2079# 0.07fF
C3780 B[4].n3 a_1596_n2079# 0.06fF $ **FLOATING
C3781 B[4].n4 a_1596_n2079# 0.02fF $ **FLOATING
C3782 B[4].t2 a_1596_n2079# 0.03fF
C3783 B[4].t10 a_1596_n2079# 0.09fF
C3784 B[4].n5 a_1596_n2079# 0.19fF $ **FLOATING
C3785 B[4].n6 a_1596_n2079# 0.22fF $ **FLOATING
C3786 B[4].n7 a_1596_n2079# 0.22fF $ **FLOATING
C3787 B[4].t7 a_1596_n2079# 0.02fF
C3788 B[4].t14 a_1596_n2079# 0.04fF
C3789 B[4].n8 a_1596_n2079# 0.04fF $ **FLOATING
C3790 B[4].t0 a_1596_n2079# 0.07fF
C3791 B[4].t11 a_1596_n2079# 0.07fF
C3792 B[4].n9 a_1596_n2079# 1.04fF $ **FLOATING
C3793 B[4].n10 a_1596_n2079# 0.22fF $ **FLOATING
C3794 carry_in.t4 a_1596_n2079# 0.02fF
C3795 carry_in.t15 a_1596_n2079# 0.04fF
C3796 carry_in.n0 a_1596_n2079# 0.05fF $ **FLOATING
C3797 carry_in.t14 a_1596_n2079# 0.08fF
C3798 carry_in.t5 a_1596_n2079# 0.08fF
C3799 carry_in.t2 a_1596_n2079# 0.04fF
C3800 carry_in.t3 a_1596_n2079# 0.05fF
C3801 carry_in.t8 a_1596_n2079# 0.05fF
C3802 carry_in.t6 a_1596_n2079# 0.07fF
C3803 carry_in.n1 a_1596_n2079# 0.07fF $ **FLOATING
C3804 carry_in.n2 a_1596_n2079# 0.07fF $ **FLOATING
C3805 carry_in.t0 a_1596_n2079# 0.06fF
C3806 carry_in.n3 a_1596_n2079# 0.06fF $ **FLOATING
C3807 carry_in.t11 a_1596_n2079# 0.04fF
C3808 carry_in.t1 a_1596_n2079# 0.03fF
C3809 carry_in.t13 a_1596_n2079# 0.10fF
C3810 carry_in.n4 a_1596_n2079# 0.21fF $ **FLOATING
C3811 carry_in.n5 a_1596_n2079# 0.19fF $ **FLOATING
C3812 carry_in.n6 a_1596_n2079# 1.99fF $ **FLOATING
C3813 carry_in.t12 a_1596_n2079# 0.02fF
C3814 carry_in.t9 a_1596_n2079# 0.04fF
C3815 carry_in.n7 a_1596_n2079# 0.05fF $ **FLOATING
C3816 carry_in.t7 a_1596_n2079# 0.08fF
C3817 carry_in.t10 a_1596_n2079# 0.08fF
C3818 carry_in.n8 a_1596_n2079# 0.83fF $ **FLOATING
C3819 a_52_n3507.t2 a_1596_n2079# 0.02fF
C3820 a_52_n3507.t0 a_1596_n2079# 0.02fF
C3821 a_52_n3507.t1 a_1596_n2079# 0.02fF
C3822 a_52_n3507.n0 a_1596_n2079# 0.26fF $ **FLOATING
C3823 a_52_n3507.t14 a_1596_n2079# 0.04fF
C3824 a_52_n3507.t13 a_1596_n2079# 0.07fF
C3825 a_52_n3507.n1 a_1596_n2079# 0.08fF $ **FLOATING
C3826 a_52_n3507.t16 a_1596_n2079# 0.13fF
C3827 a_52_n3507.t4 a_1596_n2079# 0.13fF
C3828 a_52_n3507.t9 a_1596_n2079# 0.09fF
C3829 a_52_n3507.t15 a_1596_n2079# 0.09fF
C3830 a_52_n3507.t18 a_1596_n2079# 0.12fF
C3831 a_52_n3507.n2 a_1596_n2079# 0.11fF $ **FLOATING
C3832 a_52_n3507.n3 a_1596_n2079# 0.11fF $ **FLOATING
C3833 a_52_n3507.t19 a_1596_n2079# 0.11fF
C3834 a_52_n3507.t11 a_1596_n2079# 0.07fF
C3835 a_52_n3507.n4 a_1596_n2079# 0.10fF $ **FLOATING
C3836 a_52_n3507.t12 a_1596_n2079# 0.07fF
C3837 a_52_n3507.t10 a_1596_n2079# 0.05fF
C3838 a_52_n3507.t17 a_1596_n2079# 0.18fF
C3839 a_52_n3507.n5 a_1596_n2079# 0.36fF $ **FLOATING
C3840 a_52_n3507.n6 a_1596_n2079# 0.32fF $ **FLOATING
C3841 a_52_n3507.n7 a_1596_n2079# 3.38fF $ **FLOATING
C3842 a_52_n3507.t8 a_1596_n2079# 0.04fF
C3843 a_52_n3507.t7 a_1596_n2079# 0.07fF
C3844 a_52_n3507.n8 a_1596_n2079# 0.08fF $ **FLOATING
C3845 a_52_n3507.t6 a_1596_n2079# 0.13fF
C3846 a_52_n3507.t5 a_1596_n2079# 0.14fF
C3847 a_52_n3507.n9 a_1596_n2079# 2.96fF $ **FLOATING
C3848 a_52_n3507.n10 a_1596_n2079# 1.09fF $ **FLOATING
C3849 a_52_n3507.n11 a_1596_n2079# 0.13fF $ **FLOATING
C3850 a_52_n3507.t3 a_1596_n2079# 0.02fF
C3851 A[1].t14 a_1596_n2079# 0.05fF
C3852 A[1].t3 a_1596_n2079# 0.07fF
C3853 A[1].t5 a_1596_n2079# 0.07fF
C3854 A[1].t10 a_1596_n2079# 0.09fF
C3855 A[1].n0 a_1596_n2079# 0.09fF $ **FLOATING
C3856 A[1].n1 a_1596_n2079# 0.08fF $ **FLOATING
C3857 A[1].t11 a_1596_n2079# 0.08fF
C3858 A[1].n2 a_1596_n2079# 0.08fF $ **FLOATING
C3859 A[1].t2 a_1596_n2079# 0.06fF
C3860 A[1].t0 a_1596_n2079# 0.04fF
C3861 A[1].t8 a_1596_n2079# 0.13fF
C3862 A[1].n3 a_1596_n2079# 0.28fF $ **FLOATING
C3863 A[1].n4 a_1596_n2079# 0.23fF $ **FLOATING
C3864 A[1].t4 a_1596_n2079# 0.03fF
C3865 A[1].t15 a_1596_n2079# 0.05fF
C3866 A[1].n5 a_1596_n2079# 0.06fF $ **FLOATING
C3867 A[1].t1 a_1596_n2079# 0.10fF
C3868 A[1].t12 a_1596_n2079# 0.11fF
C3869 A[1].n6 a_1596_n2079# 2.83fF $ **FLOATING
C3870 A[1].t13 a_1596_n2079# 0.03fF
C3871 A[1].t9 a_1596_n2079# 0.05fF
C3872 A[1].n7 a_1596_n2079# 0.06fF $ **FLOATING
C3873 A[1].t6 a_1596_n2079# 0.10fF
C3874 A[1].t7 a_1596_n2079# 0.10fF
C3875 A[1].n8 a_1596_n2079# 0.79fF $ **FLOATING
C3876 VSS.t4 a_1596_n2079# 0.01fF
C3877 VSS.t49 a_1596_n2079# 0.01fF
C3878 VSS.t25 a_1596_n2079# 0.01fF
C3879 VSS.n0 a_1596_n2079# 0.04fF $ **FLOATING
C3880 VSS.n1 a_1596_n2079# 0.05fF $ **FLOATING
C3881 VSS.t69 a_1596_n2079# 0.01fF
C3882 VSS.n2 a_1596_n2079# 0.06fF $ **FLOATING
C3883 VSS.t132 a_1596_n2079# 0.00fF
C3884 VSS.t80 a_1596_n2079# 0.01fF
C3885 VSS.n3 a_1596_n2079# 0.14fF $ **FLOATING
C3886 VSS.t134 a_1596_n2079# 0.00fF
C3887 VSS.t139 a_1596_n2079# 0.01fF
C3888 VSS.n4 a_1596_n2079# 0.11fF $ **FLOATING
C3889 VSS.t98 a_1596_n2079# 0.00fF
C3890 VSS.t73 a_1596_n2079# 0.01fF
C3891 VSS.n5 a_1596_n2079# 0.11fF $ **FLOATING
C3892 VSS.t61 a_1596_n2079# 0.01fF
C3893 VSS.t43 a_1596_n2079# 0.01fF
C3894 VSS.t41 a_1596_n2079# 0.01fF
C3895 VSS.t109 a_1596_n2079# 0.01fF
C3896 VSS.n6 a_1596_n2079# 0.04fF $ **FLOATING
C3897 VSS.n7 a_1596_n2079# 0.05fF $ **FLOATING
C3898 VSS.n8 a_1596_n2079# 0.06fF $ **FLOATING
C3899 VSS.n9 a_1596_n2079# 0.03fF $ **FLOATING
C3900 VSS.n10 a_1596_n2079# 0.19fF $ **FLOATING
C3901 VSS.t65 a_1596_n2079# 0.00fF
C3902 VSS.t22 a_1596_n2079# 0.00fF
C3903 VSS.t135 a_1596_n2079# 0.00fF
C3904 VSS.n11 a_1596_n2079# 0.02fF $ **FLOATING
C3905 VSS.n12 a_1596_n2079# 0.04fF $ **FLOATING
C3906 VSS.t122 a_1596_n2079# 0.00fF
C3907 VSS.t36 a_1596_n2079# 0.01fF
C3908 VSS.n13 a_1596_n2079# 0.09fF $ **FLOATING
C3909 VSS.n14 a_1596_n2079# 0.19fF $ **FLOATING
C3910 VSS.n15 a_1596_n2079# 0.01fF $ **FLOATING
C3911 VSS.n16 a_1596_n2079# 0.03fF $ **FLOATING
C3912 VSS.n17 a_1596_n2079# 0.03fF $ **FLOATING
C3913 VSS.t151 a_1596_n2079# 0.01fF
C3914 VSS.t107 a_1596_n2079# 0.01fF
C3915 VSS.t123 a_1596_n2079# 0.01fF
C3916 VSS.t145 a_1596_n2079# 0.01fF
C3917 VSS.n18 a_1596_n2079# 0.04fF $ **FLOATING
C3918 VSS.n19 a_1596_n2079# 0.05fF $ **FLOATING
C3919 VSS.n20 a_1596_n2079# 0.06fF $ **FLOATING
C3920 VSS.n21 a_1596_n2079# 0.04fF $ **FLOATING
C3921 VSS.n22 a_1596_n2079# 0.01fF $ **FLOATING
C3922 VSS.t124 a_1596_n2079# 0.00fF
C3923 VSS.t29 a_1596_n2079# 0.01fF
C3924 VSS.n23 a_1596_n2079# 0.09fF $ **FLOATING
C3925 VSS.t16 a_1596_n2079# 0.00fF
C3926 VSS.t79 a_1596_n2079# 0.00fF
C3927 VSS.t66 a_1596_n2079# 0.00fF
C3928 VSS.n24 a_1596_n2079# 0.02fF $ **FLOATING
C3929 VSS.n25 a_1596_n2079# 0.04fF $ **FLOATING
C3930 VSS.t45 a_1596_n2079# 0.00fF
C3931 VSS.t76 a_1596_n2079# 0.01fF
C3932 VSS.n26 a_1596_n2079# 0.09fF $ **FLOATING
C3933 VSS.n27 a_1596_n2079# 0.19fF $ **FLOATING
C3934 VSS.t9 a_1596_n2079# 0.01fF
C3935 VSS.t110 a_1596_n2079# 0.01fF
C3936 VSS.t81 a_1596_n2079# 0.01fF
C3937 VSS.t86 a_1596_n2079# 0.01fF
C3938 VSS.n28 a_1596_n2079# 0.04fF $ **FLOATING
C3939 VSS.n29 a_1596_n2079# 0.05fF $ **FLOATING
C3940 VSS.n30 a_1596_n2079# 0.06fF $ **FLOATING
C3941 VSS.n31 a_1596_n2079# 1.15fF $ **FLOATING
C3942 VSS.n32 a_1596_n2079# 0.22fF $ **FLOATING
C3943 VSS.t157 a_1596_n2079# 0.01fF
C3944 VSS.t72 a_1596_n2079# 0.01fF
C3945 VSS.t118 a_1596_n2079# 0.01fF
C3946 VSS.t114 a_1596_n2079# 0.01fF
C3947 VSS.n33 a_1596_n2079# 0.04fF $ **FLOATING
C3948 VSS.n34 a_1596_n2079# 0.05fF $ **FLOATING
C3949 VSS.n35 a_1596_n2079# 0.06fF $ **FLOATING
C3950 VSS.n36 a_1596_n2079# 0.05fF $ **FLOATING
C3951 VSS.t21 a_1596_n2079# 0.00fF
C3952 VSS.t100 a_1596_n2079# 0.01fF
C3953 VSS.n37 a_1596_n2079# 0.09fF $ **FLOATING
C3954 VSS.t159 a_1596_n2079# 0.00fF
C3955 VSS.t155 a_1596_n2079# 0.01fF
C3956 VSS.n38 a_1596_n2079# 0.09fF $ **FLOATING
C3957 VSS.t152 a_1596_n2079# 0.00fF
C3958 VSS.t156 a_1596_n2079# 0.01fF
C3959 VSS.n39 a_1596_n2079# 0.11fF $ **FLOATING
C3960 VSS.n40 a_1596_n2079# 6.25fF $ **FLOATING
C3961 VSS.n41 a_1596_n2079# 2.41fF $ **FLOATING
C3962 VSS.t46 a_1596_n2079# 0.00fF
C3963 VSS.t12 a_1596_n2079# 0.00fF
C3964 VSS.t51 a_1596_n2079# 0.00fF
C3965 VSS.n42 a_1596_n2079# 0.02fF $ **FLOATING
C3966 VSS.n43 a_1596_n2079# 0.04fF $ **FLOATING
C3967 VSS.n44 a_1596_n2079# 3.30fF $ **FLOATING
C3968 VSS.t19 a_1596_n2079# 0.00fF
C3969 VSS.t70 a_1596_n2079# 0.00fF
C3970 VSS.t57 a_1596_n2079# 0.00fF
C3971 VSS.n45 a_1596_n2079# 0.02fF $ **FLOATING
C3972 VSS.n46 a_1596_n2079# 0.04fF $ **FLOATING
C3973 VSS.n47 a_1596_n2079# 4.21fF $ **FLOATING
C3974 VSS.n48 a_1596_n2079# 2.72fF $ **FLOATING
C3975 VSS.n49 a_1596_n2079# 2.34fF $ **FLOATING
C3976 VSS.t50 a_1596_n2079# 0.00fF
C3977 VSS.t11 a_1596_n2079# 0.01fF
C3978 VSS.n50 a_1596_n2079# 0.09fF $ **FLOATING
C3979 VSS.t64 a_1596_n2079# 0.00fF
C3980 VSS.t6 a_1596_n2079# 0.01fF
C3981 VSS.n51 a_1596_n2079# 0.09fF $ **FLOATING
C3982 VSS.n52 a_1596_n2079# 5.21fF $ **FLOATING
C3983 VSS.t94 a_1596_n2079# 0.01fF
C3984 VSS.t62 a_1596_n2079# 0.01fF
C3985 VSS.t121 a_1596_n2079# 0.01fF
C3986 VSS.t119 a_1596_n2079# 0.01fF
C3987 VSS.n53 a_1596_n2079# 0.04fF $ **FLOATING
C3988 VSS.n54 a_1596_n2079# 0.05fF $ **FLOATING
C3989 VSS.n55 a_1596_n2079# 0.06fF $ **FLOATING
C3990 VSS.n56 a_1596_n2079# 0.26fF $ **FLOATING
C3991 VSS.n57 a_1596_n2079# 6.43fF $ **FLOATING
C3992 VSS.t67 a_1596_n2079# 0.00fF
C3993 VSS.t158 a_1596_n2079# 0.00fF
C3994 VSS.t5 a_1596_n2079# 0.00fF
C3995 VSS.n58 a_1596_n2079# 0.02fF $ **FLOATING
C3996 VSS.n59 a_1596_n2079# 0.04fF $ **FLOATING
C3997 VSS.n60 a_1596_n2079# 4.86fF $ **FLOATING
C3998 VSS.n61 a_1596_n2079# 0.83fF $ **FLOATING
C3999 VSS.t149 a_1596_n2079# 0.01fF
C4000 VSS.t63 a_1596_n2079# 0.01fF
C4001 VSS.t106 a_1596_n2079# 0.01fF
C4002 VSS.t101 a_1596_n2079# 0.01fF
C4003 VSS.n62 a_1596_n2079# 0.04fF $ **FLOATING
C4004 VSS.n63 a_1596_n2079# 0.05fF $ **FLOATING
C4005 VSS.n64 a_1596_n2079# 0.06fF $ **FLOATING
C4006 VSS.n65 a_1596_n2079# 3.14fF $ **FLOATING
C4007 VSS.t47 a_1596_n2079# 0.00fF
C4008 VSS.t140 a_1596_n2079# 0.01fF
C4009 VSS.n66 a_1596_n2079# 0.09fF $ **FLOATING
C4010 VSS.t27 a_1596_n2079# 0.00fF
C4011 VSS.t127 a_1596_n2079# 0.01fF
C4012 VSS.n67 a_1596_n2079# 0.09fF $ **FLOATING
C4013 VSS.n68 a_1596_n2079# 7.02fF $ **FLOATING
C4014 VSS.t136 a_1596_n2079# 0.01fF
C4015 VSS.t44 a_1596_n2079# 0.01fF
C4016 VSS.t95 a_1596_n2079# 0.01fF
C4017 VSS.t8 a_1596_n2079# 0.01fF
C4018 VSS.n69 a_1596_n2079# 0.04fF $ **FLOATING
C4019 VSS.n70 a_1596_n2079# 0.05fF $ **FLOATING
C4020 VSS.n71 a_1596_n2079# 0.06fF $ **FLOATING
C4021 VSS.n72 a_1596_n2079# 0.05fF $ **FLOATING
C4022 VSS.n73 a_1596_n2079# 0.03fF $ **FLOATING
C4023 VSS.n74 a_1596_n2079# 0.24fF $ **FLOATING
C4024 VSS.n75 a_1596_n2079# 0.02fF $ **FLOATING
C4025 VSS.t7 a_1596_n2079# 0.00fF
C4026 VSS.t3 a_1596_n2079# 0.00fF
C4027 VSS.t130 a_1596_n2079# 0.00fF
C4028 VSS.n76 a_1596_n2079# 0.02fF $ **FLOATING
C4029 VSS.n77 a_1596_n2079# 0.04fF $ **FLOATING
C4030 VSS.n78 a_1596_n2079# 6.35fF $ **FLOATING
C4031 VSS.t56 a_1596_n2079# 0.00fF
C4032 VSS.t142 a_1596_n2079# 0.00fF
C4033 VSS.t150 a_1596_n2079# 0.00fF
C4034 VSS.n79 a_1596_n2079# 0.02fF $ **FLOATING
C4035 VSS.n80 a_1596_n2079# 0.04fF $ **FLOATING
C4036 VSS.n81 a_1596_n2079# 4.23fF $ **FLOATING
C4037 VSS.n82 a_1596_n2079# 1.28fF $ **FLOATING
C4038 VSS.n83 a_1596_n2079# 3.10fF $ **FLOATING
C4039 VSS.t28 a_1596_n2079# 0.00fF
C4040 VSS.t146 a_1596_n2079# 0.01fF
C4041 VSS.n84 a_1596_n2079# 0.09fF $ **FLOATING
C4042 VSS.t96 a_1596_n2079# 0.00fF
C4043 VSS.t38 a_1596_n2079# 0.01fF
C4044 VSS.n85 a_1596_n2079# 0.09fF $ **FLOATING
C4045 VSS.n86 a_1596_n2079# 6.97fF $ **FLOATING
C4046 VSS.t37 a_1596_n2079# 0.01fF
C4047 VSS.t143 a_1596_n2079# 0.01fF
C4048 VSS.t138 a_1596_n2079# 0.01fF
C4049 VSS.t148 a_1596_n2079# 0.01fF
C4050 VSS.n87 a_1596_n2079# 0.04fF $ **FLOATING
C4051 VSS.n88 a_1596_n2079# 0.05fF $ **FLOATING
C4052 VSS.n89 a_1596_n2079# 0.06fF $ **FLOATING
C4053 VSS.n90 a_1596_n2079# 0.25fF $ **FLOATING
C4054 VSS.n91 a_1596_n2079# 6.43fF $ **FLOATING
C4055 VSS.t120 a_1596_n2079# 0.00fF
C4056 VSS.t75 a_1596_n2079# 0.00fF
C4057 VSS.t23 a_1596_n2079# 0.00fF
C4058 VSS.n92 a_1596_n2079# 0.02fF $ **FLOATING
C4059 VSS.n93 a_1596_n2079# 0.04fF $ **FLOATING
C4060 VSS.n94 a_1596_n2079# 4.23fF $ **FLOATING
C4061 VSS.n95 a_1596_n2079# 1.28fF $ **FLOATING
C4062 VSS.n96 a_1596_n2079# 0.89fF $ **FLOATING
C4063 VSS.n97 a_1596_n2079# 4.53fF $ **FLOATING
C4064 VSS.n98 a_1596_n2079# 4.26fF $ **FLOATING
C4065 VSS.t68 a_1596_n2079# 0.00fF
C4066 VSS.t97 a_1596_n2079# 0.00fF
C4067 VSS.n99 a_1596_n2079# 0.02fF $ **FLOATING
C4068 VSS.t74 a_1596_n2079# 0.00fF
C4069 VSS.n100 a_1596_n2079# 0.04fF $ **FLOATING
C4070 VSS.t82 a_1596_n2079# 0.00fF
C4071 VSS.t93 a_1596_n2079# 0.01fF
C4072 VSS.n101 a_1596_n2079# 0.24fF $ **FLOATING
C4073 VSS.t1 a_1596_n2079# 0.00fF
C4074 VSS.t88 a_1596_n2079# 0.00fF
C4075 VSS.n102 a_1596_n2079# 0.02fF $ **FLOATING
C4076 VSS.t55 a_1596_n2079# 0.00fF
C4077 VSS.n103 a_1596_n2079# 0.04fF $ **FLOATING
C4078 VSS.n104 a_1596_n2079# 4.22fF $ **FLOATING
C4079 VSS.t144 a_1596_n2079# 0.00fF
C4080 VSS.t92 a_1596_n2079# 0.01fF
C4081 VSS.n105 a_1596_n2079# 0.11fF $ **FLOATING
C4082 VSS.t48 a_1596_n2079# 0.00fF
C4083 VSS.t102 a_1596_n2079# 0.01fF
C4084 VSS.n106 a_1596_n2079# 0.11fF $ **FLOATING
C4085 VSS.t104 a_1596_n2079# 0.01fF
C4086 VSS.t103 a_1596_n2079# 0.01fF
C4087 VSS.t117 a_1596_n2079# 0.01fF
C4088 VSS.n107 a_1596_n2079# 0.04fF $ **FLOATING
C4089 VSS.n108 a_1596_n2079# 0.05fF $ **FLOATING
C4090 VSS.t52 a_1596_n2079# 0.01fF
C4091 VSS.n109 a_1596_n2079# 0.06fF $ **FLOATING
C4092 VSS.t153 a_1596_n2079# 0.01fF
C4093 VSS.t10 a_1596_n2079# 0.01fF
C4094 VSS.t39 a_1596_n2079# 0.01fF
C4095 VSS.n110 a_1596_n2079# 0.04fF $ **FLOATING
C4096 VSS.n111 a_1596_n2079# 0.05fF $ **FLOATING
C4097 VSS.t105 a_1596_n2079# 0.01fF
C4098 VSS.n112 a_1596_n2079# 0.06fF $ **FLOATING
C4099 VSS.n113 a_1596_n2079# 3.64fF $ **FLOATING
C4100 VSS.n114 a_1596_n2079# 5.91fF $ **FLOATING
C4101 VSS.n115 a_1596_n2079# 4.88fF $ **FLOATING
C4102 VSS.n116 a_1596_n2079# 4.21fF $ **FLOATING
C4103 VSS.n117 a_1596_n2079# 1.76fF $ **FLOATING
C4104 VSS.n118 a_1596_n2079# 5.11fF $ **FLOATING
C4105 VSS.t91 a_1596_n2079# 0.00fF
C4106 VSS.t58 a_1596_n2079# 0.00fF
C4107 VSS.n119 a_1596_n2079# 0.02fF $ **FLOATING
C4108 VSS.t90 a_1596_n2079# 0.00fF
C4109 VSS.n120 a_1596_n2079# 0.04fF $ **FLOATING
C4110 VSS.n121 a_1596_n2079# 6.69fF $ **FLOATING
C4111 VSS.t15 a_1596_n2079# 0.00fF
C4112 VSS.t128 a_1596_n2079# 0.00fF
C4113 VSS.n122 a_1596_n2079# 0.02fF $ **FLOATING
C4114 VSS.t78 a_1596_n2079# 0.00fF
C4115 VSS.n123 a_1596_n2079# 0.04fF $ **FLOATING
C4116 VSS.n124 a_1596_n2079# 4.23fF $ **FLOATING
C4117 VSS.n125 a_1596_n2079# 1.28fF $ **FLOATING
C4118 VSS.t17 a_1596_n2079# 0.01fF
C4119 VSS.t129 a_1596_n2079# 0.01fF
C4120 VSS.t85 a_1596_n2079# 0.01fF
C4121 VSS.n126 a_1596_n2079# 0.04fF $ **FLOATING
C4122 VSS.n127 a_1596_n2079# 0.05fF $ **FLOATING
C4123 VSS.t0 a_1596_n2079# 0.01fF
C4124 VSS.n128 a_1596_n2079# 0.06fF $ **FLOATING
C4125 VSS.n129 a_1596_n2079# 0.03fF $ **FLOATING
C4126 VSS.n130 a_1596_n2079# 0.19fF $ **FLOATING
C4127 VSS.n131 a_1596_n2079# 0.90fF $ **FLOATING
C4128 VSS.n132 a_1596_n2079# 0.07fF $ **FLOATING
C4129 VSS.n133 a_1596_n2079# 1.85fF $ **FLOATING
C4130 VSS.t137 a_1596_n2079# 0.00fF
C4131 VSS.t31 a_1596_n2079# 0.01fF
C4132 VSS.n134 a_1596_n2079# 0.14fF $ **FLOATING
C4133 VSS.t141 a_1596_n2079# 0.01fF
C4134 VSS.t108 a_1596_n2079# 0.01fF
C4135 VSS.t112 a_1596_n2079# 0.01fF
C4136 VSS.n135 a_1596_n2079# 0.04fF $ **FLOATING
C4137 VSS.n136 a_1596_n2079# 0.05fF $ **FLOATING
C4138 VSS.t33 a_1596_n2079# 0.01fF
C4139 VSS.n137 a_1596_n2079# 0.06fF $ **FLOATING
C4140 VSS.t99 a_1596_n2079# 0.00fF
C4141 VSS.t84 a_1596_n2079# 0.01fF
C4142 VSS.n138 a_1596_n2079# 0.14fF $ **FLOATING
C4143 VSS.t30 a_1596_n2079# 0.01fF
C4144 VSS.t147 a_1596_n2079# 0.01fF
C4145 VSS.t126 a_1596_n2079# 0.01fF
C4146 VSS.n139 a_1596_n2079# 0.04fF $ **FLOATING
C4147 VSS.n140 a_1596_n2079# 0.05fF $ **FLOATING
C4148 VSS.t14 a_1596_n2079# 0.01fF
C4149 VSS.n141 a_1596_n2079# 0.06fF $ **FLOATING
C4150 VSS.t113 a_1596_n2079# 0.00fF
C4151 VSS.t133 a_1596_n2079# 0.00fF
C4152 VSS.n142 a_1596_n2079# 0.02fF $ **FLOATING
C4153 VSS.t125 a_1596_n2079# 0.00fF
C4154 VSS.n143 a_1596_n2079# 0.06fF $ **FLOATING
C4155 VSS.t24 a_1596_n2079# 0.01fF
C4156 VSS.t35 a_1596_n2079# 0.01fF
C4157 VSS.t83 a_1596_n2079# 0.01fF
C4158 VSS.n144 a_1596_n2079# 0.04fF $ **FLOATING
C4159 VSS.n145 a_1596_n2079# 0.05fF $ **FLOATING
C4160 VSS.t87 a_1596_n2079# 0.01fF
C4161 VSS.n146 a_1596_n2079# 0.14fF $ **FLOATING
C4162 VSS.n147 a_1596_n2079# 7.20fF $ **FLOATING
C4163 VSS.t111 a_1596_n2079# 0.00fF
C4164 VSS.t53 a_1596_n2079# 0.00fF
C4165 VSS.n148 a_1596_n2079# 0.02fF $ **FLOATING
C4166 VSS.t26 a_1596_n2079# 0.00fF
C4167 VSS.n149 a_1596_n2079# 0.04fF $ **FLOATING
C4168 VSS.n150 a_1596_n2079# 6.69fF $ **FLOATING
C4169 VSS.t40 a_1596_n2079# 0.00fF
C4170 VSS.t77 a_1596_n2079# 0.01fF
C4171 VSS.n151 a_1596_n2079# 0.11fF $ **FLOATING
C4172 VSS.t154 a_1596_n2079# 0.00fF
C4173 VSS.t59 a_1596_n2079# 0.01fF
C4174 VSS.n152 a_1596_n2079# 0.09fF $ **FLOATING
C4175 VSS.n153 a_1596_n2079# 6.96fF $ **FLOATING
C4176 VSS.n154 a_1596_n2079# 2.25fF $ **FLOATING
C4177 VSS.t60 a_1596_n2079# 0.01fF
C4178 VSS.t71 a_1596_n2079# 0.01fF
C4179 VSS.t20 a_1596_n2079# 0.01fF
C4180 VSS.n155 a_1596_n2079# 0.04fF $ **FLOATING
C4181 VSS.n156 a_1596_n2079# 0.05fF $ **FLOATING
C4182 VSS.t54 a_1596_n2079# 0.01fF
C4183 VSS.n157 a_1596_n2079# 0.06fF $ **FLOATING
C4184 VSS.n158 a_1596_n2079# 0.03fF $ **FLOATING
C4185 VSS.n159 a_1596_n2079# 0.19fF $ **FLOATING
C4186 VSS.n160 a_1596_n2079# 0.90fF $ **FLOATING
C4187 VSS.n161 a_1596_n2079# 1.28fF $ **FLOATING
C4188 VSS.t42 a_1596_n2079# 0.00fF
C4189 VSS.t131 a_1596_n2079# 0.00fF
C4190 VSS.n162 a_1596_n2079# 0.02fF $ **FLOATING
C4191 VSS.t18 a_1596_n2079# 0.00fF
C4192 VSS.n163 a_1596_n2079# 0.04fF $ **FLOATING
C4193 VSS.n164 a_1596_n2079# 4.22fF $ **FLOATING
C4194 VSS.t89 a_1596_n2079# 0.00fF
C4195 VSS.t115 a_1596_n2079# 0.00fF
C4196 VSS.n165 a_1596_n2079# 0.02fF $ **FLOATING
C4197 VSS.t2 a_1596_n2079# 0.00fF
C4198 VSS.n166 a_1596_n2079# 0.04fF $ **FLOATING
C4199 VSS.n167 a_1596_n2079# 6.68fF $ **FLOATING
C4200 VSS.t116 a_1596_n2079# 0.00fF
C4201 VSS.t32 a_1596_n2079# 0.01fF
C4202 VSS.n168 a_1596_n2079# 0.11fF $ **FLOATING
C4203 VSS.t13 a_1596_n2079# 0.00fF
C4204 VSS.t34 a_1596_n2079# 0.01fF
C4205 VSS.n169 a_1596_n2079# 0.11fF $ **FLOATING
C4206 VSS.n170 a_1596_n2079# 5.11fF $ **FLOATING
C4207 VSS.n171 a_1596_n2079# 1.28fF $ **FLOATING
C4208 B[0].t13 a_1596_n2079# 0.04fF
C4209 B[0].t8 a_1596_n2079# 0.06fF
C4210 B[0].n0 a_1596_n2079# 0.07fF $ **FLOATING
C4211 B[0].t3 a_1596_n2079# 0.12fF
C4212 B[0].t6 a_1596_n2079# 0.12fF
C4213 B[0].t9 a_1596_n2079# 0.04fF
C4214 B[0].t12 a_1596_n2079# 0.08fF
C4215 B[0].t5 a_1596_n2079# 0.11fF
C4216 B[0].n1 a_1596_n2079# 0.14fF $ **FLOATING
C4217 B[0].t10 a_1596_n2079# 0.13fF
C4218 B[0].n2 a_1596_n2079# 0.10fF $ **FLOATING
C4219 B[0].t14 a_1596_n2079# 0.04fF
C4220 B[0].t4 a_1596_n2079# 0.06fF
C4221 B[0].n3 a_1596_n2079# 0.05fF $ **FLOATING
C4222 B[0].n4 a_1596_n2079# 0.03fF $ **FLOATING
C4223 B[0].t1 a_1596_n2079# 0.04fF
C4224 B[0].t11 a_1596_n2079# 0.16fF
C4225 B[0].n5 a_1596_n2079# 0.33fF $ **FLOATING
C4226 B[0].n6 a_1596_n2079# 0.38fF $ **FLOATING
C4227 B[0].n7 a_1596_n2079# 0.38fF $ **FLOATING
C4228 B[0].t7 a_1596_n2079# 0.04fF
C4229 B[0].t2 a_1596_n2079# 0.06fF
C4230 B[0].n8 a_1596_n2079# 0.07fF $ **FLOATING
C4231 B[0].t15 a_1596_n2079# 0.12fF
C4232 B[0].t0 a_1596_n2079# 0.13fF
C4233 B[0].n9 a_1596_n2079# 1.84fF $ **FLOATING
C4234 a_19657_n3503.t1 a_1596_n2079# 0.01fF
C4235 a_19657_n3503.t0 a_1596_n2079# 0.01fF
C4236 a_19657_n3503.t2 a_1596_n2079# 0.01fF
C4237 a_19657_n3503.n0 a_1596_n2079# 0.20fF $ **FLOATING
C4238 a_19657_n3503.t12 a_1596_n2079# 0.03fF
C4239 a_19657_n3503.t8 a_1596_n2079# 0.05fF
C4240 a_19657_n3503.n1 a_1596_n2079# 0.06fF $ **FLOATING
C4241 a_19657_n3503.t13 a_1596_n2079# 0.10fF
C4242 a_19657_n3503.t9 a_1596_n2079# 0.10fF
C4243 a_19657_n3503.t6 a_1596_n2079# 0.07fF
C4244 a_19657_n3503.t10 a_1596_n2079# 0.07fF
C4245 a_19657_n3503.t11 a_1596_n2079# 0.09fF
C4246 a_19657_n3503.n2 a_1596_n2079# 0.09fF $ **FLOATING
C4247 a_19657_n3503.n3 a_1596_n2079# 0.09fF $ **FLOATING
C4248 a_19657_n3503.t5 a_1596_n2079# 0.08fF
C4249 a_19657_n3503.t19 a_1596_n2079# 0.05fF
C4250 a_19657_n3503.n4 a_1596_n2079# 0.08fF $ **FLOATING
C4251 a_19657_n3503.t4 a_1596_n2079# 0.06fF
C4252 a_19657_n3503.t15 a_1596_n2079# 0.04fF
C4253 a_19657_n3503.t7 a_1596_n2079# 0.14fF
C4254 a_19657_n3503.n5 a_1596_n2079# 0.28fF $ **FLOATING
C4255 a_19657_n3503.n6 a_1596_n2079# 0.24fF $ **FLOATING
C4256 a_19657_n3503.n7 a_1596_n2079# 2.62fF $ **FLOATING
C4257 a_19657_n3503.t17 a_1596_n2079# 0.03fF
C4258 a_19657_n3503.t18 a_1596_n2079# 0.05fF
C4259 a_19657_n3503.n8 a_1596_n2079# 0.06fF $ **FLOATING
C4260 a_19657_n3503.t14 a_1596_n2079# 0.10fF
C4261 a_19657_n3503.t16 a_1596_n2079# 0.11fF
C4262 a_19657_n3503.n9 a_1596_n2079# 4.26fF $ **FLOATING
C4263 a_19657_n3503.n10 a_1596_n2079# 2.36fF $ **FLOATING
C4264 a_19657_n3503.n11 a_1596_n2079# 0.10fF $ **FLOATING
C4265 a_19657_n3503.t3 a_1596_n2079# 0.01fF
C4266 B[3].t15 a_1596_n2079# 0.04fF
C4267 B[3].t8 a_1596_n2079# 0.06fF
C4268 B[3].n0 a_1596_n2079# 0.07fF $ **FLOATING
C4269 B[3].t1 a_1596_n2079# 0.12fF
C4270 B[3].t3 a_1596_n2079# 0.12fF
C4271 B[3].t9 a_1596_n2079# 0.04fF
C4272 B[3].t7 a_1596_n2079# 0.08fF
C4273 B[3].t2 a_1596_n2079# 0.11fF
C4274 B[3].n1 a_1596_n2079# 0.14fF $ **FLOATING
C4275 B[3].t14 a_1596_n2079# 0.13fF
C4276 B[3].n2 a_1596_n2079# 0.10fF $ **FLOATING
C4277 B[3].t0 a_1596_n2079# 0.04fF
C4278 B[3].t6 a_1596_n2079# 0.06fF
C4279 B[3].n3 a_1596_n2079# 0.05fF $ **FLOATING
C4280 B[3].n4 a_1596_n2079# 0.03fF $ **FLOATING
C4281 B[3].t13 a_1596_n2079# 0.04fF
C4282 B[3].t5 a_1596_n2079# 0.16fF
C4283 B[3].n5 a_1596_n2079# 0.33fF $ **FLOATING
C4284 B[3].n6 a_1596_n2079# 0.38fF $ **FLOATING
C4285 B[3].n7 a_1596_n2079# 0.38fF $ **FLOATING
C4286 B[3].t11 a_1596_n2079# 0.04fF
C4287 B[3].t4 a_1596_n2079# 0.06fF
C4288 B[3].n8 a_1596_n2079# 0.07fF $ **FLOATING
C4289 B[3].t10 a_1596_n2079# 0.12fF
C4290 B[3].t12 a_1596_n2079# 0.13fF
C4291 B[3].n9 a_1596_n2079# 1.82fF $ **FLOATING
C4292 VDD.t213 a_1596_n2079# 0.01fF
C4293 VDD.t126 a_1596_n2079# 0.01fF
C4294 VDD.n0 a_1596_n2079# 0.05fF $ **FLOATING
C4295 VDD.t37 a_1596_n2079# 0.01fF
C4296 VDD.t147 a_1596_n2079# 0.01fF
C4297 VDD.t295 a_1596_n2079# 0.01fF
C4298 VDD.n1 a_1596_n2079# 0.05fF $ **FLOATING
C4299 VDD.n2 a_1596_n2079# 0.10fF $ **FLOATING
C4300 VDD.n3 a_1596_n2079# 0.06fF $ **FLOATING
C4301 VDD.t115 a_1596_n2079# 0.01fF
C4302 VDD.t117 a_1596_n2079# 0.01fF
C4303 VDD.n4 a_1596_n2079# 0.06fF $ **FLOATING
C4304 VDD.t116 a_1596_n2079# 0.01fF
C4305 VDD.t66 a_1596_n2079# 0.01fF
C4306 VDD.n5 a_1596_n2079# 0.05fF $ **FLOATING
C4307 VDD.n6 a_1596_n2079# 0.03fF $ **FLOATING
C4308 VDD.n7 a_1596_n2079# 0.20fF $ **FLOATING
C4309 VDD.t395 a_1596_n2079# 0.01fF
C4310 VDD.t394 a_1596_n2079# 0.01fF
C4311 VDD.n8 a_1596_n2079# 0.11fF $ **FLOATING
C4312 VDD.t393 a_1596_n2079# 0.01fF
C4313 VDD.t19 a_1596_n2079# 0.01fF
C4314 VDD.t21 a_1596_n2079# 0.01fF
C4315 VDD.t20 a_1596_n2079# 0.01fF
C4316 VDD.n9 a_1596_n2079# 0.07fF $ **FLOATING
C4317 VDD.n10 a_1596_n2079# 0.10fF $ **FLOATING
C4318 VDD.n11 a_1596_n2079# 0.13fF $ **FLOATING
C4319 VDD.n12 a_1596_n2079# 0.04fF $ **FLOATING
C4320 VDD.t478 a_1596_n2079# 0.01fF
C4321 VDD.t476 a_1596_n2079# 0.01fF
C4322 VDD.n13 a_1596_n2079# 0.11fF $ **FLOATING
C4323 VDD.t477 a_1596_n2079# 0.01fF
C4324 VDD.t453 a_1596_n2079# 0.01fF
C4325 VDD.t452 a_1596_n2079# 0.01fF
C4326 VDD.t451 a_1596_n2079# 0.01fF
C4327 VDD.n14 a_1596_n2079# 0.07fF $ **FLOATING
C4328 VDD.n15 a_1596_n2079# 0.10fF $ **FLOATING
C4329 VDD.n16 a_1596_n2079# 0.13fF $ **FLOATING
C4330 VDD.n17 a_1596_n2079# 0.04fF $ **FLOATING
C4331 VDD.t460 a_1596_n2079# 0.01fF
C4332 VDD.t143 a_1596_n2079# 0.01fF
C4333 VDD.n18 a_1596_n2079# 0.05fF $ **FLOATING
C4334 VDD.t108 a_1596_n2079# 0.01fF
C4335 VDD.t110 a_1596_n2079# 0.01fF
C4336 VDD.t33 a_1596_n2079# 0.01fF
C4337 VDD.n19 a_1596_n2079# 0.05fF $ **FLOATING
C4338 VDD.n20 a_1596_n2079# 0.10fF $ **FLOATING
C4339 VDD.n21 a_1596_n2079# 0.06fF $ **FLOATING
C4340 VDD.t157 a_1596_n2079# 0.01fF
C4341 VDD.t156 a_1596_n2079# 0.01fF
C4342 VDD.n22 a_1596_n2079# 0.06fF $ **FLOATING
C4343 VDD.t158 a_1596_n2079# 0.01fF
C4344 VDD.t144 a_1596_n2079# 0.01fF
C4345 VDD.n23 a_1596_n2079# 0.05fF $ **FLOATING
C4346 VDD.n24 a_1596_n2079# 0.03fF $ **FLOATING
C4347 VDD.n25 a_1596_n2079# 2.25fF $ **FLOATING
C4348 VDD.t214 a_1596_n2079# 0.01fF
C4349 VDD.t385 a_1596_n2079# 0.01fF
C4350 VDD.n26 a_1596_n2079# 0.05fF $ **FLOATING
C4351 VDD.t49 a_1596_n2079# 0.01fF
C4352 VDD.t430 a_1596_n2079# 0.01fF
C4353 VDD.t349 a_1596_n2079# 0.01fF
C4354 VDD.n27 a_1596_n2079# 0.05fF $ **FLOATING
C4355 VDD.n28 a_1596_n2079# 0.10fF $ **FLOATING
C4356 VDD.n29 a_1596_n2079# 0.06fF $ **FLOATING
C4357 VDD.t381 a_1596_n2079# 0.01fF
C4358 VDD.t383 a_1596_n2079# 0.01fF
C4359 VDD.n30 a_1596_n2079# 0.06fF $ **FLOATING
C4360 VDD.t382 a_1596_n2079# 0.01fF
C4361 VDD.t68 a_1596_n2079# 0.01fF
C4362 VDD.n31 a_1596_n2079# 0.05fF $ **FLOATING
C4363 VDD.n32 a_1596_n2079# 0.03fF $ **FLOATING
C4364 VDD.n33 a_1596_n2079# 0.20fF $ **FLOATING
C4365 VDD.n34 a_1596_n2079# 2.88fF $ **FLOATING
C4366 VDD.t125 a_1596_n2079# 0.01fF
C4367 VDD.t411 a_1596_n2079# 0.01fF
C4368 VDD.n35 a_1596_n2079# 0.10fF $ **FLOATING
C4369 VDD.t127 a_1596_n2079# 0.01fF
C4370 VDD.t212 a_1596_n2079# 0.01fF
C4371 VDD.n36 a_1596_n2079# 0.20fF $ **FLOATING
C4372 VDD.t67 a_1596_n2079# 0.01fF
C4373 VDD.t124 a_1596_n2079# 0.01fF
C4374 VDD.n37 a_1596_n2079# 0.08fF $ **FLOATING
C4375 VDD.n38 a_1596_n2079# 0.06fF $ **FLOATING
C4376 VDD.n39 a_1596_n2079# 0.03fF $ **FLOATING
C4377 VDD.t146 a_1596_n2079# 0.01fF
C4378 VDD.t109 a_1596_n2079# 0.01fF
C4379 VDD.n40 a_1596_n2079# 0.10fF $ **FLOATING
C4380 VDD.t36 a_1596_n2079# 0.01fF
C4381 VDD.t32 a_1596_n2079# 0.01fF
C4382 VDD.n41 a_1596_n2079# 0.20fF $ **FLOATING
C4383 VDD.t35 a_1596_n2079# 0.01fF
C4384 VDD.t34 a_1596_n2079# 0.01fF
C4385 VDD.n42 a_1596_n2079# 0.08fF $ **FLOATING
C4386 VDD.n43 a_1596_n2079# 0.06fF $ **FLOATING
C4387 VDD.n44 a_1596_n2079# 0.03fF $ **FLOATING
C4388 VDD.n45 a_1596_n2079# 0.04fF $ **FLOATING
C4389 VDD.n46 a_1596_n2079# 2.28fF $ **FLOATING
C4390 VDD.t486 a_1596_n2079# 0.01fF
C4391 VDD.t485 a_1596_n2079# 0.01fF
C4392 VDD.n47 a_1596_n2079# 0.10fF $ **FLOATING
C4393 VDD.t487 a_1596_n2079# 0.01fF
C4394 VDD.t482 a_1596_n2079# 0.01fF
C4395 VDD.n48 a_1596_n2079# 0.20fF $ **FLOATING
C4396 VDD.t484 a_1596_n2079# 0.01fF
C4397 VDD.t483 a_1596_n2079# 0.01fF
C4398 VDD.n49 a_1596_n2079# 0.08fF $ **FLOATING
C4399 VDD.n50 a_1596_n2079# 0.06fF $ **FLOATING
C4400 VDD.n51 a_1596_n2079# 0.03fF $ **FLOATING
C4401 VDD.t350 a_1596_n2079# 0.01fF
C4402 VDD.t17 a_1596_n2079# 0.01fF
C4403 VDD.n52 a_1596_n2079# 0.10fF $ **FLOATING
C4404 VDD.t142 a_1596_n2079# 0.01fF
C4405 VDD.t48 a_1596_n2079# 0.01fF
C4406 VDD.n53 a_1596_n2079# 0.20fF $ **FLOATING
C4407 VDD.t16 a_1596_n2079# 0.01fF
C4408 VDD.t431 a_1596_n2079# 0.01fF
C4409 VDD.n54 a_1596_n2079# 0.08fF $ **FLOATING
C4410 VDD.n55 a_1596_n2079# 0.06fF $ **FLOATING
C4411 VDD.n56 a_1596_n2079# 0.03fF $ **FLOATING
C4412 VDD.n57 a_1596_n2079# 0.04fF $ **FLOATING
C4413 VDD.n58 a_1596_n2079# 2.87fF $ **FLOATING
C4414 VDD.t481 a_1596_n2079# 0.01fF
C4415 VDD.t480 a_1596_n2079# 0.01fF
C4416 VDD.n59 a_1596_n2079# 0.05fF $ **FLOATING
C4417 VDD.t470 a_1596_n2079# 0.01fF
C4418 VDD.t249 a_1596_n2079# 0.01fF
C4419 VDD.t492 a_1596_n2079# 0.01fF
C4420 VDD.n60 a_1596_n2079# 0.05fF $ **FLOATING
C4421 VDD.n61 a_1596_n2079# 0.10fF $ **FLOATING
C4422 VDD.n62 a_1596_n2079# 0.06fF $ **FLOATING
C4423 VDD.t325 a_1596_n2079# 0.01fF
C4424 VDD.t323 a_1596_n2079# 0.01fF
C4425 VDD.n63 a_1596_n2079# 0.06fF $ **FLOATING
C4426 VDD.t324 a_1596_n2079# 0.01fF
C4427 VDD.t178 a_1596_n2079# 0.01fF
C4428 VDD.n64 a_1596_n2079# 0.05fF $ **FLOATING
C4429 VDD.n65 a_1596_n2079# 0.03fF $ **FLOATING
C4430 VDD.n66 a_1596_n2079# 0.20fF $ **FLOATING
C4431 VDD.t408 a_1596_n2079# 0.01fF
C4432 VDD.t410 a_1596_n2079# 0.01fF
C4433 VDD.n67 a_1596_n2079# 0.11fF $ **FLOATING
C4434 VDD.t409 a_1596_n2079# 0.01fF
C4435 VDD.t83 a_1596_n2079# 0.01fF
C4436 VDD.t82 a_1596_n2079# 0.01fF
C4437 VDD.t84 a_1596_n2079# 0.01fF
C4438 VDD.n68 a_1596_n2079# 0.07fF $ **FLOATING
C4439 VDD.n69 a_1596_n2079# 0.10fF $ **FLOATING
C4440 VDD.n70 a_1596_n2079# 0.13fF $ **FLOATING
C4441 VDD.n71 a_1596_n2079# 0.04fF $ **FLOATING
C4442 VDD.t96 a_1596_n2079# 0.01fF
C4443 VDD.t95 a_1596_n2079# 0.01fF
C4444 VDD.n72 a_1596_n2079# 0.11fF $ **FLOATING
C4445 VDD.t94 a_1596_n2079# 0.01fF
C4446 VDD.t259 a_1596_n2079# 0.01fF
C4447 VDD.t261 a_1596_n2079# 0.01fF
C4448 VDD.t260 a_1596_n2079# 0.01fF
C4449 VDD.n73 a_1596_n2079# 0.07fF $ **FLOATING
C4450 VDD.n74 a_1596_n2079# 0.10fF $ **FLOATING
C4451 VDD.n75 a_1596_n2079# 0.13fF $ **FLOATING
C4452 VDD.n76 a_1596_n2079# 0.04fF $ **FLOATING
C4453 VDD.t346 a_1596_n2079# 0.01fF
C4454 VDD.t345 a_1596_n2079# 0.01fF
C4455 VDD.n77 a_1596_n2079# 0.05fF $ **FLOATING
C4456 VDD.t148 a_1596_n2079# 0.01fF
C4457 VDD.t266 a_1596_n2079# 0.01fF
C4458 VDD.t262 a_1596_n2079# 0.01fF
C4459 VDD.n78 a_1596_n2079# 0.05fF $ **FLOATING
C4460 VDD.n79 a_1596_n2079# 0.10fF $ **FLOATING
C4461 VDD.n80 a_1596_n2079# 0.06fF $ **FLOATING
C4462 VDD.t122 a_1596_n2079# 0.01fF
C4463 VDD.t121 a_1596_n2079# 0.01fF
C4464 VDD.n81 a_1596_n2079# 0.06fF $ **FLOATING
C4465 VDD.t123 a_1596_n2079# 0.01fF
C4466 VDD.t443 a_1596_n2079# 0.01fF
C4467 VDD.n82 a_1596_n2079# 0.05fF $ **FLOATING
C4468 VDD.n83 a_1596_n2079# 0.03fF $ **FLOATING
C4469 VDD.n84 a_1596_n2079# 2.25fF $ **FLOATING
C4470 VDD.t28 a_1596_n2079# 0.01fF
C4471 VDD.t176 a_1596_n2079# 0.01fF
C4472 VDD.n85 a_1596_n2079# 0.05fF $ **FLOATING
C4473 VDD.t471 a_1596_n2079# 0.01fF
C4474 VDD.t472 a_1596_n2079# 0.01fF
C4475 VDD.t448 a_1596_n2079# 0.01fF
C4476 VDD.n86 a_1596_n2079# 0.05fF $ **FLOATING
C4477 VDD.n87 a_1596_n2079# 0.10fF $ **FLOATING
C4478 VDD.n88 a_1596_n2079# 0.06fF $ **FLOATING
C4479 VDD.t378 a_1596_n2079# 0.01fF
C4480 VDD.t377 a_1596_n2079# 0.01fF
C4481 VDD.n89 a_1596_n2079# 0.06fF $ **FLOATING
C4482 VDD.t379 a_1596_n2079# 0.01fF
C4483 VDD.t194 a_1596_n2079# 0.01fF
C4484 VDD.n90 a_1596_n2079# 0.05fF $ **FLOATING
C4485 VDD.n91 a_1596_n2079# 0.03fF $ **FLOATING
C4486 VDD.n92 a_1596_n2079# 0.20fF $ **FLOATING
C4487 VDD.n93 a_1596_n2079# 2.88fF $ **FLOATING
C4488 VDD.t177 a_1596_n2079# 0.01fF
C4489 VDD.t193 a_1596_n2079# 0.01fF
C4490 VDD.n94 a_1596_n2079# 0.10fF $ **FLOATING
C4491 VDD.t27 a_1596_n2079# 0.01fF
C4492 VDD.t479 a_1596_n2079# 0.01fF
C4493 VDD.n95 a_1596_n2079# 0.20fF $ **FLOATING
C4494 VDD.t425 a_1596_n2079# 0.01fF
C4495 VDD.t192 a_1596_n2079# 0.01fF
C4496 VDD.n96 a_1596_n2079# 0.08fF $ **FLOATING
C4497 VDD.n97 a_1596_n2079# 0.06fF $ **FLOATING
C4498 VDD.n98 a_1596_n2079# 0.03fF $ **FLOATING
C4499 VDD.t455 a_1596_n2079# 0.01fF
C4500 VDD.t265 a_1596_n2079# 0.01fF
C4501 VDD.n99 a_1596_n2079# 0.10fF $ **FLOATING
C4502 VDD.t248 a_1596_n2079# 0.01fF
C4503 VDD.t456 a_1596_n2079# 0.01fF
C4504 VDD.n100 a_1596_n2079# 0.20fF $ **FLOATING
C4505 VDD.t491 a_1596_n2079# 0.01fF
C4506 VDD.t138 a_1596_n2079# 0.01fF
C4507 VDD.n101 a_1596_n2079# 0.08fF $ **FLOATING
C4508 VDD.n102 a_1596_n2079# 0.06fF $ **FLOATING
C4509 VDD.n103 a_1596_n2079# 0.03fF $ **FLOATING
C4510 VDD.n104 a_1596_n2079# 0.04fF $ **FLOATING
C4511 VDD.n105 a_1596_n2079# 2.28fF $ **FLOATING
C4512 VDD.t221 a_1596_n2079# 0.01fF
C4513 VDD.t220 a_1596_n2079# 0.01fF
C4514 VDD.n106 a_1596_n2079# 0.10fF $ **FLOATING
C4515 VDD.t216 a_1596_n2079# 0.01fF
C4516 VDD.t219 a_1596_n2079# 0.01fF
C4517 VDD.n107 a_1596_n2079# 0.20fF $ **FLOATING
C4518 VDD.t217 a_1596_n2079# 0.01fF
C4519 VDD.t218 a_1596_n2079# 0.01fF
C4520 VDD.n108 a_1596_n2079# 0.08fF $ **FLOATING
C4521 VDD.n109 a_1596_n2079# 0.06fF $ **FLOATING
C4522 VDD.n110 a_1596_n2079# 0.03fF $ **FLOATING
C4523 VDD.t446 a_1596_n2079# 0.01fF
C4524 VDD.t444 a_1596_n2079# 0.01fF
C4525 VDD.n111 a_1596_n2079# 0.10fF $ **FLOATING
C4526 VDD.t447 a_1596_n2079# 0.01fF
C4527 VDD.t145 a_1596_n2079# 0.01fF
C4528 VDD.n112 a_1596_n2079# 0.20fF $ **FLOATING
C4529 VDD.t445 a_1596_n2079# 0.01fF
C4530 VDD.t449 a_1596_n2079# 0.01fF
C4531 VDD.n113 a_1596_n2079# 0.08fF $ **FLOATING
C4532 VDD.n114 a_1596_n2079# 0.06fF $ **FLOATING
C4533 VDD.n115 a_1596_n2079# 0.03fF $ **FLOATING
C4534 VDD.n116 a_1596_n2079# 0.04fF $ **FLOATING
C4535 VDD.n117 a_1596_n2079# 3.19fF $ **FLOATING
C4536 VDD.n118 a_1596_n2079# 3.15fF $ **FLOATING
C4537 VDD.n119 a_1596_n2079# 3.21fF $ **FLOATING
C4538 VDD.n120 a_1596_n2079# 4.34fF $ **FLOATING
C4539 VDD.n121 a_1596_n2079# 3.82fF $ **FLOATING
C4540 VDD.n122 a_1596_n2079# 1.48fF $ **FLOATING
C4541 VDD.n123 a_1596_n2079# 3.35fF $ **FLOATING
C4542 VDD.n124 a_1596_n2079# 3.69fF $ **FLOATING
C4543 VDD.t222 a_1596_n2079# 0.01fF
C4544 VDD.t269 a_1596_n2079# 0.01fF
C4545 VDD.n125 a_1596_n2079# 0.05fF $ **FLOATING
C4546 VDD.t436 a_1596_n2079# 0.01fF
C4547 VDD.t232 a_1596_n2079# 0.01fF
C4548 VDD.t235 a_1596_n2079# 0.01fF
C4549 VDD.n126 a_1596_n2079# 0.05fF $ **FLOATING
C4550 VDD.n127 a_1596_n2079# 0.10fF $ **FLOATING
C4551 VDD.n128 a_1596_n2079# 0.06fF $ **FLOATING
C4552 VDD.t173 a_1596_n2079# 0.01fF
C4553 VDD.t175 a_1596_n2079# 0.01fF
C4554 VDD.n129 a_1596_n2079# 0.06fF $ **FLOATING
C4555 VDD.t174 a_1596_n2079# 0.01fF
C4556 VDD.t338 a_1596_n2079# 0.01fF
C4557 VDD.n130 a_1596_n2079# 0.05fF $ **FLOATING
C4558 VDD.n131 a_1596_n2079# 0.03fF $ **FLOATING
C4559 VDD.n132 a_1596_n2079# 2.25fF $ **FLOATING
C4560 VDD.t344 a_1596_n2079# 0.01fF
C4561 VDD.t164 a_1596_n2079# 0.01fF
C4562 VDD.n133 a_1596_n2079# 0.05fF $ **FLOATING
C4563 VDD.t44 a_1596_n2079# 0.01fF
C4564 VDD.t296 a_1596_n2079# 0.01fF
C4565 VDD.t112 a_1596_n2079# 0.01fF
C4566 VDD.n134 a_1596_n2079# 0.05fF $ **FLOATING
C4567 VDD.n135 a_1596_n2079# 0.10fF $ **FLOATING
C4568 VDD.n136 a_1596_n2079# 0.06fF $ **FLOATING
C4569 VDD.t149 a_1596_n2079# 0.01fF
C4570 VDD.t151 a_1596_n2079# 0.01fF
C4571 VDD.n137 a_1596_n2079# 0.06fF $ **FLOATING
C4572 VDD.t150 a_1596_n2079# 0.01fF
C4573 VDD.t104 a_1596_n2079# 0.01fF
C4574 VDD.n138 a_1596_n2079# 0.05fF $ **FLOATING
C4575 VDD.n139 a_1596_n2079# 0.03fF $ **FLOATING
C4576 VDD.n140 a_1596_n2079# 0.20fF $ **FLOATING
C4577 VDD.n141 a_1596_n2079# 2.88fF $ **FLOATING
C4578 VDD.t384 a_1596_n2079# 0.01fF
C4579 VDD.t114 a_1596_n2079# 0.01fF
C4580 VDD.n142 a_1596_n2079# 0.10fF $ **FLOATING
C4581 VDD.t303 a_1596_n2079# 0.01fF
C4582 VDD.t254 a_1596_n2079# 0.01fF
C4583 VDD.n143 a_1596_n2079# 0.20fF $ **FLOATING
C4584 VDD.t134 a_1596_n2079# 0.01fF
C4585 VDD.t195 a_1596_n2079# 0.01fF
C4586 VDD.n144 a_1596_n2079# 0.08fF $ **FLOATING
C4587 VDD.n145 a_1596_n2079# 0.06fF $ **FLOATING
C4588 VDD.n146 a_1596_n2079# 0.03fF $ **FLOATING
C4589 VDD.t374 a_1596_n2079# 0.01fF
C4590 VDD.t251 a_1596_n2079# 0.01fF
C4591 VDD.n147 a_1596_n2079# 0.10fF $ **FLOATING
C4592 VDD.t234 a_1596_n2079# 0.01fF
C4593 VDD.t252 a_1596_n2079# 0.01fF
C4594 VDD.n148 a_1596_n2079# 0.20fF $ **FLOATING
C4595 VDD.t435 a_1596_n2079# 0.01fF
C4596 VDD.t233 a_1596_n2079# 0.01fF
C4597 VDD.n149 a_1596_n2079# 0.08fF $ **FLOATING
C4598 VDD.n150 a_1596_n2079# 0.06fF $ **FLOATING
C4599 VDD.n151 a_1596_n2079# 0.03fF $ **FLOATING
C4600 VDD.n152 a_1596_n2079# 0.04fF $ **FLOATING
C4601 VDD.n153 a_1596_n2079# 2.28fF $ **FLOATING
C4602 VDD.t99 a_1596_n2079# 0.01fF
C4603 VDD.t64 a_1596_n2079# 0.01fF
C4604 VDD.n154 a_1596_n2079# 0.10fF $ **FLOATING
C4605 VDD.t97 a_1596_n2079# 0.01fF
C4606 VDD.t65 a_1596_n2079# 0.01fF
C4607 VDD.n155 a_1596_n2079# 0.20fF $ **FLOATING
C4608 VDD.t473 a_1596_n2079# 0.01fF
C4609 VDD.t98 a_1596_n2079# 0.01fF
C4610 VDD.n156 a_1596_n2079# 0.08fF $ **FLOATING
C4611 VDD.n157 a_1596_n2079# 0.06fF $ **FLOATING
C4612 VDD.n158 a_1596_n2079# 0.03fF $ **FLOATING
C4613 VDD.t271 a_1596_n2079# 0.01fF
C4614 VDD.t111 a_1596_n2079# 0.01fF
C4615 VDD.n159 a_1596_n2079# 0.10fF $ **FLOATING
C4616 VDD.t43 a_1596_n2079# 0.01fF
C4617 VDD.t113 a_1596_n2079# 0.01fF
C4618 VDD.n160 a_1596_n2079# 0.20fF $ **FLOATING
C4619 VDD.t223 a_1596_n2079# 0.01fF
C4620 VDD.t270 a_1596_n2079# 0.01fF
C4621 VDD.n161 a_1596_n2079# 0.08fF $ **FLOATING
C4622 VDD.n162 a_1596_n2079# 0.06fF $ **FLOATING
C4623 VDD.n163 a_1596_n2079# 0.03fF $ **FLOATING
C4624 VDD.n164 a_1596_n2079# 0.04fF $ **FLOATING
C4625 VDD.n165 a_1596_n2079# 2.87fF $ **FLOATING
C4626 VDD.t30 a_1596_n2079# 0.01fF
C4627 VDD.t29 a_1596_n2079# 0.01fF
C4628 VDD.n166 a_1596_n2079# 0.10fF $ **FLOATING
C4629 VDD.t432 a_1596_n2079# 0.01fF
C4630 VDD.t31 a_1596_n2079# 0.01fF
C4631 VDD.n167 a_1596_n2079# 0.20fF $ **FLOATING
C4632 VDD.t38 a_1596_n2079# 0.01fF
C4633 VDD.t39 a_1596_n2079# 0.01fF
C4634 VDD.n168 a_1596_n2079# 0.08fF $ **FLOATING
C4635 VDD.n169 a_1596_n2079# 0.06fF $ **FLOATING
C4636 VDD.n170 a_1596_n2079# 0.03fF $ **FLOATING
C4637 VDD.t321 a_1596_n2079# 0.01fF
C4638 VDD.t336 a_1596_n2079# 0.01fF
C4639 VDD.n171 a_1596_n2079# 0.10fF $ **FLOATING
C4640 VDD.t363 a_1596_n2079# 0.01fF
C4641 VDD.t354 a_1596_n2079# 0.01fF
C4642 VDD.n172 a_1596_n2079# 0.20fF $ **FLOATING
C4643 VDD.t362 a_1596_n2079# 0.01fF
C4644 VDD.t283 a_1596_n2079# 0.01fF
C4645 VDD.n173 a_1596_n2079# 0.08fF $ **FLOATING
C4646 VDD.n174 a_1596_n2079# 0.06fF $ **FLOATING
C4647 VDD.n175 a_1596_n2079# 0.03fF $ **FLOATING
C4648 VDD.n176 a_1596_n2079# 0.04fF $ **FLOATING
C4649 VDD.n177 a_1596_n2079# 2.86fF $ **FLOATING
C4650 VDD.t488 a_1596_n2079# 0.01fF
C4651 VDD.t490 a_1596_n2079# 0.01fF
C4652 VDD.n178 a_1596_n2079# 0.06fF $ **FLOATING
C4653 VDD.t489 a_1596_n2079# 0.01fF
C4654 VDD.t253 a_1596_n2079# 0.01fF
C4655 VDD.n179 a_1596_n2079# 0.05fF $ **FLOATING
C4656 VDD.n180 a_1596_n2079# 0.03fF $ **FLOATING
C4657 VDD.t22 a_1596_n2079# 0.01fF
C4658 VDD.t60 a_1596_n2079# 0.01fF
C4659 VDD.n181 a_1596_n2079# 0.05fF $ **FLOATING
C4660 VDD.t454 a_1596_n2079# 0.01fF
C4661 VDD.t305 a_1596_n2079# 0.01fF
C4662 VDD.t348 a_1596_n2079# 0.01fF
C4663 VDD.n182 a_1596_n2079# 0.05fF $ **FLOATING
C4664 VDD.n183 a_1596_n2079# 0.10fF $ **FLOATING
C4665 VDD.n184 a_1596_n2079# 0.06fF $ **FLOATING
C4666 VDD.t364 a_1596_n2079# 0.01fF
C4667 VDD.t257 a_1596_n2079# 0.01fF
C4668 VDD.n185 a_1596_n2079# 0.05fF $ **FLOATING
C4669 VDD.t450 a_1596_n2079# 0.01fF
C4670 VDD.t201 a_1596_n2079# 0.01fF
C4671 VDD.t267 a_1596_n2079# 0.01fF
C4672 VDD.n186 a_1596_n2079# 0.05fF $ **FLOATING
C4673 VDD.n187 a_1596_n2079# 0.10fF $ **FLOATING
C4674 VDD.n188 a_1596_n2079# 0.06fF $ **FLOATING
C4675 VDD.t79 a_1596_n2079# 0.01fF
C4676 VDD.t81 a_1596_n2079# 0.01fF
C4677 VDD.n189 a_1596_n2079# 0.06fF $ **FLOATING
C4678 VDD.t80 a_1596_n2079# 0.01fF
C4679 VDD.t258 a_1596_n2079# 0.01fF
C4680 VDD.n190 a_1596_n2079# 0.05fF $ **FLOATING
C4681 VDD.n191 a_1596_n2079# 0.03fF $ **FLOATING
C4682 VDD.n192 a_1596_n2079# 1.05fF $ **FLOATING
C4683 VDD.t365 a_1596_n2079# 0.01fF
C4684 VDD.t366 a_1596_n2079# 0.01fF
C4685 VDD.n193 a_1596_n2079# 0.11fF $ **FLOATING
C4686 VDD.t367 a_1596_n2079# 0.01fF
C4687 VDD.t402 a_1596_n2079# 0.01fF
C4688 VDD.t404 a_1596_n2079# 0.01fF
C4689 VDD.t403 a_1596_n2079# 0.01fF
C4690 VDD.n194 a_1596_n2079# 0.07fF $ **FLOATING
C4691 VDD.n195 a_1596_n2079# 0.10fF $ **FLOATING
C4692 VDD.n196 a_1596_n2079# 0.13fF $ **FLOATING
C4693 VDD.n197 a_1596_n2079# 0.04fF $ **FLOATING
C4694 VDD.n198 a_1596_n2079# 0.25fF $ **FLOATING
C4695 VDD.t355 a_1596_n2079# 0.01fF
C4696 VDD.t356 a_1596_n2079# 0.01fF
C4697 VDD.n199 a_1596_n2079# 0.11fF $ **FLOATING
C4698 VDD.t357 a_1596_n2079# 0.01fF
C4699 VDD.t198 a_1596_n2079# 0.01fF
C4700 VDD.t196 a_1596_n2079# 0.01fF
C4701 VDD.t197 a_1596_n2079# 0.01fF
C4702 VDD.n200 a_1596_n2079# 0.07fF $ **FLOATING
C4703 VDD.n201 a_1596_n2079# 0.10fF $ **FLOATING
C4704 VDD.n202 a_1596_n2079# 0.13fF $ **FLOATING
C4705 VDD.n203 a_1596_n2079# 0.04fF $ **FLOATING
C4706 VDD.t160 a_1596_n2079# 0.01fF
C4707 VDD.t288 a_1596_n2079# 0.01fF
C4708 VDD.n204 a_1596_n2079# 0.05fF $ **FLOATING
C4709 VDD.t466 a_1596_n2079# 0.01fF
C4710 VDD.t465 a_1596_n2079# 0.01fF
C4711 VDD.t186 a_1596_n2079# 0.01fF
C4712 VDD.n205 a_1596_n2079# 0.05fF $ **FLOATING
C4713 VDD.n206 a_1596_n2079# 0.10fF $ **FLOATING
C4714 VDD.n207 a_1596_n2079# 0.06fF $ **FLOATING
C4715 VDD.t135 a_1596_n2079# 0.01fF
C4716 VDD.t137 a_1596_n2079# 0.01fF
C4717 VDD.n208 a_1596_n2079# 0.06fF $ **FLOATING
C4718 VDD.t302 a_1596_n2079# 0.01fF
C4719 VDD.t136 a_1596_n2079# 0.01fF
C4720 VDD.n209 a_1596_n2079# 0.05fF $ **FLOATING
C4721 VDD.n210 a_1596_n2079# 0.03fF $ **FLOATING
C4722 VDD.t171 a_1596_n2079# 0.01fF
C4723 VDD.t190 a_1596_n2079# 0.01fF
C4724 VDD.n211 a_1596_n2079# 0.10fF $ **FLOATING
C4725 VDD.t172 a_1596_n2079# 0.01fF
C4726 VDD.t226 a_1596_n2079# 0.01fF
C4727 VDD.n212 a_1596_n2079# 0.20fF $ **FLOATING
C4728 VDD.t319 a_1596_n2079# 0.01fF
C4729 VDD.t204 a_1596_n2079# 0.01fF
C4730 VDD.n213 a_1596_n2079# 0.08fF $ **FLOATING
C4731 VDD.n214 a_1596_n2079# 0.06fF $ **FLOATING
C4732 VDD.n215 a_1596_n2079# 0.03fF $ **FLOATING
C4733 VDD.t316 a_1596_n2079# 0.01fF
C4734 VDD.t299 a_1596_n2079# 0.01fF
C4735 VDD.n216 a_1596_n2079# 0.10fF $ **FLOATING
C4736 VDD.t312 a_1596_n2079# 0.01fF
C4737 VDD.t50 a_1596_n2079# 0.01fF
C4738 VDD.n217 a_1596_n2079# 0.20fF $ **FLOATING
C4739 VDD.t298 a_1596_n2079# 0.01fF
C4740 VDD.t102 a_1596_n2079# 0.01fF
C4741 VDD.n218 a_1596_n2079# 0.08fF $ **FLOATING
C4742 VDD.n219 a_1596_n2079# 0.06fF $ **FLOATING
C4743 VDD.n220 a_1596_n2079# 0.03fF $ **FLOATING
C4744 VDD.n221 a_1596_n2079# 0.04fF $ **FLOATING
C4745 VDD.t413 a_1596_n2079# 0.01fF
C4746 VDD.t412 a_1596_n2079# 0.01fF
C4747 VDD.n222 a_1596_n2079# 0.05fF $ **FLOATING
C4748 VDD.t77 a_1596_n2079# 0.01fF
C4749 VDD.t130 a_1596_n2079# 0.01fF
C4750 VDD.t300 a_1596_n2079# 0.01fF
C4751 VDD.n223 a_1596_n2079# 0.05fF $ **FLOATING
C4752 VDD.n224 a_1596_n2079# 0.10fF $ **FLOATING
C4753 VDD.n225 a_1596_n2079# 0.06fF $ **FLOATING
C4754 VDD.t58 a_1596_n2079# 0.01fF
C4755 VDD.t59 a_1596_n2079# 0.01fF
C4756 VDD.n226 a_1596_n2079# 0.06fF $ **FLOATING
C4757 VDD.t191 a_1596_n2079# 0.01fF
C4758 VDD.t57 a_1596_n2079# 0.01fF
C4759 VDD.n227 a_1596_n2079# 0.05fF $ **FLOATING
C4760 VDD.n228 a_1596_n2079# 0.03fF $ **FLOATING
C4761 VDD.t427 a_1596_n2079# 0.01fF
C4762 VDD.t428 a_1596_n2079# 0.01fF
C4763 VDD.n229 a_1596_n2079# 0.06fF $ **FLOATING
C4764 VDD.t341 a_1596_n2079# 0.01fF
C4765 VDD.t426 a_1596_n2079# 0.01fF
C4766 VDD.n230 a_1596_n2079# 0.05fF $ **FLOATING
C4767 VDD.n231 a_1596_n2079# 0.03fF $ **FLOATING
C4768 VDD.t203 a_1596_n2079# 0.01fF
C4769 VDD.t202 a_1596_n2079# 0.01fF
C4770 VDD.n232 a_1596_n2079# 0.05fF $ **FLOATING
C4771 VDD.t56 a_1596_n2079# 0.01fF
C4772 VDD.t55 a_1596_n2079# 0.01fF
C4773 VDD.t313 a_1596_n2079# 0.01fF
C4774 VDD.n233 a_1596_n2079# 0.05fF $ **FLOATING
C4775 VDD.n234 a_1596_n2079# 0.10fF $ **FLOATING
C4776 VDD.n235 a_1596_n2079# 0.06fF $ **FLOATING
C4777 VDD.n236 a_1596_n2079# 2.25fF $ **FLOATING
C4778 VDD.n237 a_1596_n2079# 3.06fF $ **FLOATING
C4779 VDD.n238 a_1596_n2079# 2.30fF $ **FLOATING
C4780 VDD.t118 a_1596_n2079# 0.01fF
C4781 VDD.t167 a_1596_n2079# 0.01fF
C4782 VDD.n239 a_1596_n2079# 0.10fF $ **FLOATING
C4783 VDD.t119 a_1596_n2079# 0.01fF
C4784 VDD.t120 a_1596_n2079# 0.01fF
C4785 VDD.n240 a_1596_n2079# 0.20fF $ **FLOATING
C4786 VDD.t166 a_1596_n2079# 0.01fF
C4787 VDD.t165 a_1596_n2079# 0.01fF
C4788 VDD.n241 a_1596_n2079# 0.08fF $ **FLOATING
C4789 VDD.n242 a_1596_n2079# 0.06fF $ **FLOATING
C4790 VDD.n243 a_1596_n2079# 0.03fF $ **FLOATING
C4791 VDD.t340 a_1596_n2079# 0.01fF
C4792 VDD.t475 a_1596_n2079# 0.01fF
C4793 VDD.n244 a_1596_n2079# 0.10fF $ **FLOATING
C4794 VDD.t474 a_1596_n2079# 0.01fF
C4795 VDD.t301 a_1596_n2079# 0.01fF
C4796 VDD.n245 a_1596_n2079# 0.20fF $ **FLOATING
C4797 VDD.t92 a_1596_n2079# 0.01fF
C4798 VDD.t215 a_1596_n2079# 0.01fF
C4799 VDD.n246 a_1596_n2079# 0.08fF $ **FLOATING
C4800 VDD.n247 a_1596_n2079# 0.06fF $ **FLOATING
C4801 VDD.n248 a_1596_n2079# 0.03fF $ **FLOATING
C4802 VDD.n249 a_1596_n2079# 0.04fF $ **FLOATING
C4803 VDD.n250 a_1596_n2079# 2.86fF $ **FLOATING
C4804 VDD.t139 a_1596_n2079# 0.01fF
C4805 VDD.t140 a_1596_n2079# 0.01fF
C4806 VDD.n251 a_1596_n2079# 0.11fF $ **FLOATING
C4807 VDD.t141 a_1596_n2079# 0.01fF
C4808 VDD.t398 a_1596_n2079# 0.01fF
C4809 VDD.t396 a_1596_n2079# 0.01fF
C4810 VDD.t397 a_1596_n2079# 0.01fF
C4811 VDD.n252 a_1596_n2079# 0.07fF $ **FLOATING
C4812 VDD.n253 a_1596_n2079# 0.10fF $ **FLOATING
C4813 VDD.n254 a_1596_n2079# 0.13fF $ **FLOATING
C4814 VDD.n255 a_1596_n2079# 0.04fF $ **FLOATING
C4815 VDD.t292 a_1596_n2079# 0.01fF
C4816 VDD.t293 a_1596_n2079# 0.01fF
C4817 VDD.n256 a_1596_n2079# 0.11fF $ **FLOATING
C4818 VDD.t294 a_1596_n2079# 0.01fF
C4819 VDD.t370 a_1596_n2079# 0.01fF
C4820 VDD.t368 a_1596_n2079# 0.01fF
C4821 VDD.t369 a_1596_n2079# 0.01fF
C4822 VDD.n257 a_1596_n2079# 0.07fF $ **FLOATING
C4823 VDD.n258 a_1596_n2079# 0.10fF $ **FLOATING
C4824 VDD.n259 a_1596_n2079# 0.13fF $ **FLOATING
C4825 VDD.n260 a_1596_n2079# 0.04fF $ **FLOATING
C4826 VDD.t314 a_1596_n2079# 0.01fF
C4827 VDD.t227 a_1596_n2079# 0.01fF
C4828 VDD.n261 a_1596_n2079# 0.05fF $ **FLOATING
C4829 VDD.t317 a_1596_n2079# 0.01fF
C4830 VDD.t433 a_1596_n2079# 0.01fF
C4831 VDD.t103 a_1596_n2079# 0.01fF
C4832 VDD.n262 a_1596_n2079# 0.05fF $ **FLOATING
C4833 VDD.n263 a_1596_n2079# 0.10fF $ **FLOATING
C4834 VDD.n264 a_1596_n2079# 0.06fF $ **FLOATING
C4835 VDD.t372 a_1596_n2079# 0.01fF
C4836 VDD.t371 a_1596_n2079# 0.01fF
C4837 VDD.n265 a_1596_n2079# 0.06fF $ **FLOATING
C4838 VDD.t155 a_1596_n2079# 0.01fF
C4839 VDD.t373 a_1596_n2079# 0.01fF
C4840 VDD.n266 a_1596_n2079# 0.05fF $ **FLOATING
C4841 VDD.n267 a_1596_n2079# 0.03fF $ **FLOATING
C4842 VDD.t152 a_1596_n2079# 0.01fF
C4843 VDD.t154 a_1596_n2079# 0.01fF
C4844 VDD.n268 a_1596_n2079# 0.10fF $ **FLOATING
C4845 VDD.t153 a_1596_n2079# 0.01fF
C4846 VDD.t188 a_1596_n2079# 0.01fF
C4847 VDD.n269 a_1596_n2079# 0.20fF $ **FLOATING
C4848 VDD.t243 a_1596_n2079# 0.01fF
C4849 VDD.t189 a_1596_n2079# 0.01fF
C4850 VDD.n270 a_1596_n2079# 0.08fF $ **FLOATING
C4851 VDD.n271 a_1596_n2079# 0.06fF $ **FLOATING
C4852 VDD.n272 a_1596_n2079# 0.03fF $ **FLOATING
C4853 VDD.t304 a_1596_n2079# 0.01fF
C4854 VDD.t51 a_1596_n2079# 0.01fF
C4855 VDD.n273 a_1596_n2079# 0.10fF $ **FLOATING
C4856 VDD.t236 a_1596_n2079# 0.01fF
C4857 VDD.t272 a_1596_n2079# 0.01fF
C4858 VDD.n274 a_1596_n2079# 0.20fF $ **FLOATING
C4859 VDD.t351 a_1596_n2079# 0.01fF
C4860 VDD.t429 a_1596_n2079# 0.01fF
C4861 VDD.n275 a_1596_n2079# 0.08fF $ **FLOATING
C4862 VDD.n276 a_1596_n2079# 0.06fF $ **FLOATING
C4863 VDD.n277 a_1596_n2079# 0.03fF $ **FLOATING
C4864 VDD.n278 a_1596_n2079# 0.04fF $ **FLOATING
C4865 VDD.t255 a_1596_n2079# 0.01fF
C4866 VDD.t360 a_1596_n2079# 0.01fF
C4867 VDD.n279 a_1596_n2079# 0.05fF $ **FLOATING
C4868 VDD.t85 a_1596_n2079# 0.01fF
C4869 VDD.t199 a_1596_n2079# 0.01fF
C4870 VDD.t182 a_1596_n2079# 0.01fF
C4871 VDD.n280 a_1596_n2079# 0.05fF $ **FLOATING
C4872 VDD.n281 a_1596_n2079# 0.10fF $ **FLOATING
C4873 VDD.n282 a_1596_n2079# 0.06fF $ **FLOATING
C4874 VDD.t330 a_1596_n2079# 0.01fF
C4875 VDD.t331 a_1596_n2079# 0.01fF
C4876 VDD.n283 a_1596_n2079# 0.06fF $ **FLOATING
C4877 VDD.t359 a_1596_n2079# 0.01fF
C4878 VDD.t329 a_1596_n2079# 0.01fF
C4879 VDD.n284 a_1596_n2079# 0.05fF $ **FLOATING
C4880 VDD.n285 a_1596_n2079# 0.03fF $ **FLOATING
C4881 VDD.t400 a_1596_n2079# 0.01fF
C4882 VDD.t401 a_1596_n2079# 0.01fF
C4883 VDD.n286 a_1596_n2079# 0.06fF $ **FLOATING
C4884 VDD.t76 a_1596_n2079# 0.01fF
C4885 VDD.t399 a_1596_n2079# 0.01fF
C4886 VDD.n287 a_1596_n2079# 0.05fF $ **FLOATING
C4887 VDD.n288 a_1596_n2079# 0.03fF $ **FLOATING
C4888 VDD.t105 a_1596_n2079# 0.01fF
C4889 VDD.t78 a_1596_n2079# 0.01fF
C4890 VDD.n289 a_1596_n2079# 0.05fF $ **FLOATING
C4891 VDD.t231 a_1596_n2079# 0.01fF
C4892 VDD.t87 a_1596_n2079# 0.01fF
C4893 VDD.t315 a_1596_n2079# 0.01fF
C4894 VDD.n290 a_1596_n2079# 0.05fF $ **FLOATING
C4895 VDD.n291 a_1596_n2079# 0.10fF $ **FLOATING
C4896 VDD.n292 a_1596_n2079# 0.06fF $ **FLOATING
C4897 VDD.n293 a_1596_n2079# 2.25fF $ **FLOATING
C4898 VDD.n294 a_1596_n2079# 3.06fF $ **FLOATING
C4899 VDD.n295 a_1596_n2079# 2.30fF $ **FLOATING
C4900 VDD.t6 a_1596_n2079# 0.01fF
C4901 VDD.t4 a_1596_n2079# 0.01fF
C4902 VDD.n296 a_1596_n2079# 0.10fF $ **FLOATING
C4903 VDD.t5 a_1596_n2079# 0.01fF
C4904 VDD.t3 a_1596_n2079# 0.01fF
C4905 VDD.n297 a_1596_n2079# 0.20fF $ **FLOATING
C4906 VDD.t1 a_1596_n2079# 0.01fF
C4907 VDD.t2 a_1596_n2079# 0.01fF
C4908 VDD.n298 a_1596_n2079# 0.08fF $ **FLOATING
C4909 VDD.n299 a_1596_n2079# 0.06fF $ **FLOATING
C4910 VDD.n300 a_1596_n2079# 0.03fF $ **FLOATING
C4911 VDD.t279 a_1596_n2079# 0.01fF
C4912 VDD.t380 a_1596_n2079# 0.01fF
C4913 VDD.n301 a_1596_n2079# 0.10fF $ **FLOATING
C4914 VDD.t320 a_1596_n2079# 0.01fF
C4915 VDD.t503 a_1596_n2079# 0.01fF
C4916 VDD.n302 a_1596_n2079# 0.20fF $ **FLOATING
C4917 VDD.t208 a_1596_n2079# 0.01fF
C4918 VDD.t376 a_1596_n2079# 0.01fF
C4919 VDD.n303 a_1596_n2079# 0.08fF $ **FLOATING
C4920 VDD.n304 a_1596_n2079# 0.06fF $ **FLOATING
C4921 VDD.n305 a_1596_n2079# 0.03fF $ **FLOATING
C4922 VDD.n306 a_1596_n2079# 0.04fF $ **FLOATING
C4923 VDD.n307 a_1596_n2079# 2.86fF $ **FLOATING
C4924 VDD.t73 a_1596_n2079# 0.01fF
C4925 VDD.t74 a_1596_n2079# 0.01fF
C4926 VDD.n308 a_1596_n2079# 0.11fF $ **FLOATING
C4927 VDD.t72 a_1596_n2079# 0.01fF
C4928 VDD.t390 a_1596_n2079# 0.01fF
C4929 VDD.t391 a_1596_n2079# 0.01fF
C4930 VDD.t392 a_1596_n2079# 0.01fF
C4931 VDD.n309 a_1596_n2079# 0.07fF $ **FLOATING
C4932 VDD.n310 a_1596_n2079# 0.10fF $ **FLOATING
C4933 VDD.n311 a_1596_n2079# 0.13fF $ **FLOATING
C4934 VDD.n312 a_1596_n2079# 0.04fF $ **FLOATING
C4935 VDD.t307 a_1596_n2079# 0.01fF
C4936 VDD.t308 a_1596_n2079# 0.01fF
C4937 VDD.n313 a_1596_n2079# 0.11fF $ **FLOATING
C4938 VDD.t306 a_1596_n2079# 0.01fF
C4939 VDD.t211 a_1596_n2079# 0.01fF
C4940 VDD.t209 a_1596_n2079# 0.01fF
C4941 VDD.t210 a_1596_n2079# 0.01fF
C4942 VDD.n314 a_1596_n2079# 0.07fF $ **FLOATING
C4943 VDD.n315 a_1596_n2079# 0.10fF $ **FLOATING
C4944 VDD.n316 a_1596_n2079# 0.13fF $ **FLOATING
C4945 VDD.n317 a_1596_n2079# 0.04fF $ **FLOATING
C4946 VDD.t361 a_1596_n2079# 0.01fF
C4947 VDD.t256 a_1596_n2079# 0.01fF
C4948 VDD.n318 a_1596_n2079# 0.05fF $ **FLOATING
C4949 VDD.t462 a_1596_n2079# 0.01fF
C4950 VDD.t268 a_1596_n2079# 0.01fF
C4951 VDD.t469 a_1596_n2079# 0.01fF
C4952 VDD.n319 a_1596_n2079# 0.05fF $ **FLOATING
C4953 VDD.n320 a_1596_n2079# 0.10fF $ **FLOATING
C4954 VDD.n321 a_1596_n2079# 0.06fF $ **FLOATING
C4955 VDD.t406 a_1596_n2079# 0.01fF
C4956 VDD.t407 a_1596_n2079# 0.01fF
C4957 VDD.n322 a_1596_n2079# 0.06fF $ **FLOATING
C4958 VDD.t244 a_1596_n2079# 0.01fF
C4959 VDD.t405 a_1596_n2079# 0.01fF
C4960 VDD.n323 a_1596_n2079# 0.05fF $ **FLOATING
C4961 VDD.n324 a_1596_n2079# 0.03fF $ **FLOATING
C4962 VDD.t280 a_1596_n2079# 0.01fF
C4963 VDD.t343 a_1596_n2079# 0.01fF
C4964 VDD.n325 a_1596_n2079# 0.10fF $ **FLOATING
C4965 VDD.t311 a_1596_n2079# 0.01fF
C4966 VDD.t335 a_1596_n2079# 0.01fF
C4967 VDD.n326 a_1596_n2079# 0.20fF $ **FLOATING
C4968 VDD.t440 a_1596_n2079# 0.01fF
C4969 VDD.t439 a_1596_n2079# 0.01fF
C4970 VDD.n327 a_1596_n2079# 0.08fF $ **FLOATING
C4971 VDD.n328 a_1596_n2079# 0.06fF $ **FLOATING
C4972 VDD.n329 a_1596_n2079# 0.03fF $ **FLOATING
C4973 VDD.t387 a_1596_n2079# 0.01fF
C4974 VDD.t12 a_1596_n2079# 0.01fF
C4975 VDD.n330 a_1596_n2079# 0.10fF $ **FLOATING
C4976 VDD.t183 a_1596_n2079# 0.01fF
C4977 VDD.t11 a_1596_n2079# 0.01fF
C4978 VDD.n331 a_1596_n2079# 0.20fF $ **FLOATING
C4979 VDD.t10 a_1596_n2079# 0.01fF
C4980 VDD.t86 a_1596_n2079# 0.01fF
C4981 VDD.n332 a_1596_n2079# 0.08fF $ **FLOATING
C4982 VDD.n333 a_1596_n2079# 0.06fF $ **FLOATING
C4983 VDD.n334 a_1596_n2079# 0.03fF $ **FLOATING
C4984 VDD.n335 a_1596_n2079# 0.04fF $ **FLOATING
C4985 VDD.t309 a_1596_n2079# 0.01fF
C4986 VDD.t282 a_1596_n2079# 0.01fF
C4987 VDD.n336 a_1596_n2079# 0.05fF $ **FLOATING
C4988 VDD.t423 a_1596_n2079# 0.01fF
C4989 VDD.t422 a_1596_n2079# 0.01fF
C4990 VDD.t421 a_1596_n2079# 0.01fF
C4991 VDD.n337 a_1596_n2079# 0.05fF $ **FLOATING
C4992 VDD.n338 a_1596_n2079# 0.10fF $ **FLOATING
C4993 VDD.n339 a_1596_n2079# 0.06fF $ **FLOATING
C4994 VDD.t457 a_1596_n2079# 0.01fF
C4995 VDD.t458 a_1596_n2079# 0.01fF
C4996 VDD.n340 a_1596_n2079# 0.06fF $ **FLOATING
C4997 VDD.t281 a_1596_n2079# 0.01fF
C4998 VDD.t459 a_1596_n2079# 0.01fF
C4999 VDD.n341 a_1596_n2079# 0.05fF $ **FLOATING
C5000 VDD.n342 a_1596_n2079# 0.03fF $ **FLOATING
C5001 VDD.t163 a_1596_n2079# 0.01fF
C5002 VDD.t161 a_1596_n2079# 0.01fF
C5003 VDD.n343 a_1596_n2079# 0.06fF $ **FLOATING
C5004 VDD.t416 a_1596_n2079# 0.01fF
C5005 VDD.t162 a_1596_n2079# 0.01fF
C5006 VDD.n344 a_1596_n2079# 0.05fF $ **FLOATING
C5007 VDD.n345 a_1596_n2079# 0.03fF $ **FLOATING
C5008 VDD.t420 a_1596_n2079# 0.01fF
C5009 VDD.t419 a_1596_n2079# 0.01fF
C5010 VDD.n346 a_1596_n2079# 0.05fF $ **FLOATING
C5011 VDD.t493 a_1596_n2079# 0.01fF
C5012 VDD.t42 a_1596_n2079# 0.01fF
C5013 VDD.t41 a_1596_n2079# 0.01fF
C5014 VDD.n347 a_1596_n2079# 0.05fF $ **FLOATING
C5015 VDD.n348 a_1596_n2079# 0.10fF $ **FLOATING
C5016 VDD.n349 a_1596_n2079# 0.06fF $ **FLOATING
C5017 VDD.n350 a_1596_n2079# 2.25fF $ **FLOATING
C5018 VDD.n351 a_1596_n2079# 3.06fF $ **FLOATING
C5019 VDD.n352 a_1596_n2079# 2.30fF $ **FLOATING
C5020 VDD.t75 a_1596_n2079# 0.01fF
C5021 VDD.t461 a_1596_n2079# 0.01fF
C5022 VDD.n353 a_1596_n2079# 0.10fF $ **FLOATING
C5023 VDD.t263 a_1596_n2079# 0.01fF
C5024 VDD.t318 a_1596_n2079# 0.01fF
C5025 VDD.n354 a_1596_n2079# 0.20fF $ **FLOATING
C5026 VDD.t185 a_1596_n2079# 0.01fF
C5027 VDD.t463 a_1596_n2079# 0.01fF
C5028 VDD.n355 a_1596_n2079# 0.08fF $ **FLOATING
C5029 VDD.n356 a_1596_n2079# 0.06fF $ **FLOATING
C5030 VDD.n357 a_1596_n2079# 0.03fF $ **FLOATING
C5031 VDD.t418 a_1596_n2079# 0.01fF
C5032 VDD.t417 a_1596_n2079# 0.01fF
C5033 VDD.n358 a_1596_n2079# 0.10fF $ **FLOATING
C5034 VDD.t415 a_1596_n2079# 0.01fF
C5035 VDD.t414 a_1596_n2079# 0.01fF
C5036 VDD.n359 a_1596_n2079# 0.20fF $ **FLOATING
C5037 VDD.t200 a_1596_n2079# 0.01fF
C5038 VDD.t424 a_1596_n2079# 0.01fF
C5039 VDD.n360 a_1596_n2079# 0.08fF $ **FLOATING
C5040 VDD.n361 a_1596_n2079# 0.06fF $ **FLOATING
C5041 VDD.n362 a_1596_n2079# 0.03fF $ **FLOATING
C5042 VDD.n363 a_1596_n2079# 0.04fF $ **FLOATING
C5043 VDD.n364 a_1596_n2079# 2.85fF $ **FLOATING
C5044 VDD.t8 a_1596_n2079# 0.01fF
C5045 VDD.t9 a_1596_n2079# 0.01fF
C5046 VDD.n365 a_1596_n2079# 0.11fF $ **FLOATING
C5047 VDD.t7 a_1596_n2079# 0.01fF
C5048 VDD.t290 a_1596_n2079# 0.01fF
C5049 VDD.t289 a_1596_n2079# 0.01fF
C5050 VDD.t291 a_1596_n2079# 0.01fF
C5051 VDD.n366 a_1596_n2079# 0.07fF $ **FLOATING
C5052 VDD.n367 a_1596_n2079# 0.10fF $ **FLOATING
C5053 VDD.n368 a_1596_n2079# 0.13fF $ **FLOATING
C5054 VDD.n369 a_1596_n2079# 0.04fF $ **FLOATING
C5055 VDD.t240 a_1596_n2079# 0.01fF
C5056 VDD.t241 a_1596_n2079# 0.01fF
C5057 VDD.n370 a_1596_n2079# 0.11fF $ **FLOATING
C5058 VDD.t242 a_1596_n2079# 0.01fF
C5059 VDD.t328 a_1596_n2079# 0.01fF
C5060 VDD.t326 a_1596_n2079# 0.01fF
C5061 VDD.t327 a_1596_n2079# 0.01fF
C5062 VDD.n371 a_1596_n2079# 0.07fF $ **FLOATING
C5063 VDD.n372 a_1596_n2079# 0.10fF $ **FLOATING
C5064 VDD.n373 a_1596_n2079# 0.13fF $ **FLOATING
C5065 VDD.n374 a_1596_n2079# 0.04fF $ **FLOATING
C5066 VDD.t342 a_1596_n2079# 0.01fF
C5067 VDD.t310 a_1596_n2079# 0.01fF
C5068 VDD.n375 a_1596_n2079# 0.05fF $ **FLOATING
C5069 VDD.t184 a_1596_n2079# 0.01fF
C5070 VDD.t386 a_1596_n2079# 0.01fF
C5071 VDD.t388 a_1596_n2079# 0.01fF
C5072 VDD.n376 a_1596_n2079# 0.05fF $ **FLOATING
C5073 VDD.n377 a_1596_n2079# 0.10fF $ **FLOATING
C5074 VDD.n378 a_1596_n2079# 0.06fF $ **FLOATING
C5075 VDD.t278 a_1596_n2079# 0.01fF
C5076 VDD.t277 a_1596_n2079# 0.01fF
C5077 VDD.n379 a_1596_n2079# 0.06fF $ **FLOATING
C5078 VDD.t441 a_1596_n2079# 0.01fF
C5079 VDD.t276 a_1596_n2079# 0.01fF
C5080 VDD.n380 a_1596_n2079# 0.05fF $ **FLOATING
C5081 VDD.n381 a_1596_n2079# 0.03fF $ **FLOATING
C5082 VDD.n382 a_1596_n2079# 0.96fF $ **FLOATING
C5083 VDD.n383 a_1596_n2079# 3.36fF $ **FLOATING
C5084 VDD.n384 a_1596_n2079# 1.50fF $ **FLOATING
C5085 VDD.n385 a_1596_n2079# 3.73fF $ **FLOATING
C5086 VDD.n386 a_1596_n2079# 4.52fF $ **FLOATING
C5087 VDD.n387 a_1596_n2079# 3.34fF $ **FLOATING
C5088 VDD.n388 a_1596_n2079# 1.50fF $ **FLOATING
C5089 VDD.n389 a_1596_n2079# 3.75fF $ **FLOATING
C5090 VDD.n390 a_1596_n2079# 4.54fF $ **FLOATING
C5091 VDD.n391 a_1596_n2079# 3.34fF $ **FLOATING
C5092 VDD.n392 a_1596_n2079# 1.50fF $ **FLOATING
C5093 VDD.n393 a_1596_n2079# 3.77fF $ **FLOATING
C5094 VDD.n394 a_1596_n2079# 4.55fF $ **FLOATING
C5095 VDD.n395 a_1596_n2079# 2.95fF $ **FLOATING
C5096 VDD.t169 a_1596_n2079# 0.01fF
C5097 VDD.t131 a_1596_n2079# 0.01fF
C5098 VDD.n396 a_1596_n2079# 0.10fF $ **FLOATING
C5099 VDD.t170 a_1596_n2079# 0.01fF
C5100 VDD.t285 a_1596_n2079# 0.01fF
C5101 VDD.n397 a_1596_n2079# 0.20fF $ **FLOATING
C5102 VDD.t168 a_1596_n2079# 0.01fF
C5103 VDD.t286 a_1596_n2079# 0.01fF
C5104 VDD.n398 a_1596_n2079# 0.08fF $ **FLOATING
C5105 VDD.n399 a_1596_n2079# 0.06fF $ **FLOATING
C5106 VDD.n400 a_1596_n2079# 0.03fF $ **FLOATING
C5107 VDD.t437 a_1596_n2079# 0.01fF
C5108 VDD.t132 a_1596_n2079# 0.01fF
C5109 VDD.n401 a_1596_n2079# 0.10fF $ **FLOATING
C5110 VDD.t100 a_1596_n2079# 0.01fF
C5111 VDD.t438 a_1596_n2079# 0.01fF
C5112 VDD.n402 a_1596_n2079# 0.20fF $ **FLOATING
C5113 VDD.t13 a_1596_n2079# 0.01fF
C5114 VDD.t101 a_1596_n2079# 0.01fF
C5115 VDD.n403 a_1596_n2079# 0.08fF $ **FLOATING
C5116 VDD.n404 a_1596_n2079# 0.06fF $ **FLOATING
C5117 VDD.n405 a_1596_n2079# 0.03fF $ **FLOATING
C5118 VDD.n406 a_1596_n2079# 0.04fF $ **FLOATING
C5119 VDD.t71 a_1596_n2079# 0.01fF
C5120 VDD.t70 a_1596_n2079# 0.01fF
C5121 VDD.n407 a_1596_n2079# 0.10fF $ **FLOATING
C5122 VDD.t353 a_1596_n2079# 0.01fF
C5123 VDD.t287 a_1596_n2079# 0.01fF
C5124 VDD.n408 a_1596_n2079# 0.20fF $ **FLOATING
C5125 VDD.t352 a_1596_n2079# 0.01fF
C5126 VDD.t69 a_1596_n2079# 0.01fF
C5127 VDD.n409 a_1596_n2079# 0.08fF $ **FLOATING
C5128 VDD.n410 a_1596_n2079# 0.06fF $ **FLOATING
C5129 VDD.n411 a_1596_n2079# 0.03fF $ **FLOATING
C5130 VDD.t464 a_1596_n2079# 0.01fF
C5131 VDD.t467 a_1596_n2079# 0.01fF
C5132 VDD.n412 a_1596_n2079# 0.10fF $ **FLOATING
C5133 VDD.t18 a_1596_n2079# 0.01fF
C5134 VDD.t107 a_1596_n2079# 0.01fF
C5135 VDD.n413 a_1596_n2079# 0.20fF $ **FLOATING
C5136 VDD.t106 a_1596_n2079# 0.01fF
C5137 VDD.t129 a_1596_n2079# 0.01fF
C5138 VDD.n414 a_1596_n2079# 0.08fF $ **FLOATING
C5139 VDD.n415 a_1596_n2079# 0.06fF $ **FLOATING
C5140 VDD.n416 a_1596_n2079# 0.03fF $ **FLOATING
C5141 VDD.n417 a_1596_n2079# 0.04fF $ **FLOATING
C5142 VDD.t159 a_1596_n2079# 0.01fF
C5143 VDD.t297 a_1596_n2079# 0.01fF
C5144 VDD.n418 a_1596_n2079# 0.05fF $ **FLOATING
C5145 VDD.t62 a_1596_n2079# 0.01fF
C5146 VDD.t63 a_1596_n2079# 0.01fF
C5147 VDD.t61 a_1596_n2079# 0.01fF
C5148 VDD.n419 a_1596_n2079# 0.05fF $ **FLOATING
C5149 VDD.n420 a_1596_n2079# 0.10fF $ **FLOATING
C5150 VDD.n421 a_1596_n2079# 0.06fF $ **FLOATING
C5151 VDD.t495 a_1596_n2079# 0.01fF
C5152 VDD.t496 a_1596_n2079# 0.01fF
C5153 VDD.n422 a_1596_n2079# 0.06fF $ **FLOATING
C5154 VDD.t264 a_1596_n2079# 0.01fF
C5155 VDD.t494 a_1596_n2079# 0.01fF
C5156 VDD.n423 a_1596_n2079# 0.05fF $ **FLOATING
C5157 VDD.n424 a_1596_n2079# 0.03fF $ **FLOATING
C5158 VDD.t333 a_1596_n2079# 0.01fF
C5159 VDD.t334 a_1596_n2079# 0.01fF
C5160 VDD.n425 a_1596_n2079# 0.06fF $ **FLOATING
C5161 VDD.t14 a_1596_n2079# 0.01fF
C5162 VDD.t332 a_1596_n2079# 0.01fF
C5163 VDD.n426 a_1596_n2079# 0.05fF $ **FLOATING
C5164 VDD.n427 a_1596_n2079# 0.03fF $ **FLOATING
C5165 VDD.t133 a_1596_n2079# 0.01fF
C5166 VDD.t15 a_1596_n2079# 0.01fF
C5167 VDD.n428 a_1596_n2079# 0.05fF $ **FLOATING
C5168 VDD.t187 a_1596_n2079# 0.01fF
C5169 VDD.t468 a_1596_n2079# 0.01fF
C5170 VDD.t128 a_1596_n2079# 0.01fF
C5171 VDD.n429 a_1596_n2079# 0.05fF $ **FLOATING
C5172 VDD.n430 a_1596_n2079# 0.10fF $ **FLOATING
C5173 VDD.n431 a_1596_n2079# 0.06fF $ **FLOATING
C5174 VDD.n432 a_1596_n2079# 2.25fF $ **FLOATING
C5175 VDD.n433 a_1596_n2079# 3.06fF $ **FLOATING
C5176 VDD.n434 a_1596_n2079# 2.32fF $ **FLOATING
C5177 VDD.n435 a_1596_n2079# 2.64fF $ **FLOATING
C5178 VDD.n436 a_1596_n2079# 1.45fF $ **FLOATING
C5179 VDD.n437 a_1596_n2079# 0.88fF $ **FLOATING
C5180 VDD.n438 a_1596_n2079# 2.30fF $ **FLOATING
C5181 VDD.n439 a_1596_n2079# 3.84fF $ **FLOATING
C5182 VDD.t89 a_1596_n2079# 0.01fF
C5183 VDD.t224 a_1596_n2079# 0.01fF
C5184 VDD.n440 a_1596_n2079# 0.05fF $ **FLOATING
C5185 VDD.t322 a_1596_n2079# 0.01fF
C5186 VDD.t337 a_1596_n2079# 0.01fF
C5187 VDD.t284 a_1596_n2079# 0.01fF
C5188 VDD.n441 a_1596_n2079# 0.05fF $ **FLOATING
C5189 VDD.n442 a_1596_n2079# 0.10fF $ **FLOATING
C5190 VDD.n443 a_1596_n2079# 0.06fF $ **FLOATING
C5191 VDD.t500 a_1596_n2079# 0.01fF
C5192 VDD.t502 a_1596_n2079# 0.01fF
C5193 VDD.n444 a_1596_n2079# 0.06fF $ **FLOATING
C5194 VDD.t501 a_1596_n2079# 0.01fF
C5195 VDD.t23 a_1596_n2079# 0.01fF
C5196 VDD.n445 a_1596_n2079# 0.05fF $ **FLOATING
C5197 VDD.n446 a_1596_n2079# 0.03fF $ **FLOATING
C5198 VDD.n447 a_1596_n2079# 0.51fF $ **FLOATING
C5199 VDD.t358 a_1596_n2079# 0.01fF
C5200 VDD.t88 a_1596_n2079# 0.01fF
C5201 VDD.n448 a_1596_n2079# 0.10fF $ **FLOATING
C5202 VDD.t47 a_1596_n2079# 0.01fF
C5203 VDD.t46 a_1596_n2079# 0.01fF
C5204 VDD.n449 a_1596_n2079# 0.20fF $ **FLOATING
C5205 VDD.t90 a_1596_n2079# 0.01fF
C5206 VDD.t225 a_1596_n2079# 0.01fF
C5207 VDD.n450 a_1596_n2079# 0.08fF $ **FLOATING
C5208 VDD.n451 a_1596_n2079# 0.06fF $ **FLOATING
C5209 VDD.n452 a_1596_n2079# 0.03fF $ **FLOATING
C5210 VDD.t40 a_1596_n2079# 0.01fF
C5211 VDD.t91 a_1596_n2079# 0.01fF
C5212 VDD.n453 a_1596_n2079# 0.10fF $ **FLOATING
C5213 VDD.t0 a_1596_n2079# 0.01fF
C5214 VDD.t339 a_1596_n2079# 0.01fF
C5215 VDD.n454 a_1596_n2079# 0.20fF $ **FLOATING
C5216 VDD.t45 a_1596_n2079# 0.01fF
C5217 VDD.t442 a_1596_n2079# 0.01fF
C5218 VDD.n455 a_1596_n2079# 0.08fF $ **FLOATING
C5219 VDD.n456 a_1596_n2079# 0.06fF $ **FLOATING
C5220 VDD.n457 a_1596_n2079# 0.03fF $ **FLOATING
C5221 VDD.n458 a_1596_n2079# 0.04fF $ **FLOATING
C5222 VDD.n459 a_1596_n2079# 2.36fF $ **FLOATING
C5223 VDD.n460 a_1596_n2079# 4.76fF $ **FLOATING
C5224 VDD.n461 a_1596_n2079# 5.02fF $ **FLOATING
C5225 VDD.t179 a_1596_n2079# 0.01fF
C5226 VDD.t181 a_1596_n2079# 0.01fF
C5227 VDD.n462 a_1596_n2079# 0.11fF $ **FLOATING
C5228 VDD.t180 a_1596_n2079# 0.01fF
C5229 VDD.t52 a_1596_n2079# 0.01fF
C5230 VDD.t54 a_1596_n2079# 0.01fF
C5231 VDD.t53 a_1596_n2079# 0.01fF
C5232 VDD.n463 a_1596_n2079# 0.07fF $ **FLOATING
C5233 VDD.n464 a_1596_n2079# 0.10fF $ **FLOATING
C5234 VDD.n465 a_1596_n2079# 0.13fF $ **FLOATING
C5235 VDD.n466 a_1596_n2079# 0.04fF $ **FLOATING
C5236 VDD.n467 a_1596_n2079# 3.34fF $ **FLOATING
C5237 VDD.t207 a_1596_n2079# 0.01fF
C5238 VDD.t205 a_1596_n2079# 0.01fF
C5239 VDD.n468 a_1596_n2079# 0.11fF $ **FLOATING
C5240 VDD.t206 a_1596_n2079# 0.01fF
C5241 VDD.t246 a_1596_n2079# 0.01fF
C5242 VDD.t245 a_1596_n2079# 0.01fF
C5243 VDD.t247 a_1596_n2079# 0.01fF
C5244 VDD.n469 a_1596_n2079# 0.07fF $ **FLOATING
C5245 VDD.n470 a_1596_n2079# 0.10fF $ **FLOATING
C5246 VDD.n471 a_1596_n2079# 0.13fF $ **FLOATING
C5247 VDD.n472 a_1596_n2079# 0.04fF $ **FLOATING
C5248 VDD.n473 a_1596_n2079# 1.47fF $ **FLOATING
C5249 VDD.n474 a_1596_n2079# 3.77fF $ **FLOATING
C5250 VDD.t93 a_1596_n2079# 0.01fF
C5251 VDD.t347 a_1596_n2079# 0.01fF
C5252 VDD.n475 a_1596_n2079# 0.05fF $ **FLOATING
C5253 VDD.t250 a_1596_n2079# 0.01fF
C5254 VDD.t375 a_1596_n2079# 0.01fF
C5255 VDD.t434 a_1596_n2079# 0.01fF
C5256 VDD.n476 a_1596_n2079# 0.05fF $ **FLOATING
C5257 VDD.n477 a_1596_n2079# 0.10fF $ **FLOATING
C5258 VDD.n478 a_1596_n2079# 0.06fF $ **FLOATING
C5259 VDD.t229 a_1596_n2079# 0.01fF
C5260 VDD.t228 a_1596_n2079# 0.01fF
C5261 VDD.n479 a_1596_n2079# 0.06fF $ **FLOATING
C5262 VDD.t230 a_1596_n2079# 0.01fF
C5263 VDD.t389 a_1596_n2079# 0.01fF
C5264 VDD.n480 a_1596_n2079# 0.05fF $ **FLOATING
C5265 VDD.n481 a_1596_n2079# 0.03fF $ **FLOATING
C5266 VDD.n482 a_1596_n2079# 0.20fF $ **FLOATING
C5267 VDD.n483 a_1596_n2079# 4.32fF $ **FLOATING
C5268 VDD.t239 a_1596_n2079# 0.01fF
C5269 VDD.t238 a_1596_n2079# 0.01fF
C5270 VDD.n484 a_1596_n2079# 0.11fF $ **FLOATING
C5271 VDD.t237 a_1596_n2079# 0.01fF
C5272 VDD.t274 a_1596_n2079# 0.01fF
C5273 VDD.t273 a_1596_n2079# 0.01fF
C5274 VDD.t275 a_1596_n2079# 0.01fF
C5275 VDD.n485 a_1596_n2079# 0.07fF $ **FLOATING
C5276 VDD.n486 a_1596_n2079# 0.10fF $ **FLOATING
C5277 VDD.n487 a_1596_n2079# 0.13fF $ **FLOATING
C5278 VDD.n488 a_1596_n2079# 0.04fF $ **FLOATING
C5279 VDD.n489 a_1596_n2079# 3.33fF $ **FLOATING
C5280 VDD.t26 a_1596_n2079# 0.01fF
C5281 VDD.t25 a_1596_n2079# 0.01fF
C5282 VDD.n490 a_1596_n2079# 0.11fF $ **FLOATING
C5283 VDD.t24 a_1596_n2079# 0.01fF
C5284 VDD.t499 a_1596_n2079# 0.01fF
C5285 VDD.t498 a_1596_n2079# 0.01fF
C5286 VDD.t497 a_1596_n2079# 0.01fF
C5287 VDD.n491 a_1596_n2079# 0.07fF $ **FLOATING
C5288 VDD.n492 a_1596_n2079# 0.10fF $ **FLOATING
C5289 VDD.n493 a_1596_n2079# 0.13fF $ **FLOATING
C5290 VDD.n494 a_1596_n2079# 0.04fF $ **FLOATING
C5291 VDD.n495 a_1596_n2079# 1.40fF $ **FLOATING
C5292 VDD.n496 a_1596_n2079# 1.95fF $ **FLOATING
.ends

