* NGSPICE file created from logic_xor_pex.ext - technology: sky130B

.subckt logic_xor A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3]
+ Y[4] Y[5] Y[6] Y[7] VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7]
X0 a_6543_n476.t6 a_6955_n502.t4 Y[3].t1 VDD.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1 a_4475_n478.t5 A[2].t0 VDD.t223 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2 a_692_n1210.t0 A[0].t0 Y[0].t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3 Y[3].t0 a_6955_n502.t5 a_6543_n476.t5 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4 a_2818_n502.t2 B[1].t0 VDD.t237 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 a_338_n478.t6 a_n89_215.t4 Y[0].t7 VDD.t213 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X6 a_12749_n476.t4 A[6].t0 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 Y[2].t4 a_4048_215.t4 a_4475_n478.t8 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X8 a_13161_n502.t3 B[6].t0 VSS.t12 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X9 a_14817_n474.t8 B[7].t0 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10 VDD.t231 A[4].t0 a_8612_n476.t6 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 VSS.t27 B[0].t0 a_692_n1210.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X12 a_2406_n476.t7 a_2818_n502.t4 Y[1].t4 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X13 a_n89_215.t2 A[0].t1 VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X14 a_4475_n478.t4 A[2].t1 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X15 Y[7].t7 a_14390_219.t4 a_14817_n474.t10 VDD.t184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X16 VDD.t191 A[1].t0 a_2406_n476.t11 VDD.t190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 a_6543_n476.t2 A[3].t0 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 Y[4].t5 a_8185_217.t4 a_8612_n476.t2 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_8612_n476.t1 a_9024_n502.t4 Y[4].t0 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X20 VDD.t195 B[0].t1 a_338_n478.t10 VDD.t194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X21 Y[5].t6 a_10253_219.t4 a_10680_n474.t5 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X22 Y[1].t0 a_1979_217.t4 a_2524_n1208.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X23 a_14817_n474.t5 A[7].t0 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X24 VDD.t49 B[5].t0 a_11092_n500.t2 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X25 a_13161_n502.t2 B[6].t1 VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 a_6955_n502.t3 B[3].t0 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X27 a_4475_n478.t10 a_4887_n504.t4 Y[2].t7 VDD.t171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X28 VSS.t11 A[2].t2 a_4048_215.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X29 a_4887_n504.t0 B[2].t0 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X30 VSS.t10 A[5].t0 a_10253_219.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X31 VDD.t63 A[1].t1 a_1979_217.t2 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X32 a_15229_n500.t2 B[7].t1 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X33 a_13103_n1208.t0 A[6].t1 Y[6].t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X34 a_12749_n476.t11 a_12322_217.t4 Y[6].t7 VDD.t204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X35 a_338_n478.t9 B[0].t2 VDD.t193 VDD.t192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X36 VDD.t175 A[4].t1 a_8185_217.t2 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X37 Y[6].t6 a_12322_217.t5 a_12749_n476.t6 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X38 VDD.t59 A[6].t2 a_12749_n476.t3 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 a_2406_n476.t10 A[1].t2 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X40 VDD.t23 A[2].t3 a_4475_n478.t3 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X41 VSS.t14 B[6].t2 a_13103_n1208.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X42 a_6955_n502.t0 B[3].t1 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X43 a_8612_n476.t5 A[4].t2 VDD.t225 VDD.t224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X44 a_15229_n500.t3 B[7].t2 VSS.t16 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X45 a_4593_n1210.t1 a_4887_n504.t5 VSS.t24 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X46 a_2406_n476.t8 a_1979_217.t5 Y[1].t6 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X47 a_10680_n474.t10 A[5].t1 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X48 VDD.t8 A[3].t1 a_6543_n476.t1 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X49 a_14817_n474.t1 a_15229_n500.t4 Y[7].t1 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X50 VDD.t53 A[7].t1 a_14817_n474.t3 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X51 Y[4].t4 a_8185_217.t5 a_8612_n476.t3 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X52 a_338_n478.t3 A[0].t2 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X53 VSS.t29 B[4].t0 a_8966_n1208.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X54 Y[6].t0 a_12322_217.t6 a_12867_n1208.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X55 Y[6].t5 a_13161_n502.t4 a_12749_n476.t7 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X56 Y[3].t3 a_6116_217.t4 a_6543_n476.t9 VDD.t209 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X57 VDD.t181 B[2].t1 a_4475_n478.t11 VDD.t180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X58 a_8730_n1208.t0 a_9024_n502.t5 VSS.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X59 a_10680_n474.t4 a_11092_n500.t4 Y[5].t2 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X60 VDD.t86 B[6].t3 a_13161_n502.t1 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X61 a_11092_n500.t1 B[5].t1 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X62 VDD.t133 A[2].t4 a_4048_215.t2 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 VDD.t141 B[3].t2 a_6955_n502.t2 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X64 a_8185_217.t1 A[4].t3 VDD.t229 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X65 VDD.t34 A[5].t2 a_10680_n474.t3 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X66 a_456_n1210.t1 a_750_n504.t4 VSS.t20 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X67 a_8612_n476.t11 B[4].t1 VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X68 VDD.t135 B[7].t3 a_15229_n500.t1 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X69 a_1979_217.t1 A[1].t3 VDD.t227 VDD.t226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X70 Y[3].t7 a_6116_217.t5 a_6543_n476.t11 VDD.t239 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X71 VDD.t61 B[0].t3 a_338_n478.t0 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X72 a_8966_n1208.t1 A[4].t4 Y[4].t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X73 a_12749_n476.t2 A[6].t3 VDD.t235 VDD.t234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X74 a_750_n504.t3 B[0].t4 VSS.t26 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X75 a_338_n478.t8 a_750_n504.t5 Y[0].t5 VDD.t155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X76 VDD.t13 A[0].t3 a_338_n478.t2 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X77 a_6661_n1208.t0 a_6955_n502.t6 VSS.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X78 VDD.t219 B[1].t1 a_2406_n476.t4 VDD.t218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X79 a_6543_n476.t0 A[3].t2 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X80 a_13161_n502.t0 B[6].t4 VDD.t121 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X81 VDD.t206 B[4].t2 a_8612_n476.t10 VDD.t205 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X82 a_8612_n476.t8 a_9024_n502.t6 Y[4].t6 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X83 a_4475_n478.t9 B[2].t2 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X84 VDD.t173 B[5].t2 a_10680_n474.t11 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X85 Y[3].t6 a_6116_217.t6 a_6661_n1208.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X86 Y[5].t5 a_10253_219.t5 a_10680_n474.t6 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X87 Y[7].t4 a_14390_219.t5 a_14935_n1206.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 a_338_n478.t7 a_750_n504.t6 Y[0].t2 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X89 VSS.t6 A[4].t5 a_8185_217.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X90 a_6897_n1208.t0 A[3].t3 Y[3].t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X91 a_10680_n474.t1 a_11092_n500.t5 Y[5].t1 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X92 VDD.t32 B[4].t3 a_8612_n476.t0 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X93 VDD.t40 A[5].t3 a_10253_219.t0 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X94 a_2760_n1208.t0 A[1].t4 Y[1].t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X95 a_4048_215.t1 A[2].t5 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X96 Y[2].t1 a_4887_n504.t6 a_4475_n478.t1 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X97 a_12867_n1208.t1 a_13161_n502.t5 VSS.t13 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X98 a_11092_n500.t3 B[5].t3 VSS.t9 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X99 VSS.t23 B[3].t3 a_6897_n1208.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X100 VDD.t233 A[4].t6 a_8185_217.t0 VDD.t232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X101 Y[7].t6 a_14390_219.t6 a_14817_n474.t11 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X102 VSS.t8 A[0].t4 a_n89_215.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X103 a_15229_n500.t0 B[7].t4 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X104 a_12322_217.t2 A[6].t4 VDD.t162 VDD.t161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X105 VDD.t45 A[1].t5 a_1979_217.t0 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X106 a_6116_217.t2 A[3].t4 VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X107 Y[6].t1 a_12322_217.t7 a_12749_n476.t1 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X108 a_338_n478.t1 A[0].t5 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X109 Y[1].t7 a_1979_217.t6 a_2406_n476.t9 VDD.t185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X110 VSS.t25 A[3].t5 a_6116_217.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X111 VDD.t119 B[6].t5 a_12749_n476.t8 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X112 a_2406_n476.t3 B[1].t2 VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X113 VSS.t5 A[1].t6 a_1979_217.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X114 Y[7].t2 a_15229_n500.t5 a_14817_n474.t2 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X115 VDD.t93 A[6].t5 a_12322_217.t1 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X116 VDD.t95 A[3].t6 a_6116_217.t1 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X117 Y[0].t0 a_n89_215.t5 a_338_n478.t5 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X118 a_10680_n474.t8 B[5].t4 VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X119 VDD.t179 B[3].t4 a_6543_n476.t8 VDD.t178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X120 VDD.t217 A[0].t6 a_n89_215.t1 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X121 VSS.t1 B[5].t5 a_11034_n1206.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X122 VDD.t79 A[6].t6 a_12322_217.t0 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X123 VDD.t114 A[2].t6 a_4048_215.t0 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X124 a_10253_219.t3 A[5].t4 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X125 a_4475_n478.t7 a_4048_215.t5 Y[2].t3 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X126 VDD.t21 A[7].t2 a_14390_219.t0 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X127 Y[1].t1 a_1979_217.t7 a_2406_n476.t0 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X128 a_750_n504.t2 B[0].t5 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X129 a_14817_n474.t9 A[7].t3 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X130 a_8612_n476.t7 a_8185_217.t6 Y[4].t3 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X131 Y[2].t5 a_4048_215.t6 a_4593_n1210.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X132 a_6543_n476.t10 a_6116_217.t7 Y[3].t5 VDD.t238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X133 VDD.t151 A[3].t7 a_6116_217.t0 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X134 a_750_n504.t1 B[0].t6 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X135 a_15171_n1206.t0 A[7].t4 Y[7].t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X136 a_2818_n502.t1 B[1].t3 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X137 Y[5].t3 a_10253_219.t6 a_10798_n1206.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X138 a_4887_n504.t1 B[2].t3 VSS.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X139 a_6543_n476.t4 a_6955_n502.t7 Y[3].t2 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X140 Y[0].t4 a_n89_215.t6 a_338_n478.t4 VDD.t126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X141 a_4475_n478.t0 a_4887_n504.t7 Y[2].t0 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X142 Y[1].t5 a_2818_n502.t5 a_2406_n476.t6 VDD.t220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X143 a_11034_n1206.t0 A[5].t5 Y[5].t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X144 VDD.t215 B[1].t4 a_2406_n476.t2 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X145 a_2406_n476.t5 a_2818_n502.t6 Y[1].t3 VDD.t221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X146 VSS.t19 A[6].t7 a_12322_217.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X147 a_14817_n474.t4 a_14390_219.t7 Y[7].t5 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X148 a_12749_n476.t5 B[6].t6 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X149 VSS.t31 B[1].t5 a_2760_n1208.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X150 a_6543_n476.t3 B[3].t5 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X151 Y[4].t7 a_9024_n502.t7 a_8612_n476.t9 VDD.t199 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X152 VDD.t57 A[5].t6 a_10253_219.t1 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X153 a_9024_n502.t1 B[4].t4 VSS.t28 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X154 a_2524_n1208.t1 a_2818_n502.t7 VSS.t30 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X155 VDD.t25 B[5].t6 a_10680_n474.t2 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X156 a_10680_n474.t7 a_10253_219.t7 Y[5].t4 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X157 Y[0].t6 a_750_n504.t7 a_338_n478.t11 VDD.t196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X158 VDD.t149 A[0].t7 a_n89_215.t0 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X159 a_14390_219.t2 A[7].t5 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X160 VDD.t43 B[0].t7 a_750_n504.t0 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X161 a_4887_n504.t2 B[2].t4 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X162 VDD.t203 B[4].t5 a_9024_n502.t3 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X163 VDD.t28 B[2].t5 a_4475_n478.t2 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X164 a_12749_n476.t9 a_13161_n502.t6 Y[6].t4 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X165 VDD.t128 B[1].t6 a_2818_n502.t0 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X166 a_6955_n502.t1 B[3].t6 VSS.t18 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X167 Y[5].t0 a_11092_n500.t6 a_10680_n474.t0 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X168 VDD.t212 B[7].t5 a_14817_n474.t7 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X169 a_2818_n502.t3 B[1].t7 VSS.t15 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X170 a_8612_n476.t4 A[4].t7 VDD.t187 VDD.t186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X171 a_2406_n476.t1 A[1].t7 VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X172 VDD.t183 B[6].t7 a_12749_n476.t10 VDD.t182 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X173 a_10680_n474.t9 A[5].t7 VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X174 VSS.t22 A[7].t6 a_14390_219.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X175 a_14817_n474.t0 a_15229_n500.t6 Y[7].t0 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X176 VDD.t177 B[3].t7 a_6543_n476.t7 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X177 a_9024_n502.t2 B[4].t6 VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X178 a_12749_n476.t0 a_13161_n502.t7 Y[6].t3 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X179 a_4829_n1210.t0 A[2].t7 Y[2].t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X180 VDD.t110 B[7].t6 a_14817_n474.t6 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X181 Y[2].t2 a_4048_215.t7 a_4475_n478.t6 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X182 VSS.t21 B[7].t7 a_15171_n1206.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X183 VSS.t2 B[2].t6 a_4829_n1210.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X184 VDD.t72 A[7].t7 a_14390_219.t1 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X185 a_14935_n1206.t0 a_15229_n500.t7 VSS.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X186 a_10798_n1206.t1 a_11092_n500.t7 VSS.t17 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X187 VDD.t169 B[2].t7 a_4887_n504.t3 VDD.t168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X188 a_11092_n500.t0 B[5].t7 VDD.t201 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X189 Y[4].t2 a_8185_217.t7 a_8730_n1208.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X190 Y[0].t3 a_n89_215.t7 a_456_n1210.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X191 a_9024_n502.t0 B[4].t7 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 a_6955_n502.n1 a_6955_n502.t5 318.922
R1 a_6955_n502.n0 a_6955_n502.t4 274.739
R2 a_6955_n502.n0 a_6955_n502.t7 274.739
R3 a_6955_n502.n1 a_6955_n502.t6 269.116
R4 a_6955_n502.t5 a_6955_n502.n0 179.946
R5 a_6955_n502.n2 a_6955_n502.n1 107.263
R6 a_6955_n502.n3 a_6955_n502.t3 29.444
R7 a_6955_n502.n4 a_6955_n502.t2 28.565
R8 a_6955_n502.t0 a_6955_n502.n4 28.565
R9 a_6955_n502.n2 a_6955_n502.t1 18.145
R10 a_6955_n502.n3 a_6955_n502.n2 2.878
R11 a_6955_n502.n4 a_6955_n502.n3 0.764
R12 Y[3].n7 Y[3].n6 194.965
R13 Y[3].n4 Y[3].n2 157.665
R14 Y[3].n4 Y[3].n3 122.999
R15 Y[3].n6 Y[3].n0 90.436
R16 Y[3].n5 Y[3].n1 90.416
R17 Y[3].n6 Y[3].n5 74.302
R18 Y[3].n5 Y[3].n4 50.575
R19 Y[3].n0 Y[3].t2 14.282
R20 Y[3].n0 Y[3].t0 14.282
R21 Y[3].n1 Y[3].t1 14.282
R22 Y[3].n1 Y[3].t7 14.282
R23 Y[3].n3 Y[3].t5 14.282
R24 Y[3].n3 Y[3].t3 14.282
R25 Y[3].n2 Y[3].t4 8.7
R26 Y[3].n2 Y[3].t6 8.7
R27 Y[3] Y[3].n7 0.03
R28 Y[3].n7 Y[3] 0.028
R29 a_6543_n476.n2 a_6543_n476.n0 267.767
R30 a_6543_n476.n6 a_6543_n476.t9 16.058
R31 a_6543_n476.n4 a_6543_n476.t4 16.058
R32 a_6543_n476.n5 a_6543_n476.t11 14.282
R33 a_6543_n476.n5 a_6543_n476.t10 14.282
R34 a_6543_n476.n3 a_6543_n476.t5 14.282
R35 a_6543_n476.n3 a_6543_n476.t6 14.282
R36 a_6543_n476.n1 a_6543_n476.t7 14.282
R37 a_6543_n476.n1 a_6543_n476.t2 14.282
R38 a_6543_n476.n0 a_6543_n476.t8 14.282
R39 a_6543_n476.n0 a_6543_n476.t3 14.282
R40 a_6543_n476.n9 a_6543_n476.t1 14.282
R41 a_6543_n476.t0 a_6543_n476.n9 14.282
R42 a_6543_n476.n9 a_6543_n476.n8 1.511
R43 a_6543_n476.n6 a_6543_n476.n5 0.999
R44 a_6543_n476.n4 a_6543_n476.n3 0.999
R45 a_6543_n476.n8 a_6543_n476.n2 0.669
R46 a_6543_n476.n7 a_6543_n476.n6 0.575
R47 a_6543_n476.n8 a_6543_n476.n7 0.227
R48 a_6543_n476.n7 a_6543_n476.n4 0.2
R49 a_6543_n476.n2 a_6543_n476.n1 0.001
R50 VDD.t180 VDD.t4 413.681
R51 VDD.t178 VDD.t90 413.681
R52 VDD.t172 VDD.t138 413.681
R53 VDD.t211 VDD.t111 413.681
R54 VDD.t205 VDD.t29 413.681
R55 VDD.t118 VDD.t120 413.681
R56 VDD.t218 VDD.t236 413.681
R57 VDD.t194 VDD.t87 413.681
R58 VDD.t132 VDD.t83 345.987
R59 VDD.t83 VDD.t113 345.987
R60 VDD.t168 VDD.t54 345.987
R61 VDD.t4 VDD.t168 345.987
R62 VDD.t94 VDD.t159 345.987
R63 VDD.t159 VDD.t150 345.987
R64 VDD.t140 VDD.t166 345.987
R65 VDD.t90 VDD.t140 345.987
R66 VDD.t39 VDD.t163 345.987
R67 VDD.t163 VDD.t56 345.987
R68 VDD.t48 VDD.t200 345.987
R69 VDD.t138 VDD.t48 345.987
R70 VDD.t20 VDD.t130 345.987
R71 VDD.t130 VDD.t71 345.987
R72 VDD.t134 VDD.t65 345.987
R73 VDD.t111 VDD.t134 345.987
R74 VDD.t174 VDD.t228 345.987
R75 VDD.t228 VDD.t232 345.987
R76 VDD.t202 VDD.t197 345.987
R77 VDD.t29 VDD.t202 345.987
R78 VDD.t92 VDD.t161 345.987
R79 VDD.t161 VDD.t78 345.987
R80 VDD.t85 VDD.t122 345.987
R81 VDD.t120 VDD.t85 345.987
R82 VDD.t62 VDD.t226 345.987
R83 VDD.t226 VDD.t44 345.987
R84 VDD.t127 VDD.t0 345.987
R85 VDD.t236 VDD.t127 345.987
R86 VDD.t148 VDD.t116 345.987
R87 VDD.t116 VDD.t216 345.987
R88 VDD.t42 VDD.t76 345.987
R89 VDD.t87 VDD.t42 345.987
R90 VDD.t96 VDD.t132 312.28
R91 VDD.t209 VDD.t94 312.28
R92 VDD.t165 VDD.t39 312.28
R93 VDD.t184 VDD.t20 312.28
R94 VDD.t80 VDD.t174 312.28
R95 VDD.t37 VDD.t92 312.28
R96 VDD.t185 VDD.t62 312.28
R97 VDD.t9 VDD.t148 312.28
R98 VDD.n149 VDD.t27 170.677
R99 VDD.n124 VDD.t176 170.677
R100 VDD.n45 VDD.t24 170.677
R101 VDD.n95 VDD.t109 170.677
R102 VDD.n20 VDD.t31 170.677
R103 VDD.n70 VDD.t182 170.677
R104 VDD.n174 VDD.t214 170.677
R105 VDD.n199 VDD.t60 170.677
R106 VDD.n150 VDD.n149 151.379
R107 VDD.n125 VDD.n124 151.379
R108 VDD.n46 VDD.n45 151.379
R109 VDD.n96 VDD.n95 151.379
R110 VDD.n21 VDD.n20 151.379
R111 VDD.n71 VDD.n70 151.379
R112 VDD.n175 VDD.n174 151.379
R113 VDD.n200 VDD.n199 151.379
R114 VDD.n149 VDD.n148 115.932
R115 VDD.n124 VDD.n123 115.932
R116 VDD.n45 VDD.n44 115.932
R117 VDD.n95 VDD.n94 115.932
R118 VDD.n20 VDD.n19 115.932
R119 VDD.n70 VDD.n69 115.932
R120 VDD.n174 VDD.n173 115.932
R121 VDD.n199 VDD.n198 115.932
R122 VDD.t11 VDD.t27 53.244
R123 VDD.t14 VDD.t96 53.244
R124 VDD.t75 VDD.t176 53.244
R125 VDD.t2 VDD.t209 53.244
R126 VDD.t144 VDD.t165 53.244
R127 VDD.t152 VDD.t184 53.244
R128 VDD.t224 VDD.t80 53.244
R129 VDD.t234 VDD.t37 53.244
R130 VDD.t154 VDD.t214 53.244
R131 VDD.t188 VDD.t185 53.244
R132 VDD.t155 VDD.t60 53.244
R133 VDD.t18 VDD.t9 53.244
R134 VDD.t102 VDD.n144 44.17
R135 VDD.t27 VDD.n145 44.17
R136 VDD.n147 VDD.t22 44.17
R137 VDD.n146 VDD.t14 44.17
R138 VDD.t50 VDD.n119 44.17
R139 VDD.t176 VDD.n120 44.17
R140 VDD.n122 VDD.t7 44.17
R141 VDD.n121 VDD.t2 44.17
R142 VDD.t136 VDD.n40 44.17
R143 VDD.t24 VDD.n41 44.17
R144 VDD.n43 VDD.t33 44.17
R145 VDD.n42 VDD.t144 44.17
R146 VDD.t68 VDD.n90 44.17
R147 VDD.t109 VDD.n91 44.17
R148 VDD.n93 VDD.t52 44.17
R149 VDD.n92 VDD.t152 44.17
R150 VDD.t207 VDD.n15 44.17
R151 VDD.t31 VDD.n16 44.17
R152 VDD.n18 VDD.t230 44.17
R153 VDD.n17 VDD.t224 44.17
R154 VDD.t99 VDD.n65 44.17
R155 VDD.t182 VDD.n66 44.17
R156 VDD.n68 VDD.t58 44.17
R157 VDD.n67 VDD.t234 44.17
R158 VDD.t157 VDD.n169 44.17
R159 VDD.t214 VDD.n170 44.17
R160 VDD.n172 VDD.t190 44.17
R161 VDD.n171 VDD.t188 44.17
R162 VDD.t192 VDD.n194 44.17
R163 VDD.t60 VDD.n195 44.17
R164 VDD.n197 VDD.t12 44.17
R165 VDD.n196 VDD.t18 44.17
R166 VDD.n145 VDD.t102 41.273
R167 VDD.t222 VDD.n147 41.273
R168 VDD.t22 VDD.n146 41.273
R169 VDD.n144 VDD.t180 41.273
R170 VDD.n120 VDD.t50 41.273
R171 VDD.t46 VDD.n122 41.273
R172 VDD.t7 VDD.n121 41.273
R173 VDD.n119 VDD.t178 41.273
R174 VDD.n41 VDD.t136 41.273
R175 VDD.t142 VDD.n43 41.273
R176 VDD.t33 VDD.n42 41.273
R177 VDD.n40 VDD.t172 41.273
R178 VDD.n91 VDD.t68 41.273
R179 VDD.t107 VDD.n93 41.273
R180 VDD.t52 VDD.n92 41.273
R181 VDD.n90 VDD.t211 41.273
R182 VDD.n16 VDD.t207 41.273
R183 VDD.t186 VDD.n18 41.273
R184 VDD.t230 VDD.n17 41.273
R185 VDD.n15 VDD.t205 41.273
R186 VDD.n66 VDD.t99 41.273
R187 VDD.t124 VDD.n68 41.273
R188 VDD.t58 VDD.n67 41.273
R189 VDD.n65 VDD.t118 41.273
R190 VDD.n170 VDD.t157 41.273
R191 VDD.t81 VDD.n172 41.273
R192 VDD.t190 VDD.n171 41.273
R193 VDD.n169 VDD.t218 41.273
R194 VDD.n195 VDD.t192 41.273
R195 VDD.t146 VDD.n197 41.273
R196 VDD.t12 VDD.n196 41.273
R197 VDD.n194 VDD.t194 41.273
R198 VDD.n148 VDD.t11 29.891
R199 VDD.n123 VDD.t75 29.891
R200 VDD.n44 VDD.t17 29.891
R201 VDD.n94 VDD.t6 29.891
R202 VDD.n19 VDD.t36 29.891
R203 VDD.n69 VDD.t156 29.891
R204 VDD.n173 VDD.t154 29.891
R205 VDD.n198 VDD.t155 29.891
R206 VDD.n131 VDD.t133 28.664
R207 VDD.n138 VDD.t5 28.664
R208 VDD.n106 VDD.t95 28.664
R209 VDD.n113 VDD.t91 28.664
R210 VDD.n35 VDD.t40 28.664
R211 VDD.n27 VDD.t139 28.664
R212 VDD.n85 VDD.t21 28.664
R213 VDD.n77 VDD.t112 28.664
R214 VDD.n10 VDD.t175 28.664
R215 VDD.n2 VDD.t30 28.664
R216 VDD.n60 VDD.t93 28.664
R217 VDD.n52 VDD.t121 28.664
R218 VDD.n156 VDD.t63 28.664
R219 VDD.n163 VDD.t237 28.664
R220 VDD.n181 VDD.t149 28.664
R221 VDD.n188 VDD.t88 28.664
R222 VDD.n132 VDD.t84 28.565
R223 VDD.n132 VDD.t114 28.565
R224 VDD.n139 VDD.t55 28.565
R225 VDD.n139 VDD.t169 28.565
R226 VDD.n107 VDD.t160 28.565
R227 VDD.n107 VDD.t151 28.565
R228 VDD.n114 VDD.t167 28.565
R229 VDD.n114 VDD.t141 28.565
R230 VDD.n36 VDD.t164 28.565
R231 VDD.n36 VDD.t57 28.565
R232 VDD.n28 VDD.t201 28.565
R233 VDD.n28 VDD.t49 28.565
R234 VDD.n86 VDD.t131 28.565
R235 VDD.n86 VDD.t72 28.565
R236 VDD.n78 VDD.t66 28.565
R237 VDD.n78 VDD.t135 28.565
R238 VDD.n11 VDD.t229 28.565
R239 VDD.n11 VDD.t233 28.565
R240 VDD.n3 VDD.t198 28.565
R241 VDD.n3 VDD.t203 28.565
R242 VDD.n61 VDD.t162 28.565
R243 VDD.n61 VDD.t79 28.565
R244 VDD.n53 VDD.t123 28.565
R245 VDD.n53 VDD.t86 28.565
R246 VDD.n157 VDD.t227 28.565
R247 VDD.n157 VDD.t45 28.565
R248 VDD.n164 VDD.t1 28.565
R249 VDD.n164 VDD.t128 28.565
R250 VDD.n182 VDD.t117 28.565
R251 VDD.n182 VDD.t217 28.565
R252 VDD.n189 VDD.t77 28.565
R253 VDD.n189 VDD.t43 28.565
R254 VDD.n148 VDD.t222 20.998
R255 VDD.n123 VDD.t46 20.998
R256 VDD.n44 VDD.t142 20.998
R257 VDD.n94 VDD.t107 20.998
R258 VDD.n19 VDD.t186 20.998
R259 VDD.n69 VDD.t124 20.998
R260 VDD.n173 VDD.t81 20.998
R261 VDD.n198 VDD.t146 20.998
R262 VDD.n131 VDD.t15 14.284
R263 VDD.n138 VDD.t181 14.284
R264 VDD.n106 VDD.t3 14.284
R265 VDD.n113 VDD.t179 14.284
R266 VDD.n35 VDD.t145 14.284
R267 VDD.n27 VDD.t173 14.284
R268 VDD.n85 VDD.t153 14.284
R269 VDD.n77 VDD.t212 14.284
R270 VDD.n10 VDD.t225 14.284
R271 VDD.n2 VDD.t206 14.284
R272 VDD.n60 VDD.t235 14.284
R273 VDD.n52 VDD.t119 14.284
R274 VDD.n156 VDD.t189 14.284
R275 VDD.n163 VDD.t219 14.284
R276 VDD.n181 VDD.t19 14.284
R277 VDD.n188 VDD.t195 14.284
R278 VDD.n130 VDD.t223 14.282
R279 VDD.n130 VDD.t23 14.282
R280 VDD.n137 VDD.t103 14.282
R281 VDD.n137 VDD.t28 14.282
R282 VDD.n105 VDD.t47 14.282
R283 VDD.n105 VDD.t8 14.282
R284 VDD.n112 VDD.t51 14.282
R285 VDD.n112 VDD.t177 14.282
R286 VDD.n34 VDD.t143 14.282
R287 VDD.n34 VDD.t34 14.282
R288 VDD.n26 VDD.t137 14.282
R289 VDD.n26 VDD.t25 14.282
R290 VDD.n84 VDD.t108 14.282
R291 VDD.n84 VDD.t53 14.282
R292 VDD.n76 VDD.t69 14.282
R293 VDD.n76 VDD.t110 14.282
R294 VDD.n9 VDD.t187 14.282
R295 VDD.n9 VDD.t231 14.282
R296 VDD.n1 VDD.t208 14.282
R297 VDD.n1 VDD.t32 14.282
R298 VDD.n59 VDD.t125 14.282
R299 VDD.n59 VDD.t59 14.282
R300 VDD.n51 VDD.t100 14.282
R301 VDD.n51 VDD.t183 14.282
R302 VDD.n155 VDD.t82 14.282
R303 VDD.n155 VDD.t191 14.282
R304 VDD.n162 VDD.t158 14.282
R305 VDD.n162 VDD.t215 14.282
R306 VDD.n180 VDD.t147 14.282
R307 VDD.n180 VDD.t13 14.282
R308 VDD.n187 VDD.t193 14.282
R309 VDD.n187 VDD.t61 14.282
R310 VDD.n153 VDD.n135 9.03
R311 VDD.n128 VDD.n110 9.03
R312 VDD.n178 VDD.n160 9.03
R313 VDD.n203 VDD.n185 9.03
R314 VDD.n142 VDD.n129 9
R315 VDD.n117 VDD.n104 9
R316 VDD.n167 VDD.n154 9
R317 VDD.n192 VDD.n179 9
R318 VDD.n144 VDD.t171 6.189
R319 VDD.n145 VDD.t26 6.189
R320 VDD.n147 VDD.t98 6.189
R321 VDD.n146 VDD.t97 6.189
R322 VDD.n119 VDD.t73 6.189
R323 VDD.n120 VDD.t74 6.189
R324 VDD.n122 VDD.t239 6.189
R325 VDD.n121 VDD.t238 6.189
R326 VDD.n40 VDD.t38 6.189
R327 VDD.n41 VDD.t16 6.189
R328 VDD.n43 VDD.t89 6.189
R329 VDD.n42 VDD.t129 6.189
R330 VDD.n90 VDD.t35 6.189
R331 VDD.n91 VDD.t41 6.189
R332 VDD.n93 VDD.t210 6.189
R333 VDD.n92 VDD.t67 6.189
R334 VDD.n15 VDD.t170 6.189
R335 VDD.n16 VDD.t199 6.189
R336 VDD.n18 VDD.t64 6.189
R337 VDD.n17 VDD.t104 6.189
R338 VDD.n65 VDD.t10 6.189
R339 VDD.n66 VDD.t115 6.189
R340 VDD.n68 VDD.t101 6.189
R341 VDD.n67 VDD.t204 6.189
R342 VDD.n169 VDD.t221 6.189
R343 VDD.n170 VDD.t220 6.189
R344 VDD.n172 VDD.t70 6.189
R345 VDD.n171 VDD.t106 6.189
R346 VDD.n194 VDD.t105 6.189
R347 VDD.n195 VDD.t196 6.189
R348 VDD.n197 VDD.t126 6.189
R349 VDD.n196 VDD.t213 6.189
R350 VDD.n133 VDD.n132 2.451
R351 VDD.n108 VDD.n107 2.451
R352 VDD.n37 VDD.n36 2.451
R353 VDD.n87 VDD.n86 2.451
R354 VDD.n12 VDD.n11 2.451
R355 VDD.n62 VDD.n61 2.451
R356 VDD.n158 VDD.n157 2.451
R357 VDD.n183 VDD.n182 2.451
R358 VDD.n140 VDD.n139 2.449
R359 VDD.n115 VDD.n114 2.449
R360 VDD.n29 VDD.n28 2.449
R361 VDD.n79 VDD.n78 2.449
R362 VDD.n4 VDD.n3 2.449
R363 VDD.n54 VDD.n53 2.449
R364 VDD.n165 VDD.n164 2.449
R365 VDD.n190 VDD.n189 2.449
R366 VDD.n204 VDD.n179 1.739
R367 VDD.n206 VDD.n129 1.738
R368 VDD.n207 VDD.n104 1.738
R369 VDD.n205 VDD.n154 1.738
R370 VDD.n134 VDD.n130 0.922
R371 VDD.n141 VDD.n137 0.922
R372 VDD.n109 VDD.n105 0.922
R373 VDD.n116 VDD.n112 0.922
R374 VDD.n38 VDD.n34 0.922
R375 VDD.n30 VDD.n26 0.922
R376 VDD.n88 VDD.n84 0.922
R377 VDD.n80 VDD.n76 0.922
R378 VDD.n13 VDD.n9 0.922
R379 VDD.n5 VDD.n1 0.922
R380 VDD.n63 VDD.n59 0.922
R381 VDD.n55 VDD.n51 0.922
R382 VDD.n159 VDD.n155 0.922
R383 VDD.n166 VDD.n162 0.922
R384 VDD.n184 VDD.n180 0.922
R385 VDD.n191 VDD.n187 0.922
R386 VDD.n133 VDD.n131 0.921
R387 VDD.n140 VDD.n138 0.921
R388 VDD.n108 VDD.n106 0.921
R389 VDD.n115 VDD.n113 0.921
R390 VDD.n37 VDD.n35 0.921
R391 VDD.n29 VDD.n27 0.921
R392 VDD.n87 VDD.n85 0.921
R393 VDD.n79 VDD.n77 0.921
R394 VDD.n12 VDD.n10 0.921
R395 VDD.n4 VDD.n2 0.921
R396 VDD.n62 VDD.n60 0.921
R397 VDD.n54 VDD.n52 0.921
R398 VDD.n158 VDD.n156 0.921
R399 VDD.n165 VDD.n163 0.921
R400 VDD.n183 VDD.n181 0.921
R401 VDD.n190 VDD.n188 0.921
R402 VDD.n134 VDD.n133 0.686
R403 VDD.n141 VDD.n140 0.686
R404 VDD.n109 VDD.n108 0.686
R405 VDD.n116 VDD.n115 0.686
R406 VDD.n38 VDD.n37 0.686
R407 VDD.n30 VDD.n29 0.686
R408 VDD.n88 VDD.n87 0.686
R409 VDD.n80 VDD.n79 0.686
R410 VDD.n13 VDD.n12 0.686
R411 VDD.n5 VDD.n4 0.686
R412 VDD.n63 VDD.n62 0.686
R413 VDD.n55 VDD.n54 0.686
R414 VDD.n159 VDD.n158 0.686
R415 VDD.n166 VDD.n165 0.686
R416 VDD.n184 VDD.n183 0.686
R417 VDD.n191 VDD.n190 0.686
R418 VDD.n101 VDD.n100 0.398
R419 VDD.n102 VDD.n101 0.398
R420 VDD.n103 VDD.n102 0.398
R421 VDD.n207 VDD.n206 0.398
R422 VDD.n206 VDD.n205 0.398
R423 VDD.n205 VDD.n204 0.398
R424 VDD VDD.n103 0.205
R425 VDD.n135 VDD.n134 0.193
R426 VDD.n110 VDD.n109 0.193
R427 VDD.n39 VDD.n38 0.193
R428 VDD.n89 VDD.n88 0.193
R429 VDD.n14 VDD.n13 0.193
R430 VDD.n64 VDD.n63 0.193
R431 VDD.n160 VDD.n159 0.193
R432 VDD.n185 VDD.n184 0.193
R433 VDD.n142 VDD.n141 0.189
R434 VDD.n117 VDD.n116 0.189
R435 VDD.n31 VDD.n30 0.189
R436 VDD.n81 VDD.n80 0.189
R437 VDD.n6 VDD.n5 0.189
R438 VDD.n56 VDD.n55 0.189
R439 VDD.n167 VDD.n166 0.189
R440 VDD.n192 VDD.n191 0.189
R441 VDD VDD.n207 0.154
R442 VDD.n136 VDD.n129 0.03
R443 VDD.n111 VDD.n104 0.03
R444 VDD.n33 VDD.n25 0.03
R445 VDD.n83 VDD.n75 0.03
R446 VDD.n8 VDD.n0 0.03
R447 VDD.n58 VDD.n50 0.03
R448 VDD.n161 VDD.n154 0.03
R449 VDD.n186 VDD.n179 0.03
R450 VDD.n143 VDD.n142 0.021
R451 VDD.n151 VDD.n135 0.021
R452 VDD.n118 VDD.n117 0.021
R453 VDD.n126 VDD.n110 0.021
R454 VDD.n32 VDD.n31 0.021
R455 VDD.n47 VDD.n39 0.021
R456 VDD.n82 VDD.n81 0.021
R457 VDD.n97 VDD.n89 0.021
R458 VDD.n7 VDD.n6 0.021
R459 VDD.n22 VDD.n14 0.021
R460 VDD.n57 VDD.n56 0.021
R461 VDD.n72 VDD.n64 0.021
R462 VDD.n168 VDD.n167 0.021
R463 VDD.n176 VDD.n160 0.021
R464 VDD.n193 VDD.n192 0.021
R465 VDD.n201 VDD.n185 0.021
R466 VDD.n151 VDD.n150 0.002
R467 VDD.n126 VDD.n125 0.002
R468 VDD.n47 VDD.n46 0.002
R469 VDD.n97 VDD.n96 0.002
R470 VDD.n22 VDD.n21 0.002
R471 VDD.n72 VDD.n71 0.002
R472 VDD.n176 VDD.n175 0.002
R473 VDD.n152 VDD.n136 0.002
R474 VDD.n127 VDD.n111 0.002
R475 VDD.n48 VDD.n33 0.002
R476 VDD.n98 VDD.n83 0.002
R477 VDD.n23 VDD.n8 0.002
R478 VDD.n73 VDD.n58 0.002
R479 VDD.n177 VDD.n161 0.002
R480 VDD.n202 VDD.n186 0.002
R481 VDD.n152 VDD.n151 0.002
R482 VDD.n127 VDD.n126 0.002
R483 VDD.n48 VDD.n47 0.002
R484 VDD.n98 VDD.n97 0.002
R485 VDD.n23 VDD.n22 0.002
R486 VDD.n73 VDD.n72 0.002
R487 VDD.n177 VDD.n176 0.002
R488 VDD.n201 VDD.n200 0.001
R489 VDD.n143 VDD.n136 0.001
R490 VDD.n118 VDD.n111 0.001
R491 VDD.n33 VDD.n32 0.001
R492 VDD.n83 VDD.n82 0.001
R493 VDD.n8 VDD.n7 0.001
R494 VDD.n58 VDD.n57 0.001
R495 VDD.n168 VDD.n161 0.001
R496 VDD.n193 VDD.n186 0.001
R497 VDD.n202 VDD.n201 0.001
R498 VDD.n153 VDD.n152 0.001
R499 VDD.n128 VDD.n127 0.001
R500 VDD.n49 VDD.n48 0.001
R501 VDD.n99 VDD.n98 0.001
R502 VDD.n24 VDD.n23 0.001
R503 VDD.n74 VDD.n73 0.001
R504 VDD.n178 VDD.n177 0.001
R505 VDD.n203 VDD.n202 0.001
R506 VDD.n206 VDD.n153 0.001
R507 VDD.n207 VDD.n128 0.001
R508 VDD.n102 VDD.n49 0.001
R509 VDD.n100 VDD.n99 0.001
R510 VDD.n103 VDD.n24 0.001
R511 VDD.n101 VDD.n74 0.001
R512 VDD.n205 VDD.n178 0.001
R513 VDD.n204 VDD.n203 0.001
R514 VDD.n150 VDD.n143 0.001
R515 VDD.n125 VDD.n118 0.001
R516 VDD.n175 VDD.n168 0.001
R517 VDD.n200 VDD.n193 0.001
R518 A[2].n5 A[2].n4 412.11
R519 A[2].n1 A[2].t1 394.151
R520 A[2].n4 A[2].t7 294.653
R521 A[2].n0 A[2].t0 269.523
R522 A[2].t1 A[2].n0 269.523
R523 A[2].n5 A[2].n3 224.13
R524 A[2].n2 A[2].t6 198.043
R525 A[2].n0 A[2].t3 160.666
R526 A[2] A[2].n5 138.225
R527 A[2].n4 A[2].t2 111.663
R528 A[2].n3 A[2].n1 97.816
R529 A[2].n2 A[2].t5 93.989
R530 A[2].n1 A[2].t4 80.333
R531 A[2].n3 A[2].n2 6.615
R532 a_4475_n478.n2 a_4475_n478.n0 267.767
R533 a_4475_n478.n6 a_4475_n478.t6 16.058
R534 a_4475_n478.n8 a_4475_n478.t10 16.058
R535 a_4475_n478.n1 a_4475_n478.t2 14.282
R536 a_4475_n478.n1 a_4475_n478.t5 14.282
R537 a_4475_n478.n0 a_4475_n478.t11 14.282
R538 a_4475_n478.n0 a_4475_n478.t9 14.282
R539 a_4475_n478.n3 a_4475_n478.t3 14.282
R540 a_4475_n478.n3 a_4475_n478.t4 14.282
R541 a_4475_n478.n5 a_4475_n478.t8 14.282
R542 a_4475_n478.n5 a_4475_n478.t7 14.282
R543 a_4475_n478.n9 a_4475_n478.t1 14.282
R544 a_4475_n478.t0 a_4475_n478.n9 14.282
R545 a_4475_n478.n4 a_4475_n478.n3 1.511
R546 a_4475_n478.n6 a_4475_n478.n5 0.999
R547 a_4475_n478.n9 a_4475_n478.n8 0.999
R548 a_4475_n478.n4 a_4475_n478.n2 0.669
R549 a_4475_n478.n7 a_4475_n478.n6 0.575
R550 a_4475_n478.n7 a_4475_n478.n4 0.227
R551 a_4475_n478.n8 a_4475_n478.n7 0.2
R552 a_4475_n478.n2 a_4475_n478.n1 0.001
R553 A[0].n5 A[0].n4 412.11
R554 A[0].n1 A[0].t5 394.151
R555 A[0].n4 A[0].t0 294.653
R556 A[0].n0 A[0].t2 269.523
R557 A[0].t5 A[0].n0 269.523
R558 A[0].n5 A[0].n3 224.13
R559 A[0].n2 A[0].t6 198.043
R560 A[0].n0 A[0].t3 160.666
R561 A[0] A[0].n5 138.23
R562 A[0].n4 A[0].t4 111.663
R563 A[0].n3 A[0].n1 97.816
R564 A[0].n2 A[0].t1 93.989
R565 A[0].n1 A[0].t7 80.333
R566 A[0].n3 A[0].n2 6.615
R567 Y[0].n7 Y[0].n6 194.965
R568 Y[0].n4 Y[0].n2 157.665
R569 Y[0].n4 Y[0].n3 122.999
R570 Y[0].n6 Y[0].n0 90.436
R571 Y[0].n5 Y[0].n1 90.416
R572 Y[0].n6 Y[0].n5 74.302
R573 Y[0].n5 Y[0].n4 50.575
R574 Y[0].n0 Y[0].t2 14.282
R575 Y[0].n0 Y[0].t6 14.282
R576 Y[0].n1 Y[0].t5 14.282
R577 Y[0].n1 Y[0].t4 14.282
R578 Y[0].n3 Y[0].t7 14.282
R579 Y[0].n3 Y[0].t0 14.282
R580 Y[0].n2 Y[0].t1 8.7
R581 Y[0].n2 Y[0].t3 8.7
R582 Y[0] Y[0].n7 0.034
R583 Y[0].n7 Y[0] 0.024
R584 a_692_n1210.t0 a_692_n1210.t1 17.4
R585 VSS.n16 VSS.t18 20.763
R586 VSS.n18 VSS.t3 20.763
R587 VSS.n20 VSS.t15 20.763
R588 VSS.n22 VSS.t26 20.763
R589 VSS.n1 VSS.t28 20.763
R590 VSS.n3 VSS.t9 20.763
R591 VSS.n5 VSS.t12 20.763
R592 VSS.n7 VSS.t16 20.763
R593 VSS.n23 VSS.t8 20.676
R594 VSS.n28 VSS.t25 20.676
R595 VSS.n26 VSS.t11 20.676
R596 VSS.n24 VSS.t5 20.676
R597 VSS.n14 VSS.t6 20.676
R598 VSS.n12 VSS.t10 20.676
R599 VSS.n10 VSS.t19 20.676
R600 VSS.n8 VSS.t22 20.676
R601 VSS.n15 VSS.t7 8.7
R602 VSS.n15 VSS.t23 8.7
R603 VSS.n17 VSS.t24 8.7
R604 VSS.n17 VSS.t2 8.7
R605 VSS.n19 VSS.t30 8.7
R606 VSS.n19 VSS.t31 8.7
R607 VSS.n21 VSS.t20 8.7
R608 VSS.n21 VSS.t27 8.7
R609 VSS.n0 VSS.t0 8.7
R610 VSS.n0 VSS.t29 8.7
R611 VSS.n2 VSS.t17 8.7
R612 VSS.n2 VSS.t1 8.7
R613 VSS.n4 VSS.t13 8.7
R614 VSS.n4 VSS.t14 8.7
R615 VSS.n6 VSS.t4 8.7
R616 VSS.n6 VSS.t21 8.7
R617 VSS.n16 VSS.n15 0.948
R618 VSS.n18 VSS.n17 0.948
R619 VSS.n20 VSS.n19 0.948
R620 VSS.n22 VSS.n21 0.948
R621 VSS.n1 VSS.n0 0.948
R622 VSS.n3 VSS.n2 0.948
R623 VSS.n5 VSS.n4 0.948
R624 VSS.n7 VSS.n6 0.948
R625 VSS.n26 VSS.n25 0.511
R626 VSS.n24 VSS.n23 0.51
R627 VSS.n28 VSS.n27 0.51
R628 VSS.n9 VSS.n8 0.506
R629 VSS.n13 VSS.n12 0.506
R630 VSS.n11 VSS.n10 0.506
R631 VSS VSS.n14 0.249
R632 VSS VSS.n29 0.21
R633 VSS.n8 VSS.n7 0.196
R634 VSS.n29 VSS.n16 0.196
R635 VSS.n27 VSS.n18 0.196
R636 VSS.n25 VSS.n20 0.196
R637 VSS.n23 VSS.n22 0.196
R638 VSS.n13 VSS.n1 0.196
R639 VSS.n11 VSS.n3 0.196
R640 VSS.n9 VSS.n5 0.196
R641 VSS.n25 VSS.n24 0.001
R642 VSS.n27 VSS.n26 0.001
R643 VSS.n29 VSS.n28 0.001
R644 VSS.n10 VSS.n9 0.001
R645 VSS.n14 VSS.n13 0.001
R646 VSS.n12 VSS.n11 0.001
R647 B[1].n4 B[1].n3 592.056
R648 B[1].t0 B[1].n1 313.873
R649 B[1].n3 B[1].t5 294.986
R650 B[1].n0 B[1].t4 272.288
R651 B[1].n4 B[1].t6 204.68
R652 B[1].n2 B[1].t0 190.152
R653 B[1].n2 B[1].t3 190.152
R654 B[1].n0 B[1].t2 160.666
R655 B[1].n1 B[1].t1 160.666
R656 B[1].n3 B[1].t7 110.859
R657 B[1].n1 B[1].n0 96.129
R658 B[1].t6 B[1].n2 80.333
R659 B[1] B[1].n4 42.781
R660 a_2818_n502.n1 a_2818_n502.t5 318.922
R661 a_2818_n502.n0 a_2818_n502.t4 274.739
R662 a_2818_n502.n0 a_2818_n502.t6 274.739
R663 a_2818_n502.n1 a_2818_n502.t7 269.116
R664 a_2818_n502.t5 a_2818_n502.n0 179.946
R665 a_2818_n502.n2 a_2818_n502.n1 107.263
R666 a_2818_n502.n3 a_2818_n502.t1 29.444
R667 a_2818_n502.n4 a_2818_n502.t0 28.565
R668 a_2818_n502.t2 a_2818_n502.n4 28.565
R669 a_2818_n502.n2 a_2818_n502.t3 18.145
R670 a_2818_n502.n3 a_2818_n502.n2 2.878
R671 a_2818_n502.n4 a_2818_n502.n3 0.764
R672 a_n89_215.n1 a_n89_215.t4 318.922
R673 a_n89_215.n0 a_n89_215.t5 273.935
R674 a_n89_215.n0 a_n89_215.t6 273.935
R675 a_n89_215.n1 a_n89_215.t7 269.116
R676 a_n89_215.n4 a_n89_215.n3 193.227
R677 a_n89_215.t4 a_n89_215.n0 179.142
R678 a_n89_215.n2 a_n89_215.n1 106.999
R679 a_n89_215.n3 a_n89_215.t1 28.568
R680 a_n89_215.n4 a_n89_215.t0 28.565
R681 a_n89_215.t2 a_n89_215.n4 28.565
R682 a_n89_215.n2 a_n89_215.t3 18.149
R683 a_n89_215.n3 a_n89_215.n2 3.726
R684 a_338_n478.n8 a_338_n478.n0 267.767
R685 a_338_n478.n4 a_338_n478.t5 16.058
R686 a_338_n478.n2 a_338_n478.t7 16.058
R687 a_338_n478.n3 a_338_n478.t4 14.282
R688 a_338_n478.n3 a_338_n478.t6 14.282
R689 a_338_n478.n1 a_338_n478.t11 14.282
R690 a_338_n478.n1 a_338_n478.t8 14.282
R691 a_338_n478.n6 a_338_n478.t2 14.282
R692 a_338_n478.n6 a_338_n478.t1 14.282
R693 a_338_n478.n0 a_338_n478.t10 14.282
R694 a_338_n478.n0 a_338_n478.t9 14.282
R695 a_338_n478.t0 a_338_n478.n9 14.282
R696 a_338_n478.n9 a_338_n478.t3 14.282
R697 a_338_n478.n7 a_338_n478.n6 1.511
R698 a_338_n478.n4 a_338_n478.n3 0.999
R699 a_338_n478.n2 a_338_n478.n1 0.999
R700 a_338_n478.n8 a_338_n478.n7 0.669
R701 a_338_n478.n5 a_338_n478.n4 0.575
R702 a_338_n478.n7 a_338_n478.n5 0.227
R703 a_338_n478.n5 a_338_n478.n2 0.2
R704 a_338_n478.n9 a_338_n478.n8 0.001
R705 A[6].n5 A[6].n4 412.11
R706 A[6].n1 A[6].t3 394.151
R707 A[6].n4 A[6].t1 294.653
R708 A[6].n0 A[6].t0 269.523
R709 A[6].t3 A[6].n0 269.523
R710 A[6].n5 A[6].n3 224.13
R711 A[6].n2 A[6].t6 198.043
R712 A[6].n0 A[6].t2 160.666
R713 A[6] A[6].n5 138.229
R714 A[6].n4 A[6].t7 111.663
R715 A[6].n3 A[6].n1 97.816
R716 A[6].n2 A[6].t4 93.989
R717 A[6].n1 A[6].t5 80.333
R718 A[6].n3 A[6].n2 6.615
R719 a_12749_n476.n3 a_12749_n476.n1 267.767
R720 a_12749_n476.n7 a_12749_n476.t1 16.058
R721 a_12749_n476.t0 a_12749_n476.n9 16.058
R722 a_12749_n476.n2 a_12749_n476.t10 14.282
R723 a_12749_n476.n2 a_12749_n476.t4 14.282
R724 a_12749_n476.n1 a_12749_n476.t8 14.282
R725 a_12749_n476.n1 a_12749_n476.t5 14.282
R726 a_12749_n476.n4 a_12749_n476.t3 14.282
R727 a_12749_n476.n4 a_12749_n476.t2 14.282
R728 a_12749_n476.n6 a_12749_n476.t6 14.282
R729 a_12749_n476.n6 a_12749_n476.t11 14.282
R730 a_12749_n476.n0 a_12749_n476.t7 14.282
R731 a_12749_n476.n0 a_12749_n476.t9 14.282
R732 a_12749_n476.n5 a_12749_n476.n4 1.511
R733 a_12749_n476.n7 a_12749_n476.n6 0.999
R734 a_12749_n476.n9 a_12749_n476.n0 0.999
R735 a_12749_n476.n5 a_12749_n476.n3 0.669
R736 a_12749_n476.n8 a_12749_n476.n7 0.575
R737 a_12749_n476.n8 a_12749_n476.n5 0.227
R738 a_12749_n476.n9 a_12749_n476.n8 0.2
R739 a_12749_n476.n3 a_12749_n476.n2 0.001
R740 a_4048_215.n1 a_4048_215.t5 318.922
R741 a_4048_215.n0 a_4048_215.t7 273.935
R742 a_4048_215.n0 a_4048_215.t4 273.935
R743 a_4048_215.n1 a_4048_215.t6 269.116
R744 a_4048_215.n4 a_4048_215.n3 193.227
R745 a_4048_215.t5 a_4048_215.n0 179.142
R746 a_4048_215.n2 a_4048_215.n1 106.999
R747 a_4048_215.n3 a_4048_215.t0 28.568
R748 a_4048_215.t2 a_4048_215.n4 28.565
R749 a_4048_215.n4 a_4048_215.t1 28.565
R750 a_4048_215.n2 a_4048_215.t3 18.149
R751 a_4048_215.n3 a_4048_215.n2 3.726
R752 Y[2].n7 Y[2].n6 194.965
R753 Y[2].n4 Y[2].n2 157.665
R754 Y[2].n4 Y[2].n3 122.999
R755 Y[2].n6 Y[2].n0 90.436
R756 Y[2].n5 Y[2].n1 90.416
R757 Y[2].n6 Y[2].n5 74.302
R758 Y[2].n5 Y[2].n4 50.575
R759 Y[2].n0 Y[2].t7 14.282
R760 Y[2].n0 Y[2].t1 14.282
R761 Y[2].n1 Y[2].t0 14.282
R762 Y[2].n1 Y[2].t4 14.282
R763 Y[2].n3 Y[2].t3 14.282
R764 Y[2].n3 Y[2].t2 14.282
R765 Y[2].n2 Y[2].t6 8.7
R766 Y[2].n2 Y[2].t5 8.7
R767 Y[2] Y[2].n7 0.036
R768 Y[2].n7 Y[2] 0.022
R769 B[6].n4 B[6].n3 592.056
R770 B[6].t4 B[6].n1 313.873
R771 B[6].n3 B[6].t2 294.986
R772 B[6].n0 B[6].t7 272.288
R773 B[6].n4 B[6].t3 204.68
R774 B[6].n2 B[6].t4 190.152
R775 B[6].n2 B[6].t1 190.152
R776 B[6].n0 B[6].t6 160.666
R777 B[6].n1 B[6].t5 160.666
R778 B[6].n3 B[6].t0 110.859
R779 B[6].n1 B[6].n0 96.129
R780 B[6].t3 B[6].n2 80.333
R781 B[6] B[6].n4 42.783
R782 a_13161_n502.n1 a_13161_n502.t4 318.922
R783 a_13161_n502.n0 a_13161_n502.t6 274.739
R784 a_13161_n502.n0 a_13161_n502.t7 274.739
R785 a_13161_n502.n1 a_13161_n502.t5 269.116
R786 a_13161_n502.t4 a_13161_n502.n0 179.946
R787 a_13161_n502.n2 a_13161_n502.n1 107.263
R788 a_13161_n502.t2 a_13161_n502.n4 29.444
R789 a_13161_n502.n3 a_13161_n502.t1 28.565
R790 a_13161_n502.n3 a_13161_n502.t0 28.565
R791 a_13161_n502.n2 a_13161_n502.t3 18.145
R792 a_13161_n502.n4 a_13161_n502.n2 2.878
R793 a_13161_n502.n4 a_13161_n502.n3 0.764
R794 B[7].n4 B[7].n3 592.056
R795 B[7].t4 B[7].n1 313.873
R796 B[7].n3 B[7].t7 294.986
R797 B[7].n0 B[7].t6 272.288
R798 B[7].n4 B[7].t3 204.68
R799 B[7].n2 B[7].t4 190.152
R800 B[7].n2 B[7].t1 190.152
R801 B[7].n0 B[7].t0 160.666
R802 B[7].n1 B[7].t5 160.666
R803 B[7].n3 B[7].t2 110.859
R804 B[7].n1 B[7].n0 96.129
R805 B[7].t3 B[7].n2 80.333
R806 B[7] B[7].n4 42.78
R807 a_14817_n474.n2 a_14817_n474.n0 267.767
R808 a_14817_n474.n6 a_14817_n474.t10 16.058
R809 a_14817_n474.n8 a_14817_n474.t1 16.058
R810 a_14817_n474.n1 a_14817_n474.t6 14.282
R811 a_14817_n474.n1 a_14817_n474.t5 14.282
R812 a_14817_n474.n0 a_14817_n474.t7 14.282
R813 a_14817_n474.n0 a_14817_n474.t8 14.282
R814 a_14817_n474.n3 a_14817_n474.t3 14.282
R815 a_14817_n474.n3 a_14817_n474.t9 14.282
R816 a_14817_n474.n5 a_14817_n474.t11 14.282
R817 a_14817_n474.n5 a_14817_n474.t4 14.282
R818 a_14817_n474.n9 a_14817_n474.t2 14.282
R819 a_14817_n474.t0 a_14817_n474.n9 14.282
R820 a_14817_n474.n4 a_14817_n474.n3 1.511
R821 a_14817_n474.n6 a_14817_n474.n5 0.999
R822 a_14817_n474.n9 a_14817_n474.n8 0.999
R823 a_14817_n474.n4 a_14817_n474.n2 0.669
R824 a_14817_n474.n7 a_14817_n474.n6 0.575
R825 a_14817_n474.n7 a_14817_n474.n4 0.227
R826 a_14817_n474.n8 a_14817_n474.n7 0.2
R827 a_14817_n474.n2 a_14817_n474.n1 0.001
R828 A[4].n5 A[4].n4 412.11
R829 A[4].n1 A[4].t2 394.151
R830 A[4].n4 A[4].t4 294.653
R831 A[4].n0 A[4].t7 269.523
R832 A[4].t2 A[4].n0 269.523
R833 A[4].n5 A[4].n3 224.13
R834 A[4].n2 A[4].t6 198.043
R835 A[4].n0 A[4].t0 160.666
R836 A[4] A[4].n5 138.227
R837 A[4].n4 A[4].t5 111.663
R838 A[4].n3 A[4].n1 97.816
R839 A[4].n2 A[4].t3 93.989
R840 A[4].n1 A[4].t1 80.333
R841 A[4].n3 A[4].n2 6.615
R842 a_8612_n476.n8 a_8612_n476.n0 267.767
R843 a_8612_n476.n4 a_8612_n476.t3 16.058
R844 a_8612_n476.n2 a_8612_n476.t8 16.058
R845 a_8612_n476.n3 a_8612_n476.t2 14.282
R846 a_8612_n476.n3 a_8612_n476.t7 14.282
R847 a_8612_n476.n1 a_8612_n476.t9 14.282
R848 a_8612_n476.n1 a_8612_n476.t1 14.282
R849 a_8612_n476.n6 a_8612_n476.t6 14.282
R850 a_8612_n476.n6 a_8612_n476.t5 14.282
R851 a_8612_n476.n0 a_8612_n476.t10 14.282
R852 a_8612_n476.n0 a_8612_n476.t11 14.282
R853 a_8612_n476.t0 a_8612_n476.n9 14.282
R854 a_8612_n476.n9 a_8612_n476.t4 14.282
R855 a_8612_n476.n7 a_8612_n476.n6 1.511
R856 a_8612_n476.n4 a_8612_n476.n3 0.999
R857 a_8612_n476.n2 a_8612_n476.n1 0.999
R858 a_8612_n476.n8 a_8612_n476.n7 0.669
R859 a_8612_n476.n5 a_8612_n476.n4 0.575
R860 a_8612_n476.n7 a_8612_n476.n5 0.227
R861 a_8612_n476.n5 a_8612_n476.n2 0.2
R862 a_8612_n476.n9 a_8612_n476.n8 0.001
R863 B[0].n4 B[0].n3 592.056
R864 B[0].t6 B[0].n1 313.873
R865 B[0].n3 B[0].t0 294.986
R866 B[0].n0 B[0].t3 272.288
R867 B[0].n4 B[0].t7 204.68
R868 B[0].n2 B[0].t6 190.152
R869 B[0].n2 B[0].t5 190.152
R870 B[0].n0 B[0].t2 160.666
R871 B[0].n1 B[0].t1 160.666
R872 B[0].n3 B[0].t4 110.859
R873 B[0].n1 B[0].n0 96.129
R874 B[0].t7 B[0].n2 80.333
R875 B[0] B[0].n4 42.781
R876 Y[1].n7 Y[1].n6 194.965
R877 Y[1].n4 Y[1].n2 157.665
R878 Y[1].n4 Y[1].n3 122.999
R879 Y[1].n6 Y[1].n0 90.436
R880 Y[1].n5 Y[1].n1 90.416
R881 Y[1].n6 Y[1].n5 74.302
R882 Y[1].n5 Y[1].n4 50.575
R883 Y[1].n0 Y[1].t3 14.282
R884 Y[1].n0 Y[1].t5 14.282
R885 Y[1].n1 Y[1].t4 14.282
R886 Y[1].n1 Y[1].t1 14.282
R887 Y[1].n3 Y[1].t6 14.282
R888 Y[1].n3 Y[1].t7 14.282
R889 Y[1].n2 Y[1].t2 8.7
R890 Y[1].n2 Y[1].t0 8.7
R891 Y[1] Y[1].n7 0.034
R892 Y[1].n7 Y[1] 0.024
R893 a_2406_n476.n2 a_2406_n476.n0 267.767
R894 a_2406_n476.n8 a_2406_n476.t9 16.058
R895 a_2406_n476.n6 a_2406_n476.t5 16.058
R896 a_2406_n476.n1 a_2406_n476.t2 14.282
R897 a_2406_n476.n1 a_2406_n476.t1 14.282
R898 a_2406_n476.n0 a_2406_n476.t4 14.282
R899 a_2406_n476.n0 a_2406_n476.t3 14.282
R900 a_2406_n476.n3 a_2406_n476.t11 14.282
R901 a_2406_n476.n3 a_2406_n476.t10 14.282
R902 a_2406_n476.n5 a_2406_n476.t6 14.282
R903 a_2406_n476.n5 a_2406_n476.t7 14.282
R904 a_2406_n476.t0 a_2406_n476.n9 14.282
R905 a_2406_n476.n9 a_2406_n476.t8 14.282
R906 a_2406_n476.n4 a_2406_n476.n3 1.511
R907 a_2406_n476.n6 a_2406_n476.n5 0.999
R908 a_2406_n476.n9 a_2406_n476.n8 0.999
R909 a_2406_n476.n4 a_2406_n476.n2 0.669
R910 a_2406_n476.n8 a_2406_n476.n7 0.575
R911 a_2406_n476.n7 a_2406_n476.n4 0.227
R912 a_2406_n476.n7 a_2406_n476.n6 0.2
R913 a_2406_n476.n2 a_2406_n476.n1 0.001
R914 a_14390_219.n1 a_14390_219.t7 318.922
R915 a_14390_219.n0 a_14390_219.t4 273.935
R916 a_14390_219.n0 a_14390_219.t6 273.935
R917 a_14390_219.n1 a_14390_219.t5 269.116
R918 a_14390_219.n4 a_14390_219.n3 193.227
R919 a_14390_219.t7 a_14390_219.n0 179.142
R920 a_14390_219.n2 a_14390_219.n1 106.999
R921 a_14390_219.n3 a_14390_219.t1 28.568
R922 a_14390_219.t0 a_14390_219.n4 28.565
R923 a_14390_219.n4 a_14390_219.t2 28.565
R924 a_14390_219.n2 a_14390_219.t3 18.149
R925 a_14390_219.n3 a_14390_219.n2 3.726
R926 Y[7].n7 Y[7].n6 194.965
R927 Y[7].n4 Y[7].n2 157.665
R928 Y[7].n4 Y[7].n3 122.999
R929 Y[7].n6 Y[7].n0 90.436
R930 Y[7].n5 Y[7].n1 90.416
R931 Y[7].n6 Y[7].n5 74.302
R932 Y[7].n5 Y[7].n4 50.575
R933 Y[7].n0 Y[7].t1 14.282
R934 Y[7].n0 Y[7].t2 14.282
R935 Y[7].n1 Y[7].t0 14.282
R936 Y[7].n1 Y[7].t6 14.282
R937 Y[7].n3 Y[7].t5 14.282
R938 Y[7].n3 Y[7].t7 14.282
R939 Y[7].n2 Y[7].t3 8.7
R940 Y[7].n2 Y[7].t4 8.7
R941 Y[7] Y[7].n7 0.038
R942 Y[7].n7 Y[7] 0.02
R943 A[1].n5 A[1].n4 412.11
R944 A[1].n1 A[1].t2 394.151
R945 A[1].n4 A[1].t4 294.653
R946 A[1].n0 A[1].t7 269.523
R947 A[1].t2 A[1].n0 269.523
R948 A[1].n5 A[1].n3 224.13
R949 A[1].n2 A[1].t5 198.043
R950 A[1].n0 A[1].t0 160.666
R951 A[1] A[1].n5 138.227
R952 A[1].n4 A[1].t6 111.663
R953 A[1].n3 A[1].n1 97.816
R954 A[1].n2 A[1].t3 93.989
R955 A[1].n1 A[1].t1 80.333
R956 A[1].n3 A[1].n2 6.615
R957 A[3].n5 A[3].n4 412.11
R958 A[3].n1 A[3].t2 394.151
R959 A[3].n4 A[3].t3 294.653
R960 A[3].n0 A[3].t0 269.523
R961 A[3].t2 A[3].n0 269.523
R962 A[3].n5 A[3].n3 224.13
R963 A[3].n2 A[3].t7 198.043
R964 A[3].n0 A[3].t1 160.666
R965 A[3] A[3].n5 138.229
R966 A[3].n4 A[3].t5 111.663
R967 A[3].n3 A[3].n1 97.816
R968 A[3].n2 A[3].t4 93.989
R969 A[3].n1 A[3].t6 80.333
R970 A[3].n3 A[3].n2 6.615
R971 a_8185_217.n1 a_8185_217.t6 318.922
R972 a_8185_217.n0 a_8185_217.t5 273.935
R973 a_8185_217.n0 a_8185_217.t4 273.935
R974 a_8185_217.n1 a_8185_217.t7 269.116
R975 a_8185_217.n4 a_8185_217.n3 193.227
R976 a_8185_217.t6 a_8185_217.n0 179.142
R977 a_8185_217.n2 a_8185_217.n1 106.999
R978 a_8185_217.n3 a_8185_217.t0 28.568
R979 a_8185_217.t2 a_8185_217.n4 28.565
R980 a_8185_217.n4 a_8185_217.t1 28.565
R981 a_8185_217.n2 a_8185_217.t3 18.149
R982 a_8185_217.n3 a_8185_217.n2 3.726
R983 Y[4].n7 Y[4].n6 194.965
R984 Y[4].n4 Y[4].n2 157.665
R985 Y[4].n4 Y[4].n3 122.999
R986 Y[4].n6 Y[4].n0 90.436
R987 Y[4].n5 Y[4].n1 90.416
R988 Y[4].n6 Y[4].n5 74.302
R989 Y[4].n5 Y[4].n4 50.575
R990 Y[4].n0 Y[4].t6 14.282
R991 Y[4].n0 Y[4].t7 14.282
R992 Y[4].n1 Y[4].t0 14.282
R993 Y[4].n1 Y[4].t5 14.282
R994 Y[4].n3 Y[4].t3 14.282
R995 Y[4].n3 Y[4].t4 14.282
R996 Y[4].n2 Y[4].t1 8.7
R997 Y[4].n2 Y[4].t2 8.7
R998 Y[4] Y[4].n7 0.038
R999 Y[4].n7 Y[4] 0.02
R1000 a_9024_n502.n1 a_9024_n502.t7 318.922
R1001 a_9024_n502.n0 a_9024_n502.t4 274.739
R1002 a_9024_n502.n0 a_9024_n502.t6 274.739
R1003 a_9024_n502.n1 a_9024_n502.t5 269.116
R1004 a_9024_n502.t7 a_9024_n502.n0 179.946
R1005 a_9024_n502.n2 a_9024_n502.n1 107.263
R1006 a_9024_n502.n3 a_9024_n502.t2 29.444
R1007 a_9024_n502.n4 a_9024_n502.t3 28.565
R1008 a_9024_n502.t0 a_9024_n502.n4 28.565
R1009 a_9024_n502.n2 a_9024_n502.t1 18.145
R1010 a_9024_n502.n3 a_9024_n502.n2 2.878
R1011 a_9024_n502.n4 a_9024_n502.n3 0.764
R1012 a_10253_219.n1 a_10253_219.t7 318.922
R1013 a_10253_219.n0 a_10253_219.t4 273.935
R1014 a_10253_219.n0 a_10253_219.t5 273.935
R1015 a_10253_219.n1 a_10253_219.t6 269.116
R1016 a_10253_219.n4 a_10253_219.n3 193.227
R1017 a_10253_219.t7 a_10253_219.n0 179.142
R1018 a_10253_219.n2 a_10253_219.n1 106.999
R1019 a_10253_219.n3 a_10253_219.t1 28.568
R1020 a_10253_219.t0 a_10253_219.n4 28.565
R1021 a_10253_219.n4 a_10253_219.t3 28.565
R1022 a_10253_219.n2 a_10253_219.t2 18.149
R1023 a_10253_219.n3 a_10253_219.n2 3.726
R1024 a_10680_n474.n2 a_10680_n474.n0 267.767
R1025 a_10680_n474.n6 a_10680_n474.t5 16.058
R1026 a_10680_n474.n8 a_10680_n474.t4 16.058
R1027 a_10680_n474.n1 a_10680_n474.t2 14.282
R1028 a_10680_n474.n1 a_10680_n474.t9 14.282
R1029 a_10680_n474.n0 a_10680_n474.t11 14.282
R1030 a_10680_n474.n0 a_10680_n474.t8 14.282
R1031 a_10680_n474.n3 a_10680_n474.t3 14.282
R1032 a_10680_n474.n3 a_10680_n474.t10 14.282
R1033 a_10680_n474.n5 a_10680_n474.t6 14.282
R1034 a_10680_n474.n5 a_10680_n474.t7 14.282
R1035 a_10680_n474.t0 a_10680_n474.n9 14.282
R1036 a_10680_n474.n9 a_10680_n474.t1 14.282
R1037 a_10680_n474.n4 a_10680_n474.n3 1.511
R1038 a_10680_n474.n6 a_10680_n474.n5 0.999
R1039 a_10680_n474.n9 a_10680_n474.n8 0.999
R1040 a_10680_n474.n4 a_10680_n474.n2 0.669
R1041 a_10680_n474.n7 a_10680_n474.n6 0.575
R1042 a_10680_n474.n7 a_10680_n474.n4 0.227
R1043 a_10680_n474.n8 a_10680_n474.n7 0.2
R1044 a_10680_n474.n2 a_10680_n474.n1 0.001
R1045 Y[5].n7 Y[5].n6 194.965
R1046 Y[5].n4 Y[5].n2 157.665
R1047 Y[5].n4 Y[5].n3 122.999
R1048 Y[5].n6 Y[5].n0 90.436
R1049 Y[5].n5 Y[5].n1 90.416
R1050 Y[5].n6 Y[5].n5 74.302
R1051 Y[5].n5 Y[5].n4 50.575
R1052 Y[5].n0 Y[5].t2 14.282
R1053 Y[5].n0 Y[5].t0 14.282
R1054 Y[5].n1 Y[5].t1 14.282
R1055 Y[5].n1 Y[5].t5 14.282
R1056 Y[5].n3 Y[5].t4 14.282
R1057 Y[5].n3 Y[5].t6 14.282
R1058 Y[5].n2 Y[5].t7 8.7
R1059 Y[5].n2 Y[5].t3 8.7
R1060 Y[5] Y[5].n7 0.038
R1061 Y[5].n7 Y[5] 0.02
R1062 a_1979_217.n1 a_1979_217.t5 318.922
R1063 a_1979_217.n0 a_1979_217.t6 273.935
R1064 a_1979_217.n0 a_1979_217.t7 273.935
R1065 a_1979_217.n1 a_1979_217.t4 269.116
R1066 a_1979_217.n4 a_1979_217.n3 193.227
R1067 a_1979_217.t5 a_1979_217.n0 179.142
R1068 a_1979_217.n2 a_1979_217.n1 106.999
R1069 a_1979_217.n3 a_1979_217.t0 28.568
R1070 a_1979_217.t2 a_1979_217.n4 28.565
R1071 a_1979_217.n4 a_1979_217.t1 28.565
R1072 a_1979_217.n2 a_1979_217.t3 18.149
R1073 a_1979_217.n3 a_1979_217.n2 3.726
R1074 a_2524_n1208.t0 a_2524_n1208.t1 380.209
R1075 A[7].n5 A[7].n4 412.11
R1076 A[7].n1 A[7].t3 394.151
R1077 A[7].n4 A[7].t4 294.653
R1078 A[7].n0 A[7].t0 269.523
R1079 A[7].t3 A[7].n0 269.523
R1080 A[7].n5 A[7].n3 224.13
R1081 A[7].n2 A[7].t7 198.043
R1082 A[7].n0 A[7].t1 160.666
R1083 A[7] A[7].n5 138.229
R1084 A[7].n4 A[7].t6 111.663
R1085 A[7].n3 A[7].n1 97.816
R1086 A[7].n2 A[7].t5 93.989
R1087 A[7].n1 A[7].t2 80.333
R1088 A[7].n3 A[7].n2 6.615
R1089 B[5].n4 B[5].n3 592.056
R1090 B[5].t1 B[5].n1 313.873
R1091 B[5].n3 B[5].t5 294.986
R1092 B[5].n0 B[5].t6 272.288
R1093 B[5].n4 B[5].t0 204.68
R1094 B[5].n2 B[5].t1 190.152
R1095 B[5].n2 B[5].t7 190.152
R1096 B[5].n0 B[5].t4 160.666
R1097 B[5].n1 B[5].t2 160.666
R1098 B[5].n3 B[5].t3 110.859
R1099 B[5].n1 B[5].n0 96.129
R1100 B[5].t0 B[5].n2 80.333
R1101 B[5] B[5].n4 42.781
R1102 a_11092_n500.n1 a_11092_n500.t6 318.922
R1103 a_11092_n500.n0 a_11092_n500.t5 274.739
R1104 a_11092_n500.n0 a_11092_n500.t4 274.739
R1105 a_11092_n500.n1 a_11092_n500.t7 269.116
R1106 a_11092_n500.t6 a_11092_n500.n0 179.946
R1107 a_11092_n500.n2 a_11092_n500.n1 107.263
R1108 a_11092_n500.n3 a_11092_n500.t0 29.444
R1109 a_11092_n500.t2 a_11092_n500.n4 28.565
R1110 a_11092_n500.n4 a_11092_n500.t1 28.565
R1111 a_11092_n500.n2 a_11092_n500.t3 18.145
R1112 a_11092_n500.n3 a_11092_n500.n2 2.878
R1113 a_11092_n500.n4 a_11092_n500.n3 0.764
R1114 B[3].n4 B[3].n3 592.056
R1115 B[3].t1 B[3].n1 313.873
R1116 B[3].n3 B[3].t3 294.986
R1117 B[3].n0 B[3].t7 272.288
R1118 B[3].n4 B[3].t2 204.68
R1119 B[3].n2 B[3].t1 190.152
R1120 B[3].n2 B[3].t0 190.152
R1121 B[3].n0 B[3].t5 160.666
R1122 B[3].n1 B[3].t4 160.666
R1123 B[3].n3 B[3].t6 110.859
R1124 B[3].n1 B[3].n0 96.129
R1125 B[3].t2 B[3].n2 80.333
R1126 B[3] B[3].n4 42.783
R1127 a_4887_n504.n1 a_4887_n504.t6 318.922
R1128 a_4887_n504.n0 a_4887_n504.t7 274.739
R1129 a_4887_n504.n0 a_4887_n504.t4 274.739
R1130 a_4887_n504.n1 a_4887_n504.t5 269.116
R1131 a_4887_n504.t6 a_4887_n504.n0 179.946
R1132 a_4887_n504.n2 a_4887_n504.n1 107.263
R1133 a_4887_n504.n3 a_4887_n504.t2 29.444
R1134 a_4887_n504.n4 a_4887_n504.t3 28.565
R1135 a_4887_n504.t0 a_4887_n504.n4 28.565
R1136 a_4887_n504.n2 a_4887_n504.t1 18.145
R1137 a_4887_n504.n3 a_4887_n504.n2 2.878
R1138 a_4887_n504.n4 a_4887_n504.n3 0.764
R1139 B[2].n4 B[2].n3 592.056
R1140 B[2].t0 B[2].n1 313.873
R1141 B[2].n3 B[2].t6 294.986
R1142 B[2].n0 B[2].t5 272.288
R1143 B[2].n4 B[2].t7 204.68
R1144 B[2].n2 B[2].t0 190.152
R1145 B[2].n2 B[2].t4 190.152
R1146 B[2].n0 B[2].t2 160.666
R1147 B[2].n1 B[2].t1 160.666
R1148 B[2].n3 B[2].t3 110.859
R1149 B[2].n1 B[2].n0 96.129
R1150 B[2].t7 B[2].n2 80.333
R1151 B[2] B[2].n4 42.78
R1152 A[5].n5 A[5].n4 412.11
R1153 A[5].n1 A[5].t1 394.151
R1154 A[5].n4 A[5].t5 294.653
R1155 A[5].n0 A[5].t7 269.523
R1156 A[5].t1 A[5].n0 269.523
R1157 A[5].n5 A[5].n3 224.13
R1158 A[5].n2 A[5].t6 198.043
R1159 A[5].n0 A[5].t2 160.666
R1160 A[5] A[5].n5 138.227
R1161 A[5].n4 A[5].t0 111.663
R1162 A[5].n3 A[5].n1 97.816
R1163 A[5].n2 A[5].t4 93.989
R1164 A[5].n1 A[5].t3 80.333
R1165 A[5].n3 A[5].n2 6.615
R1166 a_15229_n500.n1 a_15229_n500.t5 318.922
R1167 a_15229_n500.n0 a_15229_n500.t6 274.739
R1168 a_15229_n500.n0 a_15229_n500.t4 274.739
R1169 a_15229_n500.n1 a_15229_n500.t7 269.116
R1170 a_15229_n500.t5 a_15229_n500.n0 179.946
R1171 a_15229_n500.n2 a_15229_n500.n1 107.263
R1172 a_15229_n500.t2 a_15229_n500.n4 29.444
R1173 a_15229_n500.n3 a_15229_n500.t1 28.565
R1174 a_15229_n500.n3 a_15229_n500.t0 28.565
R1175 a_15229_n500.n2 a_15229_n500.t3 18.145
R1176 a_15229_n500.n4 a_15229_n500.n2 2.878
R1177 a_15229_n500.n4 a_15229_n500.n3 0.764
R1178 Y[6].n7 Y[6].n6 194.965
R1179 Y[6].n4 Y[6].n2 157.665
R1180 Y[6].n4 Y[6].n3 122.999
R1181 Y[6].n6 Y[6].n0 90.436
R1182 Y[6].n5 Y[6].n1 90.416
R1183 Y[6].n6 Y[6].n5 74.302
R1184 Y[6].n5 Y[6].n4 50.575
R1185 Y[6].n0 Y[6].t3 14.282
R1186 Y[6].n0 Y[6].t5 14.282
R1187 Y[6].n1 Y[6].t4 14.282
R1188 Y[6].n1 Y[6].t6 14.282
R1189 Y[6].n3 Y[6].t7 14.282
R1190 Y[6].n3 Y[6].t1 14.282
R1191 Y[6].n2 Y[6].t2 8.7
R1192 Y[6].n2 Y[6].t0 8.7
R1193 Y[6] Y[6].n7 0.034
R1194 Y[6].n7 Y[6] 0.024
R1195 a_13103_n1208.t0 a_13103_n1208.t1 17.4
R1196 a_12322_217.n1 a_12322_217.t4 318.922
R1197 a_12322_217.n0 a_12322_217.t7 273.935
R1198 a_12322_217.n0 a_12322_217.t5 273.935
R1199 a_12322_217.n1 a_12322_217.t6 269.116
R1200 a_12322_217.n4 a_12322_217.n3 193.227
R1201 a_12322_217.t4 a_12322_217.n0 179.142
R1202 a_12322_217.n2 a_12322_217.n1 106.999
R1203 a_12322_217.n3 a_12322_217.t0 28.568
R1204 a_12322_217.n4 a_12322_217.t1 28.565
R1205 a_12322_217.t2 a_12322_217.n4 28.565
R1206 a_12322_217.n2 a_12322_217.t3 18.149
R1207 a_12322_217.n3 a_12322_217.n2 3.726
R1208 a_4593_n1210.t0 a_4593_n1210.t1 380.209
R1209 B[4].n4 B[4].n3 592.056
R1210 B[4].t7 B[4].n1 313.873
R1211 B[4].n3 B[4].t0 294.986
R1212 B[4].n0 B[4].t3 272.288
R1213 B[4].n4 B[4].t5 204.68
R1214 B[4].n2 B[4].t7 190.152
R1215 B[4].n2 B[4].t6 190.152
R1216 B[4].n0 B[4].t1 160.666
R1217 B[4].n1 B[4].t2 160.666
R1218 B[4].n3 B[4].t4 110.859
R1219 B[4].n1 B[4].n0 96.129
R1220 B[4].t5 B[4].n2 80.333
R1221 B[4] B[4].n4 42.781
R1222 a_8966_n1208.t0 a_8966_n1208.t1 17.4
R1223 a_12867_n1208.t0 a_12867_n1208.t1 380.209
R1224 a_6116_217.n1 a_6116_217.t7 318.922
R1225 a_6116_217.n0 a_6116_217.t4 273.935
R1226 a_6116_217.n0 a_6116_217.t5 273.935
R1227 a_6116_217.n1 a_6116_217.t6 269.116
R1228 a_6116_217.n4 a_6116_217.n3 193.227
R1229 a_6116_217.t7 a_6116_217.n0 179.142
R1230 a_6116_217.n2 a_6116_217.n1 106.999
R1231 a_6116_217.n3 a_6116_217.t0 28.568
R1232 a_6116_217.n4 a_6116_217.t1 28.565
R1233 a_6116_217.t2 a_6116_217.n4 28.565
R1234 a_6116_217.n2 a_6116_217.t3 18.149
R1235 a_6116_217.n3 a_6116_217.n2 3.726
R1236 a_8730_n1208.t0 a_8730_n1208.t1 380.209
R1237 a_750_n504.n1 a_750_n504.t7 318.922
R1238 a_750_n504.n0 a_750_n504.t5 274.739
R1239 a_750_n504.n0 a_750_n504.t6 274.739
R1240 a_750_n504.n1 a_750_n504.t4 269.116
R1241 a_750_n504.t7 a_750_n504.n0 179.946
R1242 a_750_n504.n2 a_750_n504.n1 107.263
R1243 a_750_n504.t2 a_750_n504.n4 29.444
R1244 a_750_n504.n3 a_750_n504.t0 28.565
R1245 a_750_n504.n3 a_750_n504.t1 28.565
R1246 a_750_n504.n2 a_750_n504.t3 18.145
R1247 a_750_n504.n4 a_750_n504.n2 2.878
R1248 a_750_n504.n4 a_750_n504.n3 0.764
R1249 a_456_n1210.t0 a_456_n1210.t1 380.209
R1250 a_6661_n1208.t0 a_6661_n1208.t1 380.209
R1251 a_14935_n1206.t0 a_14935_n1206.t1 380.209
R1252 a_6897_n1208.t0 a_6897_n1208.t1 17.4
R1253 a_2760_n1208.t0 a_2760_n1208.t1 17.4
R1254 a_11034_n1206.t0 a_11034_n1206.t1 17.4
R1255 a_15171_n1206.t0 a_15171_n1206.t1 17.4
R1256 a_10798_n1206.t0 a_10798_n1206.t1 380.209
R1257 a_4829_n1210.t0 a_4829_n1210.t1 17.4
C0 A[0] VDD 0.55fF
C1 B[0] A[0] 0.21fF
C2 B[5] Y[6] 0.00fF
C3 A[5] B[4] 0.04fF
C4 A[1] VDD 0.59fF
C5 B[0] A[1] 0.04fF
C6 Y[5] B[4] 0.00fF
C7 B[6] A[7] 0.04fF
C8 A[5] VDD 0.59fF
C9 B[6] A[6] 0.21fF
C10 Y[1] A[1] 0.18fF
C11 Y[7] B[6] 0.00fF
C12 B[1] A[2] 0.03fF
C13 Y[5] VDD 0.23fF
C14 Y[2] A[3] 0.01fF
C15 B[3] Y[4] 0.00fF
C16 VDD A[3] 0.59fF
C17 A[5] A[6] 0.00fF
C18 B[4] VDD 0.81fF
C19 B[6] Y[6] 0.15fF
C20 Y[2] VDD 0.23fF
C21 A[0] Y[0] 0.18fF
C22 Y[5] A[6] 0.01fF
C23 A[2] A[1] 0.00fF
C24 B[2] A[3] 0.04fF
C25 B[7] VDD 0.76fF
C26 Y[0] A[1] 0.01fF
C27 B[0] VDD 0.81fF
C28 Y[3] Y[4] 0.01fF
C29 Y[2] B[2] 0.15fF
C30 Y[2] Y[1] 0.01fF
C31 A[4] Y[4] 0.18fF
C32 B[2] VDD 0.81fF
C33 B[3] Y[3] 0.15fF
C34 Y[1] VDD 0.23fF
C35 Y[5] Y[6] 0.01fF
C36 B[0] Y[1] 0.00fF
C37 B[7] A[7] 0.21fF
C38 B[6] B[5] 0.01fF
C39 VDD A[7] 0.59fF
C40 A[4] B[3] 0.04fF
C41 A[6] VDD 0.59fF
C42 A[2] A[3] 0.00fF
C43 Y[7] B[7] 0.15fF
C44 Y[7] VDD 0.23fF
C45 Y[2] A[2] 0.18fF
C46 A[5] Y[4] 0.01fF
C47 A[4] Y[3] 0.01fF
C48 A[5] B[5] 0.21fF
C49 A[2] VDD 0.59fF
C50 A[6] A[7] 0.00fF
C51 Y[5] Y[4] 0.01fF
C52 Y[7] A[7] 0.18fF
C53 Y[5] B[5] 0.15fF
C54 VDD Y[6] 0.23fF
C55 Y[0] VDD 0.23fF
C56 B[0] Y[0] 0.15fF
C57 A[2] B[2] 0.21fF
C58 A[2] Y[1] 0.01fF
C59 B[1] A[1] 0.21fF
C60 Y[0] Y[1] 0.01fF
C61 Y[4] B[4] 0.15fF
C62 B[5] B[4] 0.01fF
C63 Y[6] A[7] 0.01fF
C64 B[3] A[3] 0.21fF
C65 A[6] Y[6] 0.18fF
C66 A[4] A[5] 0.00fF
C67 Y[7] Y[6] 0.01fF
C68 B[3] B[4] 0.01fF
C69 A[0] A[1] 0.00fF
C70 Y[4] VDD 0.23fF
C71 B[5] VDD 0.81fF
C72 B[3] VDD 0.81fF
C73 Y[3] A[3] 0.18fF
C74 A[4] A[3] 0.00fF
C75 Y[2] Y[3] 0.01fF
C76 Y[2] B[1] 0.00fF
C77 B[3] B[2] 0.01fF
C78 A[4] B[4] 0.21fF
C79 B[5] A[6] 0.03fF
C80 Y[3] VDD 0.23fF
C81 B[1] VDD 0.81fF
C82 B[0] B[1] 0.01fF
C83 Y[5] A[5] 0.18fF
C84 A[4] VDD 0.59fF
C85 Y[3] B[2] 0.00fF
C86 B[1] B[2] 0.01fF
C87 B[7] B[6] 0.01fF
C88 B[6] VDD 0.81fF
C89 B[1] Y[1] 0.15fF
.ends

