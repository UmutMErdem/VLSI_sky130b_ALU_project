magic
tech sky130B
magscale 1 2
timestamp 1736460087
<< nwell >>
rect -471 496 1306 814
rect -484 95 -420 262
rect -476 62 -420 95
<< ndiff >>
rect 115 -1071 167 -871
rect 668 -960 735 -871
rect 667 -987 735 -960
rect 644 -1071 735 -987
<< pdiff >>
rect -484 95 -420 262
rect -476 62 -420 95
<< psubdiff >>
rect 338 -1526 524 -1502
rect 338 -1572 380 -1526
rect 484 -1572 524 -1526
rect 338 -1608 524 -1572
<< nsubdiff >>
rect 268 720 572 776
rect 268 644 322 720
rect 518 644 572 720
rect 268 630 572 644
<< psubdiffcont >>
rect 380 -1572 484 -1526
<< nsubdiffcont >>
rect 322 644 518 720
<< poly >>
rect -377 477 -81 516
rect 90 477 386 516
rect 444 477 740 516
rect 917 477 1213 516
rect -818 278 -522 317
rect 1390 278 1686 317
rect -818 -224 -758 59
rect -818 -241 -682 -224
rect -818 -296 -759 -241
rect -701 -296 -682 -241
rect -818 -311 -682 -296
rect -818 -623 -758 -311
rect -259 -356 -199 43
rect 209 -124 268 54
rect 209 -125 272 -124
rect 206 -141 272 -125
rect 206 -175 222 -141
rect 256 -175 272 -141
rect 206 -191 272 -175
rect 309 -240 404 -225
rect 309 -295 328 -240
rect 386 -263 404 -240
rect 562 -263 622 43
rect 386 -295 622 -263
rect 309 -312 622 -295
rect -259 -413 268 -356
rect 208 -512 268 -413
rect 197 -525 278 -512
rect 197 -580 210 -525
rect 268 -580 278 -525
rect 197 -591 278 -580
rect -818 -668 76 -623
rect 16 -857 76 -668
rect 208 -857 268 -591
rect 326 -857 386 -312
rect 1035 -354 1095 45
rect 1516 -87 1582 -84
rect 1626 -87 1686 59
rect 1516 -100 1686 -87
rect 1516 -134 1532 -100
rect 1566 -134 1686 -100
rect 1516 -147 1686 -134
rect 1516 -150 1582 -147
rect 557 -371 1095 -354
rect 557 -405 576 -371
rect 610 -405 1095 -371
rect 557 -411 1095 -405
rect 557 -421 626 -411
rect 557 -423 622 -421
rect 441 -761 507 -745
rect 441 -795 457 -761
rect 491 -795 507 -761
rect 441 -811 507 -795
rect 444 -855 504 -811
rect 562 -855 622 -423
rect 1626 -623 1686 -147
rect 758 -668 1686 -623
rect 758 -856 818 -668
rect 383 -1352 449 -1344
rect 758 -1352 818 -1083
rect 383 -1360 818 -1352
rect 383 -1394 399 -1360
rect 433 -1394 818 -1360
rect 383 -1403 818 -1394
rect 383 -1410 449 -1403
<< polycont >>
rect -759 -296 -701 -241
rect 222 -175 256 -141
rect 328 -295 386 -240
rect 210 -580 268 -525
rect 1532 -134 1566 -100
rect 576 -405 610 -371
rect 457 -795 491 -761
rect 399 -1394 433 -1360
<< locali >>
rect 306 720 534 738
rect 306 644 322 720
rect 518 644 534 720
rect 306 628 534 644
rect -423 503 -153 542
rect -423 431 -389 503
rect -187 431 -153 503
rect 44 502 314 541
rect 44 430 78 502
rect 280 430 314 502
rect 516 502 786 541
rect 516 430 550 502
rect 752 430 786 502
rect 989 502 1259 541
rect 989 430 1023 502
rect 1225 430 1259 502
rect -864 301 -594 340
rect -864 222 -830 301
rect -628 229 -594 301
rect 1462 300 1732 337
rect 1462 226 1496 300
rect 1698 226 1732 300
rect -746 23 -712 95
rect -510 23 -476 95
rect -746 -16 -476 23
rect -305 23 -271 95
rect -69 23 -35 95
rect 162 23 196 95
rect 398 23 432 95
rect 634 23 668 95
rect 871 23 905 95
rect 1107 23 1141 95
rect -305 -16 1141 23
rect 1344 20 1378 80
rect 1580 20 1614 92
rect 1344 -19 1614 20
rect 222 -141 256 -125
rect 1516 -134 1532 -100
rect 1566 -134 1582 -100
rect 222 -191 256 -175
rect -1007 -240 -950 -236
rect -1007 -300 -1003 -240
rect -954 -300 -950 -240
rect -1007 -304 -950 -300
rect -775 -241 -683 -224
rect -775 -296 -759 -241
rect -699 -296 -683 -241
rect -775 -309 -683 -296
rect 310 -240 402 -227
rect 310 -295 326 -240
rect 386 -295 402 -240
rect 310 -312 402 -295
rect -1007 -356 -950 -352
rect -1007 -416 -1003 -356
rect -954 -416 -950 -356
rect -1007 -420 -950 -416
rect 576 -371 610 -355
rect 576 -421 610 -405
rect -1007 -524 -950 -520
rect -1007 -584 -1003 -524
rect -954 -584 -950 -524
rect -1007 -588 -950 -584
rect 192 -525 284 -512
rect 192 -580 208 -525
rect 268 -580 284 -525
rect 192 -597 284 -580
rect 457 -761 491 -745
rect 457 -811 491 -795
rect 115 -1071 167 -871
rect 668 -960 735 -871
rect 667 -987 735 -960
rect 644 -1071 735 -987
rect 383 -1394 399 -1360
rect 433 -1394 449 -1360
rect 364 -1512 500 -1508
rect 364 -1526 402 -1512
rect 460 -1526 500 -1512
rect 364 -1572 380 -1526
rect 484 -1572 500 -1526
rect 364 -1594 500 -1572
<< viali >>
rect 388 646 460 700
rect 1532 -134 1566 -100
rect 222 -175 256 -141
rect -1003 -300 -954 -240
rect -759 -296 -701 -241
rect -701 -296 -699 -241
rect 326 -295 328 -240
rect 328 -295 386 -240
rect -1003 -416 -954 -356
rect 576 -405 610 -371
rect -1003 -584 -954 -524
rect 208 -580 210 -525
rect 210 -580 268 -525
rect 457 -795 491 -761
rect 399 -1394 433 -1360
rect 402 -1526 460 -1512
rect 402 -1558 460 -1526
<< metal1 >>
rect 374 646 384 706
rect 464 646 474 706
rect 374 606 474 646
rect -423 549 1380 606
rect -423 430 -389 549
rect 752 422 786 549
rect -865 -124 -830 110
rect -484 95 -420 262
rect 1343 234 1380 549
rect 1343 189 1364 211
rect -476 62 -420 95
rect 44 -22 78 89
rect 1225 -22 1259 90
rect 44 -64 1259 -22
rect 1225 -84 1259 -64
rect 1225 -100 1582 -84
rect -865 -141 272 -124
rect -865 -175 222 -141
rect 256 -175 272 -141
rect 1225 -134 1532 -100
rect 1566 -134 1582 -100
rect 1225 -150 1582 -134
rect -865 -191 272 -175
rect -1124 -236 -948 -228
rect -1124 -304 -1007 -236
rect -950 -304 -940 -236
rect -1124 -312 -948 -304
rect -1124 -352 -948 -344
rect -1124 -420 -1007 -352
rect -950 -420 -940 -352
rect -1124 -428 -948 -420
rect -1124 -520 -948 -512
rect -1124 -588 -1007 -520
rect -950 -588 -940 -520
rect -1124 -596 -948 -588
rect -865 -701 -830 -191
rect -775 -237 -683 -224
rect -775 -300 -763 -237
rect -692 -300 -683 -237
rect -775 -309 -683 -300
rect 310 -237 402 -227
rect 310 -299 322 -237
rect 392 -299 402 -237
rect 310 -312 402 -299
rect 1698 -292 1733 110
rect 557 -354 622 -351
rect 557 -357 626 -354
rect 557 -417 563 -357
rect 622 -417 632 -357
rect 557 -421 626 -417
rect 557 -423 622 -421
rect 1698 -438 1879 -292
rect 192 -520 284 -512
rect 192 -585 204 -520
rect 272 -585 284 -520
rect 192 -597 284 -585
rect 1698 -700 1733 -438
rect -865 -748 507 -701
rect 829 -747 1733 -700
rect -31 -950 3 -748
rect 441 -761 507 -748
rect 441 -795 457 -761
rect 491 -795 507 -761
rect 441 -811 507 -795
rect 115 -1018 167 -871
rect 668 -960 735 -871
rect 830 -950 864 -747
rect 667 -987 735 -960
rect 88 -1071 167 -1018
rect 644 -1018 735 -987
rect 644 -1071 746 -1018
rect 88 -1438 122 -1071
rect 398 -1344 432 -1242
rect 383 -1360 449 -1344
rect 383 -1394 399 -1360
rect 433 -1394 449 -1360
rect 383 -1410 449 -1394
rect 712 -1438 746 -1071
rect 88 -1490 746 -1438
rect 386 -1512 478 -1490
rect 386 -1564 398 -1512
rect 464 -1564 478 -1512
rect 386 -1568 478 -1564
<< via1 >>
rect 384 700 464 706
rect 384 646 388 700
rect 388 646 460 700
rect 460 646 464 700
rect -1007 -240 -950 -236
rect -1007 -300 -1003 -240
rect -1003 -300 -954 -240
rect -954 -300 -950 -240
rect -1007 -304 -950 -300
rect -1007 -356 -950 -352
rect -1007 -416 -1003 -356
rect -1003 -416 -954 -356
rect -954 -416 -950 -356
rect -1007 -420 -950 -416
rect -1007 -524 -950 -520
rect -1007 -584 -1003 -524
rect -1003 -584 -954 -524
rect -954 -584 -950 -524
rect -1007 -588 -950 -584
rect -763 -241 -692 -237
rect -763 -296 -759 -241
rect -759 -296 -699 -241
rect -699 -296 -692 -241
rect -763 -300 -692 -296
rect 322 -240 392 -237
rect 322 -295 326 -240
rect 326 -295 386 -240
rect 386 -295 392 -240
rect 322 -299 392 -295
rect 563 -371 622 -357
rect 563 -405 576 -371
rect 576 -405 610 -371
rect 610 -405 622 -371
rect 563 -417 622 -405
rect 204 -525 272 -520
rect 204 -580 208 -525
rect 208 -580 268 -525
rect 268 -580 272 -525
rect 204 -585 272 -580
rect 398 -1558 402 -1512
rect 402 -1558 460 -1512
rect 460 -1558 464 -1512
rect 398 -1564 464 -1558
<< metal2 >>
rect 372 734 472 744
rect 372 632 472 642
rect -1007 -227 -950 -226
rect -774 -227 -681 -225
rect -1015 -228 401 -227
rect -1124 -236 401 -228
rect -1124 -304 -1007 -236
rect -950 -237 401 -236
rect -950 -300 -763 -237
rect -692 -299 322 -237
rect 392 -299 401 -237
rect -692 -300 401 -299
rect -950 -304 401 -300
rect -1124 -311 401 -304
rect -1124 -312 -940 -311
rect -1007 -314 -950 -312
rect -1007 -344 -950 -342
rect -1124 -347 -922 -344
rect -1124 -352 622 -347
rect -1124 -420 -1007 -352
rect -950 -357 622 -352
rect -950 -417 563 -357
rect -950 -420 622 -417
rect -1124 -426 622 -420
rect -1124 -429 -922 -426
rect 563 -427 622 -426
rect -1007 -430 -950 -429
rect -1007 -511 -950 -510
rect -1124 -512 -922 -511
rect -1124 -520 283 -512
rect -1124 -588 -1007 -520
rect -950 -585 204 -520
rect 272 -585 283 -520
rect -950 -588 283 -585
rect -1124 -596 283 -588
rect -1007 -598 -950 -596
rect 392 -1510 468 -1500
rect 392 -1578 468 -1568
<< via2 >>
rect 372 706 472 734
rect 372 646 384 706
rect 384 646 464 706
rect 464 646 472 706
rect 372 642 472 646
rect 392 -1512 468 -1510
rect 392 -1564 398 -1512
rect 398 -1564 464 -1512
rect 464 -1564 468 -1512
rect 392 -1568 468 -1564
<< metal3 >>
rect 362 734 482 739
rect 362 640 372 734
rect 472 640 482 734
rect 362 637 482 640
rect 352 -1510 518 -1502
rect 352 -1578 386 -1510
rect 470 -1578 518 -1510
rect 352 -1582 518 -1578
<< via3 >>
rect 372 642 472 732
rect 372 640 472 642
rect 386 -1568 392 -1510
rect 392 -1568 468 -1510
rect 468 -1568 470 -1510
rect 386 -1578 470 -1568
<< metal4 >>
rect 136 732 710 812
rect 136 640 372 732
rect 472 640 710 732
rect 136 620 710 640
rect 238 -1510 618 -1502
rect 238 -1578 386 -1510
rect 470 -1578 618 -1510
rect 238 -1608 618 -1578
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_0
timestamp 1735665674
transform 1 0 46 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_AJ3TNB  sky130_fd_pr__nfet_01v8_AJ3TNB_1
timestamp 1735665674
transform 1 0 788 0 1 -971
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_CSZSK8  sky130_fd_pr__nfet_01v8_CSZSK8_0
timestamp 1735665674
transform 1 0 415 0 1 -1071
box -265 -226 265 226
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_0
timestamp 1735665674
transform 1 0 415 0 1 262
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_0
timestamp 1735665674
transform 1 0 1065 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_6CQCZ3  sky130_fd_pr__pfet_01v8_6CQCZ3_1
timestamp 1735665674
transform 1 0 -229 0 1 262
box -242 -262 242 262
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_0
timestamp 1735665674
transform 1 0 1538 0 1 162
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_2
timestamp 1735665674
transform 1 0 -670 0 1 162
box -242 -162 242 162
<< labels >>
flabel metal1 -1118 -590 -1020 -516 1 FreeSans 240 0 0 0 D1
port 1 n
flabel metal1 -1118 -306 -1020 -232 1 FreeSans 240 0 0 0 S
port 2 n
flabel metal1 -1118 -422 -1020 -348 1 FreeSans 240 0 0 0 D0
port 3 n
flabel metal1 1718 -428 1870 -301 1 FreeSans 240 0 0 0 OUT
port 4 n
flabel metal4 380 -1602 484 -1546 1 FreeSerif 640 0 0 0 VSS
port 8 n
flabel metal4 352 644 500 758 1 FreeSerif 640 0 0 0 VDD
port 9 n
<< end >>
