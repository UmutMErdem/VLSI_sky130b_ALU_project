** sch_path: /home/ahmet/Desktop/arithmetic_unit/logic_and_tb.sch
**.subckt logic_and_tb
x1 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] GND VDD B[0] B[1]
+ B[2] B[3] B[4] B[5] B[6] B[7] logic_and
VDD VDD GND 1.2
V1 A[2] GND pulse(0, 1.2, 40n, 0.1p, 0.1p, 20n, 80n)
V3 A[0] GND pulse(0, 1.2, 0n, 0.1p, 0.1p, 20n, 80n)
V4 A[3] GND pulse(0, 1.2, 60n, 0.1p, 0.1p, 20n, 80n)
V2 A[1] GND pulse(0, 1.2, 20n, 0.1p, 0.1p, 20n, 40n)
V5 A[6] GND pulse(0, 1.2, 40n, 0.1p, 0.1p, 20n, 80n)
V6 A[4] GND pulse(0, 1.2, 0n, 0.1p, 0.1p, 20n, 40n)
V7 A[7] GND pulse(0, 1.2, 60n, 0.1p, 0.1p, 20n, 80n)
V8 A[5] GND pulse(0, 1.2, 20n, 0.1p, 0.1p, 20n, 80n)
V9 B[2] GND pulse(0, 1.2, 40n, 0.1p, 0.1p, 20n, 80n)
V10 B[0] GND pulse(0, 1.2, 0n, 0.1p, 0.1p, 20n, 80n)
V11 B[3] GND pulse(0, 1.2, 60n, 0.1p, 0.1p, 20n, 80n)
V12 B[1] GND pulse(0, 1.2, 20n, 0.1p, 0.1p, 20n, 80n)
V13 B[6] GND pulse(0, 1.2, 40n, 0.1p, 0.1p, 20n, 80n)
V14 B[4] GND pulse(0, 1.2, 0n, 0.1p, 0.1p, 20n, 80n)
V15 B[7] GND pulse(0, 1.2, 60n, 0.1p, 0.1p, 20n, 80n)
V16 B[5] GND pulse(0, 1.2, 20n, 0.1p, 0.1p, 20n, 80n)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt_mm



.control
save all

set color0 = white
tran 1p 80n
plot "a[0]" "a[1]"+2 "a[2]"+4 "a[3]"+6 "a[4]"+8 "a[5]"+10 "a[6]"+12 "a[7]"+14
plot "b[0]" "b[1]"+2 "b[2]"+4 "b[3]"+6 "b[4]"+8 "b[5]"+10 "b[6]"+12 "b[7]"+14
plot "y[0]" "y[1]"+2 "y[2]"+4 "y[3]"+6 "y[4]"+8 "y[5]"+10 "y[6]"+12 "y[7]"+14
.endc

**** end user architecture code
**.ends

* expanding   symbol:  logic_and.sym # of pins=5
** sym_path: /home/ahmet/Desktop/arithmetic_unit/logic_and.sym
** sch_path: /home/ahmet/Desktop/arithmetic_unit/logic_and.sch
.subckt logic_and  A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
+ VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7]
*.ipin A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7]
*.opin Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7]
*.iopin VSS
*.iopin VDD
*.ipin B[0],B[1],B[2],B[3],B[4],B[5],B[6],B[7]
x1 VSS A[0] B[0] VDD Y[0] and2
x2 VSS A[1] B[1] VDD Y[1] and2
x3 VSS A[2] B[2] VDD Y[2] and2
x4 VSS A[3] B[3] VDD Y[3] and2
x5 VSS A[4] B[4] VDD Y[4] and2
x6 VSS A[5] B[5] VDD Y[5] and2
x7 VSS A[6] B[6] VDD Y[6] and2
x8 VSS A[7] B[7] VDD Y[7] and2
.ends


* expanding   symbol:  and2.sym # of pins=5
** sym_path: /home/ahmet/Desktop/arithmetic_unit/and2.sym
** sch_path: /home/ahmet/Desktop/arithmetic_unit/and2.sch
.subckt and2  VSS A B VDD OUT
*.iopin VSS
*.ipin A
*.ipin B
*.iopin VDD
*.opin OUT
XM2 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 A net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
