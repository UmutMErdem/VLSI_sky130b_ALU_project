magic
tech sky130B
magscale 1 2
timestamp 1733696680
<< poly >>
rect 95 289 391 325
rect 449 288 745 324
rect 332 -168 390 48
rect 450 -168 508 48
<< metal1 >>
rect 386 522 446 532
rect 386 452 446 462
rect 394 404 434 452
rect 50 374 790 404
rect 50 250 82 374
rect 286 250 318 374
rect 522 250 554 374
rect 758 250 790 374
rect 166 -26 202 84
rect 402 -26 438 84
rect 638 -24 674 86
rect 638 -26 836 -24
rect 166 -56 836 -26
rect 286 -194 320 -56
rect 642 -58 836 -56
rect 736 -124 836 -58
rect 694 -340 704 -332
rect 522 -380 704 -340
rect 58 -408 158 -380
rect 694 -392 704 -380
rect 764 -392 774 -332
rect 58 -456 392 -408
rect 58 -480 158 -456
rect 58 -544 158 -522
rect 450 -544 512 -408
rect 58 -592 512 -544
rect 58 -622 158 -592
<< via1 >>
rect 386 462 446 522
rect 704 -392 764 -332
<< metal2 >>
rect 366 452 376 532
rect 456 452 466 532
rect 694 -322 774 -312
rect 694 -412 774 -402
<< via2 >>
rect 376 522 456 532
rect 376 462 386 522
rect 386 462 446 522
rect 446 462 456 522
rect 376 452 456 462
rect 694 -332 774 -322
rect 694 -392 704 -332
rect 704 -392 764 -332
rect 764 -392 774 -332
rect 694 -402 774 -392
<< metal3 >>
rect 366 542 466 552
rect 366 432 466 442
rect 674 -412 684 -312
rect 784 -412 794 -312
<< via3 >>
rect 366 532 466 542
rect 366 452 376 532
rect 376 452 456 532
rect 456 452 466 532
rect 366 442 466 452
rect 684 -322 784 -312
rect 684 -402 694 -322
rect 694 -402 774 -322
rect 774 -402 784 -322
rect 684 -412 784 -402
<< metal4 >>
rect 356 638 478 640
rect 324 542 524 638
rect 324 496 366 542
rect 365 442 366 496
rect 466 496 524 542
rect 466 442 467 496
rect 365 441 467 442
rect 742 -311 910 -302
rect 683 -312 910 -311
rect 683 -412 684 -312
rect 784 -412 910 -312
rect 683 -413 910 -412
rect 742 -492 910 -413
use sky130_fd_pr__nfet_01v8_8H4MRT  sky130_fd_pr__nfet_01v8_8H4MRT_0
timestamp 1733695122
transform 1 0 480 0 1 -307
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_8H4MRT  sky130_fd_pr__nfet_01v8_8H4MRT_1
timestamp 1733695122
transform 1 0 362 0 1 -307
box -88 -157 88 157
use sky130_fd_pr__pfet_01v8_A64S85  sky130_fd_pr__pfet_01v8_A64S85_0
timestamp 1733691381
transform 1 0 420 0 1 168
box -419 -162 419 162
<< labels >>
flabel space 322 498 522 640 1 FreeSans 480 0 0 0 VDD
port 4 n
flabel metal4 760 -452 880 -348 1 FreeSans 480 0 0 0 VSS
port 1 n
flabel metal1 58 -622 158 -522 1 FreeSans 480 0 0 0 B
port 3 n
flabel metal1 58 -480 158 -380 1 FreeSans 480 0 0 0 A
port 2 n
flabel metal1 736 -124 836 -24 1 FreeSans 480 0 0 0 Y
port 5 n
<< end >>
