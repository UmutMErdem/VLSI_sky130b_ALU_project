magic
tech sky130B
magscale 1 2
timestamp 1736524280
<< nwell >>
rect 458 1226 1372 1504
rect 1626 1226 2540 1504
rect 2794 1226 3708 1504
rect 3962 1226 4876 1504
rect 5136 1228 6050 1506
rect 6304 1228 7218 1506
rect 7472 1228 8386 1506
rect 8640 1228 9554 1506
rect 888 418 1372 1226
rect 2056 418 2540 1226
rect 3224 418 3708 1226
rect 4392 418 4876 1226
rect 5566 420 6050 1228
rect 6734 420 7218 1228
rect 7902 420 8386 1228
rect 9070 420 9554 1228
<< psubdiff >>
rect 538 82 734 112
rect 538 16 578 82
rect 696 16 734 82
rect 538 -32 734 16
rect 1706 82 1902 112
rect 1706 16 1746 82
rect 1864 16 1902 82
rect 1706 -32 1902 16
rect 2874 82 3070 112
rect 2874 16 2914 82
rect 3032 16 3070 82
rect 2874 -32 3070 16
rect 4042 82 4238 112
rect 4042 16 4082 82
rect 4200 16 4238 82
rect 4042 -32 4238 16
rect 5216 84 5412 114
rect 5216 18 5256 84
rect 5374 18 5412 84
rect 5216 -30 5412 18
rect 6384 84 6580 114
rect 6384 18 6424 84
rect 6542 18 6580 84
rect 6384 -30 6580 18
rect 7552 84 7748 114
rect 7552 18 7592 84
rect 7710 18 7748 84
rect 7552 -30 7748 18
rect 8720 84 8916 114
rect 8720 18 8760 84
rect 8878 18 8916 84
rect 8720 -30 8916 18
<< nsubdiff >>
rect 978 1426 1244 1464
rect 978 1354 1034 1426
rect 1178 1354 1244 1426
rect 2146 1426 2412 1464
rect 978 1324 1244 1354
rect 2146 1354 2202 1426
rect 2346 1354 2412 1426
rect 3314 1426 3580 1464
rect 2146 1324 2412 1354
rect 3314 1354 3370 1426
rect 3514 1354 3580 1426
rect 4482 1426 4748 1464
rect 3314 1324 3580 1354
rect 4482 1354 4538 1426
rect 4682 1354 4748 1426
rect 5656 1428 5922 1466
rect 4482 1324 4748 1354
rect 5656 1356 5712 1428
rect 5856 1356 5922 1428
rect 6824 1428 7090 1466
rect 5656 1326 5922 1356
rect 6824 1356 6880 1428
rect 7024 1356 7090 1428
rect 7992 1428 8258 1466
rect 6824 1326 7090 1356
rect 7992 1356 8048 1428
rect 8192 1356 8258 1428
rect 9160 1428 9426 1466
rect 7992 1326 8258 1356
rect 9160 1356 9216 1428
rect 9360 1356 9426 1428
rect 9160 1326 9426 1356
<< psubdiffcont >>
rect 578 16 696 82
rect 1746 16 1864 82
rect 2914 16 3032 82
rect 4082 16 4200 82
rect 5256 18 5374 84
rect 6424 18 6542 84
rect 7592 18 7710 84
rect 8760 18 8878 84
<< nsubdiffcont >>
rect 1034 1354 1178 1426
rect 2202 1354 2346 1426
rect 3370 1354 3514 1426
rect 4538 1354 4682 1426
rect 5712 1356 5856 1428
rect 6880 1356 7024 1428
rect 8048 1356 8192 1428
rect 9216 1356 9360 1428
<< poly >>
rect 400 1348 466 1364
rect 400 1314 416 1348
rect 450 1344 466 1348
rect 450 1314 950 1344
rect 1568 1348 1634 1364
rect 400 1301 950 1314
rect 400 1298 466 1301
rect 400 1249 466 1256
rect 906 1249 950 1301
rect 1568 1314 1584 1348
rect 1618 1344 1634 1348
rect 1618 1314 2118 1344
rect 2736 1348 2802 1364
rect 1568 1301 2118 1314
rect 1568 1298 1634 1301
rect 1568 1249 1634 1256
rect 2074 1249 2118 1301
rect 2736 1314 2752 1348
rect 2786 1344 2802 1348
rect 2786 1314 3286 1344
rect 3904 1348 3970 1364
rect 2736 1301 3286 1314
rect 2736 1298 2802 1301
rect 2736 1249 2802 1256
rect 3242 1249 3286 1301
rect 3904 1314 3920 1348
rect 3954 1344 3970 1348
rect 3954 1314 4454 1344
rect 5078 1350 5144 1366
rect 3904 1301 4454 1314
rect 3904 1298 3970 1301
rect 3904 1249 3970 1256
rect 4410 1249 4454 1301
rect 5078 1316 5094 1350
rect 5128 1346 5144 1350
rect 5128 1316 5628 1346
rect 6246 1350 6312 1366
rect 5078 1303 5628 1316
rect 5078 1300 5144 1303
rect 5078 1251 5144 1258
rect 5584 1251 5628 1303
rect 6246 1316 6262 1350
rect 6296 1346 6312 1350
rect 6296 1316 6796 1346
rect 7414 1350 7480 1366
rect 6246 1303 6796 1316
rect 6246 1300 6312 1303
rect 6246 1251 6312 1258
rect 6752 1251 6796 1303
rect 7414 1316 7430 1350
rect 7464 1346 7480 1350
rect 7464 1316 7964 1346
rect 8582 1350 8648 1366
rect 7414 1303 7964 1316
rect 7414 1300 7480 1303
rect 7414 1251 7480 1258
rect 7920 1251 7964 1303
rect 8582 1316 8598 1350
rect 8632 1346 8648 1350
rect 8632 1316 9132 1346
rect 8582 1303 9132 1316
rect 8582 1300 8648 1303
rect 8582 1251 8648 1258
rect 9088 1251 9132 1303
rect 400 1240 848 1249
rect 400 1206 416 1240
rect 450 1208 848 1240
rect 906 1208 1202 1249
rect 1568 1240 2016 1249
rect 450 1207 584 1208
rect 450 1206 466 1207
rect 400 1190 466 1206
rect 1568 1206 1584 1240
rect 1618 1208 2016 1240
rect 2074 1208 2370 1249
rect 2736 1240 3184 1249
rect 1618 1207 1752 1208
rect 1618 1206 1634 1207
rect 1568 1190 1634 1206
rect 2736 1206 2752 1240
rect 2786 1208 3184 1240
rect 3242 1208 3538 1249
rect 3904 1240 4352 1249
rect 2786 1207 2920 1208
rect 2786 1206 2802 1207
rect 2736 1190 2802 1206
rect 3904 1206 3920 1240
rect 3954 1208 4352 1240
rect 4410 1208 4706 1249
rect 5078 1242 5526 1251
rect 5078 1208 5094 1242
rect 5128 1210 5526 1242
rect 5584 1210 5880 1251
rect 6246 1242 6694 1251
rect 5128 1209 5262 1210
rect 5128 1208 5144 1209
rect 3954 1207 4088 1208
rect 3954 1206 3970 1207
rect 3904 1190 3970 1206
rect 5078 1192 5144 1208
rect 6246 1208 6262 1242
rect 6296 1210 6694 1242
rect 6752 1210 7048 1251
rect 7414 1242 7862 1251
rect 6296 1209 6430 1210
rect 6296 1208 6312 1209
rect 6246 1192 6312 1208
rect 7414 1208 7430 1242
rect 7464 1210 7862 1242
rect 7920 1210 8216 1251
rect 8582 1242 9030 1251
rect 7464 1209 7598 1210
rect 7464 1208 7480 1209
rect 7414 1192 7480 1208
rect 8582 1208 8598 1242
rect 8632 1210 9030 1242
rect 9088 1210 9384 1251
rect 8632 1209 8766 1210
rect 8632 1208 8648 1209
rect 8582 1192 8648 1208
rect 552 681 613 770
rect 462 628 613 681
rect 462 410 522 628
rect 906 586 966 771
rect 1720 681 1781 770
rect 580 535 966 586
rect 1630 628 1781 681
rect 580 408 640 535
rect 695 477 761 493
rect 695 443 711 477
rect 745 443 761 477
rect 695 427 761 443
rect 1630 410 1690 628
rect 2074 586 2134 771
rect 2888 681 2949 770
rect 1748 535 2134 586
rect 2798 628 2949 681
rect 1748 408 1808 535
rect 1863 477 1929 493
rect 1863 443 1879 477
rect 1913 443 1929 477
rect 1863 427 1929 443
rect 2798 410 2858 628
rect 3242 586 3302 771
rect 4056 681 4117 770
rect 2916 535 3302 586
rect 3966 628 4117 681
rect 2916 408 2976 535
rect 3031 477 3097 493
rect 3031 443 3047 477
rect 3081 443 3097 477
rect 3031 427 3097 443
rect 3966 410 4026 628
rect 4410 586 4470 771
rect 5230 683 5291 772
rect 4084 535 4470 586
rect 5140 630 5291 683
rect 4084 408 4144 535
rect 4199 477 4265 493
rect 4199 443 4215 477
rect 4249 443 4265 477
rect 4199 427 4265 443
rect 5140 412 5200 630
rect 5584 588 5644 773
rect 6398 683 6459 772
rect 5258 537 5644 588
rect 6308 630 6459 683
rect 5258 410 5318 537
rect 5373 479 5439 495
rect 5373 445 5389 479
rect 5423 445 5439 479
rect 5373 429 5439 445
rect 6308 412 6368 630
rect 6752 588 6812 773
rect 7566 683 7627 772
rect 6426 537 6812 588
rect 7476 630 7627 683
rect 6426 410 6486 537
rect 6541 479 6607 495
rect 6541 445 6557 479
rect 6591 445 6607 479
rect 6541 429 6607 445
rect 7476 412 7536 630
rect 7920 588 7980 773
rect 8734 683 8795 772
rect 7594 537 7980 588
rect 8644 630 8795 683
rect 7594 410 7654 537
rect 7709 479 7775 495
rect 7709 445 7725 479
rect 7759 445 7775 479
rect 7709 429 7775 445
rect 8644 412 8704 630
rect 9088 588 9148 773
rect 8762 537 9148 588
rect 8762 410 8822 537
rect 8877 479 8943 495
rect 8877 445 8893 479
rect 8927 445 8943 479
rect 8877 429 8943 445
rect 698 172 758 194
rect 982 172 1041 194
rect 1100 172 1159 194
rect 1218 172 1277 194
rect 698 131 1277 172
rect 1866 172 1926 194
rect 2149 172 2209 194
rect 2267 172 2327 194
rect 2385 172 2445 194
rect 1866 131 2445 172
rect 3034 172 3094 194
rect 3317 172 3377 194
rect 3435 172 3495 194
rect 3553 172 3613 194
rect 3034 131 3613 172
rect 4202 172 4262 194
rect 4486 172 4546 194
rect 4604 172 4664 194
rect 4722 172 4781 194
rect 4202 131 4781 172
rect 5376 174 5436 196
rect 5659 174 5718 196
rect 5777 174 5836 196
rect 5895 174 5954 196
rect 5376 168 5954 174
rect 6544 174 6604 196
rect 6827 174 6887 196
rect 6945 174 7005 196
rect 7063 174 7123 196
rect 5376 133 5955 168
rect 6544 133 7123 174
rect 7712 174 7772 196
rect 7995 174 8055 196
rect 8113 174 8173 196
rect 8231 174 8291 196
rect 7712 133 8291 174
rect 8880 174 8940 196
rect 9163 174 9223 196
rect 9281 174 9341 196
rect 9399 174 9459 196
rect 8880 133 9459 174
<< polycont >>
rect 416 1314 450 1348
rect 1584 1314 1618 1348
rect 2752 1314 2786 1348
rect 3920 1314 3954 1348
rect 5094 1316 5128 1350
rect 6262 1316 6296 1350
rect 7430 1316 7464 1350
rect 8598 1316 8632 1350
rect 416 1206 450 1240
rect 1584 1206 1618 1240
rect 2752 1206 2786 1240
rect 3920 1206 3954 1240
rect 5094 1208 5128 1242
rect 6262 1208 6296 1242
rect 7430 1208 7464 1242
rect 8598 1208 8632 1242
rect 711 443 745 477
rect 1879 443 1913 477
rect 3047 443 3081 477
rect 4215 443 4249 477
rect 5389 445 5423 479
rect 6557 445 6591 479
rect 7725 445 7759 479
rect 8893 445 8927 479
<< locali >>
rect 1002 1426 1206 1438
rect 1002 1354 1034 1426
rect 1178 1354 1206 1426
rect 1002 1352 1064 1354
rect 1144 1352 1206 1354
rect 400 1314 416 1348
rect 450 1314 466 1348
rect 1002 1336 1206 1352
rect 2170 1426 2374 1438
rect 2170 1354 2202 1426
rect 2346 1354 2374 1426
rect 2170 1352 2232 1354
rect 2312 1352 2374 1354
rect 1568 1314 1584 1348
rect 1618 1314 1634 1348
rect 2170 1336 2374 1352
rect 3338 1426 3542 1438
rect 3338 1354 3370 1426
rect 3514 1354 3542 1426
rect 3338 1352 3400 1354
rect 3480 1352 3542 1354
rect 2736 1314 2752 1348
rect 2786 1314 2802 1348
rect 3338 1336 3542 1352
rect 4506 1426 4710 1438
rect 4506 1354 4538 1426
rect 4682 1354 4710 1426
rect 4506 1352 4568 1354
rect 4648 1352 4710 1354
rect 3904 1314 3920 1348
rect 3954 1314 3970 1348
rect 4506 1336 4710 1352
rect 5680 1428 5884 1440
rect 5680 1356 5712 1428
rect 5856 1356 5884 1428
rect 5680 1354 5742 1356
rect 5822 1354 5884 1356
rect 5078 1316 5094 1350
rect 5128 1316 5144 1350
rect 5680 1338 5884 1354
rect 6848 1428 7052 1440
rect 6848 1356 6880 1428
rect 7024 1356 7052 1428
rect 6848 1354 6910 1356
rect 6990 1354 7052 1356
rect 6246 1316 6262 1350
rect 6296 1316 6312 1350
rect 6848 1338 7052 1354
rect 8016 1428 8220 1440
rect 8016 1356 8048 1428
rect 8192 1356 8220 1428
rect 8016 1354 8078 1356
rect 8158 1354 8220 1356
rect 7414 1316 7430 1350
rect 7464 1316 7480 1350
rect 8016 1338 8220 1354
rect 9184 1428 9388 1440
rect 9184 1356 9216 1428
rect 9360 1356 9388 1428
rect 9184 1354 9246 1356
rect 9326 1354 9388 1356
rect 8582 1316 8598 1350
rect 8632 1316 8648 1350
rect 9184 1338 9388 1354
rect 400 1206 416 1240
rect 450 1206 466 1240
rect 1568 1206 1584 1240
rect 1618 1206 1634 1240
rect 2736 1206 2752 1240
rect 2786 1206 2802 1240
rect 3904 1206 3920 1240
rect 3954 1206 3970 1240
rect 5078 1208 5094 1242
rect 5128 1208 5144 1242
rect 6246 1208 6262 1242
rect 6296 1208 6312 1242
rect 7414 1208 7430 1242
rect 7464 1208 7480 1242
rect 8582 1208 8598 1242
rect 8632 1208 8648 1242
rect 695 443 711 477
rect 745 443 761 477
rect 1863 443 1879 477
rect 1913 443 1929 477
rect 3031 443 3047 477
rect 3081 443 3097 477
rect 4199 443 4215 477
rect 4249 443 4265 477
rect 5373 445 5389 479
rect 5423 445 5439 479
rect 6541 445 6557 479
rect 6591 445 6607 479
rect 7709 445 7725 479
rect 7759 445 7775 479
rect 8877 445 8893 479
rect 8927 445 8943 479
rect 560 86 702 98
rect 560 82 600 86
rect 666 82 702 86
rect 560 16 578 82
rect 696 16 702 82
rect 560 -10 702 16
rect 1728 86 1870 98
rect 1728 82 1768 86
rect 1834 82 1870 86
rect 1728 16 1746 82
rect 1864 16 1870 82
rect 1728 -10 1870 16
rect 2896 86 3038 98
rect 2896 82 2936 86
rect 3002 82 3038 86
rect 2896 16 2914 82
rect 3032 16 3038 82
rect 2896 -10 3038 16
rect 4064 86 4206 98
rect 4064 82 4104 86
rect 4170 82 4206 86
rect 4064 16 4082 82
rect 4200 16 4206 82
rect 4064 -10 4206 16
rect 5238 88 5380 100
rect 5238 84 5278 88
rect 5344 84 5380 88
rect 5238 18 5256 84
rect 5374 18 5380 84
rect 5238 -8 5380 18
rect 6406 88 6548 100
rect 6406 84 6446 88
rect 6512 84 6548 88
rect 6406 18 6424 84
rect 6542 18 6548 84
rect 6406 -8 6548 18
rect 7574 88 7716 100
rect 7574 84 7614 88
rect 7680 84 7716 88
rect 7574 18 7592 84
rect 7710 18 7716 84
rect 7574 -8 7716 18
rect 8742 88 8884 100
rect 8742 84 8782 88
rect 8848 84 8884 88
rect 8742 18 8760 84
rect 8878 18 8884 84
rect 8742 -8 8884 18
<< viali >>
rect 1064 1354 1144 1424
rect 1064 1352 1144 1354
rect 416 1314 450 1348
rect 2232 1354 2312 1424
rect 2232 1352 2312 1354
rect 1584 1314 1618 1348
rect 3400 1354 3480 1424
rect 3400 1352 3480 1354
rect 2752 1314 2786 1348
rect 4568 1354 4648 1424
rect 4568 1352 4648 1354
rect 3920 1314 3954 1348
rect 5742 1356 5822 1426
rect 5742 1354 5822 1356
rect 5094 1316 5128 1350
rect 6910 1356 6990 1426
rect 6910 1354 6990 1356
rect 6262 1316 6296 1350
rect 8078 1356 8158 1426
rect 8078 1354 8158 1356
rect 7430 1316 7464 1350
rect 9246 1356 9326 1426
rect 9246 1354 9326 1356
rect 8598 1316 8632 1350
rect 416 1206 450 1240
rect 1584 1206 1618 1240
rect 2752 1206 2786 1240
rect 3920 1206 3954 1240
rect 5094 1208 5128 1242
rect 6262 1208 6296 1242
rect 7430 1208 7464 1242
rect 8598 1208 8632 1242
rect 711 443 745 477
rect 1879 443 1913 477
rect 3047 443 3081 477
rect 4215 443 4249 477
rect 5389 445 5423 479
rect 6557 445 6591 479
rect 7725 445 7759 479
rect 8893 445 8927 479
rect 600 82 666 86
rect 600 16 666 82
rect 1768 82 1834 86
rect 1768 16 1834 82
rect 2936 82 3002 86
rect 2936 16 3002 82
rect 4104 82 4170 86
rect 4104 16 4170 82
rect 5278 84 5344 88
rect 5278 18 5344 84
rect 6446 84 6512 88
rect 6446 18 6512 84
rect 7614 84 7680 88
rect 7614 18 7680 84
rect 8782 84 8848 88
rect 8782 18 8848 84
<< metal1 >>
rect 366 1348 466 1450
rect 366 1314 416 1348
rect 450 1314 466 1348
rect 1052 1424 1156 1430
rect 1052 1352 1064 1424
rect 1144 1352 1156 1424
rect 1052 1346 1156 1352
rect 1534 1348 1634 1450
rect 366 1288 466 1314
rect 1087 1290 1122 1346
rect 1534 1314 1584 1348
rect 1618 1314 1634 1348
rect 2220 1424 2324 1430
rect 2220 1352 2232 1424
rect 2312 1352 2324 1424
rect 2220 1346 2324 1352
rect 2702 1348 2802 1450
rect 366 1240 466 1260
rect 366 1206 416 1240
rect 450 1206 466 1240
rect 366 1108 466 1206
rect 624 1249 894 1277
rect 624 1184 658 1249
rect 860 1184 894 1249
rect 978 1249 1248 1290
rect 1534 1288 1634 1314
rect 2255 1290 2290 1346
rect 2702 1314 2752 1348
rect 2786 1314 2802 1348
rect 3388 1424 3492 1430
rect 3388 1352 3400 1424
rect 3480 1352 3492 1424
rect 3388 1346 3492 1352
rect 3870 1348 3970 1450
rect 978 1180 1012 1249
rect 1214 1180 1248 1249
rect 1534 1240 1634 1260
rect 1534 1206 1584 1240
rect 1618 1206 1634 1240
rect 1534 1108 1634 1206
rect 1792 1249 2062 1277
rect 1792 1184 1826 1249
rect 2028 1184 2062 1249
rect 2146 1249 2416 1290
rect 2702 1288 2802 1314
rect 3423 1290 3458 1346
rect 3870 1314 3920 1348
rect 3954 1314 3970 1348
rect 4556 1424 4660 1430
rect 4556 1352 4568 1424
rect 4648 1352 4660 1424
rect 4556 1346 4660 1352
rect 5044 1350 5144 1452
rect 2146 1180 2180 1249
rect 2382 1180 2416 1249
rect 2702 1240 2802 1260
rect 2702 1206 2752 1240
rect 2786 1206 2802 1240
rect 2702 1108 2802 1206
rect 2960 1249 3230 1277
rect 2960 1184 2994 1249
rect 3196 1184 3230 1249
rect 3314 1249 3584 1290
rect 3870 1288 3970 1314
rect 4591 1290 4626 1346
rect 5044 1316 5094 1350
rect 5128 1316 5144 1350
rect 5730 1426 5834 1432
rect 5730 1354 5742 1426
rect 5822 1354 5834 1426
rect 5730 1348 5834 1354
rect 6212 1350 6312 1452
rect 5044 1290 5144 1316
rect 5765 1292 5800 1348
rect 6212 1316 6262 1350
rect 6296 1316 6312 1350
rect 6898 1426 7002 1432
rect 6898 1354 6910 1426
rect 6990 1354 7002 1426
rect 6898 1348 7002 1354
rect 7380 1350 7480 1452
rect 3314 1180 3348 1249
rect 3550 1180 3584 1249
rect 3870 1240 3970 1260
rect 3870 1206 3920 1240
rect 3954 1206 3970 1240
rect 3870 1108 3970 1206
rect 4128 1249 4398 1277
rect 4128 1184 4162 1249
rect 4364 1184 4398 1249
rect 4482 1249 4752 1290
rect 4482 1180 4516 1249
rect 4718 1180 4752 1249
rect 5044 1242 5144 1262
rect 5044 1208 5094 1242
rect 5128 1208 5144 1242
rect 5044 1110 5144 1208
rect 5302 1251 5572 1279
rect 5302 1186 5336 1251
rect 5538 1186 5572 1251
rect 5656 1251 5926 1292
rect 6212 1290 6312 1316
rect 6933 1292 6968 1348
rect 7380 1316 7430 1350
rect 7464 1316 7480 1350
rect 8066 1426 8170 1432
rect 8066 1354 8078 1426
rect 8158 1354 8170 1426
rect 8066 1348 8170 1354
rect 8548 1350 8648 1452
rect 5656 1182 5690 1251
rect 5892 1182 5926 1251
rect 6212 1242 6312 1262
rect 6212 1208 6262 1242
rect 6296 1208 6312 1242
rect 6212 1110 6312 1208
rect 6470 1251 6740 1279
rect 6470 1186 6504 1251
rect 6706 1186 6740 1251
rect 6824 1251 7094 1292
rect 7380 1290 7480 1316
rect 8101 1292 8136 1348
rect 8548 1316 8598 1350
rect 8632 1316 8648 1350
rect 9234 1426 9338 1432
rect 9234 1354 9246 1426
rect 9326 1354 9338 1426
rect 9234 1348 9338 1354
rect 6824 1182 6858 1251
rect 7060 1182 7094 1251
rect 7380 1242 7480 1262
rect 7380 1208 7430 1242
rect 7464 1208 7480 1242
rect 7380 1110 7480 1208
rect 7638 1251 7908 1279
rect 7638 1186 7672 1251
rect 7874 1186 7908 1251
rect 7992 1251 8262 1292
rect 8548 1290 8648 1316
rect 9269 1292 9304 1348
rect 7992 1182 8026 1251
rect 8228 1182 8262 1251
rect 8548 1242 8648 1262
rect 8548 1208 8598 1242
rect 8632 1208 8648 1242
rect 8548 1110 8648 1208
rect 8806 1251 9076 1279
rect 8806 1186 8840 1251
rect 9042 1186 9076 1251
rect 9160 1251 9430 1292
rect 9160 1182 9194 1251
rect 9396 1182 9430 1251
rect 506 745 540 816
rect 742 745 776 816
rect 506 717 776 745
rect 860 746 894 816
rect 1096 746 1130 816
rect 860 717 1130 746
rect 506 669 540 717
rect 506 639 569 669
rect 534 547 569 639
rect 1214 604 1248 788
rect 1674 745 1708 816
rect 1910 745 1944 816
rect 1674 717 1944 745
rect 2028 746 2062 816
rect 2264 746 2298 816
rect 2028 717 2298 746
rect 1674 669 1708 717
rect 1674 639 1737 669
rect 534 511 761 547
rect 534 364 569 511
rect 695 477 761 511
rect 695 443 711 477
rect 745 443 761 477
rect 1042 535 1139 586
rect 1214 550 1323 604
rect 1042 468 1099 535
rect 695 437 761 443
rect 936 432 1205 468
rect 936 394 969 432
rect 1172 397 1205 432
rect 1289 383 1323 550
rect 1702 547 1737 639
rect 2382 604 2416 788
rect 2842 745 2876 816
rect 3078 745 3112 816
rect 2842 717 3112 745
rect 3196 746 3230 816
rect 3432 746 3466 816
rect 3196 717 3466 746
rect 2842 669 2876 717
rect 2842 639 2905 669
rect 1702 511 1929 547
rect 1702 364 1737 511
rect 1863 477 1929 511
rect 1863 443 1879 477
rect 1913 443 1929 477
rect 2210 535 2307 586
rect 2382 550 2491 604
rect 2210 468 2267 535
rect 1863 437 1929 443
rect 2104 432 2373 468
rect 2104 394 2137 432
rect 2340 397 2373 432
rect 2457 383 2491 550
rect 2870 547 2905 639
rect 3550 604 3584 788
rect 4010 745 4044 816
rect 4246 745 4280 816
rect 4010 717 4280 745
rect 4364 746 4398 816
rect 4600 746 4634 816
rect 4364 717 4634 746
rect 4010 669 4044 717
rect 4010 639 4073 669
rect 2870 511 3097 547
rect 2870 364 2905 511
rect 3031 477 3097 511
rect 3031 443 3047 477
rect 3081 443 3097 477
rect 3378 535 3475 586
rect 3550 550 3659 604
rect 3378 468 3435 535
rect 3031 437 3097 443
rect 3272 432 3541 468
rect 3272 394 3305 432
rect 3508 397 3541 432
rect 3625 383 3659 550
rect 4038 547 4073 639
rect 4718 604 4752 788
rect 5184 747 5218 818
rect 5420 747 5454 818
rect 5184 719 5454 747
rect 5538 748 5572 818
rect 5774 748 5808 818
rect 5538 719 5808 748
rect 5184 671 5218 719
rect 5184 641 5247 671
rect 4038 511 4265 547
rect 4038 364 4073 511
rect 4199 477 4265 511
rect 4199 443 4215 477
rect 4249 443 4265 477
rect 4546 535 4643 586
rect 4718 550 4827 604
rect 4546 468 4603 535
rect 4199 437 4265 443
rect 4440 432 4709 468
rect 4440 394 4473 432
rect 4676 397 4709 432
rect 4793 383 4827 550
rect 5212 549 5247 641
rect 5892 606 5926 790
rect 6352 747 6386 818
rect 6588 747 6622 818
rect 6352 719 6622 747
rect 6706 748 6740 818
rect 6942 748 6976 818
rect 6706 719 6976 748
rect 6352 671 6386 719
rect 6352 641 6415 671
rect 5212 513 5439 549
rect 5212 366 5247 513
rect 5373 479 5439 513
rect 5373 445 5389 479
rect 5423 445 5439 479
rect 5720 537 5817 588
rect 5892 552 6001 606
rect 5720 470 5777 537
rect 5373 439 5439 445
rect 5614 434 5883 470
rect 5614 396 5647 434
rect 5850 399 5883 434
rect 5967 385 6001 552
rect 6380 549 6415 641
rect 7060 606 7094 790
rect 7520 747 7554 818
rect 7756 747 7790 818
rect 7520 719 7790 747
rect 7874 748 7908 818
rect 8110 748 8144 818
rect 7874 719 8144 748
rect 7520 671 7554 719
rect 7520 641 7583 671
rect 6380 513 6607 549
rect 6380 366 6415 513
rect 6541 479 6607 513
rect 6541 445 6557 479
rect 6591 445 6607 479
rect 6888 537 6985 588
rect 7060 552 7169 606
rect 6888 470 6945 537
rect 6541 439 6607 445
rect 6782 434 7051 470
rect 6782 396 6815 434
rect 7018 399 7051 434
rect 7135 385 7169 552
rect 7548 549 7583 641
rect 8228 606 8262 790
rect 8688 747 8722 818
rect 8924 747 8958 818
rect 8688 719 8958 747
rect 9042 748 9076 818
rect 9278 748 9312 818
rect 9042 719 9312 748
rect 8688 671 8722 719
rect 8688 641 8751 671
rect 7548 513 7775 549
rect 7548 366 7583 513
rect 7709 479 7775 513
rect 7709 445 7725 479
rect 7759 445 7775 479
rect 8056 537 8153 588
rect 8228 552 8337 606
rect 8056 470 8113 537
rect 7709 439 7775 445
rect 7950 434 8219 470
rect 7950 396 7983 434
rect 8186 399 8219 434
rect 8303 385 8337 552
rect 8716 549 8751 641
rect 9396 606 9430 790
rect 8716 513 8943 549
rect 8716 366 8751 513
rect 8877 479 8943 513
rect 8877 445 8893 479
rect 8927 445 8943 479
rect 9224 537 9321 588
rect 9396 552 9505 606
rect 9224 470 9281 537
rect 8877 439 8943 445
rect 9118 434 9387 470
rect 9118 396 9151 434
rect 9354 399 9387 434
rect 9471 385 9505 552
rect 787 249 952 337
rect 1955 249 2120 337
rect 3123 249 3288 337
rect 4291 249 4456 337
rect 5465 251 5630 339
rect 6633 251 6798 339
rect 7801 251 7966 339
rect 8969 251 9134 339
rect 416 165 450 218
rect 652 165 686 214
rect 416 126 686 165
rect 1053 166 1086 213
rect 1289 166 1322 213
rect 1053 130 1322 166
rect 1584 165 1618 218
rect 1820 165 1854 214
rect 1584 126 1854 165
rect 2221 166 2254 213
rect 2457 166 2490 213
rect 2221 130 2490 166
rect 2752 165 2786 218
rect 2988 165 3022 214
rect 2752 126 3022 165
rect 3389 166 3422 213
rect 3625 166 3658 213
rect 3389 130 3658 166
rect 3920 165 3954 218
rect 4156 165 4190 214
rect 3920 126 4190 165
rect 4557 166 4590 213
rect 4793 166 4826 213
rect 4557 130 4826 166
rect 5094 167 5128 220
rect 5330 167 5364 216
rect 5094 128 5364 167
rect 5731 168 5764 215
rect 5967 168 6000 215
rect 5731 132 6000 168
rect 6262 167 6296 220
rect 6498 167 6532 216
rect 6262 128 6532 167
rect 6899 168 6932 215
rect 7135 168 7168 215
rect 6899 132 7168 168
rect 7430 167 7464 220
rect 7666 167 7700 216
rect 7430 128 7700 167
rect 8067 168 8100 215
rect 8303 168 8336 215
rect 8067 132 8336 168
rect 8598 167 8632 220
rect 8834 167 8868 216
rect 8598 128 8868 167
rect 9235 168 9268 215
rect 9471 168 9504 215
rect 9235 132 9504 168
rect 616 98 650 126
rect 1784 98 1818 126
rect 2952 98 2986 126
rect 4120 98 4154 126
rect 5294 100 5328 128
rect 6462 100 6496 128
rect 7630 100 7664 128
rect 8798 100 8832 128
rect 594 86 672 98
rect 594 16 600 86
rect 666 16 672 86
rect 594 4 672 16
rect 1762 86 1840 98
rect 1762 16 1768 86
rect 1834 16 1840 86
rect 1762 4 1840 16
rect 2930 86 3008 98
rect 2930 16 2936 86
rect 3002 16 3008 86
rect 2930 4 3008 16
rect 4098 86 4176 98
rect 4098 16 4104 86
rect 4170 16 4176 86
rect 4098 4 4176 16
rect 5272 88 5350 100
rect 5272 18 5278 88
rect 5344 18 5350 88
rect 5272 6 5350 18
rect 6440 88 6518 100
rect 6440 18 6446 88
rect 6512 18 6518 88
rect 6440 6 6518 18
rect 7608 88 7686 100
rect 7608 18 7614 88
rect 7680 18 7686 88
rect 7608 6 7686 18
rect 8776 88 8854 100
rect 8776 18 8782 88
rect 8848 18 8854 88
rect 8776 6 8854 18
<< via1 >>
rect 1078 1353 1130 1405
rect 2246 1353 2298 1405
rect 3414 1353 3466 1405
rect 4582 1353 4634 1405
rect 5756 1355 5808 1407
rect 6924 1355 6976 1407
rect 8092 1355 8144 1407
rect 9260 1355 9312 1407
rect 607 29 659 81
rect 1775 29 1827 81
rect 2943 29 2995 81
rect 4111 29 4163 81
rect 5285 31 5337 83
rect 6453 31 6505 83
rect 7621 31 7673 83
rect 8789 31 8841 83
<< metal2 >>
rect 1056 1426 1146 1436
rect 1056 1325 1146 1335
rect 2224 1426 2314 1436
rect 2224 1325 2314 1335
rect 3392 1426 3482 1436
rect 3392 1325 3482 1335
rect 4560 1426 4650 1436
rect 4560 1325 4650 1335
rect 5734 1428 5824 1438
rect 5734 1327 5824 1337
rect 6902 1428 6992 1438
rect 6902 1327 6992 1337
rect 8070 1428 8160 1438
rect 8070 1327 8160 1337
rect 9238 1428 9328 1438
rect 9238 1327 9328 1337
rect 591 99 681 109
rect 591 -2 681 8
rect 1759 99 1849 109
rect 1759 -2 1849 8
rect 2927 99 3017 109
rect 2927 -2 3017 8
rect 4095 99 4185 109
rect 4095 -2 4185 8
rect 5269 101 5359 111
rect 5269 0 5359 10
rect 6437 101 6527 111
rect 6437 0 6527 10
rect 7605 101 7695 111
rect 7605 0 7695 10
rect 8773 101 8863 111
rect 8773 0 8863 10
<< via2 >>
rect 1056 1405 1146 1426
rect 1056 1353 1078 1405
rect 1078 1353 1130 1405
rect 1130 1353 1146 1405
rect 1056 1335 1146 1353
rect 2224 1405 2314 1426
rect 2224 1353 2246 1405
rect 2246 1353 2298 1405
rect 2298 1353 2314 1405
rect 2224 1335 2314 1353
rect 3392 1405 3482 1426
rect 3392 1353 3414 1405
rect 3414 1353 3466 1405
rect 3466 1353 3482 1405
rect 3392 1335 3482 1353
rect 4560 1405 4650 1426
rect 4560 1353 4582 1405
rect 4582 1353 4634 1405
rect 4634 1353 4650 1405
rect 4560 1335 4650 1353
rect 5734 1407 5824 1428
rect 5734 1355 5756 1407
rect 5756 1355 5808 1407
rect 5808 1355 5824 1407
rect 5734 1337 5824 1355
rect 6902 1407 6992 1428
rect 6902 1355 6924 1407
rect 6924 1355 6976 1407
rect 6976 1355 6992 1407
rect 6902 1337 6992 1355
rect 8070 1407 8160 1428
rect 8070 1355 8092 1407
rect 8092 1355 8144 1407
rect 8144 1355 8160 1407
rect 8070 1337 8160 1355
rect 9238 1407 9328 1428
rect 9238 1355 9260 1407
rect 9260 1355 9312 1407
rect 9312 1355 9328 1407
rect 9238 1337 9328 1355
rect 591 81 681 99
rect 591 29 607 81
rect 607 29 659 81
rect 659 29 681 81
rect 591 8 681 29
rect 1759 81 1849 99
rect 1759 29 1775 81
rect 1775 29 1827 81
rect 1827 29 1849 81
rect 1759 8 1849 29
rect 2927 81 3017 99
rect 2927 29 2943 81
rect 2943 29 2995 81
rect 2995 29 3017 81
rect 2927 8 3017 29
rect 4095 81 4185 99
rect 4095 29 4111 81
rect 4111 29 4163 81
rect 4163 29 4185 81
rect 4095 8 4185 29
rect 5269 83 5359 101
rect 5269 31 5285 83
rect 5285 31 5337 83
rect 5337 31 5359 83
rect 5269 10 5359 31
rect 6437 83 6527 101
rect 6437 31 6453 83
rect 6453 31 6505 83
rect 6505 31 6527 83
rect 6437 10 6527 31
rect 7605 83 7695 101
rect 7605 31 7621 83
rect 7621 31 7673 83
rect 7673 31 7695 83
rect 7605 10 7695 31
rect 8773 83 8863 101
rect 8773 31 8789 83
rect 8789 31 8841 83
rect 8841 31 8863 83
rect 8773 10 8863 31
<< metal3 >>
rect 1028 1320 1038 1440
rect 1160 1320 1170 1440
rect 2196 1426 2338 1440
rect 2196 1335 2224 1426
rect 2314 1335 2338 1426
rect 2196 1320 2338 1335
rect 3364 1426 3506 1440
rect 3364 1335 3392 1426
rect 3482 1335 3506 1426
rect 3364 1320 3506 1335
rect 4532 1426 4674 1440
rect 4532 1335 4560 1426
rect 4650 1335 4674 1426
rect 4532 1320 4674 1335
rect 5706 1428 5848 1442
rect 5706 1337 5734 1428
rect 5824 1337 5848 1428
rect 5706 1322 5848 1337
rect 6874 1428 7016 1442
rect 6874 1337 6902 1428
rect 6992 1337 7016 1428
rect 6874 1322 7016 1337
rect 8042 1428 8184 1442
rect 8042 1337 8070 1428
rect 8160 1337 8184 1428
rect 8042 1322 8184 1337
rect 9210 1428 9352 1442
rect 9210 1337 9238 1428
rect 9328 1337 9352 1428
rect 9210 1322 9352 1337
rect 571 -2 581 109
rect 691 -2 701 109
rect 1739 -2 1749 109
rect 1859 -2 1869 109
rect 2907 -2 2917 109
rect 3027 -2 3037 109
rect 4075 -2 4085 109
rect 4195 -2 4205 109
rect 5249 0 5259 111
rect 5369 0 5379 111
rect 6417 0 6427 111
rect 6537 0 6547 111
rect 7585 0 7595 111
rect 7705 0 7715 111
rect 8753 0 8763 111
rect 8873 0 8883 111
<< via3 >>
rect 1038 1426 1160 1440
rect 1038 1335 1056 1426
rect 1056 1335 1146 1426
rect 1146 1335 1160 1426
rect 1038 1320 1160 1335
rect 2240 1348 2304 1412
rect 3408 1348 3472 1412
rect 4578 1350 4642 1414
rect 5750 1350 5814 1414
rect 6918 1348 6982 1412
rect 8086 1350 8150 1414
rect 9254 1350 9318 1414
rect 581 99 691 109
rect 581 8 591 99
rect 591 8 681 99
rect 681 8 691 99
rect 581 -2 691 8
rect 1749 99 1859 109
rect 1749 8 1759 99
rect 1759 8 1849 99
rect 1849 8 1859 99
rect 1749 -2 1859 8
rect 2917 99 3027 109
rect 2917 8 2927 99
rect 2927 8 3017 99
rect 3017 8 3027 99
rect 2917 -2 3027 8
rect 4085 99 4195 109
rect 4085 8 4095 99
rect 4095 8 4185 99
rect 4185 8 4195 99
rect 4085 -2 4195 8
rect 5259 101 5369 111
rect 5259 10 5269 101
rect 5269 10 5359 101
rect 5359 10 5369 101
rect 5259 0 5369 10
rect 6427 101 6537 111
rect 6427 10 6437 101
rect 6437 10 6527 101
rect 6527 10 6537 101
rect 6427 0 6537 10
rect 7595 101 7705 111
rect 7595 10 7605 101
rect 7605 10 7695 101
rect 7695 10 7705 101
rect 7595 0 7705 10
rect 8763 101 8873 111
rect 8763 10 8773 101
rect 8773 10 8863 101
rect 8863 10 8873 101
rect 8763 0 8873 10
<< metal4 >>
rect 458 1440 9450 1506
rect 458 1320 1038 1440
rect 1160 1414 9450 1440
rect 1160 1412 4578 1414
rect 1160 1348 2240 1412
rect 2304 1348 3408 1412
rect 3472 1350 4578 1412
rect 4642 1350 5750 1414
rect 5814 1412 8086 1414
rect 5814 1350 6918 1412
rect 3472 1348 6918 1350
rect 6982 1350 8086 1412
rect 8150 1350 9254 1414
rect 9318 1350 9450 1414
rect 6982 1348 9450 1350
rect 1160 1320 9450 1348
rect 458 1310 9450 1320
rect 5258 111 5370 112
rect 5258 110 5259 111
rect 458 109 5259 110
rect 458 -2 581 109
rect 691 -2 1749 109
rect 1859 -2 2917 109
rect 3027 -2 4085 109
rect 4195 0 5259 109
rect 5369 110 5370 111
rect 6426 111 6538 112
rect 6426 110 6427 111
rect 5369 0 6427 110
rect 6537 110 6538 111
rect 7594 111 7706 112
rect 7594 110 7595 111
rect 6537 0 7595 110
rect 7705 110 7706 111
rect 8762 111 8874 112
rect 8762 110 8763 111
rect 7705 0 8763 110
rect 8873 110 8874 111
rect 8873 0 9556 110
rect 4195 -2 9556 0
rect 458 -86 9556 -2
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_0
timestamp 1736524280
transform 1 0 610 0 1 302
box -206 -126 206 126
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_1
timestamp 1736524280
transform 1 0 1778 0 1 304
box -206 -126 206 126
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_2
timestamp 1736524280
transform 1 0 2946 0 1 304
box -206 -126 206 126
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_3
timestamp 1736524280
transform 1 0 4114 0 1 304
box -206 -126 206 126
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_4
timestamp 1736524280
transform 1 0 5288 0 1 304
box -206 -126 206 126
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_5
timestamp 1736524280
transform 1 0 6456 0 1 304
box -206 -126 206 126
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_6
timestamp 1736524280
transform 1 0 7624 0 1 306
box -206 -126 206 126
use sky130_fd_pr__nfet_01v8_DH4BC5  sky130_fd_pr__nfet_01v8_DH4BC5_7
timestamp 1736524280
transform 1 0 8792 0 1 306
box -206 -126 206 126
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_0
timestamp 1736524280
transform 1 0 2045 0 1 988
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_1
timestamp 1736524280
transform 1 0 877 0 1 988
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_2
timestamp 1736524280
transform 1 0 3213 0 1 986
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_3
timestamp 1736524280
transform 1 0 4381 0 1 988
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_4
timestamp 1736524280
transform 1 0 5555 0 1 990
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_5
timestamp 1736524280
transform 1 0 6723 0 1 988
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_6
timestamp 1736524280
transform 1 0 7891 0 1 990
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_82VCJ4  sky130_fd_pr__pfet_01v8_82VCJ4_7
timestamp 1736524280
transform 1 0 9059 0 1 988
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_0
timestamp 1736524280
transform 1 0 4634 0 1 304
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_1
timestamp 1736524280
transform 1 0 5806 0 1 300
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_2
timestamp 1736524280
transform 1 0 1130 0 1 298
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_3
timestamp 1736524280
transform 1 0 3465 0 1 304
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_4
timestamp 1736524280
transform 1 0 2297 0 1 304
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_5
timestamp 1736524280
transform 1 0 6975 0 1 299
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_6
timestamp 1736524280
transform 1 0 8143 0 1 299
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_PCXB2D  sky130_fd_pr__pfet_01v8_PCXB2D_7
timestamp 1736524280
transform 1 0 9311 0 1 300
box -242 -162 242 162
<< labels >>
flabel metal4 4764 -86 5044 110 1 FreeSerif 800 0 0 0 VSS
port 2 n
flabel metal1 366 1368 466 1450 1 FreeSerif 480 0 0 0 B[0]
port 3 n
flabel metal1 366 1108 458 1190 1 FreeSerif 480 0 0 0 A[0]
port 4 n
flabel metal1 1534 1108 1626 1190 1 FreeSerif 480 0 0 0 A[1]
port 5 n
flabel metal1 2702 1108 2794 1190 1 FreeSerif 480 0 0 0 A[2]
port 6 n
flabel metal1 3870 1108 3962 1190 1 FreeSerif 480 0 0 0 A[3]
port 7 n
flabel metal1 5044 1110 5136 1192 1 FreeSerif 480 0 0 0 A[4]
port 8 n
flabel metal1 6212 1110 6304 1192 1 FreeSerif 480 0 0 0 A[5]
port 9 n
flabel metal1 7380 1110 7472 1192 1 FreeSerif 480 0 0 0 A[6]
port 10 n
flabel metal1 8548 1110 8640 1192 1 FreeSerif 480 0 0 0 A[7]
port 11 n
flabel metal1 9224 538 9320 588 1 FreeSerif 480 0 0 0 Y[7]
port 12 n
flabel metal1 8056 538 8152 588 1 FreeSerif 480 0 0 0 Y[6]
port 13 n
flabel metal1 6888 538 6984 588 1 FreeSerif 480 0 0 0 Y[5]
port 14 n
flabel metal1 5720 538 5816 588 1 FreeSerif 480 0 0 0 Y[4]
port 15 n
flabel metal1 4546 536 4642 586 1 FreeSerif 480 0 0 0 Y[3]
port 16 n
flabel metal1 3378 536 3474 586 1 FreeSerif 480 0 0 0 Y[2]
port 17 n
flabel metal1 2210 536 2306 586 1 FreeSerif 480 0 0 0 Y[1]
port 18 n
flabel metal1 1042 536 1138 586 1 FreeSerif 480 0 0 0 Y[0]
port 19 n
flabel metal1 1534 1368 1634 1450 1 FreeSerif 480 0 0 0 B[1]
port 20 n
flabel metal1 2702 1368 2802 1450 1 FreeSerif 480 0 0 0 B[2]
port 21 n
flabel metal1 3870 1368 3970 1450 1 FreeSerif 480 0 0 0 B[3]
port 22 n
flabel metal1 5044 1370 5144 1452 1 FreeSerif 480 0 0 0 B[4]
port 23 n
flabel metal1 6212 1370 6312 1452 1 FreeSerif 480 0 0 0 B[5]
port 24 n
flabel metal1 7380 1370 7480 1452 1 FreeSerif 480 0 0 0 B[6]
port 25 n
flabel metal1 8548 1370 8648 1452 1 FreeSerif 480 0 0 0 B[7]
port 26 n
flabel metal4 4786 1366 4910 1454 1 FreeSerif 800 0 0 0 VDD
port 27 n
<< end >>
